// Benchmark "mem_ctrl" written by ABC on Thu Sep 14 22:43:54 2023

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_,
    new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_,
    new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_,
    new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_,
    new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_,
    new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_,
    new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_,
    new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_,
    new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_,
    new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_,
    new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_,
    new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_,
    new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_,
    new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4463_, new_n4464_, new_n4465_, new_n4466_,
    new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_,
    new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_,
    new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_,
    new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_,
    new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_,
    new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_,
    new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_,
    new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_,
    new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5371_, new_n5372_,
    new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_,
    new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_,
    new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_,
    new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_,
    new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5530_,
    new_n5531_, new_n5532_, new_n5533_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_,
    new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_,
    new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_,
    new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_,
    new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_,
    new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_,
    new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_,
    new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_,
    new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_,
    new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_,
    new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_,
    new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_,
    new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_,
    new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_,
    new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_,
    new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_,
    new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5991_, new_n5992_,
    new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_,
    new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_,
    new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_,
    new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_,
    new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_,
    new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_,
    new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_,
    new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_,
    new_n6041_, new_n6042_, new_n6043_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6100_, new_n6101_, new_n6102_,
    new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_,
    new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_,
    new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_,
    new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_,
    new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_,
    new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_,
    new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_,
    new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_,
    new_n6151_, new_n6152_, new_n6153_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6209_, new_n6210_, new_n6211_, new_n6212_,
    new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_,
    new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_,
    new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_,
    new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_,
    new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_,
    new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_,
    new_n6261_, new_n6262_, new_n6263_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6302_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6339_, new_n6340_, new_n6341_, new_n6343_, new_n6345_,
    new_n6347_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6356_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6577_, new_n6581_, new_n6584_,
    new_n6595_, new_n6596_, new_n6604_, new_n6606_, new_n6643_, new_n6648_,
    new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_,
    new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_,
    new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_,
    new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6675_,
    new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_,
    new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_,
    new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_,
    new_n6695_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6742_, new_n6743_, new_n6744_,
    new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_,
    new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_,
    new_n6757_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6796_, new_n6797_, new_n6803_,
    new_n6815_, new_n6816_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6845_, new_n6878_,
    new_n6894_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6976_, new_n6977_,
    new_n6983_, new_n6989_, new_n6991_, new_n7013_, new_n7014_, new_n7015_,
    new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7082_, new_n7083_,
    new_n7084_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7110_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7132_, new_n7134_,
    new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_,
    new_n7141_, new_n7142_, new_n7143_, new_n7147_, new_n7148_, new_n7149_,
    new_n7150_, new_n7152_, new_n7153_, new_n7154_, new_n7164_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_,
    new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_,
    new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_,
    new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_,
    new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_,
    new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_,
    new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_,
    new_n7303_, new_n7304_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_,
    new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_,
    new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_,
    new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_,
    new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_,
    new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_,
    new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_,
    new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_,
    new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_,
    new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_,
    new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_,
    new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_,
    new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_,
    new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_,
    new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_,
    new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_,
    new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_,
    new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_,
    new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_,
    new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_,
    new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_,
    new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_,
    new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_,
    new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_,
    new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_,
    new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_,
    new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_,
    new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_,
    new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_,
    new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_,
    new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_,
    new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_,
    new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_,
    new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_,
    new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_,
    new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_,
    new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_,
    new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_,
    new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_,
    new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_,
    new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_,
    new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_,
    new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_,
    new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_,
    new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_,
    new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_,
    new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_,
    new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_,
    new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_,
    new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_,
    new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_,
    new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_,
    new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_,
    new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_,
    new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_,
    new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_,
    new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_,
    new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_,
    new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_,
    new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_,
    new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_,
    new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_,
    new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_,
    new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_,
    new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_,
    new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_,
    new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_,
    new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_,
    new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_,
    new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_,
    new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_,
    new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_,
    new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_,
    new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_,
    new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_,
    new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_,
    new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8274_,
    new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_,
    new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_,
    new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8318_,
    new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_,
    new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_,
    new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_,
    new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_,
    new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_,
    new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_,
    new_n8373_, new_n8374_, new_n8375_, new_n8377_, new_n8378_, new_n8379_,
    new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_,
    new_n8386_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_,
    new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_,
    new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_,
    new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8447_,
    new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_,
    new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_,
    new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_,
    new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_,
    new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_,
    new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_,
    new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_,
    new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_,
    new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8569_, new_n8570_,
    new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_,
    new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_,
    new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_,
    new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_,
    new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_,
    new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_,
    new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_,
    new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_,
    new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_,
    new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_,
    new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_,
    new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_,
    new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_,
    new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_,
    new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_,
    new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_,
    new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_,
    new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_,
    new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_,
    new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_,
    new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_,
    new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_,
    new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_,
    new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_,
    new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_,
    new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_,
    new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_,
    new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8739_,
    new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_,
    new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8875_, new_n8876_, new_n8877_, new_n8878_,
    new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_,
    new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_,
    new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_,
    new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_,
    new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_,
    new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_,
    new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_,
    new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_,
    new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_,
    new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8985_,
    new_n8986_, new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_,
    new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9148_,
    new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_,
    new_n9155_, new_n9156_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9173_, new_n9174_, new_n9176_,
    new_n9177_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9185_, new_n9186_, new_n9188_, new_n9189_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9205_, new_n9206_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9219_, new_n9221_,
    new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9279_, new_n9280_,
    new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_,
    new_n9287_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9427_, new_n9428_,
    new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_,
    new_n9435_, new_n9436_, new_n9437_, new_n9439_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_,
    new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_,
    new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_,
    new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_,
    new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_,
    new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_,
    new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_,
    new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_,
    new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_,
    new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_,
    new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_,
    new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_,
    new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_,
    new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_,
    new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_,
    new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_,
    new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_,
    new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_,
    new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_,
    new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_,
    new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_,
    new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_,
    new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_,
    new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_,
    new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_,
    new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_,
    new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_,
    new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_,
    new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_,
    new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_,
    new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_,
    new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_,
    new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_,
    new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_,
    new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_,
    new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_,
    new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_,
    new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_,
    new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_,
    new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_,
    new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_,
    new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_,
    new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_,
    new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_,
    new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_,
    new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_,
    new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_,
    new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_,
    new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_,
    new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_,
    new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_,
    new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_,
    new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_,
    new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_,
    new_n9785_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9796_, new_n9798_, new_n9799_, new_n9800_,
    new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_,
    new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_,
    new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_,
    new_n9819_, new_n9820_, new_n9825_, new_n9826_, new_n9827_, new_n9859_,
    new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_,
    new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_,
    new_n9873_, new_n9875_, new_n9876_, new_n9877_, new_n9903_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_,
    new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_,
    new_n9975_, new_n9976_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9992_, new_n9993_,
    new_n9994_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10021_, new_n10022_,
    new_n10023_, new_n10040_, new_n10046_, new_n10047_, new_n10057_,
    new_n10062_, new_n10063_, new_n10064_, new_n10065_, new_n10066_,
    new_n10067_, new_n10068_, new_n10069_, new_n10070_, new_n10071_,
    new_n10072_, new_n10073_, new_n10074_, new_n10075_, new_n10076_,
    new_n10078_, new_n10079_, new_n10080_, new_n10081_, new_n10082_,
    new_n10083_, new_n10084_, new_n10085_, new_n10086_, new_n10087_,
    new_n10088_, new_n10089_, new_n10090_, new_n10091_, new_n10092_,
    new_n10093_, new_n10094_, new_n10095_, new_n10096_, new_n10097_,
    new_n10098_, new_n10099_, new_n10100_, new_n10101_, new_n10102_,
    new_n10103_, new_n10104_, new_n10105_, new_n10106_, new_n10107_,
    new_n10108_, new_n10109_, new_n10110_, new_n10111_, new_n10112_,
    new_n10113_, new_n10114_, new_n10115_, new_n10116_, new_n10117_,
    new_n10118_, new_n10119_, new_n10120_, new_n10121_, new_n10122_,
    new_n10123_, new_n10124_, new_n10125_, new_n10126_, new_n10127_,
    new_n10128_, new_n10129_, new_n10130_, new_n10131_, new_n10132_,
    new_n10133_, new_n10134_, new_n10135_, new_n10136_, new_n10137_,
    new_n10138_, new_n10139_, new_n10140_, new_n10141_, new_n10142_,
    new_n10143_, new_n10144_, new_n10145_, new_n10146_, new_n10147_,
    new_n10148_, new_n10149_, new_n10150_, new_n10151_, new_n10152_,
    new_n10153_, new_n10154_, new_n10155_, new_n10156_, new_n10157_,
    new_n10158_, new_n10159_, new_n10160_, new_n10161_, new_n10162_,
    new_n10163_, new_n10164_, new_n10165_, new_n10166_, new_n10167_,
    new_n10168_, new_n10169_, new_n10170_, new_n10171_, new_n10172_,
    new_n10173_, new_n10174_, new_n10175_, new_n10176_, new_n10177_,
    new_n10178_, new_n10179_, new_n10180_, new_n10181_, new_n10182_,
    new_n10183_, new_n10184_, new_n10185_, new_n10186_, new_n10187_,
    new_n10188_, new_n10189_, new_n10190_, new_n10191_, new_n10192_,
    new_n10193_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10200_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10217_, new_n10218_, new_n10223_, new_n10226_,
    new_n10227_, new_n10228_, new_n10230_, new_n10231_, new_n10232_,
    new_n10233_, new_n10234_, new_n10235_, new_n10237_, new_n10238_,
    new_n10239_, new_n10240_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10258_, new_n10259_, new_n10260_, new_n10262_,
    new_n10264_, new_n10265_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10286_,
    new_n10287_, new_n10289_, new_n10290_, new_n10291_, new_n10292_,
    new_n10293_, new_n10294_, new_n10295_, new_n10297_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10304_,
    new_n10305_, new_n10306_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10321_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10331_, new_n10332_,
    new_n10333_, new_n10334_, new_n10335_, new_n10336_, new_n10338_,
    new_n10339_, new_n10340_, new_n10341_, new_n10343_, new_n10344_,
    new_n10345_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10391_,
    new_n10392_, new_n10393_, new_n10394_, new_n10395_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10405_, new_n10406_, new_n10407_, new_n10408_,
    new_n10409_, new_n10410_, new_n10411_, new_n10412_, new_n10413_,
    new_n10414_, new_n10415_, new_n10416_, new_n10417_, new_n10418_,
    new_n10419_, new_n10420_, new_n10421_, new_n10422_, new_n10423_,
    new_n10424_, new_n10425_, new_n10426_, new_n10427_, new_n10428_,
    new_n10429_, new_n10430_, new_n10431_, new_n10432_, new_n10433_,
    new_n10434_, new_n10435_, new_n10436_, new_n10437_, new_n10438_,
    new_n10439_, new_n10440_, new_n10441_, new_n10442_, new_n10443_,
    new_n10444_, new_n10445_, new_n10446_, new_n10447_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10454_, new_n10455_,
    new_n10457_, new_n10458_, new_n10459_, new_n10461_, new_n10462_,
    new_n10463_, new_n10464_, new_n10465_, new_n10466_, new_n10467_,
    new_n10468_, new_n10469_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10493_, new_n10494_, new_n10495_, new_n10496_, new_n10497_,
    new_n10499_, new_n10500_, new_n10501_, new_n10502_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10570_, new_n10571_, new_n10572_,
    new_n10573_, new_n10574_, new_n10575_, new_n10576_, new_n10577_,
    new_n10578_, new_n10579_, new_n10580_, new_n10581_, new_n10582_,
    new_n10584_, new_n10585_, new_n10586_, new_n10587_, new_n10588_,
    new_n10589_, new_n10590_, new_n10591_, new_n10592_, new_n10593_,
    new_n10594_, new_n10595_, new_n10596_, new_n10597_, new_n10598_,
    new_n10599_, new_n10600_, new_n10601_, new_n10602_, new_n10603_,
    new_n10604_, new_n10605_, new_n10606_, new_n10607_, new_n10608_,
    new_n10609_, new_n10610_, new_n10611_, new_n10612_, new_n10613_,
    new_n10614_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10628_, new_n10629_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10701_,
    new_n10702_, new_n10703_, new_n10704_, new_n10705_, new_n10706_,
    new_n10707_, new_n10708_, new_n10709_, new_n10710_, new_n10711_,
    new_n10712_, new_n10713_, new_n10714_, new_n10715_, new_n10716_,
    new_n10717_, new_n10718_, new_n10719_, new_n10720_, new_n10721_,
    new_n10722_, new_n10723_, new_n10724_, new_n10725_, new_n10726_,
    new_n10727_, new_n10728_, new_n10729_, new_n10730_, new_n10731_,
    new_n10732_, new_n10733_, new_n10734_, new_n10735_, new_n10736_,
    new_n10737_, new_n10738_, new_n10739_, new_n10740_, new_n10741_,
    new_n10742_, new_n10743_, new_n10744_, new_n10745_, new_n10746_,
    new_n10747_, new_n10748_, new_n10749_, new_n10750_, new_n10751_,
    new_n10752_, new_n10753_, new_n10754_, new_n10755_, new_n10756_,
    new_n10757_, new_n10758_, new_n10759_, new_n10760_, new_n10761_,
    new_n10762_, new_n10763_, new_n10764_, new_n10765_, new_n10766_,
    new_n10767_, new_n10768_, new_n10769_, new_n10770_, new_n10771_,
    new_n10772_, new_n10773_, new_n10774_, new_n10775_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10794_, new_n10795_, new_n10796_,
    new_n10797_, new_n10798_, new_n10799_, new_n10800_, new_n10801_,
    new_n10802_, new_n10803_, new_n10804_, new_n10805_, new_n10806_,
    new_n10807_, new_n10808_, new_n10809_, new_n10810_, new_n10811_,
    new_n10812_, new_n10813_, new_n10814_, new_n10815_, new_n10816_,
    new_n10817_, new_n10818_, new_n10819_, new_n10820_, new_n10821_,
    new_n10822_, new_n10823_, new_n10824_, new_n10825_, new_n10826_,
    new_n10827_, new_n10828_, new_n10829_, new_n10830_, new_n10831_,
    new_n10832_, new_n10833_, new_n10834_, new_n10835_, new_n10836_,
    new_n10837_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10858_, new_n10859_, new_n10860_, new_n10861_, new_n10862_,
    new_n10863_, new_n10864_, new_n10865_, new_n10866_, new_n10867_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10873_,
    new_n10874_, new_n10875_, new_n10876_, new_n10877_, new_n10878_,
    new_n10879_, new_n10880_, new_n10881_, new_n10882_, new_n10883_,
    new_n10884_, new_n10885_, new_n10886_, new_n10887_, new_n10888_,
    new_n10889_, new_n10890_, new_n10891_, new_n10892_, new_n10893_,
    new_n10894_, new_n10895_, new_n10896_, new_n10897_, new_n10898_,
    new_n10899_, new_n10900_, new_n10901_, new_n10902_, new_n10903_,
    new_n10904_, new_n10905_, new_n10906_, new_n10907_, new_n10908_,
    new_n10909_, new_n10910_, new_n10911_, new_n10912_, new_n10913_,
    new_n10914_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10921_, new_n10922_, new_n10923_,
    new_n10924_, new_n10925_, new_n10926_, new_n10927_, new_n10928_,
    new_n10929_, new_n10930_, new_n10931_, new_n10932_, new_n10933_,
    new_n10934_, new_n10935_, new_n10936_, new_n10937_, new_n10938_,
    new_n10939_, new_n10940_, new_n10941_, new_n10942_, new_n10943_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10958_, new_n10961_, new_n10962_, new_n10963_,
    new_n10964_, new_n10965_, new_n10966_, new_n10967_, new_n10968_,
    new_n10969_, new_n10970_, new_n10971_, new_n10972_, new_n10973_,
    new_n10974_, new_n10975_, new_n10976_, new_n10977_, new_n10978_,
    new_n10979_, new_n10980_, new_n10981_, new_n10982_, new_n10983_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11005_, new_n11006_, new_n11007_, new_n11008_,
    new_n11009_, new_n11010_, new_n11011_, new_n11012_, new_n11013_,
    new_n11014_, new_n11015_, new_n11016_, new_n11017_, new_n11018_,
    new_n11019_, new_n11020_, new_n11021_, new_n11022_, new_n11023_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11030_, new_n11031_, new_n11032_, new_n11033_,
    new_n11034_, new_n11035_, new_n11036_, new_n11037_, new_n11038_,
    new_n11039_, new_n11040_, new_n11041_, new_n11042_, new_n11043_,
    new_n11044_, new_n11045_, new_n11046_, new_n11047_, new_n11048_,
    new_n11049_, new_n11050_, new_n11051_, new_n11052_, new_n11053_,
    new_n11054_, new_n11055_, new_n11056_, new_n11057_, new_n11058_,
    new_n11059_, new_n11060_, new_n11061_, new_n11062_, new_n11063_,
    new_n11064_, new_n11065_, new_n11066_, new_n11067_, new_n11068_,
    new_n11069_, new_n11070_, new_n11071_, new_n11072_, new_n11073_,
    new_n11074_, new_n11075_, new_n11076_, new_n11077_, new_n11078_,
    new_n11079_, new_n11080_, new_n11081_, new_n11082_, new_n11083_,
    new_n11084_, new_n11085_, new_n11086_, new_n11087_, new_n11088_,
    new_n11089_, new_n11090_, new_n11091_, new_n11092_, new_n11093_,
    new_n11094_, new_n11095_, new_n11096_, new_n11097_, new_n11098_,
    new_n11099_, new_n11100_, new_n11101_, new_n11102_, new_n11103_,
    new_n11104_, new_n11105_, new_n11106_, new_n11107_, new_n11108_,
    new_n11109_, new_n11110_, new_n11111_, new_n11112_, new_n11113_,
    new_n11114_, new_n11115_, new_n11116_, new_n11117_, new_n11118_,
    new_n11119_, new_n11120_, new_n11121_, new_n11122_, new_n11123_,
    new_n11124_, new_n11125_, new_n11126_, new_n11127_, new_n11128_,
    new_n11129_, new_n11130_, new_n11131_, new_n11132_, new_n11133_,
    new_n11134_, new_n11135_, new_n11136_, new_n11137_, new_n11138_,
    new_n11139_, new_n11140_, new_n11141_, new_n11142_, new_n11143_,
    new_n11144_, new_n11145_, new_n11146_, new_n11147_, new_n11148_,
    new_n11149_, new_n11150_, new_n11151_, new_n11152_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11509_, new_n11510_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11555_, new_n11556_, new_n11557_, new_n11558_,
    new_n11559_, new_n11560_, new_n11561_, new_n11562_, new_n11563_,
    new_n11564_, new_n11565_, new_n11566_, new_n11567_, new_n11568_,
    new_n11569_, new_n11570_, new_n11571_, new_n11572_, new_n11573_,
    new_n11574_, new_n11575_, new_n11576_, new_n11577_, new_n11578_,
    new_n11579_, new_n11580_, new_n11581_, new_n11582_, new_n11583_,
    new_n11584_, new_n11585_, new_n11586_, new_n11587_, new_n11588_,
    new_n11589_, new_n11590_, new_n11591_, new_n11592_, new_n11593_,
    new_n11594_, new_n11595_, new_n11596_, new_n11597_, new_n11598_,
    new_n11599_, new_n11600_, new_n11601_, new_n11602_, new_n11603_,
    new_n11604_, new_n11605_, new_n11606_, new_n11607_, new_n11608_,
    new_n11609_, new_n11610_, new_n11611_, new_n11612_, new_n11613_,
    new_n11614_, new_n11615_, new_n11616_, new_n11617_, new_n11618_,
    new_n11619_, new_n11620_, new_n11621_, new_n11622_, new_n11623_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11631_, new_n11632_, new_n11633_,
    new_n11634_, new_n11635_, new_n11636_, new_n11637_, new_n11638_,
    new_n11639_, new_n11640_, new_n11641_, new_n11642_, new_n11643_,
    new_n11644_, new_n11645_, new_n11646_, new_n11647_, new_n11648_,
    new_n11649_, new_n11650_, new_n11651_, new_n11652_, new_n11653_,
    new_n11654_, new_n11655_, new_n11656_, new_n11657_, new_n11658_,
    new_n11659_, new_n11660_, new_n11661_, new_n11662_, new_n11663_,
    new_n11664_, new_n11665_, new_n11666_, new_n11667_, new_n11668_,
    new_n11669_, new_n11670_, new_n11671_, new_n11672_, new_n11673_,
    new_n11674_, new_n11675_, new_n11676_, new_n11677_, new_n11678_,
    new_n11679_, new_n11680_, new_n11681_, new_n11682_, new_n11683_,
    new_n11684_, new_n11685_, new_n11686_, new_n11687_, new_n11688_,
    new_n11689_, new_n11690_, new_n11691_, new_n11692_, new_n11693_,
    new_n11694_, new_n11695_, new_n11696_, new_n11697_, new_n11698_,
    new_n11699_, new_n11700_, new_n11701_, new_n11702_, new_n11703_,
    new_n11704_, new_n11705_, new_n11706_, new_n11707_, new_n11708_,
    new_n11709_, new_n11710_, new_n11711_, new_n11712_, new_n11713_,
    new_n11714_, new_n11715_, new_n11716_, new_n11717_, new_n11718_,
    new_n11719_, new_n11720_, new_n11721_, new_n11722_, new_n11723_,
    new_n11724_, new_n11725_, new_n11726_, new_n11727_, new_n11728_,
    new_n11729_, new_n11730_, new_n11731_, new_n11732_, new_n11733_,
    new_n11734_, new_n11735_, new_n11736_, new_n11737_, new_n11738_,
    new_n11739_, new_n11740_, new_n11741_, new_n11742_, new_n11743_,
    new_n11744_, new_n11745_, new_n11746_, new_n11747_, new_n11748_,
    new_n11749_, new_n11750_, new_n11751_, new_n11752_, new_n11753_,
    new_n11754_, new_n11755_, new_n11756_, new_n11757_, new_n11758_,
    new_n11759_, new_n11760_, new_n11761_, new_n11762_, new_n11763_,
    new_n11764_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11771_, new_n11772_, new_n11773_,
    new_n11774_, new_n11775_, new_n11776_, new_n11777_, new_n11778_,
    new_n11779_, new_n11780_, new_n11781_, new_n11782_, new_n11783_,
    new_n11784_, new_n11785_, new_n11786_, new_n11787_, new_n11788_,
    new_n11789_, new_n11790_, new_n11791_, new_n11792_, new_n11793_,
    new_n11794_, new_n11795_, new_n11796_, new_n11797_, new_n11798_,
    new_n11799_, new_n11800_, new_n11801_, new_n11802_, new_n11803_,
    new_n11804_, new_n11805_, new_n11806_, new_n11807_, new_n11808_,
    new_n11809_, new_n11810_, new_n11811_, new_n11812_, new_n11813_,
    new_n11814_, new_n11815_, new_n11816_, new_n11817_, new_n11818_,
    new_n11819_, new_n11820_, new_n11821_, new_n11822_, new_n11823_,
    new_n11824_, new_n11825_, new_n11826_, new_n11827_, new_n11828_,
    new_n11829_, new_n11830_, new_n11831_, new_n11832_, new_n11833_,
    new_n11834_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11856_, new_n11857_, new_n11858_, new_n11859_,
    new_n11860_, new_n11861_, new_n11862_, new_n11863_, new_n11864_,
    new_n11865_, new_n11866_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11903_, new_n11904_,
    new_n11905_, new_n11906_, new_n11907_, new_n11908_, new_n11909_,
    new_n11910_, new_n11911_, new_n11912_, new_n11913_, new_n11914_,
    new_n11915_, new_n11916_, new_n11917_, new_n11918_, new_n11919_,
    new_n11920_, new_n11921_, new_n11922_, new_n11923_, new_n11924_,
    new_n11925_, new_n11926_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11932_, new_n11933_, new_n11934_,
    new_n11935_, new_n11936_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11947_, new_n11948_, new_n11949_,
    new_n11950_, new_n11951_, new_n11952_, new_n11953_, new_n11954_,
    new_n11955_, new_n11956_, new_n11957_, new_n11958_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11970_, new_n11971_, new_n11972_, new_n11973_, new_n11974_,
    new_n11975_, new_n11976_, new_n11977_, new_n11978_, new_n11979_,
    new_n11980_, new_n11981_, new_n11982_, new_n11983_, new_n11984_,
    new_n11985_, new_n11986_, new_n11987_, new_n11988_, new_n11989_,
    new_n11990_, new_n11991_, new_n11992_, new_n11993_, new_n11994_,
    new_n11995_, new_n11996_, new_n11997_, new_n11998_, new_n11999_,
    new_n12000_, new_n12001_, new_n12002_, new_n12003_, new_n12004_,
    new_n12005_, new_n12006_, new_n12007_, new_n12008_, new_n12009_,
    new_n12010_, new_n12011_, new_n12012_, new_n12013_, new_n12014_,
    new_n12015_, new_n12016_, new_n12017_, new_n12018_, new_n12019_,
    new_n12020_, new_n12021_, new_n12022_, new_n12023_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12074_, new_n12105_, new_n12106_,
    new_n12107_, new_n12108_, new_n12109_, new_n12110_, new_n12111_,
    new_n12112_, new_n12113_, new_n12114_, new_n12115_, new_n12116_,
    new_n12117_, new_n12118_, new_n12119_, new_n12120_, new_n12121_,
    new_n12122_, new_n12123_, new_n12124_, new_n12125_, new_n12126_,
    new_n12127_, new_n12128_, new_n12129_, new_n12130_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12161_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12327_, new_n12328_, new_n12329_, new_n12330_, new_n12331_,
    new_n12332_, new_n12333_, new_n12334_, new_n12335_, new_n12336_,
    new_n12337_, new_n12338_, new_n12339_, new_n12340_, new_n12341_,
    new_n12342_, new_n12343_, new_n12344_, new_n12345_, new_n12346_,
    new_n12347_, new_n12348_, new_n12349_, new_n12350_, new_n12351_,
    new_n12352_, new_n12353_, new_n12354_, new_n12355_, new_n12356_,
    new_n12357_, new_n12358_, new_n12359_, new_n12360_, new_n12361_,
    new_n12362_, new_n12363_, new_n12364_, new_n12365_, new_n12366_,
    new_n12367_, new_n12368_, new_n12369_, new_n12370_, new_n12371_,
    new_n12372_, new_n12373_, new_n12374_, new_n12375_, new_n12376_,
    new_n12377_, new_n12378_, new_n12379_, new_n12380_, new_n12381_,
    new_n12382_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12519_, new_n12520_, new_n12521_,
    new_n12522_, new_n12523_, new_n12524_, new_n12525_, new_n12526_,
    new_n12527_, new_n12528_, new_n12529_, new_n12530_, new_n12531_,
    new_n12532_, new_n12533_, new_n12534_, new_n12535_, new_n12536_,
    new_n12537_, new_n12538_, new_n12539_, new_n12540_, new_n12541_,
    new_n12542_, new_n12543_, new_n12544_, new_n12545_, new_n12546_,
    new_n12547_, new_n12548_, new_n12549_, new_n12550_, new_n12551_,
    new_n12552_, new_n12553_, new_n12554_, new_n12555_, new_n12556_,
    new_n12557_, new_n12558_, new_n12559_, new_n12560_, new_n12562_,
    new_n12563_, new_n12564_, new_n12565_, new_n12566_, new_n12567_,
    new_n12568_, new_n12569_, new_n12570_, new_n12571_, new_n12572_,
    new_n12573_, new_n12574_, new_n12575_, new_n12576_, new_n12577_,
    new_n12578_, new_n12579_, new_n12580_, new_n12581_, new_n12582_,
    new_n12583_, new_n12584_, new_n12585_, new_n12586_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12593_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12617_, new_n12618_,
    new_n12619_, new_n12620_, new_n12621_, new_n12622_, new_n12623_,
    new_n12624_, new_n12625_, new_n12626_, new_n12627_, new_n12628_,
    new_n12629_, new_n12630_, new_n12631_, new_n12632_, new_n12633_,
    new_n12634_, new_n12635_, new_n12636_, new_n12637_, new_n12638_,
    new_n12639_, new_n12640_, new_n12641_, new_n12642_, new_n12643_,
    new_n12644_, new_n12645_, new_n12646_, new_n12647_, new_n12648_,
    new_n12649_, new_n12650_, new_n12651_, new_n12652_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12683_,
    new_n12684_, new_n12685_, new_n12686_, new_n12687_, new_n12688_,
    new_n12689_, new_n12690_, new_n12691_, new_n12692_, new_n12693_,
    new_n12694_, new_n12695_, new_n12696_, new_n12697_, new_n12698_,
    new_n12699_, new_n12700_, new_n12701_, new_n12702_, new_n12703_,
    new_n12704_, new_n12705_, new_n12706_, new_n12707_, new_n12708_,
    new_n12709_, new_n12710_, new_n12711_, new_n12712_, new_n12713_,
    new_n12714_, new_n12715_, new_n12716_, new_n12717_, new_n12718_,
    new_n12719_, new_n12720_, new_n12721_, new_n12722_, new_n12723_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13010_, new_n13011_,
    new_n13012_, new_n13013_, new_n13014_, new_n13015_, new_n13016_,
    new_n13017_, new_n13018_, new_n13019_, new_n13020_, new_n13021_,
    new_n13022_, new_n13023_, new_n13024_, new_n13025_, new_n13026_,
    new_n13027_, new_n13028_, new_n13029_, new_n13030_, new_n13031_,
    new_n13032_, new_n13033_, new_n13034_, new_n13035_, new_n13036_,
    new_n13037_, new_n13038_, new_n13039_, new_n13040_, new_n13041_,
    new_n13043_, new_n13044_, new_n13045_, new_n13046_, new_n13047_,
    new_n13048_, new_n13049_, new_n13050_, new_n13051_, new_n13052_,
    new_n13053_, new_n13054_, new_n13055_, new_n13056_, new_n13057_,
    new_n13058_, new_n13059_, new_n13060_, new_n13061_, new_n13062_,
    new_n13063_, new_n13064_, new_n13065_, new_n13066_, new_n13067_,
    new_n13068_, new_n13069_, new_n13070_, new_n13071_, new_n13072_,
    new_n13073_, new_n13074_, new_n13075_, new_n13076_, new_n13077_,
    new_n13078_, new_n13079_, new_n13080_, new_n13081_, new_n13082_,
    new_n13083_, new_n13084_, new_n13085_, new_n13086_, new_n13087_,
    new_n13088_, new_n13089_, new_n13090_, new_n13091_, new_n13092_,
    new_n13093_, new_n13094_, new_n13095_, new_n13096_, new_n13097_,
    new_n13098_, new_n13099_, new_n13100_, new_n13101_, new_n13102_,
    new_n13103_, new_n13104_, new_n13105_, new_n13106_, new_n13107_,
    new_n13108_, new_n13109_, new_n13110_, new_n13111_, new_n13112_,
    new_n13113_, new_n13114_, new_n13115_, new_n13116_, new_n13117_,
    new_n13118_, new_n13119_, new_n13120_, new_n13121_, new_n13122_,
    new_n13123_, new_n13124_, new_n13125_, new_n13126_, new_n13127_,
    new_n13128_, new_n13129_, new_n13130_, new_n13131_, new_n13132_,
    new_n13133_, new_n13134_, new_n13135_, new_n13136_, new_n13137_,
    new_n13138_, new_n13139_, new_n13140_, new_n13141_, new_n13142_,
    new_n13143_, new_n13144_, new_n13145_, new_n13146_, new_n13147_,
    new_n13148_, new_n13149_, new_n13150_, new_n13151_, new_n13152_,
    new_n13153_, new_n13154_, new_n13155_, new_n13156_, new_n13157_,
    new_n13158_, new_n13159_, new_n13160_, new_n13161_, new_n13162_,
    new_n13163_, new_n13164_, new_n13165_, new_n13166_, new_n13167_,
    new_n13168_, new_n13169_, new_n13170_, new_n13171_, new_n13172_,
    new_n13173_, new_n13174_, new_n13175_, new_n13176_, new_n13177_,
    new_n13178_, new_n13179_, new_n13180_, new_n13181_, new_n13182_,
    new_n13183_, new_n13184_, new_n13185_, new_n13186_, new_n13187_,
    new_n13188_, new_n13189_, new_n13190_, new_n13191_, new_n13192_,
    new_n13193_, new_n13194_, new_n13195_, new_n13196_, new_n13197_,
    new_n13198_, new_n13199_, new_n13200_, new_n13201_, new_n13202_,
    new_n13203_, new_n13204_, new_n13205_, new_n13206_, new_n13207_,
    new_n13208_, new_n13209_, new_n13210_, new_n13211_, new_n13212_,
    new_n13213_, new_n13218_, new_n13219_, new_n13220_, new_n13221_,
    new_n13222_, new_n13223_, new_n13224_, new_n13225_, new_n13226_,
    new_n13227_, new_n13228_, new_n13229_, new_n13230_, new_n13231_,
    new_n13232_, new_n13233_, new_n13234_, new_n13235_, new_n13236_,
    new_n13237_, new_n13238_, new_n13239_, new_n13240_, new_n13241_,
    new_n13242_, new_n13243_, new_n13244_, new_n13245_, new_n13246_,
    new_n13247_, new_n13248_, new_n13249_, new_n13250_, new_n13251_,
    new_n13252_, new_n13253_, new_n13254_, new_n13255_, new_n13256_,
    new_n13257_, new_n13258_, new_n13259_, new_n13260_, new_n13261_,
    new_n13262_, new_n13263_, new_n13264_, new_n13265_, new_n13266_,
    new_n13267_, new_n13268_, new_n13269_, new_n13270_, new_n13271_,
    new_n13272_, new_n13273_, new_n13274_, new_n13275_, new_n13276_,
    new_n13277_, new_n13278_, new_n13279_, new_n13280_, new_n13281_,
    new_n13282_, new_n13283_, new_n13284_, new_n13285_, new_n13286_,
    new_n13287_, new_n13288_, new_n13289_, new_n13290_, new_n13291_,
    new_n13292_, new_n13293_, new_n13294_, new_n13295_, new_n13296_,
    new_n13297_, new_n13298_, new_n13299_, new_n13300_, new_n13301_,
    new_n13302_, new_n13303_, new_n13304_, new_n13305_, new_n13306_,
    new_n13307_, new_n13308_, new_n13309_, new_n13310_, new_n13311_,
    new_n13312_, new_n13313_, new_n13314_, new_n13315_, new_n13316_,
    new_n13317_, new_n13318_, new_n13319_, new_n13320_, new_n13321_,
    new_n13322_, new_n13323_, new_n13324_, new_n13325_, new_n13326_,
    new_n13327_, new_n13328_, new_n13329_, new_n13330_, new_n13331_,
    new_n13332_, new_n13333_, new_n13334_, new_n13335_, new_n13336_,
    new_n13337_, new_n13338_, new_n13339_, new_n13340_, new_n13341_,
    new_n13342_, new_n13343_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13350_, new_n13351_,
    new_n13352_, new_n13353_, new_n13354_, new_n13355_, new_n13356_,
    new_n13357_, new_n13358_, new_n13359_, new_n13360_, new_n13361_,
    new_n13362_, new_n13363_, new_n13364_, new_n13365_, new_n13366_,
    new_n13367_, new_n13368_, new_n13369_, new_n13370_, new_n13371_,
    new_n13372_, new_n13373_, new_n13374_, new_n13375_, new_n13376_,
    new_n13377_, new_n13378_, new_n13379_, new_n13380_, new_n13381_,
    new_n13382_, new_n13383_, new_n13384_, new_n13385_, new_n13386_,
    new_n13387_, new_n13388_, new_n13389_, new_n13390_, new_n13391_,
    new_n13392_, new_n13393_, new_n13394_, new_n13395_, new_n13396_,
    new_n13397_, new_n13398_, new_n13399_, new_n13400_, new_n13401_,
    new_n13402_, new_n13403_, new_n13404_, new_n13405_, new_n13406_,
    new_n13407_, new_n13408_, new_n13409_, new_n13410_, new_n13411_,
    new_n13412_, new_n13413_, new_n13414_, new_n13415_, new_n13416_,
    new_n13417_, new_n13418_, new_n13419_, new_n13420_, new_n13421_,
    new_n13422_, new_n13423_, new_n13424_, new_n13425_, new_n13426_,
    new_n13427_, new_n13428_, new_n13429_, new_n13430_, new_n13431_,
    new_n13432_, new_n13433_, new_n13434_, new_n13435_, new_n13436_,
    new_n13437_, new_n13438_, new_n13439_, new_n13440_, new_n13441_,
    new_n13442_, new_n13443_, new_n13444_, new_n13445_, new_n13446_,
    new_n13447_, new_n13448_, new_n13449_, new_n13450_, new_n13451_,
    new_n13452_, new_n13453_, new_n13454_, new_n13455_, new_n13456_,
    new_n13457_, new_n13458_, new_n13459_, new_n13460_, new_n13461_,
    new_n13462_, new_n13463_, new_n13464_, new_n13465_, new_n13466_,
    new_n13467_, new_n13468_, new_n13469_, new_n13470_, new_n13471_,
    new_n13472_, new_n13473_, new_n13474_, new_n13475_, new_n13476_,
    new_n13477_, new_n13478_, new_n13479_, new_n13480_, new_n13481_,
    new_n13482_, new_n13483_, new_n13484_, new_n13485_, new_n13486_,
    new_n13487_, new_n13488_, new_n13489_, new_n13490_, new_n13491_,
    new_n13492_, new_n13493_, new_n13494_, new_n13495_, new_n13496_,
    new_n13497_, new_n13498_, new_n13499_, new_n13500_, new_n13501_,
    new_n13502_, new_n13503_, new_n13504_, new_n13505_, new_n13506_,
    new_n13507_, new_n13508_, new_n13509_, new_n13510_, new_n13511_,
    new_n13512_, new_n13513_, new_n13514_, new_n13515_, new_n13516_,
    new_n13517_, new_n13518_, new_n13519_, new_n13520_, new_n13521_,
    new_n13522_, new_n13523_, new_n13524_, new_n13525_, new_n13526_,
    new_n13527_, new_n13528_, new_n13529_, new_n13530_, new_n13531_,
    new_n13532_, new_n13533_, new_n13534_, new_n13535_, new_n13536_,
    new_n13537_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13963_, new_n13964_,
    new_n13965_, new_n13966_, new_n13967_, new_n13968_, new_n13969_,
    new_n13970_, new_n13971_, new_n13972_, new_n13973_, new_n13974_,
    new_n13975_, new_n13976_, new_n13977_, new_n13978_, new_n13979_,
    new_n13980_, new_n13981_, new_n13982_, new_n13983_, new_n13984_,
    new_n13985_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14302_,
    new_n14303_, new_n14304_, new_n14305_, new_n14306_, new_n14307_,
    new_n14308_, new_n14309_, new_n14310_, new_n14311_, new_n14312_,
    new_n14313_, new_n14314_, new_n14315_, new_n14316_, new_n14317_,
    new_n14318_, new_n14319_, new_n14320_, new_n14321_, new_n14322_,
    new_n14323_, new_n14324_, new_n14325_, new_n14326_, new_n14327_,
    new_n14328_, new_n14329_, new_n14330_, new_n14331_, new_n14332_,
    new_n14333_, new_n14334_, new_n14335_, new_n14336_, new_n14337_,
    new_n14338_, new_n14339_, new_n14340_, new_n14341_, new_n14342_,
    new_n14343_, new_n14344_, new_n14345_, new_n14346_, new_n14347_,
    new_n14348_, new_n14349_, new_n14350_, new_n14351_, new_n14352_,
    new_n14353_, new_n14354_, new_n14355_, new_n14356_, new_n14357_,
    new_n14358_, new_n14359_, new_n14360_, new_n14361_, new_n14362_,
    new_n14363_, new_n14364_, new_n14365_, new_n14366_, new_n14367_,
    new_n14368_, new_n14369_, new_n14370_, new_n14371_, new_n14372_,
    new_n14373_, new_n14374_, new_n14375_, new_n14376_, new_n14377_,
    new_n14378_, new_n14379_, new_n14380_, new_n14381_, new_n14382_,
    new_n14383_, new_n14384_, new_n14385_, new_n14386_, new_n14387_,
    new_n14388_, new_n14389_, new_n14390_, new_n14391_, new_n14392_,
    new_n14393_, new_n14394_, new_n14395_, new_n14396_, new_n14397_,
    new_n14398_, new_n14399_, new_n14400_, new_n14401_, new_n14402_,
    new_n14403_, new_n14404_, new_n14405_, new_n14406_, new_n14407_,
    new_n14408_, new_n14409_, new_n14410_, new_n14411_, new_n14412_,
    new_n14413_, new_n14414_, new_n14415_, new_n14416_, new_n14417_,
    new_n14418_, new_n14419_, new_n14420_, new_n14421_, new_n14422_,
    new_n14423_, new_n14424_, new_n14425_, new_n14426_, new_n14427_,
    new_n14428_, new_n14429_, new_n14430_, new_n14431_, new_n14432_,
    new_n14433_, new_n14434_, new_n14435_, new_n14436_, new_n14437_,
    new_n14438_, new_n14439_, new_n14441_, new_n14442_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14456_,
    new_n14457_, new_n14458_, new_n14459_, new_n14460_, new_n14461_,
    new_n14462_, new_n14463_, new_n14464_, new_n14465_, new_n14466_,
    new_n14467_, new_n14468_, new_n14469_, new_n14470_, new_n14471_,
    new_n14472_, new_n14473_, new_n14474_, new_n14475_, new_n14476_,
    new_n14477_, new_n14478_, new_n14479_, new_n14480_, new_n14481_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14487_, new_n14488_, new_n14489_, new_n14490_, new_n14491_,
    new_n14492_, new_n14493_, new_n14494_, new_n14495_, new_n14496_,
    new_n14497_, new_n14498_, new_n14499_, new_n14500_, new_n14501_,
    new_n14502_, new_n14503_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14522_, new_n14523_, new_n14524_, new_n14525_, new_n14526_,
    new_n14527_, new_n14528_, new_n14529_, new_n14530_, new_n14531_,
    new_n14532_, new_n14533_, new_n14534_, new_n14535_, new_n14536_,
    new_n14537_, new_n14538_, new_n14539_, new_n14540_, new_n14541_,
    new_n14542_, new_n14543_, new_n14544_, new_n14545_, new_n14546_,
    new_n14547_, new_n14548_, new_n14549_, new_n14550_, new_n14551_,
    new_n14552_, new_n14553_, new_n14554_, new_n14555_, new_n14556_,
    new_n14557_, new_n14558_, new_n14559_, new_n14560_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14575_, new_n14576_, new_n14577_, new_n14578_, new_n14579_,
    new_n14580_, new_n14581_, new_n14582_, new_n14583_, new_n14584_,
    new_n14585_, new_n14586_, new_n14587_, new_n14588_, new_n14589_,
    new_n14590_, new_n14591_, new_n14592_, new_n14593_, new_n14594_,
    new_n14595_, new_n14596_, new_n14597_, new_n14598_, new_n14599_,
    new_n14600_, new_n14601_, new_n14602_, new_n14603_, new_n14604_,
    new_n14605_, new_n14606_, new_n14607_, new_n14608_, new_n14609_,
    new_n14613_, new_n14614_, new_n14615_, new_n14616_, new_n14617_,
    new_n14618_, new_n14619_, new_n14620_, new_n14621_, new_n14622_,
    new_n14623_, new_n14624_, new_n14625_, new_n14626_, new_n14627_,
    new_n14628_, new_n14629_, new_n14630_, new_n14631_, new_n14632_,
    new_n14633_, new_n14634_, new_n14635_, new_n14636_, new_n14637_,
    new_n14638_, new_n14639_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14676_, new_n14677_,
    new_n14678_, new_n14679_, new_n14680_, new_n14681_, new_n14682_,
    new_n14683_, new_n14684_, new_n14685_, new_n14686_, new_n14687_,
    new_n14688_, new_n14689_, new_n14690_, new_n14691_, new_n14692_,
    new_n14693_, new_n14694_, new_n14695_, new_n14696_, new_n14697_,
    new_n14698_, new_n14699_, new_n14700_, new_n14701_, new_n14702_,
    new_n14703_, new_n14704_, new_n14705_, new_n14706_, new_n14707_,
    new_n14708_, new_n14709_, new_n14710_, new_n14711_, new_n14712_,
    new_n14713_, new_n14714_, new_n14715_, new_n14716_, new_n14717_,
    new_n14718_, new_n14719_, new_n14720_, new_n14721_, new_n14722_,
    new_n14723_, new_n14724_, new_n14725_, new_n14726_, new_n14727_,
    new_n14728_, new_n14729_, new_n14730_, new_n14731_, new_n14732_,
    new_n14733_, new_n14734_, new_n14735_, new_n14736_, new_n14737_,
    new_n14738_, new_n14739_, new_n14740_, new_n14741_, new_n14742_,
    new_n14743_, new_n14744_, new_n14745_, new_n14746_, new_n14747_,
    new_n14748_, new_n14749_, new_n14750_, new_n14751_, new_n14752_,
    new_n14753_, new_n14754_, new_n14755_, new_n14756_, new_n14757_,
    new_n14758_, new_n14759_, new_n14760_, new_n14761_, new_n14762_,
    new_n14763_, new_n14764_, new_n14765_, new_n14766_, new_n14767_,
    new_n14768_, new_n14769_, new_n14770_, new_n14771_, new_n14772_,
    new_n14773_, new_n14774_, new_n14775_, new_n14776_, new_n14777_,
    new_n14778_, new_n14779_, new_n14780_, new_n14781_, new_n14782_,
    new_n14783_, new_n14784_, new_n14785_, new_n14786_, new_n14787_,
    new_n14788_, new_n14789_, new_n14790_, new_n14791_, new_n14792_,
    new_n14793_, new_n14794_, new_n14795_, new_n14796_, new_n14797_,
    new_n14798_, new_n14799_, new_n14800_, new_n14801_, new_n14802_,
    new_n14803_, new_n14804_, new_n14805_, new_n14806_, new_n14807_,
    new_n14808_, new_n14809_, new_n14810_, new_n14811_, new_n14812_,
    new_n14813_, new_n14814_, new_n14815_, new_n14816_, new_n14817_,
    new_n14818_, new_n14819_, new_n14820_, new_n14821_, new_n14822_,
    new_n14823_, new_n14824_, new_n14825_, new_n14826_, new_n14827_,
    new_n14828_, new_n14829_, new_n14830_, new_n14832_, new_n14833_,
    new_n14834_, new_n14835_, new_n14836_, new_n14837_, new_n14838_,
    new_n14839_, new_n14840_, new_n14841_, new_n14842_, new_n14843_,
    new_n14844_, new_n14845_, new_n14846_, new_n14847_, new_n14848_,
    new_n14849_, new_n14850_, new_n14851_, new_n14852_, new_n14853_,
    new_n14854_, new_n14855_, new_n14856_, new_n14857_, new_n14858_,
    new_n14859_, new_n14860_, new_n14861_, new_n14862_, new_n14863_,
    new_n14864_, new_n14865_, new_n14866_, new_n14867_, new_n14868_,
    new_n14869_, new_n14870_, new_n14871_, new_n14872_, new_n14873_,
    new_n14874_, new_n14875_, new_n14876_, new_n14877_, new_n14878_,
    new_n14879_, new_n14880_, new_n14881_, new_n14882_, new_n14883_,
    new_n14884_, new_n14885_, new_n14886_, new_n14887_, new_n14888_,
    new_n14889_, new_n14890_, new_n14891_, new_n14892_, new_n14893_,
    new_n14894_, new_n14895_, new_n14896_, new_n14897_, new_n14898_,
    new_n14899_, new_n14900_, new_n14901_, new_n14902_, new_n14903_,
    new_n14904_, new_n14905_, new_n14906_, new_n14907_, new_n14908_,
    new_n14909_, new_n14910_, new_n14911_, new_n14912_, new_n14913_,
    new_n14914_, new_n14915_, new_n14916_, new_n14917_, new_n14918_,
    new_n14919_, new_n14920_, new_n14921_, new_n14922_, new_n14923_,
    new_n14924_, new_n14925_, new_n14926_, new_n14927_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14951_, new_n14952_, new_n14953_,
    new_n14954_, new_n14955_, new_n14956_, new_n14957_, new_n14958_,
    new_n14959_, new_n14960_, new_n14961_, new_n14962_, new_n14963_,
    new_n14964_, new_n14965_, new_n14966_, new_n14967_, new_n14968_,
    new_n14969_, new_n14970_, new_n14971_, new_n14972_, new_n14973_,
    new_n14974_, new_n14975_, new_n14976_, new_n14977_, new_n14978_,
    new_n14979_, new_n14980_, new_n14981_, new_n14982_, new_n14983_,
    new_n14984_, new_n14985_, new_n14986_, new_n14987_, new_n14988_,
    new_n14989_, new_n14990_, new_n14991_, new_n14992_, new_n14993_,
    new_n14994_, new_n14995_, new_n14996_, new_n14997_, new_n14998_,
    new_n14999_, new_n15000_, new_n15001_, new_n15002_, new_n15003_,
    new_n15004_, new_n15005_, new_n15006_, new_n15007_, new_n15008_,
    new_n15009_, new_n15010_, new_n15011_, new_n15012_, new_n15013_,
    new_n15014_, new_n15015_, new_n15016_, new_n15017_, new_n15018_,
    new_n15019_, new_n15020_, new_n15021_, new_n15022_, new_n15023_,
    new_n15024_, new_n15025_, new_n15026_, new_n15027_, new_n15028_,
    new_n15029_, new_n15030_, new_n15031_, new_n15032_, new_n15033_,
    new_n15034_, new_n15035_, new_n15036_, new_n15037_, new_n15038_,
    new_n15039_, new_n15040_, new_n15041_, new_n15042_, new_n15043_,
    new_n15044_, new_n15045_, new_n15046_, new_n15047_, new_n15048_,
    new_n15049_, new_n15050_, new_n15051_, new_n15052_, new_n15053_,
    new_n15054_, new_n15055_, new_n15056_, new_n15057_, new_n15058_,
    new_n15059_, new_n15060_, new_n15061_, new_n15062_, new_n15063_,
    new_n15064_, new_n15065_, new_n15066_, new_n15067_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15087_, new_n15088_,
    new_n15089_, new_n15090_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15097_, new_n15098_,
    new_n15099_, new_n15100_, new_n15101_, new_n15102_, new_n15103_,
    new_n15104_, new_n15105_, new_n15106_, new_n15107_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15112_, new_n15113_,
    new_n15114_, new_n15115_, new_n15116_, new_n15117_, new_n15118_,
    new_n15119_, new_n15120_, new_n15121_, new_n15122_, new_n15123_,
    new_n15124_, new_n15125_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15138_,
    new_n15139_, new_n15140_, new_n15141_, new_n15142_, new_n15143_,
    new_n15144_, new_n15145_, new_n15146_, new_n15147_, new_n15148_,
    new_n15149_, new_n15150_, new_n15151_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15157_, new_n15158_,
    new_n15159_, new_n15160_, new_n15161_, new_n15162_, new_n15163_,
    new_n15164_, new_n15165_, new_n15166_, new_n15167_, new_n15168_,
    new_n15169_, new_n15170_, new_n15171_, new_n15172_, new_n15173_,
    new_n15174_, new_n15175_, new_n15176_, new_n15177_, new_n15178_,
    new_n15179_, new_n15180_, new_n15181_, new_n15182_, new_n15183_,
    new_n15184_, new_n15185_, new_n15186_, new_n15187_, new_n15188_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15199_, new_n15200_, new_n15201_, new_n15202_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15214_, new_n15215_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15232_, new_n15233_,
    new_n15234_, new_n15235_, new_n15236_, new_n15237_, new_n15238_,
    new_n15239_, new_n15240_, new_n15241_, new_n15242_, new_n15243_,
    new_n15244_, new_n15245_, new_n15246_, new_n15247_, new_n15248_,
    new_n15249_, new_n15251_, new_n15252_, new_n15253_, new_n15256_,
    new_n15257_, new_n15258_, new_n15259_, new_n15260_, new_n15261_,
    new_n15262_, new_n15263_, new_n15264_, new_n15265_, new_n15266_,
    new_n15267_, new_n15268_, new_n15269_, new_n15270_, new_n15271_,
    new_n15272_, new_n15273_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15280_, new_n15281_,
    new_n15282_, new_n15283_, new_n15284_, new_n15285_, new_n15286_,
    new_n15287_, new_n15288_, new_n15289_, new_n15290_, new_n15291_,
    new_n15294_, new_n15295_, new_n15296_, new_n15297_, new_n15298_,
    new_n15299_, new_n15300_, new_n15301_, new_n15302_, new_n15303_,
    new_n15304_, new_n15305_, new_n15306_, new_n15307_, new_n15308_,
    new_n15309_, new_n15310_, new_n15311_, new_n15312_, new_n15313_,
    new_n15314_, new_n15315_, new_n15316_, new_n15317_, new_n15318_,
    new_n15319_, new_n15320_, new_n15321_, new_n15322_, new_n15323_,
    new_n15324_, new_n15325_, new_n15326_, new_n15327_, new_n15328_,
    new_n15329_, new_n15330_, new_n15331_, new_n15332_, new_n15333_,
    new_n15334_, new_n15335_, new_n15336_, new_n15337_, new_n15338_,
    new_n15339_, new_n15340_, new_n15341_, new_n15342_, new_n15343_,
    new_n15344_, new_n15345_, new_n15346_, new_n15347_, new_n15348_,
    new_n15349_, new_n15350_, new_n15351_, new_n15352_, new_n15353_,
    new_n15354_, new_n15355_, new_n15356_, new_n15357_, new_n15358_,
    new_n15359_, new_n15360_, new_n15361_, new_n15362_, new_n15363_,
    new_n15364_, new_n15365_, new_n15366_, new_n15367_, new_n15368_,
    new_n15369_, new_n15370_, new_n15371_, new_n15372_, new_n15373_,
    new_n15374_, new_n15375_, new_n15376_, new_n15377_, new_n15378_,
    new_n15379_, new_n15380_, new_n15381_, new_n15382_, new_n15383_,
    new_n15384_, new_n15385_, new_n15386_, new_n15387_, new_n15388_,
    new_n15389_, new_n15390_, new_n15391_, new_n15392_, new_n15393_,
    new_n15394_, new_n15395_, new_n15396_, new_n15397_, new_n15398_,
    new_n15399_, new_n15400_, new_n15401_, new_n15402_, new_n15403_,
    new_n15404_, new_n15405_, new_n15406_, new_n15407_, new_n15408_,
    new_n15409_, new_n15410_, new_n15411_, new_n15412_, new_n15413_,
    new_n15414_, new_n15415_, new_n15416_, new_n15417_, new_n15418_,
    new_n15419_, new_n15420_, new_n15421_, new_n15422_, new_n15423_,
    new_n15424_, new_n15425_, new_n15426_, new_n15427_, new_n15428_,
    new_n15429_, new_n15430_, new_n15431_, new_n15432_, new_n15433_,
    new_n15434_, new_n15435_, new_n15436_, new_n15437_, new_n15438_,
    new_n15439_, new_n15440_, new_n15441_, new_n15442_, new_n15443_,
    new_n15444_, new_n15445_, new_n15446_, new_n15447_, new_n15448_,
    new_n15449_, new_n15450_, new_n15451_, new_n15452_, new_n15453_,
    new_n15454_, new_n15455_, new_n15456_, new_n15457_, new_n15458_,
    new_n15459_, new_n15460_, new_n15461_, new_n15462_, new_n15463_,
    new_n15464_, new_n15465_, new_n15466_, new_n15467_, new_n15468_,
    new_n15469_, new_n15470_, new_n15471_, new_n15472_, new_n15473_,
    new_n15474_, new_n15475_, new_n15476_, new_n15477_, new_n15478_,
    new_n15479_, new_n15480_, new_n15481_, new_n15482_, new_n15483_,
    new_n15484_, new_n15485_, new_n15486_, new_n15487_, new_n15488_,
    new_n15489_, new_n15490_, new_n15491_, new_n15492_, new_n15493_,
    new_n15494_, new_n15495_, new_n15496_, new_n15497_, new_n15498_,
    new_n15499_, new_n15500_, new_n15501_, new_n15502_, new_n15503_,
    new_n15504_, new_n15505_, new_n15506_, new_n15507_, new_n15508_,
    new_n15509_, new_n15510_, new_n15511_, new_n15512_, new_n15513_,
    new_n15514_, new_n15515_, new_n15516_, new_n15517_, new_n15518_,
    new_n15519_, new_n15520_, new_n15521_, new_n15522_, new_n15523_,
    new_n15524_, new_n15525_, new_n15526_, new_n15527_, new_n15528_,
    new_n15529_, new_n15530_, new_n15531_, new_n15532_, new_n15533_,
    new_n15534_, new_n15535_, new_n15536_, new_n15537_, new_n15538_,
    new_n15539_, new_n15540_, new_n15541_, new_n15542_, new_n15543_,
    new_n15544_, new_n15545_, new_n15546_, new_n15547_, new_n15548_,
    new_n15549_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15562_, new_n15563_, new_n15564_,
    new_n15565_, new_n15566_, new_n15567_, new_n15568_, new_n15569_,
    new_n15570_, new_n15571_, new_n15572_, new_n15573_, new_n15574_,
    new_n15575_, new_n15576_, new_n15577_, new_n15578_, new_n15579_,
    new_n15580_, new_n15581_, new_n15582_, new_n15583_, new_n15584_,
    new_n15585_, new_n15586_, new_n15587_, new_n15588_, new_n15589_,
    new_n15590_, new_n15591_, new_n15592_, new_n15593_, new_n15594_,
    new_n15595_, new_n15596_, new_n15597_, new_n15598_, new_n15599_,
    new_n15600_, new_n15601_, new_n15602_, new_n15603_, new_n15604_,
    new_n15605_, new_n15606_, new_n15607_, new_n15608_, new_n15609_,
    new_n15610_, new_n15611_, new_n15612_, new_n15613_, new_n15614_,
    new_n15615_, new_n15616_, new_n15617_, new_n15618_, new_n15619_,
    new_n15620_, new_n15621_, new_n15622_, new_n15623_, new_n15624_,
    new_n15625_, new_n15626_, new_n15627_, new_n15628_, new_n15629_,
    new_n15630_, new_n15631_, new_n15632_, new_n15633_, new_n15634_,
    new_n15635_, new_n15636_, new_n15637_, new_n15638_, new_n15639_,
    new_n15640_, new_n15641_, new_n15642_, new_n15643_, new_n15644_,
    new_n15645_, new_n15646_, new_n15647_, new_n15648_, new_n15649_,
    new_n15650_, new_n15651_, new_n15652_, new_n15653_, new_n15654_,
    new_n15655_, new_n15656_, new_n15657_, new_n15658_, new_n15659_,
    new_n15660_, new_n15661_, new_n15662_, new_n15663_, new_n15664_,
    new_n15665_, new_n15666_, new_n15667_, new_n15668_, new_n15669_,
    new_n15670_, new_n15671_, new_n15672_, new_n15673_, new_n15674_,
    new_n15675_, new_n15676_, new_n15677_, new_n15678_, new_n15679_,
    new_n15680_, new_n15681_, new_n15682_, new_n15683_, new_n15684_,
    new_n15685_, new_n15686_, new_n15687_, new_n15688_, new_n15689_,
    new_n15690_, new_n15691_, new_n15692_, new_n15693_, new_n15694_,
    new_n15695_, new_n15696_, new_n15697_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15832_,
    new_n15833_, new_n15834_, new_n15835_, new_n15836_, new_n15837_,
    new_n15838_, new_n15839_, new_n15840_, new_n15841_, new_n15842_,
    new_n15843_, new_n15844_, new_n15845_, new_n15846_, new_n15847_,
    new_n15848_, new_n15849_, new_n15850_, new_n15851_, new_n15852_,
    new_n15853_, new_n15854_, new_n15855_, new_n15856_, new_n15857_,
    new_n15858_, new_n15859_, new_n15860_, new_n15861_, new_n15862_,
    new_n15863_, new_n15864_, new_n15865_, new_n15868_, new_n15869_,
    new_n15870_, new_n15871_, new_n15872_, new_n15873_, new_n15874_,
    new_n15875_, new_n15876_, new_n15877_, new_n15878_, new_n15879_,
    new_n15880_, new_n15881_, new_n15882_, new_n15883_, new_n15884_,
    new_n15885_, new_n15886_, new_n15887_, new_n15888_, new_n15889_,
    new_n15890_, new_n15891_, new_n15892_, new_n15893_, new_n15894_,
    new_n15895_, new_n15896_, new_n15897_, new_n15898_, new_n15899_,
    new_n15900_, new_n15901_, new_n15902_, new_n15903_, new_n15904_,
    new_n15905_, new_n15906_, new_n15907_, new_n15908_, new_n15909_,
    new_n15910_, new_n15911_, new_n15912_, new_n15913_, new_n15914_,
    new_n15915_, new_n15916_, new_n15917_, new_n15918_, new_n15919_,
    new_n15920_, new_n15921_, new_n15922_, new_n15923_, new_n15924_,
    new_n15925_, new_n15926_, new_n15927_, new_n15928_, new_n15929_,
    new_n15930_, new_n15931_, new_n15932_, new_n15933_, new_n15934_,
    new_n15935_, new_n15936_, new_n15937_, new_n15938_, new_n15939_,
    new_n15940_, new_n15941_, new_n15942_, new_n15943_, new_n15944_,
    new_n15945_, new_n15946_, new_n15947_, new_n15948_, new_n15949_,
    new_n15950_, new_n15951_, new_n15952_, new_n15953_, new_n15954_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16067_, new_n16068_, new_n16069_,
    new_n16070_, new_n16071_, new_n16072_, new_n16073_, new_n16074_,
    new_n16075_, new_n16076_, new_n16077_, new_n16078_, new_n16079_,
    new_n16080_, new_n16081_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16166_, new_n16167_, new_n16168_, new_n16169_, new_n16170_,
    new_n16171_, new_n16172_, new_n16173_, new_n16174_, new_n16175_,
    new_n16176_, new_n16177_, new_n16178_, new_n16179_, new_n16180_,
    new_n16181_, new_n16182_, new_n16183_, new_n16184_, new_n16185_,
    new_n16186_, new_n16187_, new_n16188_, new_n16189_, new_n16190_,
    new_n16191_, new_n16192_, new_n16193_, new_n16194_, new_n16195_,
    new_n16196_, new_n16197_, new_n16198_, new_n16199_, new_n16200_,
    new_n16201_, new_n16202_, new_n16203_, new_n16204_, new_n16205_,
    new_n16206_, new_n16207_, new_n16208_, new_n16209_, new_n16210_,
    new_n16211_, new_n16212_, new_n16213_, new_n16214_, new_n16215_,
    new_n16216_, new_n16217_, new_n16218_, new_n16219_, new_n16220_,
    new_n16221_, new_n16222_, new_n16223_, new_n16224_, new_n16225_,
    new_n16226_, new_n16227_, new_n16228_, new_n16229_, new_n16230_,
    new_n16231_, new_n16232_, new_n16233_, new_n16234_, new_n16235_,
    new_n16236_, new_n16237_, new_n16238_, new_n16239_, new_n16240_,
    new_n16241_, new_n16242_, new_n16243_, new_n16244_, new_n16245_,
    new_n16246_, new_n16247_, new_n16248_, new_n16249_, new_n16250_,
    new_n16251_, new_n16252_, new_n16253_, new_n16254_, new_n16255_,
    new_n16256_, new_n16257_, new_n16258_, new_n16259_, new_n16260_,
    new_n16261_, new_n16262_, new_n16263_, new_n16264_, new_n16265_,
    new_n16266_, new_n16267_, new_n16268_, new_n16269_, new_n16270_,
    new_n16271_, new_n16272_, new_n16273_, new_n16276_, new_n16277_,
    new_n16278_, new_n16279_, new_n16280_, new_n16281_, new_n16282_,
    new_n16283_, new_n16284_, new_n16285_, new_n16286_, new_n16287_,
    new_n16288_, new_n16289_, new_n16290_, new_n16291_, new_n16292_,
    new_n16293_, new_n16294_, new_n16295_, new_n16296_, new_n16297_,
    new_n16298_, new_n16299_, new_n16300_, new_n16301_, new_n16304_,
    new_n16305_, new_n16306_, new_n16307_, new_n16308_, new_n16309_,
    new_n16310_, new_n16311_, new_n16312_, new_n16313_, new_n16314_,
    new_n16315_, new_n16316_, new_n16317_, new_n16318_, new_n16319_,
    new_n16320_, new_n16321_, new_n16322_, new_n16323_, new_n16324_,
    new_n16325_, new_n16326_, new_n16327_, new_n16328_, new_n16329_,
    new_n16330_, new_n16331_, new_n16332_, new_n16333_, new_n16334_,
    new_n16335_, new_n16336_, new_n16337_, new_n16338_, new_n16339_,
    new_n16340_, new_n16341_, new_n16342_, new_n16343_, new_n16344_,
    new_n16345_, new_n16346_, new_n16347_, new_n16348_, new_n16349_,
    new_n16350_, new_n16351_, new_n16352_, new_n16353_, new_n16354_,
    new_n16355_, new_n16356_, new_n16357_, new_n16358_, new_n16359_,
    new_n16360_, new_n16361_, new_n16362_, new_n16363_, new_n16365_,
    new_n16366_, new_n16367_, new_n16368_, new_n16369_, new_n16370_,
    new_n16371_, new_n16372_, new_n16373_, new_n16374_, new_n16375_,
    new_n16376_, new_n16377_, new_n16378_, new_n16379_, new_n16380_,
    new_n16381_, new_n16382_, new_n16383_, new_n16384_, new_n16385_,
    new_n16386_, new_n16387_, new_n16388_, new_n16389_, new_n16390_,
    new_n16391_, new_n16392_, new_n16393_, new_n16394_, new_n16395_,
    new_n16396_, new_n16397_, new_n16398_, new_n16399_, new_n16400_,
    new_n16401_, new_n16402_, new_n16403_, new_n16404_, new_n16405_,
    new_n16406_, new_n16407_, new_n16408_, new_n16409_, new_n16410_,
    new_n16411_, new_n16412_, new_n16413_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16494_, new_n16495_, new_n16496_, new_n16497_,
    new_n16498_, new_n16499_, new_n16500_, new_n16501_, new_n16502_,
    new_n16503_, new_n16504_, new_n16505_, new_n16506_, new_n16507_,
    new_n16508_, new_n16509_, new_n16510_, new_n16511_, new_n16512_,
    new_n16513_, new_n16514_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16523_,
    new_n16524_, new_n16525_, new_n16526_, new_n16527_, new_n16528_,
    new_n16529_, new_n16530_, new_n16531_, new_n16532_, new_n16533_,
    new_n16534_, new_n16535_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16590_, new_n16591_, new_n16592_, new_n16593_,
    new_n16594_, new_n16595_, new_n16596_, new_n16597_, new_n16598_,
    new_n16599_, new_n16600_, new_n16601_, new_n16602_, new_n16603_,
    new_n16604_, new_n16605_, new_n16606_, new_n16607_, new_n16608_,
    new_n16609_, new_n16610_, new_n16611_, new_n16612_, new_n16613_,
    new_n16614_, new_n16615_, new_n16616_, new_n16617_, new_n16618_,
    new_n16619_, new_n16620_, new_n16621_, new_n16622_, new_n16623_,
    new_n16624_, new_n16625_, new_n16626_, new_n16627_, new_n16628_,
    new_n16629_, new_n16630_, new_n16631_, new_n16632_, new_n16633_,
    new_n16634_, new_n16635_, new_n16636_, new_n16637_, new_n16638_,
    new_n16639_, new_n16640_, new_n16641_, new_n16642_, new_n16643_,
    new_n16644_, new_n16645_, new_n16646_, new_n16647_, new_n16648_,
    new_n16649_, new_n16650_, new_n16651_, new_n16652_, new_n16653_,
    new_n16654_, new_n16655_, new_n16656_, new_n16657_, new_n16658_,
    new_n16659_, new_n16660_, new_n16661_, new_n16662_, new_n16663_,
    new_n16664_, new_n16665_, new_n16666_, new_n16667_, new_n16668_,
    new_n16669_, new_n16670_, new_n16671_, new_n16672_, new_n16673_,
    new_n16674_, new_n16675_, new_n16676_, new_n16677_, new_n16678_,
    new_n16679_, new_n16680_, new_n16681_, new_n16682_, new_n16683_,
    new_n16684_, new_n16685_, new_n16686_, new_n16687_, new_n16688_,
    new_n16689_, new_n16690_, new_n16691_, new_n16692_, new_n16693_,
    new_n16694_, new_n16695_, new_n16696_, new_n16697_, new_n16698_,
    new_n16699_, new_n16700_, new_n16701_, new_n16702_, new_n16703_,
    new_n16704_, new_n16705_, new_n16706_, new_n16707_, new_n16708_,
    new_n16709_, new_n16710_, new_n16711_, new_n16712_, new_n16713_,
    new_n16714_, new_n16715_, new_n16716_, new_n16717_, new_n16718_,
    new_n16719_, new_n16720_, new_n16721_, new_n16722_, new_n16723_,
    new_n16724_, new_n16725_, new_n16726_, new_n16727_, new_n16728_,
    new_n16729_, new_n16730_, new_n16731_, new_n16732_, new_n16733_,
    new_n16734_, new_n16735_, new_n16736_, new_n16737_, new_n16738_,
    new_n16739_, new_n16740_, new_n16741_, new_n16742_, new_n16743_,
    new_n16744_, new_n16745_, new_n16746_, new_n16747_, new_n16748_,
    new_n16749_, new_n16750_, new_n16751_, new_n16752_, new_n16753_,
    new_n16754_, new_n16755_, new_n16756_, new_n16757_, new_n16758_,
    new_n16759_, new_n16760_, new_n16761_, new_n16762_, new_n16763_,
    new_n16764_, new_n16765_, new_n16766_, new_n16767_, new_n16768_,
    new_n16769_, new_n16770_, new_n16771_, new_n16772_, new_n16773_,
    new_n16774_, new_n16775_, new_n16776_, new_n16777_, new_n16778_,
    new_n16779_, new_n16780_, new_n16781_, new_n16782_, new_n16783_,
    new_n16784_, new_n16785_, new_n16786_, new_n16787_, new_n16788_,
    new_n16789_, new_n16790_, new_n16791_, new_n16792_, new_n16793_,
    new_n16794_, new_n16795_, new_n16796_, new_n16797_, new_n16798_,
    new_n16799_, new_n16800_, new_n16801_, new_n16802_, new_n16803_,
    new_n16804_, new_n16805_, new_n16806_, new_n16807_, new_n16808_,
    new_n16809_, new_n16810_, new_n16811_, new_n16812_, new_n16813_,
    new_n16814_, new_n16815_, new_n16816_, new_n16817_, new_n16818_,
    new_n16819_, new_n16820_, new_n16821_, new_n16822_, new_n16823_,
    new_n16824_, new_n16825_, new_n16826_, new_n16827_, new_n16828_,
    new_n16829_, new_n16830_, new_n16831_, new_n16832_, new_n16833_,
    new_n16834_, new_n16835_, new_n16836_, new_n16837_, new_n16838_,
    new_n16839_, new_n16840_, new_n16841_, new_n16842_, new_n16843_,
    new_n16844_, new_n16845_, new_n16846_, new_n16847_, new_n16848_,
    new_n16849_, new_n16850_, new_n16851_, new_n16852_, new_n16853_,
    new_n16854_, new_n16855_, new_n16856_, new_n16857_, new_n16858_,
    new_n16859_, new_n16860_, new_n16861_, new_n16862_, new_n16863_,
    new_n16864_, new_n16865_, new_n16866_, new_n16867_, new_n16868_,
    new_n16869_, new_n16870_, new_n16871_, new_n16872_, new_n16873_,
    new_n16874_, new_n16875_, new_n16876_, new_n16877_, new_n16878_,
    new_n16879_, new_n16880_, new_n16881_, new_n16882_, new_n16883_,
    new_n16884_, new_n16885_, new_n16886_, new_n16887_, new_n16888_,
    new_n16889_, new_n16890_, new_n16891_, new_n16892_, new_n16893_,
    new_n16894_, new_n16895_, new_n16896_, new_n16897_, new_n16898_,
    new_n16899_, new_n16900_, new_n16901_, new_n16902_, new_n16903_,
    new_n16904_, new_n16905_, new_n16906_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16954_, new_n16955_,
    new_n16956_, new_n16957_, new_n16958_, new_n16959_, new_n16961_,
    new_n16962_, new_n16963_, new_n16964_, new_n16965_, new_n16966_,
    new_n16967_, new_n16968_, new_n16969_, new_n16970_, new_n16971_,
    new_n16972_, new_n16973_, new_n16974_, new_n16975_, new_n16976_,
    new_n16977_, new_n16978_, new_n16979_, new_n16980_, new_n16981_,
    new_n16982_, new_n16983_, new_n16984_, new_n16985_, new_n16986_,
    new_n16987_, new_n16988_, new_n16989_, new_n16990_, new_n16991_,
    new_n16992_, new_n16993_, new_n16994_, new_n16995_, new_n16996_,
    new_n16997_, new_n16998_, new_n16999_, new_n17000_, new_n17001_,
    new_n17002_, new_n17003_, new_n17004_, new_n17005_, new_n17006_,
    new_n17007_, new_n17008_, new_n17009_, new_n17010_, new_n17011_,
    new_n17012_, new_n17013_, new_n17014_, new_n17015_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17148_,
    new_n17149_, new_n17150_, new_n17151_, new_n17152_, new_n17153_,
    new_n17154_, new_n17155_, new_n17156_, new_n17157_, new_n17158_,
    new_n17159_, new_n17160_, new_n17161_, new_n17162_, new_n17163_,
    new_n17164_, new_n17165_, new_n17166_, new_n17167_, new_n17168_,
    new_n17169_, new_n17170_, new_n17171_, new_n17172_, new_n17173_,
    new_n17174_, new_n17175_, new_n17176_, new_n17177_, new_n17178_,
    new_n17179_, new_n17180_, new_n17181_, new_n17182_, new_n17183_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17190_, new_n17191_, new_n17192_, new_n17193_, new_n17194_,
    new_n17195_, new_n17196_, new_n17197_, new_n17198_, new_n17199_,
    new_n17200_, new_n17201_, new_n17202_, new_n17203_, new_n17204_,
    new_n17205_, new_n17206_, new_n17207_, new_n17208_, new_n17209_,
    new_n17210_, new_n17211_, new_n17212_, new_n17213_, new_n17214_,
    new_n17215_, new_n17216_, new_n17217_, new_n17218_, new_n17219_,
    new_n17220_, new_n17221_, new_n17222_, new_n17223_, new_n17224_,
    new_n17225_, new_n17227_, new_n17228_, new_n17229_, new_n17230_,
    new_n17231_, new_n17232_, new_n17233_, new_n17234_, new_n17235_,
    new_n17236_, new_n17237_, new_n17238_, new_n17239_, new_n17240_,
    new_n17241_, new_n17242_, new_n17243_, new_n17244_, new_n17245_,
    new_n17246_, new_n17247_, new_n17248_, new_n17249_, new_n17250_,
    new_n17251_, new_n17252_, new_n17253_, new_n17254_, new_n17255_,
    new_n17256_, new_n17257_, new_n17258_, new_n17259_, new_n17260_,
    new_n17261_, new_n17262_, new_n17263_, new_n17264_, new_n17265_,
    new_n17266_, new_n17267_, new_n17268_, new_n17269_, new_n17270_,
    new_n17271_, new_n17272_, new_n17273_, new_n17274_, new_n17275_,
    new_n17276_, new_n17277_, new_n17278_, new_n17279_, new_n17280_,
    new_n17281_, new_n17282_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17330_, new_n17331_, new_n17332_, new_n17333_,
    new_n17334_, new_n17335_, new_n17336_, new_n17337_, new_n17338_,
    new_n17339_, new_n17340_, new_n17341_, new_n17342_, new_n17343_,
    new_n17344_, new_n17345_, new_n17346_, new_n17347_, new_n17348_,
    new_n17349_, new_n17350_, new_n17351_, new_n17352_, new_n17353_,
    new_n17355_, new_n17356_, new_n17357_, new_n17358_, new_n17359_,
    new_n17360_, new_n17361_, new_n17362_, new_n17363_, new_n17364_,
    new_n17365_, new_n17366_, new_n17367_, new_n17368_, new_n17369_,
    new_n17370_, new_n17371_, new_n17372_, new_n17373_, new_n17374_,
    new_n17375_, new_n17376_, new_n17377_, new_n17378_, new_n17379_,
    new_n17380_, new_n17381_, new_n17382_, new_n17383_, new_n17384_,
    new_n17385_, new_n17386_, new_n17387_, new_n17388_, new_n17389_,
    new_n17390_, new_n17391_, new_n17392_, new_n17393_, new_n17394_,
    new_n17395_, new_n17396_, new_n17397_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17406_, new_n17407_, new_n17408_,
    new_n17409_, new_n17410_, new_n17411_, new_n17412_, new_n17413_,
    new_n17414_, new_n17415_, new_n17416_, new_n17417_, new_n17418_,
    new_n17419_, new_n17420_, new_n17421_, new_n17422_, new_n17423_,
    new_n17424_, new_n17425_, new_n17426_, new_n17427_, new_n17428_,
    new_n17429_, new_n17430_, new_n17431_, new_n17432_, new_n17433_,
    new_n17434_, new_n17435_, new_n17436_, new_n17437_, new_n17438_,
    new_n17440_, new_n17441_, new_n17442_, new_n17443_, new_n17444_,
    new_n17445_, new_n17446_, new_n17447_, new_n17448_, new_n17449_,
    new_n17450_, new_n17451_, new_n17452_, new_n17453_, new_n17454_,
    new_n17455_, new_n17456_, new_n17457_, new_n17458_, new_n17459_,
    new_n17460_, new_n17461_, new_n17462_, new_n17463_, new_n17464_,
    new_n17465_, new_n17466_, new_n17467_, new_n17468_, new_n17469_,
    new_n17470_, new_n17472_, new_n17473_, new_n17474_, new_n17475_,
    new_n17476_, new_n17477_, new_n17478_, new_n17479_, new_n17480_,
    new_n17481_, new_n17482_, new_n17483_, new_n17484_, new_n17485_,
    new_n17486_, new_n17487_, new_n17488_, new_n17489_, new_n17490_,
    new_n17491_, new_n17492_, new_n17493_, new_n17495_, new_n17496_,
    new_n17497_, new_n17498_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17504_, new_n17505_, new_n17506_,
    new_n17507_, new_n17508_, new_n17509_, new_n17510_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17516_,
    new_n17517_, new_n17518_, new_n17519_, new_n17520_, new_n17521_,
    new_n17522_, new_n17523_, new_n17524_, new_n17525_, new_n17526_,
    new_n17527_, new_n17528_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17567_, new_n17568_,
    new_n17569_, new_n17570_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17576_, new_n17577_, new_n17578_,
    new_n17579_, new_n17580_, new_n17581_, new_n17582_, new_n17583_,
    new_n17584_, new_n17585_, new_n17586_, new_n17587_, new_n17588_,
    new_n17589_, new_n17590_, new_n17591_, new_n17592_, new_n17593_,
    new_n17594_, new_n17595_, new_n17596_, new_n17597_, new_n17598_,
    new_n17599_, new_n17600_, new_n17601_, new_n17602_, new_n17604_,
    new_n17605_, new_n17606_, new_n17607_, new_n17608_, new_n17609_,
    new_n17610_, new_n17611_, new_n17612_, new_n17613_, new_n17614_,
    new_n17615_, new_n17616_, new_n17617_, new_n17618_, new_n17619_,
    new_n17620_, new_n17621_, new_n17622_, new_n17623_, new_n17624_,
    new_n17625_, new_n17626_, new_n17627_, new_n17628_, new_n17629_,
    new_n17630_, new_n17631_, new_n17632_, new_n17633_, new_n17634_,
    new_n17635_, new_n17636_, new_n17637_, new_n17638_, new_n17639_,
    new_n17640_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17700_, new_n17701_, new_n17702_, new_n17703_,
    new_n17704_, new_n17705_, new_n17706_, new_n17707_, new_n17708_,
    new_n17709_, new_n17710_, new_n17711_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17730_, new_n17731_, new_n17732_, new_n17733_, new_n17734_,
    new_n17735_, new_n17736_, new_n17737_, new_n17738_, new_n17739_,
    new_n17740_, new_n17741_, new_n17742_, new_n17743_, new_n17744_,
    new_n17745_, new_n17746_, new_n17747_, new_n17748_, new_n17749_,
    new_n17750_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17766_, new_n17767_, new_n17768_, new_n17769_, new_n17770_,
    new_n17771_, new_n17772_, new_n17773_, new_n17774_, new_n17775_,
    new_n17776_, new_n17777_, new_n17778_, new_n17779_, new_n17780_,
    new_n17781_, new_n17782_, new_n17783_, new_n17784_, new_n17785_,
    new_n17786_, new_n17787_, new_n17788_, new_n17789_, new_n17790_,
    new_n17792_, new_n17793_, new_n17794_, new_n17795_, new_n17796_,
    new_n17797_, new_n17798_, new_n17799_, new_n17800_, new_n17801_,
    new_n17802_, new_n17803_, new_n17804_, new_n17805_, new_n17806_,
    new_n17807_, new_n17808_, new_n17809_, new_n17810_, new_n17811_,
    new_n17812_, new_n17814_, new_n17815_, new_n17816_, new_n17817_,
    new_n17818_, new_n17819_, new_n17820_, new_n17821_, new_n17822_,
    new_n17823_, new_n17824_, new_n17825_, new_n17826_, new_n17827_,
    new_n17828_, new_n17829_, new_n17830_, new_n17831_, new_n17832_,
    new_n17833_, new_n17834_, new_n17835_, new_n17836_, new_n17837_,
    new_n17838_, new_n17839_, new_n17840_, new_n17841_, new_n17842_,
    new_n17843_, new_n17844_, new_n17845_, new_n17846_, new_n17847_,
    new_n17848_, new_n17849_, new_n17850_, new_n17851_, new_n17852_,
    new_n17853_, new_n17854_, new_n17855_, new_n17856_, new_n17857_,
    new_n17858_, new_n17859_, new_n17860_, new_n17861_, new_n17862_,
    new_n17863_, new_n17864_, new_n17865_, new_n17866_, new_n17867_,
    new_n17868_, new_n17869_, new_n17870_, new_n17871_, new_n17872_,
    new_n17873_, new_n17874_, new_n17875_, new_n17876_, new_n17877_,
    new_n17878_, new_n17880_, new_n17881_, new_n17882_, new_n17883_,
    new_n17884_, new_n17885_, new_n17886_, new_n17887_, new_n17888_,
    new_n17889_, new_n17890_, new_n17891_, new_n17892_, new_n17893_,
    new_n17894_, new_n17895_, new_n17896_, new_n17897_, new_n17898_,
    new_n17899_, new_n17900_, new_n17901_, new_n17902_, new_n17903_,
    new_n17904_, new_n17905_, new_n17906_, new_n17907_, new_n17908_,
    new_n17909_, new_n17910_, new_n17912_, new_n17913_, new_n17914_,
    new_n17915_, new_n17916_, new_n17917_, new_n17918_, new_n17919_,
    new_n17920_, new_n17921_, new_n17922_, new_n17923_, new_n17924_,
    new_n17925_, new_n17926_, new_n17927_, new_n17928_, new_n17929_,
    new_n17930_, new_n17931_, new_n17932_, new_n17933_, new_n17934_,
    new_n17935_, new_n17936_, new_n17937_, new_n17938_, new_n17939_,
    new_n17940_, new_n17941_, new_n17942_, new_n17943_, new_n17944_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17952_,
    new_n17953_, new_n17954_, new_n17956_, new_n17957_, new_n17958_,
    new_n17959_, new_n17960_, new_n17961_, new_n17962_, new_n17963_,
    new_n17964_, new_n17965_, new_n17966_, new_n17967_, new_n17968_,
    new_n17969_, new_n17970_, new_n17971_, new_n17972_, new_n17973_,
    new_n17974_, new_n17975_, new_n17976_, new_n17977_, new_n17978_,
    new_n17979_, new_n17980_, new_n17981_, new_n17982_, new_n17983_,
    new_n17984_, new_n17985_, new_n17986_, new_n17987_, new_n17988_,
    new_n17989_, new_n17990_, new_n17991_, new_n17992_, new_n17996_,
    new_n17997_, new_n17998_, new_n18000_, new_n18001_, new_n18002_,
    new_n18003_, new_n18004_, new_n18005_, new_n18006_, new_n18007_,
    new_n18008_, new_n18009_, new_n18010_, new_n18011_, new_n18012_,
    new_n18013_, new_n18014_, new_n18015_, new_n18016_, new_n18017_,
    new_n18018_, new_n18019_, new_n18020_, new_n18021_, new_n18022_,
    new_n18023_, new_n18024_, new_n18025_, new_n18026_, new_n18027_,
    new_n18028_, new_n18029_, new_n18030_, new_n18031_, new_n18032_,
    new_n18033_, new_n18034_, new_n18035_, new_n18036_, new_n18037_,
    new_n18038_, new_n18039_, new_n18040_, new_n18041_, new_n18042_,
    new_n18043_, new_n18044_, new_n18045_, new_n18046_, new_n18047_,
    new_n18048_, new_n18049_, new_n18051_, new_n18052_, new_n18053_,
    new_n18054_, new_n18055_, new_n18056_, new_n18057_, new_n18058_,
    new_n18059_, new_n18060_, new_n18061_, new_n18062_, new_n18063_,
    new_n18064_, new_n18065_, new_n18066_, new_n18067_, new_n18068_,
    new_n18069_, new_n18070_, new_n18071_, new_n18072_, new_n18073_,
    new_n18074_, new_n18075_, new_n18076_, new_n18077_, new_n18078_,
    new_n18079_, new_n18080_, new_n18081_, new_n18082_, new_n18083_,
    new_n18084_, new_n18085_, new_n18086_, new_n18087_, new_n18091_,
    new_n18092_, new_n18093_, new_n18095_, new_n18096_, new_n18097_,
    new_n18098_, new_n18099_, new_n18100_, new_n18101_, new_n18102_,
    new_n18103_, new_n18104_, new_n18105_, new_n18106_, new_n18107_,
    new_n18108_, new_n18109_, new_n18110_, new_n18111_, new_n18112_,
    new_n18113_, new_n18114_, new_n18115_, new_n18116_, new_n18117_,
    new_n18118_, new_n18119_, new_n18120_, new_n18121_, new_n18122_,
    new_n18123_, new_n18124_, new_n18125_, new_n18126_, new_n18127_,
    new_n18128_, new_n18129_, new_n18130_, new_n18131_, new_n18132_,
    new_n18133_, new_n18134_, new_n18139_, new_n18140_, new_n18142_,
    new_n18143_, new_n18144_, new_n18145_, new_n18146_, new_n18147_,
    new_n18148_, new_n18149_, new_n18150_, new_n18151_, new_n18152_,
    new_n18153_, new_n18154_, new_n18155_, new_n18156_, new_n18157_,
    new_n18158_, new_n18159_, new_n18160_, new_n18161_, new_n18162_,
    new_n18163_, new_n18164_, new_n18165_, new_n18166_, new_n18167_,
    new_n18168_, new_n18169_, new_n18170_, new_n18171_, new_n18172_,
    new_n18173_, new_n18174_, new_n18175_, new_n18176_, new_n18177_,
    new_n18178_, new_n18179_, new_n18180_, new_n18181_, new_n18182_,
    new_n18183_, new_n18184_, new_n18185_, new_n18186_, new_n18187_,
    new_n18188_, new_n18189_, new_n18190_, new_n18191_, new_n18192_,
    new_n18193_, new_n18194_, new_n18195_, new_n18196_, new_n18197_,
    new_n18198_, new_n18199_, new_n18200_, new_n18201_, new_n18202_,
    new_n18203_, new_n18204_, new_n18205_, new_n18206_, new_n18207_,
    new_n18208_, new_n18209_, new_n18210_, new_n18211_, new_n18212_,
    new_n18213_, new_n18214_, new_n18215_, new_n18216_, new_n18217_,
    new_n18218_, new_n18219_, new_n18220_, new_n18221_, new_n18222_,
    new_n18223_, new_n18224_, new_n18225_, new_n18226_, new_n18227_,
    new_n18228_, new_n18229_, new_n18230_, new_n18231_, new_n18232_,
    new_n18233_, new_n18234_, new_n18235_, new_n18236_, new_n18237_,
    new_n18238_, new_n18239_, new_n18240_, new_n18241_, new_n18242_,
    new_n18243_, new_n18244_, new_n18245_, new_n18246_, new_n18247_,
    new_n18248_, new_n18249_, new_n18250_, new_n18251_, new_n18252_,
    new_n18253_, new_n18254_, new_n18255_, new_n18256_, new_n18257_,
    new_n18258_, new_n18259_, new_n18260_, new_n18261_, new_n18262_,
    new_n18263_, new_n18264_, new_n18265_, new_n18266_, new_n18267_,
    new_n18268_, new_n18269_, new_n18270_, new_n18271_, new_n18272_,
    new_n18273_, new_n18274_, new_n18275_, new_n18276_, new_n18277_,
    new_n18278_, new_n18279_, new_n18280_, new_n18281_, new_n18282_,
    new_n18283_, new_n18284_, new_n18285_, new_n18286_, new_n18287_,
    new_n18288_, new_n18289_, new_n18290_, new_n18291_, new_n18292_,
    new_n18293_, new_n18294_, new_n18295_, new_n18296_, new_n18297_,
    new_n18298_, new_n18299_, new_n18300_, new_n18301_, new_n18302_,
    new_n18303_, new_n18304_, new_n18305_, new_n18306_, new_n18307_,
    new_n18308_, new_n18309_, new_n18310_, new_n18311_, new_n18312_,
    new_n18313_, new_n18314_, new_n18315_, new_n18316_, new_n18317_,
    new_n18318_, new_n18319_, new_n18320_, new_n18321_, new_n18322_,
    new_n18323_, new_n18324_, new_n18325_, new_n18326_, new_n18327_,
    new_n18328_, new_n18329_, new_n18330_, new_n18331_, new_n18332_,
    new_n18333_, new_n18334_, new_n18335_, new_n18336_, new_n18337_,
    new_n18338_, new_n18339_, new_n18340_, new_n18341_, new_n18342_,
    new_n18343_, new_n18344_, new_n18345_, new_n18346_, new_n18347_,
    new_n18348_, new_n18349_, new_n18350_, new_n18351_, new_n18352_,
    new_n18353_, new_n18354_, new_n18355_, new_n18356_, new_n18357_,
    new_n18358_, new_n18359_, new_n18360_, new_n18361_, new_n18362_,
    new_n18363_, new_n18364_, new_n18365_, new_n18366_, new_n18367_,
    new_n18368_, new_n18369_, new_n18370_, new_n18371_, new_n18372_,
    new_n18373_, new_n18374_, new_n18375_, new_n18376_, new_n18377_,
    new_n18378_, new_n18379_, new_n18380_, new_n18381_, new_n18382_,
    new_n18383_, new_n18384_, new_n18385_, new_n18386_, new_n18387_,
    new_n18388_, new_n18389_, new_n18390_, new_n18391_, new_n18392_,
    new_n18393_, new_n18394_, new_n18395_, new_n18396_, new_n18397_,
    new_n18398_, new_n18399_, new_n18400_, new_n18401_, new_n18402_,
    new_n18403_, new_n18404_, new_n18405_, new_n18406_, new_n18407_,
    new_n18408_, new_n18409_, new_n18410_, new_n18411_, new_n18412_,
    new_n18413_, new_n18414_, new_n18415_, new_n18416_, new_n18417_,
    new_n18418_, new_n18419_, new_n18420_, new_n18421_, new_n18422_,
    new_n18423_, new_n18424_, new_n18425_, new_n18426_, new_n18427_,
    new_n18428_, new_n18429_, new_n18430_, new_n18431_, new_n18432_,
    new_n18433_, new_n18434_, new_n18435_, new_n18436_, new_n18437_,
    new_n18438_, new_n18439_, new_n18440_, new_n18441_, new_n18442_,
    new_n18443_, new_n18444_, new_n18445_, new_n18446_, new_n18447_,
    new_n18448_, new_n18449_, new_n18450_, new_n18451_, new_n18452_,
    new_n18453_, new_n18454_, new_n18455_, new_n18456_, new_n18457_,
    new_n18458_, new_n18459_, new_n18460_, new_n18461_, new_n18462_,
    new_n18463_, new_n18464_, new_n18465_, new_n18466_, new_n18467_,
    new_n18468_, new_n18469_, new_n18470_, new_n18471_, new_n18472_,
    new_n18473_, new_n18474_, new_n18475_, new_n18476_, new_n18477_,
    new_n18478_, new_n18479_, new_n18480_, new_n18481_, new_n18482_,
    new_n18483_, new_n18484_, new_n18485_, new_n18486_, new_n18487_,
    new_n18488_, new_n18489_, new_n18490_, new_n18491_, new_n18492_,
    new_n18493_, new_n18494_, new_n18495_, new_n18496_, new_n18497_,
    new_n18498_, new_n18499_, new_n18500_, new_n18501_, new_n18502_,
    new_n18503_, new_n18504_, new_n18505_, new_n18506_, new_n18507_,
    new_n18508_, new_n18509_, new_n18510_, new_n18511_, new_n18513_,
    new_n18514_, new_n18515_, new_n18516_, new_n18517_, new_n18518_,
    new_n18519_, new_n18520_, new_n18521_, new_n18522_, new_n18523_,
    new_n18524_, new_n18525_, new_n18526_, new_n18527_, new_n18528_,
    new_n18529_, new_n18530_, new_n18531_, new_n18532_, new_n18533_,
    new_n18534_, new_n18535_, new_n18536_, new_n18537_, new_n18538_,
    new_n18544_, new_n18545_, new_n18546_, new_n18547_, new_n18548_,
    new_n18549_, new_n18550_, new_n18551_, new_n18552_, new_n18553_,
    new_n18554_, new_n18555_, new_n18556_, new_n18557_, new_n18558_,
    new_n18559_, new_n18560_, new_n18561_, new_n18562_, new_n18563_,
    new_n18564_, new_n18565_, new_n18566_, new_n18567_, new_n18568_,
    new_n18569_, new_n18570_, new_n18571_, new_n18572_, new_n18573_,
    new_n18574_, new_n18575_, new_n18576_, new_n18577_, new_n18578_,
    new_n18579_, new_n18580_, new_n18581_, new_n18582_, new_n18583_,
    new_n18584_, new_n18585_, new_n18586_, new_n18587_, new_n18588_,
    new_n18589_, new_n18590_, new_n18591_, new_n18592_, new_n18593_,
    new_n18594_, new_n18595_, new_n18596_, new_n18597_, new_n18598_,
    new_n18599_, new_n18600_, new_n18601_, new_n18602_, new_n18603_,
    new_n18604_, new_n18605_, new_n18606_, new_n18607_, new_n18608_,
    new_n18609_, new_n18610_, new_n18611_, new_n18612_, new_n18613_,
    new_n18614_, new_n18615_, new_n18616_, new_n18617_, new_n18618_,
    new_n18619_, new_n18620_, new_n18621_, new_n18622_, new_n18623_,
    new_n18624_, new_n18625_, new_n18626_, new_n18627_, new_n18628_,
    new_n18629_, new_n18630_, new_n18631_, new_n18632_, new_n18633_,
    new_n18634_, new_n18635_, new_n18636_, new_n18637_, new_n18638_,
    new_n18639_, new_n18640_, new_n18641_, new_n18642_, new_n18643_,
    new_n18644_, new_n18645_, new_n18646_, new_n18647_, new_n18648_,
    new_n18649_, new_n18650_, new_n18651_, new_n18652_, new_n18653_,
    new_n18654_, new_n18655_, new_n18656_, new_n18657_, new_n18658_,
    new_n18659_, new_n18660_, new_n18661_, new_n18662_, new_n18663_,
    new_n18664_, new_n18665_, new_n18666_, new_n18667_, new_n18668_,
    new_n18669_, new_n18670_, new_n18671_, new_n18672_, new_n18676_,
    new_n18677_, new_n18678_, new_n18679_, new_n18680_, new_n18681_,
    new_n18682_, new_n18683_, new_n18684_, new_n18685_, new_n18686_,
    new_n18687_, new_n18688_, new_n18689_, new_n18690_, new_n18691_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18703_, new_n18704_,
    new_n18705_, new_n18708_, new_n18709_, new_n18710_, new_n18711_,
    new_n18712_, new_n18713_, new_n18714_, new_n18715_, new_n18716_,
    new_n18717_, new_n18718_, new_n18719_, new_n18720_, new_n18721_,
    new_n18722_, new_n18723_, new_n18724_, new_n18725_, new_n18726_,
    new_n18727_, new_n18728_, new_n18729_, new_n18730_, new_n18731_,
    new_n18732_, new_n18733_, new_n18734_, new_n18735_, new_n18736_,
    new_n18737_, new_n18738_, new_n18739_, new_n18740_, new_n18741_,
    new_n18742_, new_n18743_, new_n18744_, new_n18745_, new_n18746_,
    new_n18747_, new_n18748_, new_n18749_, new_n18750_, new_n18751_,
    new_n18752_, new_n18753_, new_n18754_, new_n18755_, new_n18756_,
    new_n18757_, new_n18758_, new_n18759_, new_n18760_, new_n18761_,
    new_n18762_, new_n18763_, new_n18764_, new_n18765_, new_n18766_,
    new_n18767_, new_n18768_, new_n18769_, new_n18770_, new_n18771_,
    new_n18772_, new_n18773_, new_n18774_, new_n18775_, new_n18776_,
    new_n18777_, new_n18778_, new_n18779_, new_n18780_, new_n18781_,
    new_n18782_, new_n18783_, new_n18784_, new_n18785_, new_n18786_,
    new_n18787_, new_n18788_, new_n18789_, new_n18790_, new_n18791_,
    new_n18792_, new_n18793_, new_n18794_, new_n18795_, new_n18796_,
    new_n18797_, new_n18798_, new_n18799_, new_n18800_, new_n18801_,
    new_n18802_, new_n18803_, new_n18804_, new_n18805_, new_n18806_,
    new_n18807_, new_n18808_, new_n18809_, new_n18810_, new_n18811_,
    new_n18812_, new_n18813_, new_n18814_, new_n18815_, new_n18816_,
    new_n18817_, new_n18818_, new_n18819_, new_n18820_, new_n18821_,
    new_n18822_, new_n18823_, new_n18824_, new_n18825_, new_n18826_,
    new_n18827_, new_n18828_, new_n18829_, new_n18830_, new_n18831_,
    new_n18832_, new_n18833_, new_n18834_, new_n18835_, new_n18836_,
    new_n18837_, new_n18838_, new_n18839_, new_n18840_, new_n18841_,
    new_n18842_, new_n18843_, new_n18844_, new_n18845_, new_n18846_,
    new_n18847_, new_n18848_, new_n18849_, new_n18850_, new_n18851_,
    new_n18852_, new_n18853_, new_n18854_, new_n18855_, new_n18856_,
    new_n18857_, new_n18858_, new_n18859_, new_n18860_, new_n18861_,
    new_n18862_, new_n18863_, new_n18864_, new_n18865_, new_n18866_,
    new_n18867_, new_n18868_, new_n18869_, new_n18870_, new_n18871_,
    new_n18872_, new_n18873_, new_n18874_, new_n18875_, new_n18876_,
    new_n18877_, new_n18878_, new_n18879_, new_n18880_, new_n18881_,
    new_n18882_, new_n18883_, new_n18884_, new_n18885_, new_n18886_,
    new_n18887_, new_n18888_, new_n18889_, new_n18890_, new_n18891_,
    new_n18892_, new_n18893_, new_n18894_, new_n18895_, new_n18896_,
    new_n18897_, new_n18898_, new_n18899_, new_n18900_, new_n18901_,
    new_n18902_, new_n18903_, new_n18904_, new_n18905_, new_n18906_,
    new_n18907_, new_n18908_, new_n18909_, new_n18911_, new_n18912_,
    new_n18913_, new_n18914_, new_n18915_, new_n18916_, new_n18917_,
    new_n18918_, new_n18919_, new_n18920_, new_n18921_, new_n18922_,
    new_n18923_, new_n18924_, new_n18925_, new_n18926_, new_n18927_,
    new_n18928_, new_n18929_, new_n18930_, new_n18931_, new_n18932_,
    new_n18933_, new_n18934_, new_n18935_, new_n18936_, new_n18937_,
    new_n18938_, new_n18939_, new_n18940_, new_n18941_, new_n18942_,
    new_n18943_, new_n18944_, new_n18945_, new_n18946_, new_n18947_,
    new_n18948_, new_n18949_, new_n18950_, new_n18951_, new_n18952_,
    new_n18953_, new_n18954_, new_n18955_, new_n18956_, new_n18957_,
    new_n18958_, new_n18959_, new_n18960_, new_n18961_, new_n18962_,
    new_n18963_, new_n18964_, new_n18965_, new_n18966_, new_n18967_,
    new_n18968_, new_n18969_, new_n18970_, new_n18971_, new_n18972_,
    new_n18973_, new_n18974_, new_n18975_, new_n18976_, new_n18977_,
    new_n18978_, new_n18979_, new_n18980_, new_n18981_, new_n18982_,
    new_n18983_, new_n18984_, new_n18985_, new_n18986_, new_n18987_,
    new_n18988_, new_n18989_, new_n18992_, new_n18993_, new_n18994_,
    new_n18995_, new_n18996_, new_n18997_, new_n18998_, new_n18999_,
    new_n19000_, new_n19001_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19007_, new_n19008_, new_n19009_,
    new_n19010_, new_n19011_, new_n19012_, new_n19013_, new_n19014_,
    new_n19015_, new_n19016_, new_n19017_, new_n19018_, new_n19019_,
    new_n19020_, new_n19021_, new_n19022_, new_n19023_, new_n19024_,
    new_n19025_, new_n19026_, new_n19027_, new_n19028_, new_n19029_,
    new_n19030_, new_n19031_, new_n19032_, new_n19033_, new_n19034_,
    new_n19035_, new_n19036_, new_n19037_, new_n19038_, new_n19039_,
    new_n19040_, new_n19041_, new_n19042_, new_n19043_, new_n19044_,
    new_n19045_, new_n19046_, new_n19047_, new_n19048_, new_n19049_,
    new_n19050_, new_n19051_, new_n19052_, new_n19053_, new_n19054_,
    new_n19055_, new_n19056_, new_n19057_, new_n19058_, new_n19059_,
    new_n19060_, new_n19061_, new_n19062_, new_n19063_, new_n19064_,
    new_n19065_, new_n19066_, new_n19067_, new_n19068_, new_n19069_,
    new_n19070_, new_n19071_, new_n19072_, new_n19073_, new_n19074_,
    new_n19075_, new_n19076_, new_n19077_, new_n19078_, new_n19079_,
    new_n19080_, new_n19081_, new_n19082_, new_n19083_, new_n19084_,
    new_n19085_, new_n19086_, new_n19087_, new_n19088_, new_n19089_,
    new_n19090_, new_n19091_, new_n19092_, new_n19093_, new_n19094_,
    new_n19095_, new_n19096_, new_n19097_, new_n19098_, new_n19099_,
    new_n19100_, new_n19101_, new_n19102_, new_n19103_, new_n19104_,
    new_n19105_, new_n19106_, new_n19107_, new_n19108_, new_n19109_,
    new_n19110_, new_n19111_, new_n19112_, new_n19113_, new_n19114_,
    new_n19115_, new_n19116_, new_n19117_, new_n19118_, new_n19119_,
    new_n19120_, new_n19121_, new_n19122_, new_n19123_, new_n19124_,
    new_n19125_, new_n19126_, new_n19127_, new_n19128_, new_n19129_,
    new_n19130_, new_n19131_, new_n19132_, new_n19133_, new_n19134_,
    new_n19135_, new_n19136_, new_n19137_, new_n19138_, new_n19139_,
    new_n19140_, new_n19141_, new_n19142_, new_n19143_, new_n19144_,
    new_n19145_, new_n19146_, new_n19147_, new_n19148_, new_n19149_,
    new_n19150_, new_n19151_, new_n19152_, new_n19153_, new_n19154_,
    new_n19155_, new_n19156_, new_n19157_, new_n19158_, new_n19159_,
    new_n19160_, new_n19161_, new_n19162_, new_n19163_, new_n19164_,
    new_n19165_, new_n19166_, new_n19167_, new_n19168_, new_n19169_,
    new_n19170_, new_n19171_, new_n19172_, new_n19173_, new_n19174_,
    new_n19175_, new_n19176_, new_n19177_, new_n19178_, new_n19179_,
    new_n19180_, new_n19181_, new_n19182_, new_n19183_, new_n19184_,
    new_n19185_, new_n19186_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19278_, new_n19279_, new_n19280_,
    new_n19281_, new_n19282_, new_n19283_, new_n19284_, new_n19285_,
    new_n19286_, new_n19287_, new_n19288_, new_n19289_, new_n19290_,
    new_n19291_, new_n19292_, new_n19293_, new_n19294_, new_n19295_,
    new_n19296_, new_n19297_, new_n19298_, new_n19299_, new_n19300_,
    new_n19301_, new_n19302_, new_n19303_, new_n19304_, new_n19305_,
    new_n19306_, new_n19307_, new_n19308_, new_n19309_, new_n19310_,
    new_n19311_, new_n19312_, new_n19313_, new_n19314_, new_n19315_,
    new_n19316_, new_n19317_, new_n19318_, new_n19319_, new_n19320_,
    new_n19321_, new_n19322_, new_n19323_, new_n19324_, new_n19325_,
    new_n19326_, new_n19327_, new_n19328_, new_n19329_, new_n19330_,
    new_n19331_, new_n19332_, new_n19333_, new_n19334_, new_n19335_,
    new_n19336_, new_n19337_, new_n19338_, new_n19339_, new_n19340_,
    new_n19341_, new_n19342_, new_n19343_, new_n19344_, new_n19345_,
    new_n19346_, new_n19347_, new_n19348_, new_n19349_, new_n19350_,
    new_n19351_, new_n19352_, new_n19353_, new_n19354_, new_n19355_,
    new_n19356_, new_n19357_, new_n19358_, new_n19359_, new_n19360_,
    new_n19361_, new_n19362_, new_n19363_, new_n19364_, new_n19365_,
    new_n19366_, new_n19367_, new_n19368_, new_n19369_, new_n19370_,
    new_n19371_, new_n19372_, new_n19373_, new_n19374_, new_n19375_,
    new_n19376_, new_n19377_, new_n19378_, new_n19379_, new_n19380_,
    new_n19381_, new_n19382_, new_n19383_, new_n19384_, new_n19385_,
    new_n19386_, new_n19387_, new_n19388_, new_n19389_, new_n19390_,
    new_n19391_, new_n19392_, new_n19393_, new_n19394_, new_n19395_,
    new_n19396_, new_n19397_, new_n19398_, new_n19399_, new_n19400_,
    new_n19401_, new_n19402_, new_n19403_, new_n19404_, new_n19405_,
    new_n19406_, new_n19407_, new_n19408_, new_n19409_, new_n19410_,
    new_n19411_, new_n19412_, new_n19413_, new_n19414_, new_n19415_,
    new_n19416_, new_n19417_, new_n19418_, new_n19419_, new_n19420_,
    new_n19421_, new_n19422_, new_n19423_, new_n19424_, new_n19425_,
    new_n19426_, new_n19427_, new_n19428_, new_n19429_, new_n19430_,
    new_n19431_, new_n19432_, new_n19433_, new_n19434_, new_n19435_,
    new_n19436_, new_n19437_, new_n19438_, new_n19439_, new_n19440_,
    new_n19441_, new_n19442_, new_n19443_, new_n19444_, new_n19445_,
    new_n19446_, new_n19447_, new_n19448_, new_n19449_, new_n19450_,
    new_n19451_, new_n19452_, new_n19453_, new_n19454_, new_n19455_,
    new_n19456_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19637_, new_n19638_, new_n19639_, new_n19640_, new_n19641_,
    new_n19642_, new_n19645_, new_n19646_, new_n19647_, new_n19648_,
    new_n19649_, new_n19650_, new_n19651_, new_n19652_, new_n19653_,
    new_n19654_, new_n19655_, new_n19656_, new_n19657_, new_n19658_,
    new_n19659_, new_n19660_, new_n19661_, new_n19662_, new_n19663_,
    new_n19664_, new_n19665_, new_n19666_, new_n19667_, new_n19668_,
    new_n19669_, new_n19670_, new_n19671_, new_n19672_, new_n19673_,
    new_n19674_, new_n19675_, new_n19676_, new_n19677_, new_n19678_,
    new_n19679_, new_n19680_, new_n19681_, new_n19682_, new_n19683_,
    new_n19684_, new_n19689_, new_n19690_, new_n19691_, new_n19692_,
    new_n19693_, new_n19694_, new_n19695_, new_n19696_, new_n19697_,
    new_n19698_, new_n19699_, new_n19700_, new_n19701_, new_n19702_,
    new_n19703_, new_n19704_, new_n19705_, new_n19706_, new_n19707_,
    new_n19708_, new_n19709_, new_n19710_, new_n19711_, new_n19712_,
    new_n19713_, new_n19714_, new_n19715_, new_n19716_, new_n19717_,
    new_n19718_, new_n19719_, new_n19720_, new_n19721_, new_n19722_,
    new_n19723_, new_n19724_, new_n19725_, new_n19726_, new_n19727_,
    new_n19728_, new_n19729_, new_n19730_, new_n19731_, new_n19732_,
    new_n19733_, new_n19734_, new_n19735_, new_n19736_, new_n19737_,
    new_n19738_, new_n19739_, new_n19740_, new_n19741_, new_n19742_,
    new_n19743_, new_n19744_, new_n19745_, new_n19746_, new_n19747_,
    new_n19748_, new_n19749_, new_n19750_, new_n19751_, new_n19752_,
    new_n19753_, new_n19754_, new_n19755_, new_n19756_, new_n19757_,
    new_n19758_, new_n19759_, new_n19760_, new_n19761_, new_n19762_,
    new_n19763_, new_n19764_, new_n19765_, new_n19766_, new_n19767_,
    new_n19768_, new_n19769_, new_n19770_, new_n19771_, new_n19772_,
    new_n19773_, new_n19774_, new_n19775_, new_n19776_, new_n19777_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19800_, new_n19801_, new_n19802_,
    new_n19805_, new_n19806_, new_n19807_, new_n19808_, new_n19809_,
    new_n19810_, new_n19811_, new_n19812_, new_n19813_, new_n19814_,
    new_n19815_, new_n19816_, new_n19817_, new_n19818_, new_n19819_,
    new_n19820_, new_n19821_, new_n19822_, new_n19823_, new_n19824_,
    new_n19825_, new_n19826_, new_n19827_, new_n19828_, new_n19829_,
    new_n19830_, new_n19831_, new_n19832_, new_n19833_, new_n19834_,
    new_n19835_, new_n19836_, new_n19837_, new_n19838_, new_n19839_,
    new_n19840_, new_n19841_, new_n19842_, new_n19843_, new_n19844_,
    new_n19845_, new_n19846_, new_n19847_, new_n19848_, new_n19849_,
    new_n19850_, new_n19851_, new_n19852_, new_n19853_, new_n19854_,
    new_n19855_, new_n19856_, new_n19857_, new_n19858_, new_n19859_,
    new_n19860_, new_n19861_, new_n19862_, new_n19863_, new_n19864_,
    new_n19865_, new_n19866_, new_n19867_, new_n19868_, new_n19869_,
    new_n19870_, new_n19871_, new_n19872_, new_n19873_, new_n19874_,
    new_n19875_, new_n19876_, new_n19877_, new_n19878_, new_n19879_,
    new_n19880_, new_n19881_, new_n19882_, new_n19883_, new_n19884_,
    new_n19885_, new_n19886_, new_n19887_, new_n19888_, new_n19889_,
    new_n19890_, new_n19891_, new_n19892_, new_n19893_, new_n19894_,
    new_n19895_, new_n19896_, new_n19897_, new_n19898_, new_n19899_,
    new_n19900_, new_n19901_, new_n19902_, new_n19903_, new_n19904_,
    new_n19905_, new_n19906_, new_n19907_, new_n19908_, new_n19909_,
    new_n19910_, new_n19911_, new_n19912_, new_n19913_, new_n19914_,
    new_n19915_, new_n19916_, new_n19917_, new_n19918_, new_n19919_,
    new_n19920_, new_n19921_, new_n19922_, new_n19923_, new_n19924_,
    new_n19925_, new_n19926_, new_n19927_, new_n19928_, new_n19929_,
    new_n19930_, new_n19931_, new_n19932_, new_n19933_, new_n19934_,
    new_n19935_, new_n19936_, new_n19937_, new_n19938_, new_n19939_,
    new_n19940_, new_n19941_, new_n19942_, new_n19943_, new_n19944_,
    new_n19945_, new_n19946_, new_n19947_, new_n19948_, new_n19949_,
    new_n19950_, new_n19951_, new_n19952_, new_n19953_, new_n19954_,
    new_n19955_, new_n19956_, new_n19957_, new_n19958_, new_n19959_,
    new_n19960_, new_n19961_, new_n19962_, new_n19963_, new_n19964_,
    new_n19965_, new_n19966_, new_n19967_, new_n19968_, new_n19969_,
    new_n19970_, new_n19971_, new_n19972_, new_n19973_, new_n19974_,
    new_n19975_, new_n19976_, new_n19977_, new_n19978_, new_n19979_,
    new_n19980_, new_n19981_, new_n19982_, new_n19983_, new_n19984_,
    new_n19985_, new_n19986_, new_n19987_, new_n19988_, new_n19989_,
    new_n19990_, new_n19991_, new_n19992_, new_n19993_, new_n19994_,
    new_n19995_, new_n19996_, new_n19997_, new_n19998_, new_n19999_,
    new_n20000_, new_n20001_, new_n20003_, new_n20004_, new_n20005_,
    new_n20006_, new_n20007_, new_n20008_, new_n20009_, new_n20010_,
    new_n20011_, new_n20012_, new_n20013_, new_n20014_, new_n20015_,
    new_n20016_, new_n20017_, new_n20018_, new_n20019_, new_n20020_,
    new_n20021_, new_n20022_, new_n20023_, new_n20024_, new_n20025_,
    new_n20026_, new_n20027_, new_n20028_, new_n20029_, new_n20030_,
    new_n20031_, new_n20032_, new_n20033_, new_n20034_, new_n20035_,
    new_n20036_, new_n20037_, new_n20038_, new_n20039_, new_n20040_,
    new_n20041_, new_n20042_, new_n20043_, new_n20044_, new_n20045_,
    new_n20046_, new_n20047_, new_n20048_, new_n20049_, new_n20050_,
    new_n20051_, new_n20052_, new_n20053_, new_n20054_, new_n20055_,
    new_n20056_, new_n20057_, new_n20058_, new_n20059_, new_n20060_,
    new_n20061_, new_n20062_, new_n20063_, new_n20064_, new_n20065_,
    new_n20066_, new_n20067_, new_n20068_, new_n20069_, new_n20070_,
    new_n20071_, new_n20072_, new_n20073_, new_n20074_, new_n20075_,
    new_n20076_, new_n20077_, new_n20078_, new_n20079_, new_n20080_,
    new_n20081_, new_n20082_, new_n20083_, new_n20084_, new_n20085_,
    new_n20086_, new_n20087_, new_n20088_, new_n20089_, new_n20090_,
    new_n20091_, new_n20092_, new_n20093_, new_n20094_, new_n20095_,
    new_n20096_, new_n20097_, new_n20098_, new_n20099_, new_n20100_,
    new_n20101_, new_n20102_, new_n20103_, new_n20104_, new_n20105_,
    new_n20106_, new_n20107_, new_n20108_, new_n20109_, new_n20110_,
    new_n20111_, new_n20112_, new_n20113_, new_n20114_, new_n20115_,
    new_n20116_, new_n20117_, new_n20118_, new_n20119_, new_n20120_,
    new_n20121_, new_n20122_, new_n20123_, new_n20124_, new_n20125_,
    new_n20126_, new_n20127_, new_n20128_, new_n20129_, new_n20130_,
    new_n20131_, new_n20132_, new_n20133_, new_n20134_, new_n20135_,
    new_n20136_, new_n20137_, new_n20138_, new_n20139_, new_n20140_,
    new_n20141_, new_n20142_, new_n20143_, new_n20144_, new_n20145_,
    new_n20146_, new_n20147_, new_n20148_, new_n20149_, new_n20150_,
    new_n20151_, new_n20152_, new_n20153_, new_n20154_, new_n20155_,
    new_n20156_, new_n20157_, new_n20158_, new_n20159_, new_n20160_,
    new_n20161_, new_n20162_, new_n20163_, new_n20164_, new_n20165_,
    new_n20166_, new_n20167_, new_n20168_, new_n20169_, new_n20170_,
    new_n20171_, new_n20172_, new_n20173_, new_n20174_, new_n20175_,
    new_n20176_, new_n20177_, new_n20178_, new_n20179_, new_n20180_,
    new_n20181_, new_n20182_, new_n20183_, new_n20184_, new_n20185_,
    new_n20186_, new_n20187_, new_n20188_, new_n20189_, new_n20190_,
    new_n20191_, new_n20192_, new_n20193_, new_n20194_, new_n20195_,
    new_n20196_, new_n20197_, new_n20198_, new_n20199_, new_n20200_,
    new_n20201_, new_n20202_, new_n20203_, new_n20204_, new_n20205_,
    new_n20206_, new_n20207_, new_n20208_, new_n20209_, new_n20210_,
    new_n20211_, new_n20212_, new_n20213_, new_n20214_, new_n20215_,
    new_n20216_, new_n20217_, new_n20218_, new_n20219_, new_n20220_,
    new_n20221_, new_n20222_, new_n20223_, new_n20224_, new_n20225_,
    new_n20226_, new_n20227_, new_n20228_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20305_, new_n20306_, new_n20307_, new_n20308_, new_n20309_,
    new_n20310_, new_n20311_, new_n20312_, new_n20313_, new_n20314_,
    new_n20315_, new_n20316_, new_n20317_, new_n20318_, new_n20319_,
    new_n20320_, new_n20321_, new_n20322_, new_n20323_, new_n20324_,
    new_n20325_, new_n20326_, new_n20327_, new_n20328_, new_n20329_,
    new_n20330_, new_n20331_, new_n20332_, new_n20333_, new_n20334_,
    new_n20335_, new_n20336_, new_n20337_, new_n20338_, new_n20339_,
    new_n20340_, new_n20341_, new_n20342_, new_n20343_, new_n20344_,
    new_n20345_, new_n20346_, new_n20347_, new_n20348_, new_n20349_,
    new_n20350_, new_n20351_, new_n20352_, new_n20353_, new_n20354_,
    new_n20355_, new_n20356_, new_n20357_, new_n20358_, new_n20359_,
    new_n20360_, new_n20361_, new_n20362_, new_n20363_, new_n20364_,
    new_n20365_, new_n20366_, new_n20367_, new_n20368_, new_n20369_,
    new_n20370_, new_n20371_, new_n20373_, new_n20374_, new_n20375_,
    new_n20376_, new_n20377_, new_n20378_, new_n20379_, new_n20380_,
    new_n20381_, new_n20382_, new_n20383_, new_n20384_, new_n20385_,
    new_n20386_, new_n20387_, new_n20388_, new_n20389_, new_n20390_,
    new_n20391_, new_n20392_, new_n20393_, new_n20397_, new_n20398_,
    new_n20399_, new_n20400_, new_n20401_, new_n20402_, new_n20403_,
    new_n20404_, new_n20405_, new_n20406_, new_n20407_, new_n20408_,
    new_n20409_, new_n20412_, new_n20413_, new_n20414_, new_n20415_,
    new_n20416_, new_n20417_, new_n20418_, new_n20419_, new_n20420_,
    new_n20421_, new_n20422_, new_n20423_, new_n20424_, new_n20425_,
    new_n20426_, new_n20427_, new_n20428_, new_n20429_, new_n20430_,
    new_n20431_, new_n20432_, new_n20433_, new_n20434_, new_n20435_,
    new_n20436_, new_n20437_, new_n20438_, new_n20439_, new_n20440_,
    new_n20441_, new_n20442_, new_n20443_, new_n20444_, new_n20445_,
    new_n20446_, new_n20447_, new_n20448_, new_n20449_, new_n20450_,
    new_n20451_, new_n20452_, new_n20453_, new_n20454_, new_n20455_,
    new_n20456_, new_n20457_, new_n20458_, new_n20459_, new_n20460_,
    new_n20461_, new_n20462_, new_n20463_, new_n20464_, new_n20465_,
    new_n20466_, new_n20467_, new_n20468_, new_n20469_, new_n20470_,
    new_n20471_, new_n20472_, new_n20473_, new_n20474_, new_n20475_,
    new_n20476_, new_n20477_, new_n20478_, new_n20479_, new_n20480_,
    new_n20481_, new_n20482_, new_n20483_, new_n20484_, new_n20485_,
    new_n20486_, new_n20487_, new_n20488_, new_n20489_, new_n20490_,
    new_n20491_, new_n20492_, new_n20493_, new_n20494_, new_n20495_,
    new_n20496_, new_n20497_, new_n20502_, new_n20503_, new_n20504_,
    new_n20505_, new_n20506_, new_n20507_, new_n20508_, new_n20509_,
    new_n20510_, new_n20511_, new_n20512_, new_n20513_, new_n20514_,
    new_n20515_, new_n20516_, new_n20517_, new_n20518_, new_n20519_,
    new_n20520_, new_n20523_, new_n20524_, new_n20525_, new_n20526_,
    new_n20527_, new_n20528_, new_n20529_, new_n20530_, new_n20531_,
    new_n20532_, new_n20533_, new_n20534_, new_n20535_, new_n20536_,
    new_n20537_, new_n20538_, new_n20539_, new_n20540_, new_n20541_,
    new_n20542_, new_n20543_, new_n20544_, new_n20545_, new_n20546_,
    new_n20547_, new_n20548_, new_n20549_, new_n20550_, new_n20551_,
    new_n20552_, new_n20553_, new_n20554_, new_n20555_, new_n20556_,
    new_n20557_, new_n20558_, new_n20559_, new_n20560_, new_n20561_,
    new_n20562_, new_n20563_, new_n20564_, new_n20565_, new_n20566_,
    new_n20567_, new_n20568_, new_n20569_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20679_, new_n20680_, new_n20681_,
    new_n20682_, new_n20683_, new_n20684_, new_n20685_, new_n20686_,
    new_n20687_, new_n20688_, new_n20689_, new_n20690_, new_n20691_,
    new_n20692_, new_n20693_, new_n20694_, new_n20695_, new_n20696_,
    new_n20697_, new_n20698_, new_n20699_, new_n20700_, new_n20701_,
    new_n20702_, new_n20703_, new_n20704_, new_n20705_, new_n20706_,
    new_n20707_, new_n20708_, new_n20709_, new_n20710_, new_n20711_,
    new_n20712_, new_n20713_, new_n20714_, new_n20715_, new_n20716_,
    new_n20717_, new_n20718_, new_n20720_, new_n20721_, new_n20722_,
    new_n20723_, new_n20724_, new_n20725_, new_n20726_, new_n20727_,
    new_n20728_, new_n20729_, new_n20730_, new_n20731_, new_n20732_,
    new_n20733_, new_n20734_, new_n20735_, new_n20736_, new_n20737_,
    new_n20738_, new_n20739_, new_n20740_, new_n20741_, new_n20742_,
    new_n20743_, new_n20744_, new_n20745_, new_n20746_, new_n20747_,
    new_n20748_, new_n20749_, new_n20750_, new_n20751_, new_n20752_,
    new_n20753_, new_n20754_, new_n20755_, new_n20756_, new_n20757_,
    new_n20758_, new_n20759_, new_n20760_, new_n20761_, new_n20762_,
    new_n20763_, new_n20764_, new_n20765_, new_n20766_, new_n20767_,
    new_n20768_, new_n20769_, new_n20770_, new_n20771_, new_n20772_,
    new_n20773_, new_n20774_, new_n20775_, new_n20776_, new_n20777_,
    new_n20778_, new_n20779_, new_n20780_, new_n20781_, new_n20782_,
    new_n20783_, new_n20784_, new_n20785_, new_n20786_, new_n20787_,
    new_n20788_, new_n20789_, new_n20790_, new_n20791_, new_n20792_,
    new_n20793_, new_n20794_, new_n20795_, new_n20796_, new_n20797_,
    new_n20798_, new_n20799_, new_n20800_, new_n20801_, new_n20802_,
    new_n20803_, new_n20804_, new_n20805_, new_n20806_, new_n20807_,
    new_n20808_, new_n20809_, new_n20810_, new_n20811_, new_n20812_,
    new_n20813_, new_n20814_, new_n20815_, new_n20816_, new_n20817_,
    new_n20818_, new_n20819_, new_n20820_, new_n20821_, new_n20822_,
    new_n20823_, new_n20824_, new_n20825_, new_n20826_, new_n20827_,
    new_n20828_, new_n20829_, new_n20830_, new_n20831_, new_n20832_,
    new_n20833_, new_n20834_, new_n20835_, new_n20836_, new_n20837_,
    new_n20838_, new_n20839_, new_n20840_, new_n20841_, new_n20842_,
    new_n20843_, new_n20844_, new_n20845_, new_n20846_, new_n20847_,
    new_n20848_, new_n20849_, new_n20850_, new_n20851_, new_n20852_,
    new_n20853_, new_n20854_, new_n20855_, new_n20856_, new_n20857_,
    new_n20858_, new_n20859_, new_n20860_, new_n20861_, new_n20862_,
    new_n20863_, new_n20864_, new_n20865_, new_n20866_, new_n20867_,
    new_n20868_, new_n20869_, new_n20870_, new_n20871_, new_n20872_,
    new_n20873_, new_n20874_, new_n20875_, new_n20876_, new_n20877_,
    new_n20878_, new_n20879_, new_n20880_, new_n20881_, new_n20882_,
    new_n20883_, new_n20884_, new_n20885_, new_n20886_, new_n20887_,
    new_n20888_, new_n20889_, new_n20890_, new_n20891_, new_n20892_,
    new_n20893_, new_n20894_, new_n20895_, new_n20896_, new_n20897_,
    new_n20898_, new_n20899_, new_n20900_, new_n20901_, new_n20902_,
    new_n20903_, new_n20904_, new_n20905_, new_n20906_, new_n20907_,
    new_n20908_, new_n20909_, new_n20910_, new_n20911_, new_n20912_,
    new_n20913_, new_n20914_, new_n20915_, new_n20916_, new_n20917_,
    new_n20918_, new_n20919_, new_n20920_, new_n20921_, new_n20922_,
    new_n20923_, new_n20924_, new_n20925_, new_n20926_, new_n20927_,
    new_n20928_, new_n20929_, new_n20930_, new_n20931_, new_n20932_,
    new_n20933_, new_n20934_, new_n20935_, new_n20936_, new_n20937_,
    new_n20938_, new_n20939_, new_n20940_, new_n20941_, new_n20942_,
    new_n20943_, new_n20944_, new_n20945_, new_n20946_, new_n20947_,
    new_n20948_, new_n20949_, new_n20950_, new_n20951_, new_n20952_,
    new_n20953_, new_n20954_, new_n20955_, new_n20956_, new_n20957_,
    new_n20958_, new_n20959_, new_n20960_, new_n20961_, new_n20962_,
    new_n20963_, new_n20964_, new_n20965_, new_n20966_, new_n20967_,
    new_n20968_, new_n20969_, new_n20970_, new_n20971_, new_n20972_,
    new_n20973_, new_n20974_, new_n20975_, new_n20976_, new_n20977_,
    new_n20978_, new_n20979_, new_n20980_, new_n20981_, new_n20982_,
    new_n20983_, new_n20984_, new_n20985_, new_n20986_, new_n20987_,
    new_n20988_, new_n20989_, new_n20990_, new_n20991_, new_n20992_,
    new_n20993_, new_n20994_, new_n20995_, new_n20996_, new_n20997_,
    new_n20998_, new_n20999_, new_n21000_, new_n21001_, new_n21002_,
    new_n21003_, new_n21004_, new_n21005_, new_n21006_, new_n21007_,
    new_n21008_, new_n21009_, new_n21010_, new_n21011_, new_n21012_,
    new_n21013_, new_n21014_, new_n21015_, new_n21016_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21074_, new_n21075_,
    new_n21076_, new_n21077_, new_n21078_, new_n21079_, new_n21080_,
    new_n21081_, new_n21082_, new_n21083_, new_n21084_, new_n21085_,
    new_n21086_, new_n21087_, new_n21088_, new_n21089_, new_n21090_,
    new_n21091_, new_n21092_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21101_,
    new_n21102_, new_n21103_, new_n21104_, new_n21105_, new_n21106_,
    new_n21107_, new_n21108_, new_n21109_, new_n21110_, new_n21111_,
    new_n21112_, new_n21113_, new_n21114_, new_n21115_, new_n21116_,
    new_n21117_, new_n21118_, new_n21119_, new_n21120_, new_n21121_,
    new_n21122_, new_n21123_, new_n21124_, new_n21125_, new_n21126_,
    new_n21127_, new_n21128_, new_n21129_, new_n21130_, new_n21131_,
    new_n21132_, new_n21133_, new_n21134_, new_n21135_, new_n21136_,
    new_n21137_, new_n21138_, new_n21139_, new_n21140_, new_n21141_,
    new_n21142_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21178_, new_n21179_, new_n21180_, new_n21181_,
    new_n21182_, new_n21183_, new_n21184_, new_n21185_, new_n21186_,
    new_n21187_, new_n21188_, new_n21189_, new_n21190_, new_n21191_,
    new_n21192_, new_n21193_, new_n21194_, new_n21195_, new_n21196_,
    new_n21197_, new_n21198_, new_n21199_, new_n21200_, new_n21201_,
    new_n21202_, new_n21203_, new_n21204_, new_n21205_, new_n21206_,
    new_n21207_, new_n21208_, new_n21209_, new_n21210_, new_n21211_,
    new_n21212_, new_n21213_, new_n21214_, new_n21215_, new_n21216_,
    new_n21217_, new_n21218_, new_n21219_, new_n21220_, new_n21221_,
    new_n21222_, new_n21223_, new_n21224_, new_n21225_, new_n21226_,
    new_n21227_, new_n21228_, new_n21229_, new_n21230_, new_n21231_,
    new_n21232_, new_n21233_, new_n21234_, new_n21235_, new_n21236_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21377_, new_n21378_, new_n21379_, new_n21380_, new_n21381_,
    new_n21382_, new_n21383_, new_n21384_, new_n21385_, new_n21386_,
    new_n21387_, new_n21388_, new_n21389_, new_n21390_, new_n21391_,
    new_n21392_, new_n21393_, new_n21394_, new_n21395_, new_n21399_,
    new_n21400_, new_n21401_, new_n21402_, new_n21403_, new_n21404_,
    new_n21405_, new_n21406_, new_n21407_, new_n21408_, new_n21409_,
    new_n21410_, new_n21411_, new_n21412_, new_n21413_, new_n21414_,
    new_n21415_, new_n21416_, new_n21417_, new_n21418_, new_n21419_,
    new_n21420_, new_n21421_, new_n21422_, new_n21423_, new_n21424_,
    new_n21425_, new_n21426_, new_n21427_, new_n21428_, new_n21429_,
    new_n21430_, new_n21431_, new_n21432_, new_n21433_, new_n21434_,
    new_n21435_, new_n21436_, new_n21437_, new_n21438_, new_n21439_,
    new_n21440_, new_n21441_, new_n21442_, new_n21443_, new_n21444_,
    new_n21445_, new_n21446_, new_n21447_, new_n21448_, new_n21449_,
    new_n21450_, new_n21451_, new_n21452_, new_n21453_, new_n21454_,
    new_n21455_, new_n21456_, new_n21457_, new_n21458_, new_n21459_,
    new_n21460_, new_n21461_, new_n21462_, new_n21463_, new_n21464_,
    new_n21465_, new_n21466_, new_n21467_, new_n21468_, new_n21469_,
    new_n21470_, new_n21471_, new_n21472_, new_n21473_, new_n21474_,
    new_n21475_, new_n21476_, new_n21477_, new_n21478_, new_n21480_,
    new_n21481_, new_n21482_, new_n21483_, new_n21484_, new_n21485_,
    new_n21486_, new_n21487_, new_n21488_, new_n21489_, new_n21490_,
    new_n21491_, new_n21492_, new_n21493_, new_n21494_, new_n21495_,
    new_n21496_, new_n21497_, new_n21498_, new_n21499_, new_n21500_,
    new_n21501_, new_n21502_, new_n21503_, new_n21504_, new_n21505_,
    new_n21506_, new_n21507_, new_n21508_, new_n21509_, new_n21510_,
    new_n21511_, new_n21512_, new_n21513_, new_n21514_, new_n21515_,
    new_n21516_, new_n21517_, new_n21518_, new_n21519_, new_n21520_,
    new_n21521_, new_n21522_, new_n21523_, new_n21524_, new_n21525_,
    new_n21526_, new_n21527_, new_n21528_, new_n21529_, new_n21530_,
    new_n21531_, new_n21532_, new_n21533_, new_n21534_, new_n21535_,
    new_n21536_, new_n21537_, new_n21538_, new_n21539_, new_n21540_,
    new_n21541_, new_n21542_, new_n21543_, new_n21544_, new_n21545_,
    new_n21546_, new_n21547_, new_n21548_, new_n21549_, new_n21550_,
    new_n21551_, new_n21552_, new_n21553_, new_n21554_, new_n21555_,
    new_n21556_, new_n21557_, new_n21558_, new_n21559_, new_n21560_,
    new_n21561_, new_n21562_, new_n21563_, new_n21564_, new_n21565_,
    new_n21566_, new_n21567_, new_n21568_, new_n21569_, new_n21570_,
    new_n21571_, new_n21572_, new_n21573_, new_n21574_, new_n21575_,
    new_n21576_, new_n21577_, new_n21578_, new_n21579_, new_n21580_,
    new_n21581_, new_n21582_, new_n21583_, new_n21584_, new_n21585_,
    new_n21586_, new_n21587_, new_n21588_, new_n21589_, new_n21590_,
    new_n21591_, new_n21592_, new_n21593_, new_n21594_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21602_, new_n21603_, new_n21604_, new_n21605_,
    new_n21606_, new_n21607_, new_n21608_, new_n21609_, new_n21610_,
    new_n21611_, new_n21612_, new_n21613_, new_n21614_, new_n21615_,
    new_n21616_, new_n21617_, new_n21618_, new_n21619_, new_n21620_,
    new_n21621_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21630_,
    new_n21631_, new_n21632_, new_n21633_, new_n21634_, new_n21635_,
    new_n21636_, new_n21637_, new_n21638_, new_n21639_, new_n21640_,
    new_n21641_, new_n21642_, new_n21643_, new_n21644_, new_n21645_,
    new_n21646_, new_n21647_, new_n21648_, new_n21649_, new_n21650_,
    new_n21651_, new_n21652_, new_n21653_, new_n21654_, new_n21655_,
    new_n21656_, new_n21657_, new_n21658_, new_n21659_, new_n21660_,
    new_n21661_, new_n21662_, new_n21663_, new_n21664_, new_n21665_,
    new_n21666_, new_n21667_, new_n21668_, new_n21669_, new_n21670_,
    new_n21671_, new_n21672_, new_n21673_, new_n21674_, new_n21675_,
    new_n21676_, new_n21677_, new_n21678_, new_n21679_, new_n21680_,
    new_n21681_, new_n21682_, new_n21683_, new_n21684_, new_n21685_,
    new_n21686_, new_n21687_, new_n21688_, new_n21689_, new_n21690_,
    new_n21691_, new_n21692_, new_n21693_, new_n21694_, new_n21695_,
    new_n21696_, new_n21697_, new_n21698_, new_n21699_, new_n21700_,
    new_n21701_, new_n21702_, new_n21704_, new_n21705_, new_n21706_,
    new_n21707_, new_n21708_, new_n21709_, new_n21710_, new_n21711_,
    new_n21712_, new_n21713_, new_n21714_, new_n21715_, new_n21716_,
    new_n21717_, new_n21718_, new_n21719_, new_n21720_, new_n21721_,
    new_n21722_, new_n21723_, new_n21724_, new_n21725_, new_n21726_,
    new_n21727_, new_n21728_, new_n21729_, new_n21730_, new_n21731_,
    new_n21732_, new_n21733_, new_n21734_, new_n21735_, new_n21736_,
    new_n21737_, new_n21738_, new_n21739_, new_n21740_, new_n21741_,
    new_n21742_, new_n21743_, new_n21744_, new_n21745_, new_n21746_,
    new_n21747_, new_n21748_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21779_,
    new_n21780_, new_n21781_, new_n21782_, new_n21783_, new_n21784_,
    new_n21785_, new_n21786_, new_n21787_, new_n21788_, new_n21789_,
    new_n21790_, new_n21791_, new_n21792_, new_n21793_, new_n21794_,
    new_n21795_, new_n21796_, new_n21797_, new_n21798_, new_n21799_,
    new_n21800_, new_n21801_, new_n21802_, new_n21803_, new_n21804_,
    new_n21805_, new_n21806_, new_n21807_, new_n21808_, new_n21809_,
    new_n21810_, new_n21811_, new_n21812_, new_n21813_, new_n21814_,
    new_n21815_, new_n21816_, new_n21817_, new_n21818_, new_n21819_,
    new_n21820_, new_n21821_, new_n21822_, new_n21823_, new_n21824_,
    new_n21825_, new_n21826_, new_n21827_, new_n21828_, new_n21829_,
    new_n21830_, new_n21831_, new_n21832_, new_n21833_, new_n21834_,
    new_n21835_, new_n21836_, new_n21837_, new_n21838_, new_n21839_,
    new_n21840_, new_n21841_, new_n21842_, new_n21843_, new_n21844_,
    new_n21845_, new_n21847_, new_n21848_, new_n21849_, new_n21850_,
    new_n21851_, new_n21852_, new_n21853_, new_n21854_, new_n21855_,
    new_n21856_, new_n21857_, new_n21858_, new_n21859_, new_n21860_,
    new_n21861_, new_n21862_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21880_,
    new_n21881_, new_n21882_, new_n21883_, new_n21884_, new_n21885_,
    new_n21886_, new_n21887_, new_n21888_, new_n21889_, new_n21890_,
    new_n21891_, new_n21892_, new_n21893_, new_n21894_, new_n21895_,
    new_n21896_, new_n21897_, new_n21898_, new_n21899_, new_n21900_,
    new_n21901_, new_n21902_, new_n21903_, new_n21904_, new_n21905_,
    new_n21906_, new_n21907_, new_n21908_, new_n21909_, new_n21910_,
    new_n21911_, new_n21912_, new_n21913_, new_n21914_, new_n21915_,
    new_n21916_, new_n21917_, new_n21918_, new_n21919_, new_n21920_,
    new_n21921_, new_n21922_, new_n21923_, new_n21924_, new_n21925_,
    new_n21926_, new_n21927_, new_n21928_, new_n21929_, new_n21930_,
    new_n21931_, new_n21932_, new_n21933_, new_n21934_, new_n21935_,
    new_n21936_, new_n21937_, new_n21938_, new_n21939_, new_n21940_,
    new_n21941_, new_n21942_, new_n21943_, new_n21944_, new_n21945_,
    new_n21946_, new_n21947_, new_n21948_, new_n21949_, new_n21950_,
    new_n21951_, new_n21952_, new_n21953_, new_n21954_, new_n21955_,
    new_n21956_, new_n21957_, new_n21958_, new_n21959_, new_n21960_,
    new_n21961_, new_n21962_, new_n21963_, new_n21964_, new_n21965_,
    new_n21966_, new_n21967_, new_n21968_, new_n21969_, new_n21970_,
    new_n21971_, new_n21972_, new_n21973_, new_n21974_, new_n21975_,
    new_n21976_, new_n21977_, new_n21978_, new_n21979_, new_n21980_,
    new_n21981_, new_n21982_, new_n21983_, new_n21984_, new_n21985_,
    new_n21986_, new_n21987_, new_n21988_, new_n21989_, new_n21990_,
    new_n21991_, new_n21992_, new_n21993_, new_n21994_, new_n21995_,
    new_n21996_, new_n21997_, new_n21998_, new_n21999_, new_n22000_,
    new_n22001_, new_n22002_, new_n22003_, new_n22004_, new_n22005_,
    new_n22006_, new_n22007_, new_n22008_, new_n22009_, new_n22010_,
    new_n22011_, new_n22012_, new_n22013_, new_n22014_, new_n22015_,
    new_n22016_, new_n22017_, new_n22018_, new_n22019_, new_n22020_,
    new_n22021_, new_n22022_, new_n22023_, new_n22024_, new_n22025_,
    new_n22026_, new_n22027_, new_n22028_, new_n22029_, new_n22030_,
    new_n22031_, new_n22032_, new_n22033_, new_n22034_, new_n22035_,
    new_n22036_, new_n22037_, new_n22038_, new_n22039_, new_n22040_,
    new_n22041_, new_n22042_, new_n22043_, new_n22044_, new_n22045_,
    new_n22046_, new_n22047_, new_n22048_, new_n22049_, new_n22050_,
    new_n22051_, new_n22052_, new_n22053_, new_n22054_, new_n22055_,
    new_n22056_, new_n22057_, new_n22058_, new_n22059_, new_n22060_,
    new_n22061_, new_n22062_, new_n22063_, new_n22064_, new_n22065_,
    new_n22066_, new_n22067_, new_n22068_, new_n22069_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22138_, new_n22139_, new_n22140_, new_n22141_,
    new_n22142_, new_n22146_, new_n22147_, new_n22148_, new_n22149_,
    new_n22150_, new_n22151_, new_n22152_, new_n22153_, new_n22154_,
    new_n22155_, new_n22156_, new_n22157_, new_n22158_, new_n22159_,
    new_n22160_, new_n22161_, new_n22162_, new_n22163_, new_n22164_,
    new_n22165_, new_n22166_, new_n22167_, new_n22168_, new_n22169_,
    new_n22170_, new_n22171_, new_n22172_, new_n22173_, new_n22174_,
    new_n22175_, new_n22176_, new_n22177_, new_n22178_, new_n22179_,
    new_n22180_, new_n22181_, new_n22182_, new_n22183_, new_n22184_,
    new_n22185_, new_n22186_, new_n22187_, new_n22188_, new_n22189_,
    new_n22190_, new_n22191_, new_n22192_, new_n22193_, new_n22194_,
    new_n22195_, new_n22196_, new_n22197_, new_n22198_, new_n22199_,
    new_n22200_, new_n22201_, new_n22202_, new_n22203_, new_n22204_,
    new_n22205_, new_n22206_, new_n22207_, new_n22208_, new_n22209_,
    new_n22210_, new_n22211_, new_n22212_, new_n22214_, new_n22215_,
    new_n22216_, new_n22217_, new_n22218_, new_n22219_, new_n22220_,
    new_n22221_, new_n22222_, new_n22223_, new_n22224_, new_n22225_,
    new_n22226_, new_n22227_, new_n22228_, new_n22229_, new_n22230_,
    new_n22231_, new_n22232_, new_n22233_, new_n22234_, new_n22235_,
    new_n22236_, new_n22237_, new_n22238_, new_n22239_, new_n22240_,
    new_n22241_, new_n22242_, new_n22243_, new_n22244_, new_n22245_,
    new_n22246_, new_n22247_, new_n22248_, new_n22249_, new_n22250_,
    new_n22251_, new_n22252_, new_n22253_, new_n22254_, new_n22255_,
    new_n22256_, new_n22257_, new_n22258_, new_n22259_, new_n22260_,
    new_n22261_, new_n22262_, new_n22263_, new_n22264_, new_n22265_,
    new_n22266_, new_n22267_, new_n22268_, new_n22269_, new_n22270_,
    new_n22271_, new_n22272_, new_n22273_, new_n22274_, new_n22275_,
    new_n22276_, new_n22277_, new_n22278_, new_n22279_, new_n22280_,
    new_n22281_, new_n22282_, new_n22283_, new_n22284_, new_n22285_,
    new_n22286_, new_n22287_, new_n22288_, new_n22289_, new_n22290_,
    new_n22291_, new_n22292_, new_n22293_, new_n22294_, new_n22295_,
    new_n22296_, new_n22297_, new_n22298_, new_n22299_, new_n22300_,
    new_n22301_, new_n22302_, new_n22303_, new_n22304_, new_n22305_,
    new_n22306_, new_n22307_, new_n22308_, new_n22309_, new_n22310_,
    new_n22311_, new_n22312_, new_n22313_, new_n22314_, new_n22315_,
    new_n22316_, new_n22317_, new_n22318_, new_n22319_, new_n22320_,
    new_n22321_, new_n22322_, new_n22323_, new_n22324_, new_n22325_,
    new_n22326_, new_n22327_, new_n22328_, new_n22329_, new_n22330_,
    new_n22331_, new_n22332_, new_n22333_, new_n22334_, new_n22335_,
    new_n22336_, new_n22337_, new_n22338_, new_n22339_, new_n22340_,
    new_n22341_, new_n22342_, new_n22343_, new_n22344_, new_n22345_,
    new_n22346_, new_n22347_, new_n22348_, new_n22349_, new_n22350_,
    new_n22351_, new_n22352_, new_n22353_, new_n22354_, new_n22355_,
    new_n22356_, new_n22357_, new_n22358_, new_n22359_, new_n22360_,
    new_n22361_, new_n22362_, new_n22363_, new_n22364_, new_n22365_,
    new_n22366_, new_n22367_, new_n22368_, new_n22369_, new_n22370_,
    new_n22371_, new_n22372_, new_n22373_, new_n22374_, new_n22375_,
    new_n22376_, new_n22377_, new_n22378_, new_n22379_, new_n22380_,
    new_n22381_, new_n22382_, new_n22383_, new_n22384_, new_n22385_,
    new_n22386_, new_n22387_, new_n22388_, new_n22389_, new_n22390_,
    new_n22391_, new_n22392_, new_n22393_, new_n22394_, new_n22395_,
    new_n22396_, new_n22397_, new_n22398_, new_n22399_, new_n22400_,
    new_n22401_, new_n22402_, new_n22403_, new_n22404_, new_n22405_,
    new_n22406_, new_n22407_, new_n22408_, new_n22409_, new_n22410_,
    new_n22411_, new_n22412_, new_n22413_, new_n22414_, new_n22415_,
    new_n22416_, new_n22417_, new_n22418_, new_n22419_, new_n22420_,
    new_n22421_, new_n22422_, new_n22423_, new_n22424_, new_n22425_,
    new_n22426_, new_n22427_, new_n22428_, new_n22429_, new_n22430_,
    new_n22431_, new_n22432_, new_n22433_, new_n22434_, new_n22435_,
    new_n22436_, new_n22438_, new_n22439_, new_n22440_, new_n22441_,
    new_n22442_, new_n22443_, new_n22444_, new_n22445_, new_n22446_,
    new_n22447_, new_n22448_, new_n22449_, new_n22450_, new_n22451_,
    new_n22452_, new_n22453_, new_n22454_, new_n22455_, new_n22456_,
    new_n22457_, new_n22458_, new_n22459_, new_n22460_, new_n22461_,
    new_n22462_, new_n22463_, new_n22464_, new_n22465_, new_n22466_,
    new_n22467_, new_n22468_, new_n22469_, new_n22470_, new_n22471_,
    new_n22472_, new_n22473_, new_n22474_, new_n22475_, new_n22476_,
    new_n22477_, new_n22478_, new_n22479_, new_n22480_, new_n22481_,
    new_n22482_, new_n22483_, new_n22484_, new_n22485_, new_n22486_,
    new_n22487_, new_n22488_, new_n22489_, new_n22490_, new_n22491_,
    new_n22492_, new_n22493_, new_n22494_, new_n22495_, new_n22496_,
    new_n22497_, new_n22498_, new_n22499_, new_n22500_, new_n22501_,
    new_n22502_, new_n22503_, new_n22504_, new_n22505_, new_n22506_,
    new_n22507_, new_n22508_, new_n22509_, new_n22513_, new_n22514_,
    new_n22515_, new_n22516_, new_n22517_, new_n22518_, new_n22519_,
    new_n22520_, new_n22521_, new_n22522_, new_n22523_, new_n22524_,
    new_n22525_, new_n22526_, new_n22527_, new_n22528_, new_n22529_,
    new_n22530_, new_n22531_, new_n22532_, new_n22533_, new_n22534_,
    new_n22535_, new_n22536_, new_n22537_, new_n22538_, new_n22539_,
    new_n22540_, new_n22541_, new_n22542_, new_n22543_, new_n22544_,
    new_n22545_, new_n22546_, new_n22547_, new_n22548_, new_n22549_,
    new_n22550_, new_n22551_, new_n22552_, new_n22553_, new_n22554_,
    new_n22555_, new_n22556_, new_n22557_, new_n22558_, new_n22559_,
    new_n22560_, new_n22561_, new_n22562_, new_n22563_, new_n22564_,
    new_n22565_, new_n22566_, new_n22567_, new_n22568_, new_n22569_,
    new_n22570_, new_n22571_, new_n22572_, new_n22573_, new_n22574_,
    new_n22575_, new_n22576_, new_n22577_, new_n22578_, new_n22579_,
    new_n22581_, new_n22582_, new_n22583_, new_n22584_, new_n22585_,
    new_n22586_, new_n22587_, new_n22588_, new_n22589_, new_n22590_,
    new_n22591_, new_n22592_, new_n22593_, new_n22594_, new_n22595_,
    new_n22596_, new_n22597_, new_n22598_, new_n22599_, new_n22600_,
    new_n22601_, new_n22602_, new_n22603_, new_n22604_, new_n22605_,
    new_n22606_, new_n22607_, new_n22608_, new_n22609_, new_n22610_,
    new_n22611_, new_n22612_, new_n22613_, new_n22614_, new_n22615_,
    new_n22616_, new_n22617_, new_n22618_, new_n22619_, new_n22620_,
    new_n22621_, new_n22622_, new_n22623_, new_n22624_, new_n22625_,
    new_n22626_, new_n22627_, new_n22628_, new_n22629_, new_n22630_,
    new_n22631_, new_n22632_, new_n22633_, new_n22634_, new_n22635_,
    new_n22636_, new_n22637_, new_n22638_, new_n22639_, new_n22640_,
    new_n22641_, new_n22642_, new_n22643_, new_n22644_, new_n22645_,
    new_n22646_, new_n22647_, new_n22648_, new_n22649_, new_n22650_,
    new_n22651_, new_n22652_, new_n22653_, new_n22654_, new_n22655_,
    new_n22656_, new_n22657_, new_n22658_, new_n22659_, new_n22660_,
    new_n22661_, new_n22662_, new_n22663_, new_n22664_, new_n22665_,
    new_n22666_, new_n22667_, new_n22668_, new_n22669_, new_n22670_,
    new_n22671_, new_n22672_, new_n22673_, new_n22674_, new_n22675_,
    new_n22676_, new_n22677_, new_n22678_, new_n22679_, new_n22680_,
    new_n22681_, new_n22682_, new_n22683_, new_n22684_, new_n22685_,
    new_n22686_, new_n22687_, new_n22688_, new_n22689_, new_n22690_,
    new_n22691_, new_n22692_, new_n22693_, new_n22694_, new_n22695_,
    new_n22696_, new_n22697_, new_n22698_, new_n22699_, new_n22700_,
    new_n22701_, new_n22702_, new_n22703_, new_n22704_, new_n22705_,
    new_n22706_, new_n22707_, new_n22708_, new_n22709_, new_n22710_,
    new_n22711_, new_n22712_, new_n22713_, new_n22714_, new_n22715_,
    new_n22716_, new_n22717_, new_n22718_, new_n22719_, new_n22720_,
    new_n22721_, new_n22722_, new_n22723_, new_n22724_, new_n22725_,
    new_n22726_, new_n22727_, new_n22728_, new_n22729_, new_n22730_,
    new_n22731_, new_n22732_, new_n22733_, new_n22734_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22744_, new_n22745_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22879_, new_n22880_, new_n22881_, new_n22882_, new_n22883_,
    new_n22884_, new_n22885_, new_n22886_, new_n22887_, new_n22888_,
    new_n22889_, new_n22890_, new_n22891_, new_n22892_, new_n22893_,
    new_n22894_, new_n22895_, new_n22896_, new_n22897_, new_n22898_,
    new_n22899_, new_n22900_, new_n22901_, new_n22902_, new_n22903_,
    new_n22904_, new_n22905_, new_n22906_, new_n22907_, new_n22908_,
    new_n22909_, new_n22910_, new_n22911_, new_n22912_, new_n22913_,
    new_n22914_, new_n22915_, new_n22916_, new_n22917_, new_n22918_,
    new_n22919_, new_n22920_, new_n22921_, new_n22922_, new_n22923_,
    new_n22924_, new_n22925_, new_n22926_, new_n22927_, new_n22928_,
    new_n22929_, new_n22930_, new_n22931_, new_n22932_, new_n22933_,
    new_n22934_, new_n22935_, new_n22936_, new_n22937_, new_n22938_,
    new_n22939_, new_n22940_, new_n22941_, new_n22942_, new_n22943_,
    new_n22944_, new_n22945_, new_n22946_, new_n22947_, new_n22948_,
    new_n22949_, new_n22950_, new_n22951_, new_n22952_, new_n22953_,
    new_n22954_, new_n22955_, new_n22956_, new_n22957_, new_n22958_,
    new_n22960_, new_n22961_, new_n22962_, new_n22963_, new_n22964_,
    new_n22965_, new_n22966_, new_n22967_, new_n22968_, new_n22969_,
    new_n22970_, new_n22971_, new_n22972_, new_n22973_, new_n22974_,
    new_n22975_, new_n22976_, new_n22977_, new_n22978_, new_n22979_,
    new_n22980_, new_n22981_, new_n22982_, new_n22983_, new_n22984_,
    new_n22985_, new_n22986_, new_n22987_, new_n22988_, new_n22989_,
    new_n22990_, new_n22991_, new_n22992_, new_n22993_, new_n22994_,
    new_n22995_, new_n22996_, new_n22997_, new_n22998_, new_n22999_,
    new_n23000_, new_n23001_, new_n23002_, new_n23003_, new_n23004_,
    new_n23005_, new_n23006_, new_n23007_, new_n23008_, new_n23009_,
    new_n23010_, new_n23011_, new_n23012_, new_n23013_, new_n23014_,
    new_n23015_, new_n23016_, new_n23017_, new_n23018_, new_n23019_,
    new_n23020_, new_n23021_, new_n23022_, new_n23023_, new_n23024_,
    new_n23025_, new_n23026_, new_n23027_, new_n23028_, new_n23029_,
    new_n23030_, new_n23031_, new_n23032_, new_n23033_, new_n23034_,
    new_n23035_, new_n23036_, new_n23037_, new_n23038_, new_n23039_,
    new_n23041_, new_n23042_, new_n23043_, new_n23044_, new_n23045_,
    new_n23046_, new_n23047_, new_n23048_, new_n23049_, new_n23050_,
    new_n23051_, new_n23052_, new_n23053_, new_n23054_, new_n23055_,
    new_n23056_, new_n23057_, new_n23058_, new_n23059_, new_n23060_,
    new_n23061_, new_n23062_, new_n23063_, new_n23064_, new_n23065_,
    new_n23066_, new_n23067_, new_n23068_, new_n23069_, new_n23070_,
    new_n23071_, new_n23072_, new_n23073_, new_n23074_, new_n23075_,
    new_n23076_, new_n23077_, new_n23078_, new_n23079_, new_n23080_,
    new_n23081_, new_n23082_, new_n23083_, new_n23084_, new_n23085_,
    new_n23086_, new_n23087_, new_n23088_, new_n23089_, new_n23090_,
    new_n23091_, new_n23092_, new_n23093_, new_n23094_, new_n23095_,
    new_n23096_, new_n23097_, new_n23098_, new_n23099_, new_n23100_,
    new_n23101_, new_n23102_, new_n23103_, new_n23104_, new_n23105_,
    new_n23106_, new_n23107_, new_n23108_, new_n23109_, new_n23110_,
    new_n23111_, new_n23112_, new_n23113_, new_n23114_, new_n23115_,
    new_n23116_, new_n23117_, new_n23118_, new_n23119_, new_n23120_,
    new_n23121_, new_n23122_, new_n23123_, new_n23124_, new_n23125_,
    new_n23126_, new_n23127_, new_n23128_, new_n23129_, new_n23134_,
    new_n23135_, new_n23136_, new_n23137_, new_n23138_, new_n23139_,
    new_n23140_, new_n23141_, new_n23142_, new_n23143_, new_n23144_,
    new_n23145_, new_n23146_, new_n23147_, new_n23148_, new_n23149_,
    new_n23150_, new_n23151_, new_n23153_, new_n23154_, new_n23155_,
    new_n23156_, new_n23157_, new_n23158_, new_n23159_, new_n23162_,
    new_n23163_, new_n23164_, new_n23165_, new_n23169_, new_n23170_,
    new_n23171_, new_n23172_, new_n23173_, new_n23174_, new_n23175_,
    new_n23176_, new_n23177_, new_n23178_, new_n23179_, new_n23180_,
    new_n23181_, new_n23182_, new_n23183_, new_n23184_, new_n23185_,
    new_n23186_, new_n23187_, new_n23188_, new_n23189_, new_n23190_,
    new_n23191_, new_n23192_, new_n23193_, new_n23194_, new_n23195_,
    new_n23196_, new_n23197_, new_n23198_, new_n23199_, new_n23200_,
    new_n23201_, new_n23202_, new_n23203_, new_n23204_, new_n23205_,
    new_n23206_, new_n23207_, new_n23208_, new_n23209_, new_n23210_,
    new_n23211_, new_n23212_, new_n23213_, new_n23214_, new_n23215_,
    new_n23216_, new_n23217_, new_n23218_, new_n23219_, new_n23220_,
    new_n23221_, new_n23222_, new_n23223_, new_n23224_, new_n23225_,
    new_n23226_, new_n23227_, new_n23228_, new_n23229_, new_n23230_,
    new_n23231_, new_n23232_, new_n23233_, new_n23234_, new_n23235_,
    new_n23236_, new_n23237_, new_n23238_, new_n23239_, new_n23240_,
    new_n23241_, new_n23242_, new_n23243_, new_n23244_, new_n23245_,
    new_n23246_, new_n23247_, new_n23248_, new_n23249_, new_n23250_,
    new_n23251_, new_n23252_, new_n23253_, new_n23254_, new_n23255_,
    new_n23256_, new_n23257_, new_n23258_, new_n23259_, new_n23260_,
    new_n23261_, new_n23262_, new_n23263_, new_n23264_, new_n23265_,
    new_n23266_, new_n23267_, new_n23268_, new_n23269_, new_n23270_,
    new_n23271_, new_n23272_, new_n23273_, new_n23274_, new_n23275_,
    new_n23276_, new_n23277_, new_n23278_, new_n23279_, new_n23280_,
    new_n23281_, new_n23282_, new_n23283_, new_n23284_, new_n23285_,
    new_n23286_, new_n23287_, new_n23288_, new_n23289_, new_n23290_,
    new_n23291_, new_n23292_, new_n23293_, new_n23294_, new_n23295_,
    new_n23296_, new_n23297_, new_n23298_, new_n23299_, new_n23300_,
    new_n23301_, new_n23302_, new_n23303_, new_n23304_, new_n23305_,
    new_n23306_, new_n23307_, new_n23308_, new_n23309_, new_n23310_,
    new_n23311_, new_n23312_, new_n23313_, new_n23314_, new_n23315_,
    new_n23316_, new_n23317_, new_n23318_, new_n23319_, new_n23320_,
    new_n23321_, new_n23322_, new_n23323_, new_n23324_, new_n23325_,
    new_n23326_, new_n23327_, new_n23328_, new_n23329_, new_n23330_,
    new_n23331_, new_n23332_, new_n23333_, new_n23334_, new_n23335_,
    new_n23336_, new_n23337_, new_n23338_, new_n23339_, new_n23340_,
    new_n23341_, new_n23342_, new_n23343_, new_n23344_, new_n23345_,
    new_n23346_, new_n23347_, new_n23348_, new_n23349_, new_n23350_,
    new_n23351_, new_n23352_, new_n23353_, new_n23354_, new_n23355_,
    new_n23356_, new_n23357_, new_n23358_, new_n23359_, new_n23360_,
    new_n23361_, new_n23362_, new_n23363_, new_n23364_, new_n23365_,
    new_n23366_, new_n23367_, new_n23368_, new_n23369_, new_n23370_,
    new_n23371_, new_n23372_, new_n23373_, new_n23374_, new_n23375_,
    new_n23376_, new_n23377_, new_n23378_, new_n23379_, new_n23380_,
    new_n23381_, new_n23382_, new_n23383_, new_n23384_, new_n23385_,
    new_n23386_, new_n23387_, new_n23388_, new_n23389_, new_n23390_,
    new_n23391_, new_n23392_, new_n23393_, new_n23394_, new_n23395_,
    new_n23396_, new_n23397_, new_n23398_, new_n23400_, new_n23401_,
    new_n23402_, new_n23404_, new_n23405_, new_n23406_, new_n23407_,
    new_n23408_, new_n23409_, new_n23410_, new_n23411_, new_n23412_,
    new_n23413_, new_n23414_, new_n23415_, new_n23416_, new_n23417_,
    new_n23418_, new_n23419_, new_n23420_, new_n23421_, new_n23422_,
    new_n23423_, new_n23427_, new_n23428_, new_n23429_, new_n23430_,
    new_n23431_, new_n23432_, new_n23433_, new_n23434_, new_n23435_,
    new_n23436_, new_n23437_, new_n23438_, new_n23439_, new_n23440_,
    new_n23441_, new_n23442_, new_n23443_, new_n23444_, new_n23445_,
    new_n23446_, new_n23447_, new_n23448_, new_n23449_, new_n23450_,
    new_n23451_, new_n23452_, new_n23453_, new_n23454_, new_n23455_,
    new_n23456_, new_n23457_, new_n23458_, new_n23459_, new_n23460_,
    new_n23461_, new_n23462_, new_n23463_, new_n23464_, new_n23465_,
    new_n23466_, new_n23467_, new_n23468_, new_n23469_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23501_, new_n23502_, new_n23503_, new_n23504_, new_n23505_,
    new_n23506_, new_n23507_, new_n23508_, new_n23509_, new_n23510_,
    new_n23511_, new_n23512_, new_n23513_, new_n23514_, new_n23515_,
    new_n23520_, new_n23521_, new_n23522_, new_n23523_, new_n23524_,
    new_n23525_, new_n23526_, new_n23527_, new_n23528_, new_n23529_,
    new_n23530_, new_n23531_, new_n23532_, new_n23533_, new_n23534_,
    new_n23535_, new_n23536_, new_n23538_, new_n23539_, new_n23540_,
    new_n23543_, new_n23544_, new_n23545_, new_n23546_, new_n23547_,
    new_n23548_, new_n23549_, new_n23550_, new_n23551_, new_n23552_,
    new_n23553_, new_n23554_, new_n23555_, new_n23556_, new_n23557_,
    new_n23558_, new_n23559_, new_n23560_, new_n23561_, new_n23562_,
    new_n23563_, new_n23564_, new_n23565_, new_n23566_, new_n23567_,
    new_n23568_, new_n23569_, new_n23570_, new_n23571_, new_n23572_,
    new_n23573_, new_n23574_, new_n23575_, new_n23576_, new_n23577_,
    new_n23578_, new_n23579_, new_n23580_, new_n23581_, new_n23582_,
    new_n23583_, new_n23584_, new_n23585_, new_n23586_, new_n23587_,
    new_n23588_, new_n23589_, new_n23590_, new_n23591_, new_n23592_,
    new_n23593_, new_n23594_, new_n23595_, new_n23596_, new_n23597_,
    new_n23598_, new_n23599_, new_n23600_, new_n23601_, new_n23602_,
    new_n23603_, new_n23604_, new_n23605_, new_n23606_, new_n23607_,
    new_n23608_, new_n23609_, new_n23610_, new_n23611_, new_n23612_,
    new_n23613_, new_n23614_, new_n23615_, new_n23616_, new_n23617_,
    new_n23618_, new_n23619_, new_n23620_, new_n23621_, new_n23622_,
    new_n23623_, new_n23624_, new_n23625_, new_n23626_, new_n23627_,
    new_n23628_, new_n23629_, new_n23630_, new_n23631_, new_n23632_,
    new_n23633_, new_n23634_, new_n23635_, new_n23636_, new_n23637_,
    new_n23638_, new_n23639_, new_n23640_, new_n23641_, new_n23642_,
    new_n23643_, new_n23644_, new_n23645_, new_n23646_, new_n23647_,
    new_n23648_, new_n23649_, new_n23650_, new_n23651_, new_n23652_,
    new_n23653_, new_n23654_, new_n23655_, new_n23656_, new_n23657_,
    new_n23658_, new_n23659_, new_n23660_, new_n23661_, new_n23662_,
    new_n23663_, new_n23664_, new_n23665_, new_n23666_, new_n23667_,
    new_n23668_, new_n23669_, new_n23670_, new_n23671_, new_n23672_,
    new_n23673_, new_n23674_, new_n23675_, new_n23676_, new_n23677_,
    new_n23678_, new_n23679_, new_n23680_, new_n23681_, new_n23682_,
    new_n23683_, new_n23684_, new_n23685_, new_n23686_, new_n23687_,
    new_n23688_, new_n23689_, new_n23690_, new_n23691_, new_n23692_,
    new_n23693_, new_n23694_, new_n23695_, new_n23696_, new_n23697_,
    new_n23698_, new_n23699_, new_n23700_, new_n23701_, new_n23702_,
    new_n23703_, new_n23704_, new_n23705_, new_n23706_, new_n23707_,
    new_n23708_, new_n23709_, new_n23710_, new_n23711_, new_n23712_,
    new_n23713_, new_n23714_, new_n23715_, new_n23716_, new_n23717_,
    new_n23718_, new_n23719_, new_n23720_, new_n23721_, new_n23722_,
    new_n23723_, new_n23724_, new_n23725_, new_n23726_, new_n23727_,
    new_n23728_, new_n23729_, new_n23730_, new_n23731_, new_n23732_,
    new_n23733_, new_n23734_, new_n23735_, new_n23736_, new_n23737_,
    new_n23738_, new_n23739_, new_n23740_, new_n23741_, new_n23742_,
    new_n23743_, new_n23744_, new_n23745_, new_n23746_, new_n23749_,
    new_n23750_, new_n23751_, new_n23752_, new_n23753_, new_n23754_,
    new_n23755_, new_n23756_, new_n23757_, new_n23758_, new_n23759_,
    new_n23760_, new_n23761_, new_n23762_, new_n23763_, new_n23764_,
    new_n23765_, new_n23766_, new_n23767_, new_n23768_, new_n23772_,
    new_n23773_, new_n23774_, new_n23775_, new_n23776_, new_n23777_,
    new_n23778_, new_n23779_, new_n23780_, new_n23781_, new_n23782_,
    new_n23783_, new_n23784_, new_n23785_, new_n23786_, new_n23787_,
    new_n23788_, new_n23789_, new_n23790_, new_n23791_, new_n23792_,
    new_n23793_, new_n23794_, new_n23795_, new_n23796_, new_n23797_,
    new_n23798_, new_n23799_, new_n23800_, new_n23801_, new_n23802_,
    new_n23803_, new_n23804_, new_n23805_, new_n23806_, new_n23807_,
    new_n23808_, new_n23809_, new_n23810_, new_n23811_, new_n23812_,
    new_n23813_, new_n23814_, new_n23815_, new_n23816_, new_n23817_,
    new_n23818_, new_n23819_, new_n23820_, new_n23821_, new_n23822_,
    new_n23823_, new_n23824_, new_n23825_, new_n23826_, new_n23827_,
    new_n23828_, new_n23829_, new_n23830_, new_n23831_, new_n23832_,
    new_n23833_, new_n23834_, new_n23835_, new_n23836_, new_n23837_,
    new_n23838_, new_n23839_, new_n23840_, new_n23841_, new_n23842_,
    new_n23843_, new_n23844_, new_n23845_, new_n23846_, new_n23847_,
    new_n23848_, new_n23849_, new_n23850_, new_n23851_, new_n23852_,
    new_n23853_, new_n23854_, new_n23855_, new_n23856_, new_n23857_,
    new_n23858_, new_n23859_, new_n23860_, new_n23865_, new_n23866_,
    new_n23867_, new_n23868_, new_n23869_, new_n23870_, new_n23871_,
    new_n23872_, new_n23873_, new_n23874_, new_n23875_, new_n23876_,
    new_n23877_, new_n23878_, new_n23879_, new_n23880_, new_n23881_,
    new_n23883_, new_n23884_, new_n23885_, new_n23888_, new_n23889_,
    new_n23890_, new_n23891_, new_n23892_, new_n23893_, new_n23894_,
    new_n23895_, new_n23896_, new_n23897_, new_n23898_, new_n23899_,
    new_n23900_, new_n23901_, new_n23902_, new_n23903_, new_n23904_,
    new_n23905_, new_n23906_, new_n23907_, new_n23908_, new_n23909_,
    new_n23910_, new_n23911_, new_n23912_, new_n23913_, new_n23914_,
    new_n23915_, new_n23916_, new_n23917_, new_n23918_, new_n23919_,
    new_n23920_, new_n23921_, new_n23922_, new_n23923_, new_n23924_,
    new_n23925_, new_n23926_, new_n23927_, new_n23928_, new_n23929_,
    new_n23930_, new_n23931_, new_n23932_, new_n23933_, new_n23934_,
    new_n23935_, new_n23936_, new_n23937_, new_n23938_, new_n23939_,
    new_n23940_, new_n23941_, new_n23942_, new_n23943_, new_n23944_,
    new_n23945_, new_n23946_, new_n23947_, new_n23948_, new_n23949_,
    new_n23950_, new_n23951_, new_n23952_, new_n23953_, new_n23954_,
    new_n23955_, new_n23956_, new_n23957_, new_n23958_, new_n23959_,
    new_n23960_, new_n23961_, new_n23962_, new_n23963_, new_n23964_,
    new_n23965_, new_n23966_, new_n23967_, new_n23968_, new_n23969_,
    new_n23970_, new_n23971_, new_n23972_, new_n23973_, new_n23974_,
    new_n23975_, new_n23976_, new_n23977_, new_n23978_, new_n23979_,
    new_n23980_, new_n23981_, new_n23982_, new_n23983_, new_n23984_,
    new_n23985_, new_n23986_, new_n23987_, new_n23988_, new_n23989_,
    new_n23990_, new_n23991_, new_n23992_, new_n23993_, new_n23994_,
    new_n23995_, new_n23996_, new_n23997_, new_n23998_, new_n23999_,
    new_n24000_, new_n24001_, new_n24002_, new_n24003_, new_n24004_,
    new_n24005_, new_n24006_, new_n24007_, new_n24008_, new_n24009_,
    new_n24010_, new_n24011_, new_n24012_, new_n24013_, new_n24014_,
    new_n24015_, new_n24016_, new_n24017_, new_n24018_, new_n24019_,
    new_n24020_, new_n24021_, new_n24022_, new_n24023_, new_n24024_,
    new_n24025_, new_n24026_, new_n24027_, new_n24028_, new_n24029_,
    new_n24030_, new_n24031_, new_n24032_, new_n24033_, new_n24034_,
    new_n24035_, new_n24036_, new_n24037_, new_n24038_, new_n24039_,
    new_n24040_, new_n24041_, new_n24042_, new_n24043_, new_n24044_,
    new_n24045_, new_n24046_, new_n24047_, new_n24048_, new_n24049_,
    new_n24050_, new_n24051_, new_n24052_, new_n24053_, new_n24054_,
    new_n24055_, new_n24056_, new_n24057_, new_n24058_, new_n24059_,
    new_n24060_, new_n24061_, new_n24062_, new_n24063_, new_n24064_,
    new_n24065_, new_n24066_, new_n24067_, new_n24068_, new_n24069_,
    new_n24070_, new_n24071_, new_n24072_, new_n24073_, new_n24074_,
    new_n24075_, new_n24076_, new_n24077_, new_n24078_, new_n24079_,
    new_n24080_, new_n24081_, new_n24082_, new_n24083_, new_n24084_,
    new_n24085_, new_n24086_, new_n24087_, new_n24088_, new_n24089_,
    new_n24090_, new_n24091_, new_n24093_, new_n24094_, new_n24095_,
    new_n24096_, new_n24097_, new_n24098_, new_n24099_, new_n24100_,
    new_n24101_, new_n24102_, new_n24103_, new_n24104_, new_n24105_,
    new_n24106_, new_n24107_, new_n24108_, new_n24109_, new_n24110_,
    new_n24111_, new_n24112_, new_n24113_, new_n24114_, new_n24115_,
    new_n24116_, new_n24117_, new_n24122_, new_n24123_, new_n24124_,
    new_n24125_, new_n24126_, new_n24127_, new_n24128_, new_n24129_,
    new_n24130_, new_n24131_, new_n24132_, new_n24133_, new_n24134_,
    new_n24135_, new_n24136_, new_n24137_, new_n24138_, new_n24139_,
    new_n24140_, new_n24141_, new_n24142_, new_n24143_, new_n24144_,
    new_n24145_, new_n24146_, new_n24147_, new_n24148_, new_n24149_,
    new_n24150_, new_n24151_, new_n24152_, new_n24153_, new_n24154_,
    new_n24155_, new_n24156_, new_n24157_, new_n24158_, new_n24159_,
    new_n24160_, new_n24161_, new_n24162_, new_n24163_, new_n24164_,
    new_n24165_, new_n24166_, new_n24167_, new_n24168_, new_n24169_,
    new_n24170_, new_n24171_, new_n24172_, new_n24173_, new_n24174_,
    new_n24175_, new_n24176_, new_n24177_, new_n24178_, new_n24179_,
    new_n24180_, new_n24181_, new_n24182_, new_n24183_, new_n24184_,
    new_n24185_, new_n24186_, new_n24187_, new_n24188_, new_n24189_,
    new_n24190_, new_n24191_, new_n24192_, new_n24193_, new_n24194_,
    new_n24195_, new_n24196_, new_n24197_, new_n24198_, new_n24199_,
    new_n24200_, new_n24201_, new_n24202_, new_n24203_, new_n24204_,
    new_n24205_, new_n24206_, new_n24207_, new_n24208_, new_n24209_,
    new_n24210_, new_n24211_, new_n24212_, new_n24213_, new_n24214_,
    new_n24215_, new_n24216_, new_n24217_, new_n24218_, new_n24219_,
    new_n24220_, new_n24221_, new_n24222_, new_n24223_, new_n24224_,
    new_n24225_, new_n24226_, new_n24227_, new_n24228_, new_n24229_,
    new_n24230_, new_n24231_, new_n24232_, new_n24233_, new_n24234_,
    new_n24235_, new_n24236_, new_n24237_, new_n24238_, new_n24239_,
    new_n24240_, new_n24241_, new_n24242_, new_n24243_, new_n24244_,
    new_n24245_, new_n24246_, new_n24247_, new_n24248_, new_n24249_,
    new_n24250_, new_n24254_, new_n24255_, new_n24256_, new_n24257_,
    new_n24258_, new_n24259_, new_n24260_, new_n24261_, new_n24262_,
    new_n24263_, new_n24264_, new_n24265_, new_n24266_, new_n24267_,
    new_n24268_, new_n24269_, new_n24271_, new_n24272_, new_n24273_,
    new_n24274_, new_n24275_, new_n24276_, new_n24277_, new_n24278_,
    new_n24281_, new_n24282_, new_n24283_, new_n24286_, new_n24287_,
    new_n24288_, new_n24289_, new_n24290_, new_n24291_, new_n24292_,
    new_n24293_, new_n24294_, new_n24295_, new_n24296_, new_n24297_,
    new_n24298_, new_n24299_, new_n24300_, new_n24301_, new_n24302_,
    new_n24303_, new_n24304_, new_n24305_, new_n24306_, new_n24307_,
    new_n24308_, new_n24309_, new_n24310_, new_n24311_, new_n24312_,
    new_n24313_, new_n24314_, new_n24315_, new_n24316_, new_n24317_,
    new_n24318_, new_n24319_, new_n24320_, new_n24321_, new_n24322_,
    new_n24323_, new_n24324_, new_n24325_, new_n24326_, new_n24327_,
    new_n24328_, new_n24329_, new_n24330_, new_n24331_, new_n24332_,
    new_n24333_, new_n24334_, new_n24335_, new_n24336_, new_n24337_,
    new_n24338_, new_n24339_, new_n24340_, new_n24341_, new_n24342_,
    new_n24343_, new_n24344_, new_n24345_, new_n24346_, new_n24347_,
    new_n24348_, new_n24349_, new_n24350_, new_n24351_, new_n24352_,
    new_n24353_, new_n24354_, new_n24355_, new_n24356_, new_n24357_,
    new_n24358_, new_n24359_, new_n24360_, new_n24361_, new_n24362_,
    new_n24363_, new_n24364_, new_n24365_, new_n24366_, new_n24367_,
    new_n24368_, new_n24369_, new_n24370_, new_n24371_, new_n24372_,
    new_n24373_, new_n24374_, new_n24375_, new_n24376_, new_n24377_,
    new_n24378_, new_n24379_, new_n24380_, new_n24381_, new_n24382_,
    new_n24383_, new_n24384_, new_n24385_, new_n24386_, new_n24387_,
    new_n24388_, new_n24389_, new_n24390_, new_n24391_, new_n24392_,
    new_n24393_, new_n24394_, new_n24395_, new_n24396_, new_n24397_,
    new_n24398_, new_n24399_, new_n24400_, new_n24401_, new_n24402_,
    new_n24403_, new_n24404_, new_n24405_, new_n24406_, new_n24407_,
    new_n24408_, new_n24409_, new_n24410_, new_n24411_, new_n24412_,
    new_n24413_, new_n24414_, new_n24415_, new_n24416_, new_n24417_,
    new_n24418_, new_n24419_, new_n24420_, new_n24421_, new_n24422_,
    new_n24423_, new_n24424_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24463_, new_n24464_, new_n24465_, new_n24466_, new_n24467_,
    new_n24468_, new_n24469_, new_n24470_, new_n24471_, new_n24472_,
    new_n24473_, new_n24474_, new_n24475_, new_n24477_, new_n24478_,
    new_n24479_, new_n24480_, new_n24481_, new_n24482_, new_n24483_,
    new_n24484_, new_n24485_, new_n24486_, new_n24487_, new_n24488_,
    new_n24489_, new_n24490_, new_n24491_, new_n24492_, new_n24493_,
    new_n24494_, new_n24495_, new_n24496_, new_n24497_, new_n24498_,
    new_n24499_, new_n24500_, new_n24501_, new_n24502_, new_n24503_,
    new_n24504_, new_n24505_, new_n24506_, new_n24507_, new_n24508_,
    new_n24509_, new_n24510_, new_n24511_, new_n24512_, new_n24513_,
    new_n24514_, new_n24515_, new_n24516_, new_n24517_, new_n24518_,
    new_n24519_, new_n24520_, new_n24521_, new_n24522_, new_n24523_,
    new_n24524_, new_n24525_, new_n24526_, new_n24527_, new_n24528_,
    new_n24529_, new_n24530_, new_n24531_, new_n24532_, new_n24533_,
    new_n24534_, new_n24535_, new_n24536_, new_n24537_, new_n24538_,
    new_n24539_, new_n24540_, new_n24541_, new_n24542_, new_n24543_,
    new_n24544_, new_n24545_, new_n24546_, new_n24547_, new_n24548_,
    new_n24551_, new_n24552_, new_n24553_, new_n24554_, new_n24555_,
    new_n24556_, new_n24557_, new_n24558_, new_n24559_, new_n24560_,
    new_n24561_, new_n24562_, new_n24563_, new_n24564_, new_n24565_,
    new_n24566_, new_n24567_, new_n24568_, new_n24569_, new_n24570_,
    new_n24571_, new_n24572_, new_n24573_, new_n24574_, new_n24575_,
    new_n24576_, new_n24577_, new_n24578_, new_n24579_, new_n24580_,
    new_n24581_, new_n24582_, new_n24583_, new_n24584_, new_n24585_,
    new_n24586_, new_n24587_, new_n24588_, new_n24589_, new_n24590_,
    new_n24591_, new_n24592_, new_n24593_, new_n24594_, new_n24595_,
    new_n24596_, new_n24597_, new_n24598_, new_n24599_, new_n24600_,
    new_n24601_, new_n24602_, new_n24603_, new_n24604_, new_n24605_,
    new_n24606_, new_n24607_, new_n24608_, new_n24609_, new_n24610_,
    new_n24611_, new_n24612_, new_n24613_, new_n24614_, new_n24615_,
    new_n24616_, new_n24617_, new_n24618_, new_n24619_, new_n24620_,
    new_n24621_, new_n24622_, new_n24623_, new_n24624_, new_n24625_,
    new_n24626_, new_n24627_, new_n24628_, new_n24629_, new_n24630_,
    new_n24631_, new_n24632_, new_n24633_, new_n24634_, new_n24635_,
    new_n24636_, new_n24637_, new_n24638_, new_n24639_, new_n24640_,
    new_n24641_, new_n24642_, new_n24643_, new_n24644_, new_n24645_,
    new_n24646_, new_n24647_, new_n24648_, new_n24649_, new_n24650_,
    new_n24651_, new_n24652_, new_n24653_, new_n24654_, new_n24655_,
    new_n24656_, new_n24657_, new_n24658_, new_n24659_, new_n24660_,
    new_n24661_, new_n24662_, new_n24663_, new_n24664_, new_n24665_,
    new_n24666_, new_n24667_, new_n24668_, new_n24669_, new_n24670_,
    new_n24671_, new_n24672_, new_n24673_, new_n24674_, new_n24675_,
    new_n24676_, new_n24677_, new_n24678_, new_n24679_, new_n24680_,
    new_n24681_, new_n24682_, new_n24683_, new_n24684_, new_n24685_,
    new_n24686_, new_n24687_, new_n24688_, new_n24689_, new_n24690_,
    new_n24691_, new_n24692_, new_n24693_, new_n24694_, new_n24695_,
    new_n24696_, new_n24697_, new_n24698_, new_n24699_, new_n24700_,
    new_n24701_, new_n24702_, new_n24703_, new_n24704_, new_n24705_,
    new_n24706_, new_n24707_, new_n24708_, new_n24709_, new_n24710_,
    new_n24711_, new_n24712_, new_n24713_, new_n24714_, new_n24715_,
    new_n24716_, new_n24717_, new_n24718_, new_n24719_, new_n24720_,
    new_n24721_, new_n24722_, new_n24723_, new_n24724_, new_n24725_,
    new_n24726_, new_n24727_, new_n24728_, new_n24729_, new_n24730_,
    new_n24731_, new_n24732_, new_n24733_, new_n24734_, new_n24735_,
    new_n24736_, new_n24737_, new_n24738_, new_n24739_, new_n24740_,
    new_n24741_, new_n24742_, new_n24743_, new_n24744_, new_n24745_,
    new_n24746_, new_n24747_, new_n24748_, new_n24749_, new_n24750_,
    new_n24751_, new_n24752_, new_n24753_, new_n24754_, new_n24755_,
    new_n24756_, new_n24757_, new_n24758_, new_n24759_, new_n24760_,
    new_n24761_, new_n24762_, new_n24763_, new_n24764_, new_n24765_,
    new_n24766_, new_n24767_, new_n24768_, new_n24769_, new_n24770_,
    new_n24771_, new_n24772_, new_n24773_, new_n24774_, new_n24775_,
    new_n24776_, new_n24777_, new_n24778_, new_n24779_, new_n24780_,
    new_n24781_, new_n24782_, new_n24783_, new_n24784_, new_n24785_,
    new_n24786_, new_n24787_, new_n24788_, new_n24789_, new_n24790_,
    new_n24791_, new_n24792_, new_n24793_, new_n24794_, new_n24795_,
    new_n24796_, new_n24797_, new_n24798_, new_n24799_, new_n24800_,
    new_n24801_, new_n24802_, new_n24803_, new_n24804_, new_n24805_,
    new_n24806_, new_n24807_, new_n24808_, new_n24809_, new_n24810_,
    new_n24811_, new_n24812_, new_n24813_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24820_,
    new_n24821_, new_n24822_, new_n24824_, new_n24825_, new_n24826_,
    new_n24827_, new_n24828_, new_n24829_, new_n24830_, new_n24831_,
    new_n24832_, new_n24833_, new_n24834_, new_n24835_, new_n24836_,
    new_n24837_, new_n24838_, new_n24839_, new_n24840_, new_n24841_,
    new_n24842_, new_n24843_, new_n24844_, new_n24845_, new_n24846_,
    new_n24847_, new_n24848_, new_n24849_, new_n24850_, new_n24851_,
    new_n24852_, new_n24853_, new_n24854_, new_n24855_, new_n24856_,
    new_n24857_, new_n24858_, new_n24859_, new_n24860_, new_n24861_,
    new_n24862_, new_n24863_, new_n24864_, new_n24865_, new_n24866_,
    new_n24867_, new_n24868_, new_n24869_, new_n24870_, new_n24871_,
    new_n24872_, new_n24873_, new_n24874_, new_n24875_, new_n24876_,
    new_n24877_, new_n24878_, new_n24879_, new_n24880_, new_n24881_,
    new_n24882_, new_n24883_, new_n24884_, new_n24885_, new_n24886_,
    new_n24887_, new_n24888_, new_n24889_, new_n24890_, new_n24891_,
    new_n24892_, new_n24893_, new_n24894_, new_n24895_, new_n24898_,
    new_n24899_, new_n24900_, new_n24901_, new_n24902_, new_n24903_,
    new_n24904_, new_n24905_, new_n24906_, new_n24907_, new_n24908_,
    new_n24909_, new_n24910_, new_n24911_, new_n24912_, new_n24913_,
    new_n24914_, new_n24915_, new_n24916_, new_n24917_, new_n24918_,
    new_n24919_, new_n24920_, new_n24921_, new_n24922_, new_n24923_,
    new_n24924_, new_n24925_, new_n24926_, new_n24927_, new_n24928_,
    new_n24929_, new_n24930_, new_n24931_, new_n24932_, new_n24933_,
    new_n24934_, new_n24935_, new_n24936_, new_n24937_, new_n24938_,
    new_n24939_, new_n24940_, new_n24941_, new_n24942_, new_n24943_,
    new_n24944_, new_n24945_, new_n24946_, new_n24947_, new_n24948_,
    new_n24949_, new_n24950_, new_n24951_, new_n24952_, new_n24953_,
    new_n24954_, new_n24955_, new_n24956_, new_n24957_, new_n24958_,
    new_n24959_, new_n24960_, new_n24961_, new_n24962_, new_n24963_,
    new_n24964_, new_n24965_, new_n24966_, new_n24967_, new_n24968_,
    new_n24969_, new_n24970_, new_n24971_, new_n24972_, new_n24973_,
    new_n24974_, new_n24975_, new_n24976_, new_n24977_, new_n24978_,
    new_n24979_, new_n24980_, new_n24981_, new_n24982_, new_n24983_,
    new_n24984_, new_n24985_, new_n24986_, new_n24987_, new_n24988_,
    new_n24989_, new_n24990_, new_n24991_, new_n24992_, new_n24993_,
    new_n24994_, new_n24995_, new_n24996_, new_n24997_, new_n24998_,
    new_n24999_, new_n25000_, new_n25001_, new_n25002_, new_n25003_,
    new_n25004_, new_n25005_, new_n25006_, new_n25007_, new_n25008_,
    new_n25009_, new_n25010_, new_n25011_, new_n25012_, new_n25013_,
    new_n25014_, new_n25015_, new_n25016_, new_n25017_, new_n25018_,
    new_n25019_, new_n25020_, new_n25021_, new_n25022_, new_n25023_,
    new_n25024_, new_n25025_, new_n25026_, new_n25027_, new_n25028_,
    new_n25029_, new_n25030_, new_n25031_, new_n25032_, new_n25033_,
    new_n25034_, new_n25035_, new_n25036_, new_n25037_, new_n25038_,
    new_n25039_, new_n25040_, new_n25041_, new_n25042_, new_n25043_,
    new_n25044_, new_n25045_, new_n25046_, new_n25047_, new_n25048_,
    new_n25049_, new_n25050_, new_n25051_, new_n25052_, new_n25053_,
    new_n25054_, new_n25055_, new_n25056_, new_n25057_, new_n25058_,
    new_n25059_, new_n25060_, new_n25061_, new_n25062_, new_n25063_,
    new_n25064_, new_n25065_, new_n25066_, new_n25067_, new_n25068_,
    new_n25069_, new_n25070_, new_n25071_, new_n25072_, new_n25073_,
    new_n25074_, new_n25075_, new_n25076_, new_n25077_, new_n25078_,
    new_n25079_, new_n25080_, new_n25081_, new_n25082_, new_n25083_,
    new_n25084_, new_n25085_, new_n25086_, new_n25087_, new_n25088_,
    new_n25089_, new_n25090_, new_n25091_, new_n25092_, new_n25093_,
    new_n25094_, new_n25095_, new_n25096_, new_n25097_, new_n25098_,
    new_n25099_, new_n25100_, new_n25101_, new_n25102_, new_n25103_,
    new_n25104_, new_n25105_, new_n25106_, new_n25107_, new_n25108_,
    new_n25109_, new_n25110_, new_n25111_, new_n25112_, new_n25113_,
    new_n25114_, new_n25115_, new_n25116_, new_n25117_, new_n25118_,
    new_n25119_, new_n25120_, new_n25121_, new_n25122_, new_n25123_,
    new_n25124_, new_n25125_, new_n25126_, new_n25127_, new_n25128_,
    new_n25129_, new_n25130_, new_n25131_, new_n25132_, new_n25133_,
    new_n25134_, new_n25135_, new_n25136_, new_n25137_, new_n25138_,
    new_n25139_, new_n25140_, new_n25141_, new_n25142_, new_n25143_,
    new_n25144_, new_n25145_, new_n25146_, new_n25147_, new_n25148_,
    new_n25149_, new_n25150_, new_n25151_, new_n25152_, new_n25153_,
    new_n25154_, new_n25155_, new_n25156_, new_n25157_, new_n25158_,
    new_n25159_, new_n25160_, new_n25161_, new_n25162_, new_n25163_,
    new_n25164_, new_n25165_, new_n25166_, new_n25167_, new_n25168_,
    new_n25169_, new_n25171_, new_n25172_, new_n25173_, new_n25174_,
    new_n25175_, new_n25176_, new_n25177_, new_n25178_, new_n25179_,
    new_n25180_, new_n25181_, new_n25182_, new_n25183_, new_n25184_,
    new_n25185_, new_n25186_, new_n25187_, new_n25188_, new_n25189_,
    new_n25190_, new_n25191_, new_n25192_, new_n25193_, new_n25194_,
    new_n25195_, new_n25196_, new_n25197_, new_n25198_, new_n25199_,
    new_n25200_, new_n25201_, new_n25202_, new_n25203_, new_n25204_,
    new_n25205_, new_n25206_, new_n25207_, new_n25208_, new_n25209_,
    new_n25210_, new_n25211_, new_n25212_, new_n25213_, new_n25214_,
    new_n25215_, new_n25216_, new_n25217_, new_n25218_, new_n25219_,
    new_n25220_, new_n25221_, new_n25222_, new_n25223_, new_n25224_,
    new_n25225_, new_n25226_, new_n25227_, new_n25228_, new_n25229_,
    new_n25230_, new_n25231_, new_n25232_, new_n25233_, new_n25234_,
    new_n25235_, new_n25236_, new_n25237_, new_n25238_, new_n25239_,
    new_n25240_, new_n25241_, new_n25242_, new_n25245_, new_n25246_,
    new_n25247_, new_n25248_, new_n25249_, new_n25250_, new_n25251_,
    new_n25252_, new_n25253_, new_n25254_, new_n25255_, new_n25256_,
    new_n25257_, new_n25258_, new_n25259_, new_n25260_, new_n25261_,
    new_n25262_, new_n25263_, new_n25264_, new_n25265_, new_n25266_,
    new_n25267_, new_n25268_, new_n25269_, new_n25270_, new_n25271_,
    new_n25272_, new_n25273_, new_n25274_, new_n25275_, new_n25276_,
    new_n25277_, new_n25278_, new_n25279_, new_n25280_, new_n25281_,
    new_n25282_, new_n25283_, new_n25284_, new_n25285_, new_n25286_,
    new_n25287_, new_n25288_, new_n25289_, new_n25290_, new_n25291_,
    new_n25292_, new_n25293_, new_n25294_, new_n25295_, new_n25296_,
    new_n25297_, new_n25298_, new_n25299_, new_n25300_, new_n25301_,
    new_n25302_, new_n25303_, new_n25304_, new_n25305_, new_n25306_,
    new_n25307_, new_n25308_, new_n25309_, new_n25310_, new_n25311_,
    new_n25312_, new_n25313_, new_n25314_, new_n25315_, new_n25316_,
    new_n25317_, new_n25318_, new_n25319_, new_n25320_, new_n25321_,
    new_n25322_, new_n25323_, new_n25324_, new_n25325_, new_n25326_,
    new_n25327_, new_n25328_, new_n25329_, new_n25330_, new_n25331_,
    new_n25332_, new_n25333_, new_n25334_, new_n25335_, new_n25336_,
    new_n25337_, new_n25338_, new_n25339_, new_n25340_, new_n25341_,
    new_n25342_, new_n25343_, new_n25344_, new_n25345_, new_n25346_,
    new_n25347_, new_n25348_, new_n25349_, new_n25350_, new_n25351_,
    new_n25352_, new_n25353_, new_n25354_, new_n25355_, new_n25356_,
    new_n25357_, new_n25358_, new_n25359_, new_n25360_, new_n25361_,
    new_n25362_, new_n25363_, new_n25364_, new_n25365_, new_n25366_,
    new_n25367_, new_n25368_, new_n25369_, new_n25370_, new_n25371_,
    new_n25372_, new_n25373_, new_n25374_, new_n25375_, new_n25376_,
    new_n25377_, new_n25378_, new_n25379_, new_n25380_, new_n25381_,
    new_n25382_, new_n25383_, new_n25384_, new_n25385_, new_n25386_,
    new_n25387_, new_n25388_, new_n25389_, new_n25390_, new_n25391_,
    new_n25392_, new_n25393_, new_n25394_, new_n25395_, new_n25396_,
    new_n25397_, new_n25398_, new_n25399_, new_n25400_, new_n25401_,
    new_n25402_, new_n25403_, new_n25404_, new_n25405_, new_n25406_,
    new_n25407_, new_n25408_, new_n25409_, new_n25410_, new_n25411_,
    new_n25412_, new_n25413_, new_n25414_, new_n25415_, new_n25416_,
    new_n25417_, new_n25418_, new_n25419_, new_n25420_, new_n25421_,
    new_n25422_, new_n25423_, new_n25424_, new_n25425_, new_n25426_,
    new_n25427_, new_n25428_, new_n25429_, new_n25430_, new_n25431_,
    new_n25432_, new_n25433_, new_n25434_, new_n25435_, new_n25436_,
    new_n25437_, new_n25438_, new_n25439_, new_n25440_, new_n25441_,
    new_n25442_, new_n25443_, new_n25444_, new_n25445_, new_n25446_,
    new_n25447_, new_n25448_, new_n25449_, new_n25450_, new_n25451_,
    new_n25452_, new_n25453_, new_n25454_, new_n25455_, new_n25456_,
    new_n25457_, new_n25458_, new_n25459_, new_n25460_, new_n25461_,
    new_n25462_, new_n25463_, new_n25464_, new_n25465_, new_n25466_,
    new_n25467_, new_n25468_, new_n25469_, new_n25470_, new_n25471_,
    new_n25472_, new_n25473_, new_n25474_, new_n25475_, new_n25476_,
    new_n25477_, new_n25478_, new_n25479_, new_n25480_, new_n25481_,
    new_n25482_, new_n25483_, new_n25484_, new_n25485_, new_n25486_,
    new_n25487_, new_n25488_, new_n25489_, new_n25490_, new_n25491_,
    new_n25492_, new_n25493_, new_n25494_, new_n25495_, new_n25496_,
    new_n25497_, new_n25498_, new_n25499_, new_n25500_, new_n25501_,
    new_n25502_, new_n25503_, new_n25504_, new_n25505_, new_n25506_,
    new_n25507_, new_n25508_, new_n25509_, new_n25510_, new_n25511_,
    new_n25512_, new_n25513_, new_n25514_, new_n25515_, new_n25516_,
    new_n25518_, new_n25519_, new_n25520_, new_n25521_, new_n25522_,
    new_n25523_, new_n25524_, new_n25525_, new_n25526_, new_n25527_,
    new_n25528_, new_n25529_, new_n25530_, new_n25531_, new_n25532_,
    new_n25533_, new_n25534_, new_n25535_, new_n25536_, new_n25537_,
    new_n25538_, new_n25539_, new_n25540_, new_n25541_, new_n25542_,
    new_n25543_, new_n25544_, new_n25545_, new_n25546_, new_n25547_,
    new_n25548_, new_n25549_, new_n25550_, new_n25551_, new_n25552_,
    new_n25553_, new_n25554_, new_n25555_, new_n25556_, new_n25557_,
    new_n25558_, new_n25559_, new_n25560_, new_n25561_, new_n25562_,
    new_n25563_, new_n25564_, new_n25565_, new_n25566_, new_n25567_,
    new_n25568_, new_n25569_, new_n25570_, new_n25571_, new_n25572_,
    new_n25573_, new_n25574_, new_n25575_, new_n25576_, new_n25577_,
    new_n25578_, new_n25579_, new_n25580_, new_n25581_, new_n25582_,
    new_n25583_, new_n25584_, new_n25585_, new_n25586_, new_n25587_,
    new_n25588_, new_n25589_, new_n25590_, new_n25591_, new_n25592_,
    new_n25593_, new_n25594_, new_n25595_, new_n25596_, new_n25597_,
    new_n25598_, new_n25599_, new_n25600_, new_n25601_, new_n25602_,
    new_n25603_, new_n25604_, new_n25605_, new_n25606_, new_n25607_,
    new_n25608_, new_n25609_, new_n25610_, new_n25611_, new_n25612_,
    new_n25613_, new_n25614_, new_n25615_, new_n25616_, new_n25617_,
    new_n25618_, new_n25619_, new_n25620_, new_n25621_, new_n25622_,
    new_n25623_, new_n25624_, new_n25625_, new_n25626_, new_n25627_,
    new_n25628_, new_n25629_, new_n25630_, new_n25631_, new_n25632_,
    new_n25634_, new_n25635_, new_n25636_, new_n25637_, new_n25638_,
    new_n25639_, new_n25640_, new_n25641_, new_n25642_, new_n25643_,
    new_n25644_, new_n25645_, new_n25646_, new_n25647_, new_n25648_,
    new_n25649_, new_n25650_, new_n25651_, new_n25652_, new_n25653_,
    new_n25654_, new_n25655_, new_n25656_, new_n25657_, new_n25658_,
    new_n25659_, new_n25660_, new_n25661_, new_n25662_, new_n25663_,
    new_n25664_, new_n25665_, new_n25666_, new_n25667_, new_n25668_,
    new_n25669_, new_n25670_, new_n25671_, new_n25672_, new_n25673_,
    new_n25674_, new_n25675_, new_n25676_, new_n25677_, new_n25678_,
    new_n25679_, new_n25680_, new_n25681_, new_n25682_, new_n25683_,
    new_n25684_, new_n25685_, new_n25686_, new_n25687_, new_n25688_,
    new_n25689_, new_n25690_, new_n25691_, new_n25692_, new_n25693_,
    new_n25694_, new_n25695_, new_n25696_, new_n25697_, new_n25698_,
    new_n25699_, new_n25700_, new_n25701_, new_n25702_, new_n25703_,
    new_n25704_, new_n25705_, new_n25706_, new_n25707_, new_n25708_,
    new_n25709_, new_n25710_, new_n25711_, new_n25712_, new_n25713_,
    new_n25714_, new_n25715_, new_n25716_, new_n25717_, new_n25718_,
    new_n25719_, new_n25720_, new_n25721_, new_n25722_, new_n25723_,
    new_n25724_, new_n25725_, new_n25726_, new_n25727_, new_n25728_,
    new_n25729_, new_n25730_, new_n25731_, new_n25732_, new_n25733_,
    new_n25734_, new_n25735_, new_n25736_, new_n25737_, new_n25738_,
    new_n25739_, new_n25740_, new_n25741_, new_n25742_, new_n25743_,
    new_n25744_, new_n25745_, new_n25746_, new_n25747_, new_n25748_,
    new_n25749_, new_n25750_, new_n25751_, new_n25752_, new_n25753_,
    new_n25754_, new_n25755_, new_n25756_, new_n25757_, new_n25758_,
    new_n25759_, new_n25760_, new_n25761_, new_n25762_, new_n25763_,
    new_n25764_, new_n25765_, new_n25766_, new_n25767_, new_n25768_,
    new_n25769_, new_n25770_, new_n25771_, new_n25772_, new_n25773_,
    new_n25774_, new_n25775_, new_n25776_, new_n25777_, new_n25778_,
    new_n25779_, new_n25780_, new_n25781_, new_n25782_, new_n25783_,
    new_n25784_, new_n25785_, new_n25786_, new_n25787_, new_n25788_,
    new_n25789_, new_n25790_, new_n25791_, new_n25792_, new_n25793_,
    new_n25794_, new_n25795_, new_n25796_, new_n25797_, new_n25798_,
    new_n25799_, new_n25800_, new_n25801_, new_n25802_, new_n25803_,
    new_n25804_, new_n25805_, new_n25806_, new_n25810_, new_n25811_,
    new_n25812_, new_n25813_, new_n25814_, new_n25815_, new_n25816_,
    new_n25817_, new_n25818_, new_n25819_, new_n25820_, new_n25821_,
    new_n25822_, new_n25823_, new_n25824_, new_n25825_, new_n25826_,
    new_n25827_, new_n25828_, new_n25829_, new_n25830_, new_n25831_,
    new_n25832_, new_n25833_, new_n25834_, new_n25835_, new_n25836_,
    new_n25837_, new_n25838_, new_n25839_, new_n25840_, new_n25841_,
    new_n25842_, new_n25843_, new_n25844_, new_n25845_, new_n25846_,
    new_n25847_, new_n25848_, new_n25849_, new_n25850_, new_n25851_,
    new_n25852_, new_n25853_, new_n25854_, new_n25855_, new_n25856_,
    new_n25857_, new_n25858_, new_n25859_, new_n25860_, new_n25861_,
    new_n25862_, new_n25863_, new_n25864_, new_n25865_, new_n25866_,
    new_n25867_, new_n25868_, new_n25869_, new_n25870_, new_n25871_,
    new_n25872_, new_n25873_, new_n25874_, new_n25875_, new_n25876_,
    new_n25878_, new_n25879_, new_n25880_, new_n25881_, new_n25882_,
    new_n25883_, new_n25884_, new_n25885_, new_n25886_, new_n25887_,
    new_n25888_, new_n25889_, new_n25890_, new_n25891_, new_n25892_,
    new_n25893_, new_n25894_, new_n25895_, new_n25896_, new_n25897_,
    new_n25898_, new_n25899_, new_n25900_, new_n25901_, new_n25902_,
    new_n25903_, new_n25904_, new_n25905_, new_n25906_, new_n25907_,
    new_n25908_, new_n25909_, new_n25910_, new_n25911_, new_n25912_,
    new_n25913_, new_n25914_, new_n25915_, new_n25916_, new_n25917_,
    new_n25918_, new_n25919_, new_n25920_, new_n25921_, new_n25922_,
    new_n25923_, new_n25924_, new_n25925_, new_n25926_, new_n25927_,
    new_n25928_, new_n25929_, new_n25930_, new_n25931_, new_n25932_,
    new_n25933_, new_n25934_, new_n25935_, new_n25936_, new_n25937_,
    new_n25938_, new_n25939_, new_n25940_, new_n25941_, new_n25942_,
    new_n25943_, new_n25944_, new_n25945_, new_n25946_, new_n25947_,
    new_n25948_, new_n25949_, new_n25951_, new_n25952_, new_n25953_,
    new_n25954_, new_n25955_, new_n25956_, new_n25957_, new_n25958_,
    new_n25959_, new_n25960_, new_n25961_, new_n25962_, new_n25963_,
    new_n25964_, new_n25965_, new_n25966_, new_n25967_, new_n25968_,
    new_n25969_, new_n25970_, new_n25971_, new_n25972_, new_n25973_,
    new_n25974_, new_n25975_, new_n25976_, new_n25977_, new_n25978_,
    new_n25979_, new_n25980_, new_n25981_, new_n25982_, new_n25983_,
    new_n25984_, new_n25985_, new_n25986_, new_n25987_, new_n25988_,
    new_n25989_, new_n25990_, new_n25991_, new_n25992_, new_n25993_,
    new_n25994_, new_n25995_, new_n25996_, new_n25997_, new_n25998_,
    new_n25999_, new_n26000_, new_n26001_, new_n26002_, new_n26003_,
    new_n26004_, new_n26005_, new_n26006_, new_n26007_, new_n26008_,
    new_n26009_, new_n26010_, new_n26011_, new_n26012_, new_n26013_,
    new_n26014_, new_n26015_, new_n26016_, new_n26017_, new_n26018_,
    new_n26019_, new_n26020_, new_n26021_, new_n26022_, new_n26023_,
    new_n26024_, new_n26025_, new_n26026_, new_n26027_, new_n26028_,
    new_n26029_, new_n26030_, new_n26031_, new_n26032_, new_n26033_,
    new_n26034_, new_n26035_, new_n26036_, new_n26037_, new_n26038_,
    new_n26039_, new_n26040_, new_n26041_, new_n26042_, new_n26043_,
    new_n26044_, new_n26045_, new_n26046_, new_n26047_, new_n26048_,
    new_n26049_, new_n26050_, new_n26051_, new_n26052_, new_n26053_,
    new_n26054_, new_n26055_, new_n26056_, new_n26057_, new_n26058_,
    new_n26059_, new_n26060_, new_n26061_, new_n26062_, new_n26063_,
    new_n26064_, new_n26065_, new_n26066_, new_n26067_, new_n26068_,
    new_n26069_, new_n26070_, new_n26071_, new_n26072_, new_n26073_,
    new_n26077_, new_n26078_, new_n26079_, new_n26080_, new_n26081_,
    new_n26082_, new_n26083_, new_n26084_, new_n26085_, new_n26086_,
    new_n26087_, new_n26088_, new_n26089_, new_n26090_, new_n26091_,
    new_n26092_, new_n26093_, new_n26094_, new_n26095_, new_n26096_,
    new_n26097_, new_n26098_, new_n26099_, new_n26100_, new_n26101_,
    new_n26102_, new_n26104_, new_n26105_, new_n26106_, new_n26108_,
    new_n26109_, new_n26110_, new_n26112_, new_n26113_, new_n26114_,
    new_n26115_, new_n26116_, new_n26117_, new_n26118_, new_n26119_,
    new_n26120_, new_n26121_, new_n26122_, new_n26123_, new_n26124_,
    new_n26125_, new_n26126_, new_n26127_, new_n26128_, new_n26129_,
    new_n26130_, new_n26131_, new_n26132_, new_n26133_, new_n26134_,
    new_n26135_, new_n26136_, new_n26137_, new_n26138_, new_n26139_,
    new_n26140_, new_n26141_, new_n26142_, new_n26143_, new_n26144_,
    new_n26145_, new_n26146_, new_n26147_, new_n26148_, new_n26149_,
    new_n26150_, new_n26151_, new_n26152_, new_n26153_, new_n26154_,
    new_n26155_, new_n26156_, new_n26157_, new_n26158_, new_n26159_,
    new_n26160_, new_n26161_, new_n26162_, new_n26163_, new_n26164_,
    new_n26165_, new_n26166_, new_n26167_, new_n26168_, new_n26169_,
    new_n26170_, new_n26171_, new_n26172_, new_n26173_, new_n26174_,
    new_n26175_, new_n26176_, new_n26177_, new_n26178_, new_n26179_,
    new_n26180_, new_n26181_, new_n26182_, new_n26183_, new_n26184_,
    new_n26185_, new_n26186_, new_n26187_, new_n26188_, new_n26189_,
    new_n26190_, new_n26191_, new_n26192_, new_n26193_, new_n26194_,
    new_n26195_, new_n26196_, new_n26197_, new_n26198_, new_n26199_,
    new_n26200_, new_n26201_, new_n26202_, new_n26203_, new_n26204_,
    new_n26205_, new_n26206_, new_n26207_, new_n26208_, new_n26209_,
    new_n26210_, new_n26211_, new_n26212_, new_n26213_, new_n26214_,
    new_n26215_, new_n26216_, new_n26217_, new_n26218_, new_n26219_,
    new_n26220_, new_n26221_, new_n26222_, new_n26223_, new_n26224_,
    new_n26225_, new_n26226_, new_n26227_, new_n26228_, new_n26229_,
    new_n26230_, new_n26231_, new_n26232_, new_n26233_, new_n26234_,
    new_n26235_, new_n26236_, new_n26237_, new_n26238_, new_n26239_,
    new_n26240_, new_n26241_, new_n26242_, new_n26243_, new_n26244_,
    new_n26245_, new_n26246_, new_n26247_, new_n26248_, new_n26249_,
    new_n26250_, new_n26251_, new_n26252_, new_n26253_, new_n26254_,
    new_n26255_, new_n26256_, new_n26257_, new_n26258_, new_n26259_,
    new_n26260_, new_n26261_, new_n26262_, new_n26263_, new_n26264_,
    new_n26265_, new_n26266_, new_n26267_, new_n26268_, new_n26269_,
    new_n26270_, new_n26271_, new_n26272_, new_n26273_, new_n26274_,
    new_n26275_, new_n26276_, new_n26277_, new_n26278_, new_n26279_,
    new_n26280_, new_n26281_, new_n26282_, new_n26283_, new_n26284_,
    new_n26285_, new_n26286_, new_n26287_, new_n26288_, new_n26289_,
    new_n26290_, new_n26291_, new_n26292_, new_n26293_, new_n26294_,
    new_n26295_, new_n26296_, new_n26297_, new_n26298_, new_n26299_,
    new_n26300_, new_n26301_, new_n26302_, new_n26303_, new_n26304_,
    new_n26305_, new_n26306_, new_n26307_, new_n26308_, new_n26309_,
    new_n26310_, new_n26311_, new_n26312_, new_n26313_, new_n26314_,
    new_n26315_, new_n26316_, new_n26318_, new_n26319_, new_n26320_,
    new_n26321_, new_n26322_, new_n26323_, new_n26324_, new_n26325_,
    new_n26326_, new_n26327_, new_n26328_, new_n26329_, new_n26330_,
    new_n26331_, new_n26332_, new_n26333_, new_n26334_, new_n26335_,
    new_n26336_, new_n26337_, new_n26338_, new_n26339_, new_n26340_,
    new_n26341_, new_n26342_, new_n26343_, new_n26344_, new_n26345_,
    new_n26347_, new_n26348_, new_n26349_, new_n26350_, new_n26351_,
    new_n26352_, new_n26353_, new_n26354_, new_n26355_, new_n26356_,
    new_n26357_, new_n26358_, new_n26359_, new_n26360_, new_n26361_,
    new_n26362_, new_n26363_, new_n26364_, new_n26365_, new_n26366_,
    new_n26367_, new_n26368_, new_n26369_, new_n26370_, new_n26371_,
    new_n26372_, new_n26373_, new_n26374_, new_n26375_, new_n26376_,
    new_n26377_, new_n26378_, new_n26379_, new_n26380_, new_n26381_,
    new_n26382_, new_n26383_, new_n26384_, new_n26385_, new_n26386_,
    new_n26387_, new_n26388_, new_n26389_, new_n26391_, new_n26392_,
    new_n26393_, new_n26394_, new_n26395_, new_n26396_, new_n26397_,
    new_n26398_, new_n26399_, new_n26400_, new_n26401_, new_n26402_,
    new_n26403_, new_n26404_, new_n26405_, new_n26406_, new_n26407_,
    new_n26408_, new_n26409_, new_n26410_, new_n26411_, new_n26412_,
    new_n26413_, new_n26414_, new_n26415_, new_n26416_, new_n26417_,
    new_n26418_, new_n26419_, new_n26420_, new_n26421_, new_n26422_,
    new_n26423_, new_n26424_, new_n26425_, new_n26427_, new_n26428_,
    new_n26429_, new_n26430_, new_n26431_, new_n26432_, new_n26433_,
    new_n26434_, new_n26435_, new_n26436_, new_n26437_, new_n26438_,
    new_n26439_, new_n26440_, new_n26441_, new_n26442_, new_n26443_,
    new_n26444_, new_n26445_, new_n26446_, new_n26447_, new_n26448_,
    new_n26449_, new_n26450_, new_n26451_, new_n26452_, new_n26453_,
    new_n26454_, new_n26455_, new_n26456_, new_n26457_, new_n26458_,
    new_n26459_, new_n26460_, new_n26461_, new_n26462_, new_n26463_,
    new_n26464_, new_n26465_, new_n26466_, new_n26467_, new_n26468_,
    new_n26469_, new_n26470_, new_n26471_, new_n26472_, new_n26473_,
    new_n26474_, new_n26475_, new_n26476_, new_n26477_, new_n26478_,
    new_n26479_, new_n26480_, new_n26482_, new_n26483_, new_n26484_,
    new_n26485_, new_n26486_, new_n26487_, new_n26488_, new_n26489_,
    new_n26490_, new_n26491_, new_n26492_, new_n26493_, new_n26494_,
    new_n26495_, new_n26496_, new_n26497_, new_n26498_, new_n26499_,
    new_n26500_, new_n26501_, new_n26502_, new_n26503_, new_n26504_,
    new_n26505_, new_n26506_, new_n26507_, new_n26508_, new_n26509_,
    new_n26510_, new_n26511_, new_n26512_, new_n26513_, new_n26514_,
    new_n26515_, new_n26516_, new_n26517_, new_n26518_, new_n26519_,
    new_n26520_, new_n26521_, new_n26522_, new_n26523_, new_n26524_,
    new_n26525_, new_n26526_, new_n26527_, new_n26528_, new_n26529_,
    new_n26530_, new_n26531_, new_n26532_, new_n26533_, new_n26534_,
    new_n26535_, new_n26536_, new_n26537_, new_n26538_, new_n26539_,
    new_n26540_, new_n26541_, new_n26542_, new_n26543_, new_n26544_,
    new_n26545_, new_n26546_, new_n26547_, new_n26548_, new_n26549_,
    new_n26550_, new_n26551_, new_n26552_, new_n26553_, new_n26554_,
    new_n26555_, new_n26556_, new_n26557_, new_n26558_, new_n26559_,
    new_n26560_, new_n26561_, new_n26562_, new_n26563_, new_n26564_,
    new_n26565_, new_n26566_, new_n26567_, new_n26568_, new_n26569_,
    new_n26570_, new_n26571_, new_n26572_, new_n26573_, new_n26574_,
    new_n26575_, new_n26576_, new_n26577_, new_n26578_, new_n26579_,
    new_n26580_, new_n26581_, new_n26582_, new_n26583_, new_n26584_,
    new_n26585_, new_n26586_, new_n26587_, new_n26588_, new_n26589_,
    new_n26590_, new_n26591_, new_n26592_, new_n26593_, new_n26594_,
    new_n26595_, new_n26596_, new_n26597_, new_n26598_, new_n26599_,
    new_n26600_, new_n26601_, new_n26602_, new_n26603_, new_n26604_,
    new_n26605_, new_n26606_, new_n26607_, new_n26608_, new_n26609_,
    new_n26610_, new_n26611_, new_n26612_, new_n26613_, new_n26614_,
    new_n26615_, new_n26616_, new_n26617_, new_n26618_, new_n26619_,
    new_n26620_, new_n26621_, new_n26622_, new_n26623_, new_n26624_,
    new_n26625_, new_n26626_, new_n26627_, new_n26628_, new_n26629_,
    new_n26630_, new_n26631_, new_n26632_, new_n26633_, new_n26634_,
    new_n26635_, new_n26636_, new_n26637_, new_n26638_, new_n26639_,
    new_n26640_, new_n26641_, new_n26642_, new_n26643_, new_n26644_,
    new_n26645_, new_n26646_, new_n26647_, new_n26648_, new_n26649_,
    new_n26650_, new_n26651_, new_n26652_, new_n26653_, new_n26654_,
    new_n26655_, new_n26656_, new_n26657_, new_n26658_, new_n26659_,
    new_n26660_, new_n26661_, new_n26662_, new_n26663_, new_n26664_,
    new_n26665_, new_n26666_, new_n26667_, new_n26668_, new_n26669_,
    new_n26670_, new_n26671_, new_n26672_, new_n26673_, new_n26674_,
    new_n26675_, new_n26676_, new_n26677_, new_n26678_, new_n26679_,
    new_n26680_, new_n26681_, new_n26682_, new_n26683_, new_n26684_,
    new_n26685_, new_n26686_, new_n26687_, new_n26688_, new_n26689_,
    new_n26690_, new_n26691_, new_n26692_, new_n26693_, new_n26694_,
    new_n26695_, new_n26696_, new_n26697_, new_n26698_, new_n26699_,
    new_n26700_, new_n26701_, new_n26702_, new_n26703_, new_n26704_,
    new_n26705_, new_n26706_, new_n26707_, new_n26708_, new_n26709_,
    new_n26710_, new_n26711_, new_n26712_, new_n26713_, new_n26714_,
    new_n26715_, new_n26716_, new_n26717_, new_n26718_, new_n26719_,
    new_n26720_, new_n26721_, new_n26722_, new_n26723_, new_n26724_,
    new_n26725_, new_n26726_, new_n26727_, new_n26728_, new_n26729_,
    new_n26730_, new_n26731_, new_n26732_, new_n26733_, new_n26734_,
    new_n26735_, new_n26736_, new_n26737_, new_n26738_, new_n26739_,
    new_n26740_, new_n26741_, new_n26742_, new_n26743_, new_n26744_,
    new_n26745_, new_n26746_, new_n26747_, new_n26748_, new_n26749_,
    new_n26750_, new_n26751_, new_n26754_, new_n26755_, new_n26756_,
    new_n26757_, new_n26758_, new_n26759_, new_n26760_, new_n26761_,
    new_n26762_, new_n26763_, new_n26764_, new_n26765_, new_n26766_,
    new_n26767_, new_n26768_, new_n26769_, new_n26770_, new_n26771_,
    new_n26772_, new_n26773_, new_n26774_, new_n26775_, new_n26776_,
    new_n26777_, new_n26778_, new_n26779_, new_n26780_, new_n26781_,
    new_n26782_, new_n26783_, new_n26784_, new_n26785_, new_n26786_,
    new_n26787_, new_n26788_, new_n26789_, new_n26790_, new_n26791_,
    new_n26792_, new_n26793_, new_n26794_, new_n26795_, new_n26796_,
    new_n26797_, new_n26798_, new_n26799_, new_n26800_, new_n26801_,
    new_n26802_, new_n26803_, new_n26804_, new_n26805_, new_n26806_,
    new_n26807_, new_n26808_, new_n26809_, new_n26810_, new_n26811_,
    new_n26812_, new_n26813_, new_n26814_, new_n26815_, new_n26816_,
    new_n26817_, new_n26818_, new_n26819_, new_n26820_, new_n26821_,
    new_n26822_, new_n26823_, new_n26824_, new_n26825_, new_n26826_,
    new_n26827_, new_n26828_, new_n26829_, new_n26830_, new_n26831_,
    new_n26833_, new_n26834_, new_n26835_, new_n26836_, new_n26837_,
    new_n26838_, new_n26839_, new_n26840_, new_n26841_, new_n26842_,
    new_n26843_, new_n26844_, new_n26845_, new_n26846_, new_n26847_,
    new_n26848_, new_n26849_, new_n26850_, new_n26851_, new_n26852_,
    new_n26853_, new_n26854_, new_n26855_, new_n26856_, new_n26857_,
    new_n26858_, new_n26859_, new_n26860_, new_n26861_, new_n26862_,
    new_n26863_, new_n26864_, new_n26865_, new_n26866_, new_n26867_,
    new_n26868_, new_n26869_, new_n26870_, new_n26871_, new_n26872_,
    new_n26873_, new_n26874_, new_n26875_, new_n26876_, new_n26877_,
    new_n26878_, new_n26879_, new_n26880_, new_n26881_, new_n26882_,
    new_n26883_, new_n26884_, new_n26885_, new_n26886_, new_n26887_,
    new_n26888_, new_n26889_, new_n26890_, new_n26891_, new_n26892_,
    new_n26893_, new_n26894_, new_n26895_, new_n26896_, new_n26897_,
    new_n26898_, new_n26899_, new_n26900_, new_n26901_, new_n26902_,
    new_n26903_, new_n26904_, new_n26905_, new_n26906_, new_n26907_,
    new_n26908_, new_n26909_, new_n26910_, new_n26911_, new_n26912_,
    new_n26913_, new_n26914_, new_n26915_, new_n26916_, new_n26917_,
    new_n26918_, new_n26919_, new_n26920_, new_n26921_, new_n26922_,
    new_n26923_, new_n26924_, new_n26925_, new_n26926_, new_n26927_,
    new_n26928_, new_n26929_, new_n26930_, new_n26931_, new_n26932_,
    new_n26933_, new_n26934_, new_n26935_, new_n26936_, new_n26937_,
    new_n26938_, new_n26939_, new_n26940_, new_n26941_, new_n26942_,
    new_n26943_, new_n26944_, new_n26945_, new_n26946_, new_n26947_,
    new_n26948_, new_n26949_, new_n26950_, new_n26951_, new_n26952_,
    new_n26953_, new_n26954_, new_n26955_, new_n26958_, new_n26959_,
    new_n26960_, new_n26962_, new_n26963_, new_n26964_, new_n26965_,
    new_n26966_, new_n26967_, new_n26968_, new_n26969_, new_n26970_,
    new_n26971_, new_n26972_, new_n26973_, new_n26974_, new_n26975_,
    new_n26976_, new_n26977_, new_n26978_, new_n26979_, new_n26980_,
    new_n26981_, new_n26982_, new_n26983_, new_n26984_, new_n26985_,
    new_n26986_, new_n26987_, new_n26988_, new_n26989_, new_n26990_,
    new_n26991_, new_n26992_, new_n26993_, new_n26994_, new_n26995_,
    new_n26996_, new_n26997_, new_n26998_, new_n26999_, new_n27000_,
    new_n27001_, new_n27002_, new_n27003_, new_n27004_, new_n27005_,
    new_n27006_, new_n27007_, new_n27008_, new_n27009_, new_n27010_,
    new_n27011_, new_n27012_, new_n27013_, new_n27014_, new_n27015_,
    new_n27016_, new_n27017_, new_n27018_, new_n27019_, new_n27020_,
    new_n27021_, new_n27022_, new_n27023_, new_n27024_, new_n27025_,
    new_n27026_, new_n27027_, new_n27028_, new_n27029_, new_n27030_,
    new_n27031_, new_n27032_, new_n27033_, new_n27034_, new_n27035_,
    new_n27036_, new_n27037_, new_n27038_, new_n27039_, new_n27040_,
    new_n27041_, new_n27042_, new_n27043_, new_n27044_, new_n27045_,
    new_n27046_, new_n27047_, new_n27048_, new_n27049_, new_n27050_,
    new_n27051_, new_n27052_, new_n27053_, new_n27054_, new_n27055_,
    new_n27056_, new_n27057_, new_n27058_, new_n27059_, new_n27060_,
    new_n27061_, new_n27062_, new_n27063_, new_n27064_, new_n27065_,
    new_n27066_, new_n27067_, new_n27068_, new_n27069_, new_n27070_,
    new_n27071_, new_n27072_, new_n27073_, new_n27074_, new_n27075_,
    new_n27076_, new_n27077_, new_n27078_, new_n27079_, new_n27080_,
    new_n27081_, new_n27082_, new_n27083_, new_n27084_, new_n27085_,
    new_n27086_, new_n27087_, new_n27088_, new_n27089_, new_n27090_,
    new_n27091_, new_n27092_, new_n27093_, new_n27094_, new_n27095_,
    new_n27096_, new_n27097_, new_n27098_, new_n27099_, new_n27100_,
    new_n27101_, new_n27102_, new_n27103_, new_n27104_, new_n27105_,
    new_n27106_, new_n27107_, new_n27108_, new_n27109_, new_n27110_,
    new_n27111_, new_n27112_, new_n27113_, new_n27114_, new_n27115_,
    new_n27116_, new_n27117_, new_n27118_, new_n27119_, new_n27120_,
    new_n27121_, new_n27122_, new_n27123_, new_n27124_, new_n27125_,
    new_n27126_, new_n27127_, new_n27128_, new_n27129_, new_n27130_,
    new_n27131_, new_n27132_, new_n27133_, new_n27134_, new_n27135_,
    new_n27136_, new_n27137_, new_n27138_, new_n27139_, new_n27143_,
    new_n27144_, new_n27145_, new_n27146_, new_n27147_, new_n27148_,
    new_n27149_, new_n27150_, new_n27151_, new_n27152_, new_n27153_,
    new_n27154_, new_n27155_, new_n27156_, new_n27157_, new_n27158_,
    new_n27159_, new_n27160_, new_n27161_, new_n27162_, new_n27163_,
    new_n27164_, new_n27165_, new_n27166_, new_n27167_, new_n27168_,
    new_n27169_, new_n27170_, new_n27171_, new_n27172_, new_n27173_,
    new_n27174_, new_n27175_, new_n27176_, new_n27177_, new_n27179_,
    new_n27180_, new_n27182_, new_n27183_, new_n27184_, new_n27186_,
    new_n27187_, new_n27188_, new_n27189_, new_n27190_, new_n27191_,
    new_n27192_, new_n27193_, new_n27194_, new_n27195_, new_n27196_,
    new_n27197_, new_n27198_, new_n27199_, new_n27200_, new_n27201_,
    new_n27202_, new_n27203_, new_n27204_, new_n27205_, new_n27206_,
    new_n27207_, new_n27208_, new_n27209_, new_n27210_, new_n27211_,
    new_n27212_, new_n27213_, new_n27214_, new_n27215_, new_n27216_,
    new_n27217_, new_n27218_, new_n27219_, new_n27220_, new_n27221_,
    new_n27222_, new_n27223_, new_n27224_, new_n27225_, new_n27226_,
    new_n27227_, new_n27228_, new_n27229_, new_n27230_, new_n27231_,
    new_n27232_, new_n27233_, new_n27234_, new_n27235_, new_n27236_,
    new_n27237_, new_n27238_, new_n27239_, new_n27240_, new_n27241_,
    new_n27244_, new_n27245_, new_n27246_, new_n27247_, new_n27248_,
    new_n27249_, new_n27250_, new_n27251_, new_n27252_, new_n27254_,
    new_n27255_, new_n27256_, new_n27257_, new_n27258_, new_n27259_,
    new_n27260_, new_n27261_, new_n27262_, new_n27263_, new_n27264_,
    new_n27265_, new_n27266_, new_n27267_, new_n27268_, new_n27269_,
    new_n27270_, new_n27271_, new_n27272_, new_n27273_, new_n27274_,
    new_n27275_, new_n27276_, new_n27277_, new_n27278_, new_n27279_,
    new_n27280_, new_n27281_, new_n27282_, new_n27283_, new_n27284_,
    new_n27285_, new_n27286_, new_n27287_, new_n27288_, new_n27289_,
    new_n27290_, new_n27291_, new_n27292_, new_n27293_, new_n27294_,
    new_n27295_, new_n27296_, new_n27297_, new_n27298_, new_n27299_,
    new_n27300_, new_n27301_, new_n27302_, new_n27303_, new_n27304_,
    new_n27305_, new_n27306_, new_n27307_, new_n27308_, new_n27309_,
    new_n27310_, new_n27311_, new_n27312_, new_n27313_, new_n27314_,
    new_n27315_, new_n27316_, new_n27317_, new_n27318_, new_n27319_,
    new_n27320_, new_n27321_, new_n27322_, new_n27323_, new_n27324_,
    new_n27325_, new_n27326_, new_n27327_, new_n27328_, new_n27329_,
    new_n27330_, new_n27331_, new_n27332_, new_n27333_, new_n27334_,
    new_n27335_, new_n27336_, new_n27337_, new_n27338_, new_n27339_,
    new_n27340_, new_n27341_, new_n27342_, new_n27343_, new_n27344_,
    new_n27345_, new_n27346_, new_n27347_, new_n27348_, new_n27349_,
    new_n27350_, new_n27351_, new_n27352_, new_n27353_, new_n27354_,
    new_n27355_, new_n27356_, new_n27357_, new_n27358_, new_n27359_,
    new_n27360_, new_n27361_, new_n27362_, new_n27363_, new_n27364_,
    new_n27365_, new_n27366_, new_n27367_, new_n27368_, new_n27369_,
    new_n27370_, new_n27371_, new_n27372_, new_n27373_, new_n27374_,
    new_n27375_, new_n27376_, new_n27377_, new_n27378_, new_n27379_,
    new_n27380_, new_n27381_, new_n27382_, new_n27383_, new_n27384_,
    new_n27385_, new_n27386_, new_n27387_, new_n27388_, new_n27389_,
    new_n27390_, new_n27391_, new_n27392_, new_n27393_, new_n27394_,
    new_n27395_, new_n27396_, new_n27397_, new_n27398_, new_n27399_,
    new_n27400_, new_n27401_, new_n27402_, new_n27403_, new_n27404_,
    new_n27405_, new_n27406_, new_n27407_, new_n27408_, new_n27409_,
    new_n27410_, new_n27411_, new_n27412_, new_n27413_, new_n27414_,
    new_n27415_, new_n27416_, new_n27417_, new_n27418_, new_n27419_,
    new_n27420_, new_n27421_, new_n27422_, new_n27423_, new_n27424_,
    new_n27425_, new_n27426_, new_n27427_, new_n27428_, new_n27429_,
    new_n27430_, new_n27431_, new_n27432_, new_n27433_, new_n27434_,
    new_n27435_, new_n27436_, new_n27437_, new_n27438_, new_n27439_,
    new_n27440_, new_n27441_, new_n27442_, new_n27443_, new_n27444_,
    new_n27445_, new_n27446_, new_n27447_, new_n27448_, new_n27449_,
    new_n27450_, new_n27451_, new_n27452_, new_n27453_, new_n27454_,
    new_n27455_, new_n27456_, new_n27457_, new_n27458_, new_n27459_,
    new_n27460_, new_n27461_, new_n27462_, new_n27463_, new_n27464_,
    new_n27465_, new_n27466_, new_n27467_, new_n27468_, new_n27469_,
    new_n27470_, new_n27471_, new_n27472_, new_n27473_, new_n27474_,
    new_n27475_, new_n27476_, new_n27477_, new_n27478_, new_n27479_,
    new_n27480_, new_n27481_, new_n27482_, new_n27483_, new_n27484_,
    new_n27485_, new_n27486_, new_n27487_, new_n27488_, new_n27489_,
    new_n27490_, new_n27491_, new_n27492_, new_n27493_, new_n27494_,
    new_n27495_, new_n27496_, new_n27497_, new_n27498_, new_n27499_,
    new_n27500_, new_n27501_, new_n27502_, new_n27503_, new_n27504_,
    new_n27505_, new_n27506_, new_n27507_, new_n27508_, new_n27509_,
    new_n27510_, new_n27511_, new_n27512_, new_n27513_, new_n27514_,
    new_n27515_, new_n27516_, new_n27517_, new_n27518_, new_n27519_,
    new_n27520_, new_n27521_, new_n27522_, new_n27527_, new_n27528_,
    new_n27529_, new_n27530_, new_n27531_, new_n27532_, new_n27533_,
    new_n27535_, new_n27536_, new_n27537_, new_n27538_, new_n27539_,
    new_n27540_, new_n27541_, new_n27542_, new_n27543_, new_n27544_,
    new_n27545_, new_n27546_, new_n27547_, new_n27548_, new_n27549_,
    new_n27550_, new_n27551_, new_n27552_, new_n27553_, new_n27554_,
    new_n27555_, new_n27556_, new_n27557_, new_n27558_, new_n27559_,
    new_n27560_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27599_, new_n27600_, new_n27601_, new_n27602_, new_n27603_,
    new_n27604_, new_n27605_, new_n27606_, new_n27607_, new_n27608_,
    new_n27609_, new_n27610_, new_n27611_, new_n27612_, new_n27613_,
    new_n27614_, new_n27615_, new_n27616_, new_n27617_, new_n27618_,
    new_n27619_, new_n27620_, new_n27621_, new_n27622_, new_n27623_,
    new_n27624_, new_n27625_, new_n27626_, new_n27627_, new_n27628_,
    new_n27629_, new_n27632_, new_n27633_, new_n27634_, new_n27635_,
    new_n27636_, new_n27637_, new_n27638_, new_n27639_, new_n27640_,
    new_n27641_, new_n27642_, new_n27643_, new_n27644_, new_n27645_,
    new_n27646_, new_n27647_, new_n27648_, new_n27649_, new_n27650_,
    new_n27651_, new_n27652_, new_n27653_, new_n27654_, new_n27655_,
    new_n27656_, new_n27657_, new_n27658_, new_n27659_, new_n27660_,
    new_n27661_, new_n27662_, new_n27663_, new_n27664_, new_n27665_,
    new_n27666_, new_n27667_, new_n27668_, new_n27669_, new_n27670_,
    new_n27672_, new_n27673_, new_n27674_, new_n27675_, new_n27677_,
    new_n27678_, new_n27679_, new_n27680_, new_n27681_, new_n27683_,
    new_n27684_, new_n27686_, new_n27687_, new_n27688_, new_n27689_,
    new_n27690_, new_n27691_, new_n27692_, new_n27693_, new_n27694_,
    new_n27695_, new_n27696_, new_n27697_, new_n27698_, new_n27699_,
    new_n27700_, new_n27701_, new_n27702_, new_n27703_, new_n27704_,
    new_n27705_, new_n27706_, new_n27707_, new_n27708_, new_n27709_,
    new_n27710_, new_n27711_, new_n27712_, new_n27713_, new_n27714_,
    new_n27715_, new_n27716_, new_n27717_, new_n27718_, new_n27719_,
    new_n27720_, new_n27721_, new_n27722_, new_n27723_, new_n27724_,
    new_n27725_, new_n27726_, new_n27727_, new_n27728_, new_n27729_,
    new_n27730_, new_n27731_, new_n27732_, new_n27733_, new_n27734_,
    new_n27735_, new_n27736_, new_n27737_, new_n27738_, new_n27739_,
    new_n27740_, new_n27741_, new_n27742_, new_n27743_, new_n27744_,
    new_n27745_, new_n27746_, new_n27747_, new_n27748_, new_n27749_,
    new_n27750_, new_n27751_, new_n27752_, new_n27753_, new_n27754_,
    new_n27755_, new_n27756_, new_n27757_, new_n27758_, new_n27759_,
    new_n27760_, new_n27761_, new_n27763_, new_n27764_, new_n27766_,
    new_n27767_, new_n27769_, new_n27770_, new_n27771_, new_n27772_,
    new_n27773_, new_n27774_, new_n27775_, new_n27776_, new_n27777_,
    new_n27778_, new_n27779_, new_n27780_, new_n27781_, new_n27782_,
    new_n27783_, new_n27784_, new_n27785_, new_n27786_, new_n27787_,
    new_n27788_, new_n27789_, new_n27790_, new_n27791_, new_n27792_,
    new_n27793_, new_n27794_, new_n27795_, new_n27796_, new_n27797_,
    new_n27798_, new_n27799_, new_n27800_, new_n27801_, new_n27802_,
    new_n27803_, new_n27804_, new_n27805_, new_n27806_, new_n27807_,
    new_n27808_, new_n27809_, new_n27810_, new_n27811_, new_n27812_,
    new_n27813_, new_n27814_, new_n27815_, new_n27816_, new_n27817_,
    new_n27818_, new_n27819_, new_n27820_, new_n27821_, new_n27822_,
    new_n27823_, new_n27824_, new_n27825_, new_n27826_, new_n27827_,
    new_n27828_, new_n27829_, new_n27830_, new_n27831_, new_n27832_,
    new_n27833_, new_n27834_, new_n27835_, new_n27836_, new_n27837_,
    new_n27838_, new_n27839_, new_n27840_, new_n27841_, new_n27842_,
    new_n27843_, new_n27844_, new_n27845_, new_n27846_, new_n27847_,
    new_n27848_, new_n27849_, new_n27850_, new_n27851_, new_n27852_,
    new_n27853_, new_n27854_, new_n27855_, new_n27856_, new_n27857_,
    new_n27858_, new_n27859_, new_n27860_, new_n27861_, new_n27862_,
    new_n27863_, new_n27864_, new_n27865_, new_n27866_, new_n27867_,
    new_n27868_, new_n27869_, new_n27870_, new_n27871_, new_n27872_,
    new_n27873_, new_n27874_, new_n27875_, new_n27876_, new_n27877_,
    new_n27878_, new_n27879_, new_n27880_, new_n27883_, new_n27884_,
    new_n27885_, new_n27886_, new_n27887_, new_n27888_, new_n27889_,
    new_n27890_, new_n27891_, new_n27892_, new_n27893_, new_n27894_,
    new_n27895_, new_n27896_, new_n27897_, new_n27898_, new_n27899_,
    new_n27900_, new_n27901_, new_n27902_, new_n27903_, new_n27904_,
    new_n27905_, new_n27906_, new_n27907_, new_n27908_, new_n27909_,
    new_n27910_, new_n27913_, new_n27914_, new_n27915_, new_n27916_,
    new_n27917_, new_n27918_, new_n27919_, new_n27920_, new_n27921_,
    new_n27922_, new_n27923_, new_n27924_, new_n27925_, new_n27926_,
    new_n27927_, new_n27928_, new_n27929_, new_n27930_, new_n27931_,
    new_n27932_, new_n27933_, new_n27934_, new_n27935_, new_n27936_,
    new_n27937_, new_n27938_, new_n27939_, new_n27940_, new_n27941_,
    new_n27942_, new_n27943_, new_n27944_, new_n27945_, new_n27946_,
    new_n27947_, new_n27948_, new_n27949_, new_n27950_, new_n27951_,
    new_n27952_, new_n27953_, new_n27954_, new_n27955_, new_n27956_,
    new_n27957_, new_n27958_, new_n27959_, new_n27960_, new_n27961_,
    new_n27962_, new_n27963_, new_n27964_, new_n27965_, new_n27966_,
    new_n27967_, new_n27968_, new_n27969_, new_n27970_, new_n27971_,
    new_n27972_, new_n27973_, new_n27974_, new_n27975_, new_n27976_,
    new_n27977_, new_n27978_, new_n27979_, new_n27980_, new_n27981_,
    new_n27982_, new_n27983_, new_n27984_, new_n27985_, new_n27986_,
    new_n27987_, new_n27988_, new_n27989_, new_n27990_, new_n27991_,
    new_n27992_, new_n27993_, new_n27994_, new_n27995_, new_n27996_,
    new_n27997_, new_n27998_, new_n27999_, new_n28000_, new_n28001_,
    new_n28002_, new_n28003_, new_n28004_, new_n28005_, new_n28006_,
    new_n28007_, new_n28008_, new_n28009_, new_n28010_, new_n28011_,
    new_n28012_, new_n28013_, new_n28014_, new_n28015_, new_n28016_,
    new_n28017_, new_n28018_, new_n28019_, new_n28020_, new_n28021_,
    new_n28022_, new_n28023_, new_n28024_, new_n28025_, new_n28026_,
    new_n28027_, new_n28028_, new_n28029_, new_n28030_, new_n28031_,
    new_n28032_, new_n28033_, new_n28034_, new_n28035_, new_n28036_,
    new_n28037_, new_n28038_, new_n28039_, new_n28040_, new_n28041_,
    new_n28042_, new_n28043_, new_n28044_, new_n28045_, new_n28046_,
    new_n28047_, new_n28048_, new_n28049_, new_n28050_, new_n28051_,
    new_n28052_, new_n28053_, new_n28054_, new_n28055_, new_n28056_,
    new_n28057_, new_n28058_, new_n28059_, new_n28060_, new_n28061_,
    new_n28062_, new_n28063_, new_n28064_, new_n28065_, new_n28066_,
    new_n28067_, new_n28068_, new_n28069_, new_n28070_, new_n28071_,
    new_n28072_, new_n28073_, new_n28074_, new_n28075_, new_n28076_,
    new_n28077_, new_n28078_, new_n28079_, new_n28080_, new_n28081_,
    new_n28082_, new_n28083_, new_n28084_, new_n28085_, new_n28086_,
    new_n28088_, new_n28089_, new_n28091_, new_n28092_, new_n28093_,
    new_n28094_, new_n28095_, new_n28096_, new_n28097_, new_n28098_,
    new_n28099_, new_n28100_, new_n28101_, new_n28102_, new_n28103_,
    new_n28104_, new_n28105_, new_n28106_, new_n28107_, new_n28108_,
    new_n28109_, new_n28110_, new_n28111_, new_n28112_, new_n28113_,
    new_n28114_, new_n28115_, new_n28116_, new_n28117_, new_n28118_,
    new_n28119_, new_n28120_, new_n28121_, new_n28122_, new_n28123_,
    new_n28124_, new_n28125_, new_n28126_, new_n28127_, new_n28128_,
    new_n28129_, new_n28130_, new_n28131_, new_n28132_, new_n28133_,
    new_n28134_, new_n28135_, new_n28136_, new_n28137_, new_n28138_,
    new_n28139_, new_n28140_, new_n28141_, new_n28142_, new_n28143_,
    new_n28144_, new_n28145_, new_n28146_, new_n28147_, new_n28148_,
    new_n28149_, new_n28150_, new_n28151_, new_n28152_, new_n28153_,
    new_n28154_, new_n28155_, new_n28156_, new_n28157_, new_n28158_,
    new_n28159_, new_n28160_, new_n28161_, new_n28162_, new_n28163_,
    new_n28164_, new_n28165_, new_n28166_, new_n28167_, new_n28168_,
    new_n28169_, new_n28170_, new_n28171_, new_n28172_, new_n28173_,
    new_n28174_, new_n28175_, new_n28176_, new_n28177_, new_n28178_,
    new_n28179_, new_n28180_, new_n28181_, new_n28182_, new_n28183_,
    new_n28184_, new_n28185_, new_n28186_, new_n28187_, new_n28188_,
    new_n28189_, new_n28190_, new_n28191_, new_n28192_, new_n28193_,
    new_n28194_, new_n28195_, new_n28196_, new_n28197_, new_n28198_,
    new_n28199_, new_n28200_, new_n28201_, new_n28202_, new_n28203_,
    new_n28204_, new_n28205_, new_n28206_, new_n28207_, new_n28208_,
    new_n28209_, new_n28210_, new_n28211_, new_n28212_, new_n28213_,
    new_n28214_, new_n28215_, new_n28216_, new_n28217_, new_n28218_,
    new_n28219_, new_n28220_, new_n28221_, new_n28222_, new_n28223_,
    new_n28224_, new_n28225_, new_n28226_, new_n28227_, new_n28229_,
    new_n28230_, new_n28232_, new_n28233_, new_n28234_, new_n28235_,
    new_n28236_, new_n28237_, new_n28238_, new_n28239_, new_n28240_,
    new_n28241_, new_n28242_, new_n28243_, new_n28244_, new_n28245_,
    new_n28246_, new_n28247_, new_n28248_, new_n28249_, new_n28250_,
    new_n28251_, new_n28252_, new_n28253_, new_n28254_, new_n28255_,
    new_n28256_, new_n28257_, new_n28258_, new_n28259_, new_n28260_,
    new_n28261_, new_n28262_, new_n28263_, new_n28264_, new_n28265_,
    new_n28266_, new_n28267_, new_n28268_, new_n28269_, new_n28270_,
    new_n28271_, new_n28272_, new_n28273_, new_n28274_, new_n28275_,
    new_n28276_, new_n28277_, new_n28278_, new_n28279_, new_n28280_,
    new_n28281_, new_n28282_, new_n28283_, new_n28284_, new_n28285_,
    new_n28286_, new_n28287_, new_n28288_, new_n28289_, new_n28290_,
    new_n28292_, new_n28293_, new_n28295_, new_n28296_, new_n28297_,
    new_n28298_, new_n28299_, new_n28300_, new_n28301_, new_n28302_,
    new_n28303_, new_n28304_, new_n28305_, new_n28306_, new_n28307_,
    new_n28308_, new_n28309_, new_n28310_, new_n28311_, new_n28312_,
    new_n28313_, new_n28314_, new_n28315_, new_n28316_, new_n28317_,
    new_n28318_, new_n28319_, new_n28320_, new_n28321_, new_n28322_,
    new_n28323_, new_n28324_, new_n28325_, new_n28326_, new_n28327_,
    new_n28328_, new_n28329_, new_n28330_, new_n28331_, new_n28332_,
    new_n28333_, new_n28334_, new_n28335_, new_n28336_, new_n28337_,
    new_n28338_, new_n28339_, new_n28340_, new_n28341_, new_n28342_,
    new_n28343_, new_n28344_, new_n28345_, new_n28346_, new_n28347_,
    new_n28348_, new_n28349_, new_n28350_, new_n28351_, new_n28352_,
    new_n28353_, new_n28354_, new_n28355_, new_n28356_, new_n28357_,
    new_n28358_, new_n28359_, new_n28360_, new_n28361_, new_n28362_,
    new_n28363_, new_n28364_, new_n28365_, new_n28366_, new_n28367_,
    new_n28368_, new_n28369_, new_n28370_, new_n28371_, new_n28372_,
    new_n28373_, new_n28374_, new_n28375_, new_n28376_, new_n28377_,
    new_n28378_, new_n28379_, new_n28380_, new_n28381_, new_n28382_,
    new_n28383_, new_n28384_, new_n28385_, new_n28386_, new_n28387_,
    new_n28388_, new_n28389_, new_n28390_, new_n28391_, new_n28392_,
    new_n28393_, new_n28394_, new_n28395_, new_n28396_, new_n28398_,
    new_n28399_, new_n28400_, new_n28401_, new_n28402_, new_n28403_,
    new_n28404_, new_n28405_, new_n28406_, new_n28407_, new_n28408_,
    new_n28409_, new_n28410_, new_n28411_, new_n28412_, new_n28413_,
    new_n28414_, new_n28415_, new_n28416_, new_n28417_, new_n28418_,
    new_n28419_, new_n28420_, new_n28422_, new_n28423_, new_n28424_,
    new_n28425_, new_n28426_, new_n28427_, new_n28428_, new_n28429_,
    new_n28430_, new_n28431_, new_n28432_, new_n28433_, new_n28434_,
    new_n28435_, new_n28436_, new_n28437_, new_n28438_, new_n28439_,
    new_n28440_, new_n28441_, new_n28442_, new_n28443_, new_n28444_,
    new_n28445_, new_n28446_, new_n28447_, new_n28448_, new_n28449_,
    new_n28450_, new_n28451_, new_n28452_, new_n28453_, new_n28454_,
    new_n28455_, new_n28456_, new_n28457_, new_n28458_, new_n28459_,
    new_n28460_, new_n28461_, new_n28462_, new_n28463_, new_n28464_,
    new_n28465_, new_n28466_, new_n28467_, new_n28468_, new_n28469_,
    new_n28470_, new_n28471_, new_n28472_, new_n28473_, new_n28474_,
    new_n28475_, new_n28476_, new_n28477_, new_n28478_, new_n28479_,
    new_n28480_, new_n28481_, new_n28482_, new_n28483_, new_n28484_,
    new_n28485_, new_n28486_, new_n28487_, new_n28488_, new_n28489_,
    new_n28490_, new_n28491_, new_n28492_, new_n28493_, new_n28494_,
    new_n28495_, new_n28496_, new_n28497_, new_n28498_, new_n28499_,
    new_n28500_, new_n28501_, new_n28502_, new_n28503_, new_n28504_,
    new_n28505_, new_n28506_, new_n28507_, new_n28508_, new_n28509_,
    new_n28510_, new_n28511_, new_n28512_, new_n28513_, new_n28515_,
    new_n28516_, new_n28517_, new_n28518_, new_n28519_, new_n28520_,
    new_n28521_, new_n28522_, new_n28524_, new_n28525_, new_n28526_,
    new_n28527_, new_n28529_, new_n28530_, new_n28531_, new_n28532_,
    new_n28533_, new_n28535_, new_n28536_, new_n28537_, new_n28538_,
    new_n28540_, new_n28541_, new_n28542_, new_n28543_, new_n28544_,
    new_n28545_, new_n28546_, new_n28547_, new_n28548_, new_n28549_,
    new_n28550_, new_n28551_, new_n28552_, new_n28553_, new_n28554_,
    new_n28555_, new_n28556_, new_n28557_, new_n28558_, new_n28559_,
    new_n28560_, new_n28561_, new_n28562_, new_n28563_, new_n28564_,
    new_n28565_, new_n28566_, new_n28567_, new_n28568_, new_n28569_,
    new_n28570_, new_n28571_, new_n28572_, new_n28573_, new_n28574_,
    new_n28575_, new_n28576_, new_n28577_, new_n28578_, new_n28579_,
    new_n28580_, new_n28581_, new_n28582_, new_n28583_, new_n28584_,
    new_n28585_, new_n28586_, new_n28587_, new_n28588_, new_n28589_,
    new_n28590_, new_n28591_, new_n28592_, new_n28593_, new_n28594_,
    new_n28595_, new_n28596_, new_n28597_, new_n28598_, new_n28599_,
    new_n28600_, new_n28601_, new_n28602_, new_n28603_, new_n28604_,
    new_n28605_, new_n28606_, new_n28607_, new_n28609_, new_n28610_,
    new_n28611_, new_n28612_, new_n28613_, new_n28614_, new_n28615_,
    new_n28616_, new_n28617_, new_n28618_, new_n28619_, new_n28620_,
    new_n28621_, new_n28622_, new_n28623_, new_n28624_, new_n28625_,
    new_n28626_, new_n28627_, new_n28628_, new_n28629_, new_n28630_,
    new_n28631_, new_n28632_, new_n28633_, new_n28634_, new_n28635_,
    new_n28636_, new_n28637_, new_n28638_, new_n28639_, new_n28640_,
    new_n28641_, new_n28642_, new_n28643_, new_n28644_, new_n28645_,
    new_n28646_, new_n28647_, new_n28648_, new_n28649_, new_n28650_,
    new_n28651_, new_n28652_, new_n28653_, new_n28654_, new_n28655_,
    new_n28656_, new_n28657_, new_n28658_, new_n28659_, new_n28660_,
    new_n28661_, new_n28662_, new_n28663_, new_n28664_, new_n28665_,
    new_n28666_, new_n28667_, new_n28668_, new_n28669_, new_n28670_,
    new_n28671_, new_n28672_, new_n28673_, new_n28674_, new_n28675_,
    new_n28676_, new_n28677_, new_n28678_, new_n28679_, new_n28680_,
    new_n28682_, new_n28683_, new_n28684_, new_n28685_, new_n28686_,
    new_n28687_, new_n28688_, new_n28689_, new_n28690_, new_n28691_,
    new_n28692_, new_n28693_, new_n28694_, new_n28695_, new_n28696_,
    new_n28698_, new_n28699_, new_n28701_, new_n28702_, new_n28703_,
    new_n28704_, new_n28706_, new_n28708_, new_n28709_, new_n28710_,
    new_n28711_, new_n28712_, new_n28713_, new_n28714_, new_n28715_,
    new_n28716_, new_n28717_, new_n28718_, new_n28719_, new_n28720_,
    new_n28721_, new_n28722_, new_n28723_, new_n28724_, new_n28725_,
    new_n28726_, new_n28727_, new_n28728_, new_n28729_, new_n28730_,
    new_n28731_, new_n28732_, new_n28733_, new_n28734_, new_n28735_,
    new_n28736_, new_n28737_, new_n28738_, new_n28739_, new_n28740_,
    new_n28741_, new_n28742_, new_n28743_, new_n28744_, new_n28745_,
    new_n28746_, new_n28747_, new_n28748_, new_n28749_, new_n28750_,
    new_n28751_, new_n28752_, new_n28753_, new_n28754_, new_n28755_,
    new_n28756_, new_n28757_, new_n28758_, new_n28759_, new_n28760_,
    new_n28761_, new_n28762_, new_n28763_, new_n28764_, new_n28765_,
    new_n28766_, new_n28767_, new_n28768_, new_n28769_, new_n28770_,
    new_n28771_, new_n28772_, new_n28773_, new_n28774_, new_n28775_,
    new_n28776_, new_n28777_, new_n28778_, new_n28779_, new_n28780_,
    new_n28782_, new_n28783_, new_n28784_, new_n28785_, new_n28786_,
    new_n28787_, new_n28788_, new_n28789_, new_n28790_, new_n28791_,
    new_n28792_, new_n28793_, new_n28794_, new_n28795_, new_n28796_,
    new_n28797_, new_n28798_, new_n28799_, new_n28800_, new_n28801_,
    new_n28802_, new_n28803_, new_n28804_, new_n28805_, new_n28806_,
    new_n28807_, new_n28808_, new_n28809_, new_n28810_, new_n28811_,
    new_n28812_, new_n28813_, new_n28814_, new_n28815_, new_n28816_,
    new_n28818_, new_n28819_, new_n28820_, new_n28821_, new_n28822_,
    new_n28823_, new_n28824_, new_n28825_, new_n28826_, new_n28827_,
    new_n28828_, new_n28829_, new_n28830_, new_n28831_, new_n28832_,
    new_n28833_, new_n28834_, new_n28835_, new_n28836_, new_n28837_,
    new_n28838_, new_n28839_, new_n28840_, new_n28841_, new_n28842_,
    new_n28843_, new_n28844_, new_n28845_, new_n28846_, new_n28847_,
    new_n28848_, new_n28849_, new_n28850_, new_n28851_, new_n28852_,
    new_n28853_, new_n28854_, new_n28855_, new_n28856_, new_n28857_,
    new_n28858_, new_n28859_, new_n28860_, new_n28861_, new_n28862_,
    new_n28863_, new_n28864_, new_n28865_, new_n28866_, new_n28867_,
    new_n28868_, new_n28869_, new_n28870_, new_n28871_, new_n28872_,
    new_n28873_, new_n28874_, new_n28875_, new_n28876_, new_n28877_,
    new_n28878_, new_n28879_, new_n28880_, new_n28881_, new_n28882_,
    new_n28883_, new_n28884_, new_n28885_, new_n28886_, new_n28887_,
    new_n28888_, new_n28889_, new_n28890_, new_n28891_, new_n28892_,
    new_n28893_, new_n28894_, new_n28895_, new_n28896_, new_n28897_,
    new_n28898_, new_n28899_, new_n28900_, new_n28901_, new_n28902_,
    new_n28903_, new_n28904_, new_n28905_, new_n28906_, new_n28907_,
    new_n28908_, new_n28909_, new_n28910_, new_n28911_, new_n28912_,
    new_n28913_, new_n28914_, new_n28915_, new_n28916_, new_n28917_,
    new_n28918_, new_n28919_, new_n28920_, new_n28921_, new_n28922_,
    new_n28923_, new_n28924_, new_n28925_, new_n28926_, new_n28927_,
    new_n28928_, new_n28929_, new_n28930_, new_n28931_, new_n28932_,
    new_n28933_, new_n28934_, new_n28935_, new_n28936_, new_n28937_,
    new_n28938_, new_n28939_, new_n28940_, new_n28941_, new_n28942_,
    new_n28943_, new_n28944_, new_n28945_, new_n28946_, new_n28947_,
    new_n28948_, new_n28949_, new_n28950_, new_n28951_, new_n28952_,
    new_n28953_, new_n28954_, new_n28955_, new_n28956_, new_n28957_,
    new_n28958_, new_n28959_, new_n28960_, new_n28961_, new_n28962_,
    new_n28963_, new_n28964_, new_n28965_, new_n28966_, new_n28967_,
    new_n28968_, new_n28969_, new_n28970_, new_n28971_, new_n28972_,
    new_n28973_, new_n28974_, new_n28975_, new_n28976_, new_n28977_,
    new_n28978_, new_n28979_, new_n28980_, new_n28981_, new_n28982_,
    new_n28983_, new_n28984_, new_n28985_, new_n28986_, new_n28987_,
    new_n28988_, new_n28989_, new_n28990_, new_n28991_, new_n28992_,
    new_n28993_, new_n28994_, new_n28995_, new_n28996_, new_n28997_,
    new_n28998_, new_n28999_, new_n29000_, new_n29001_, new_n29002_,
    new_n29003_, new_n29004_, new_n29005_, new_n29006_, new_n29007_,
    new_n29008_, new_n29009_, new_n29010_, new_n29011_, new_n29012_,
    new_n29013_, new_n29014_, new_n29015_, new_n29016_, new_n29017_,
    new_n29018_, new_n29019_, new_n29020_, new_n29021_, new_n29022_,
    new_n29023_, new_n29024_, new_n29025_, new_n29026_, new_n29027_,
    new_n29028_, new_n29029_, new_n29030_, new_n29031_, new_n29032_,
    new_n29033_, new_n29034_, new_n29035_, new_n29036_, new_n29037_,
    new_n29038_, new_n29039_, new_n29040_, new_n29041_, new_n29042_,
    new_n29043_, new_n29044_, new_n29045_, new_n29046_, new_n29047_,
    new_n29048_, new_n29049_, new_n29050_, new_n29051_, new_n29052_,
    new_n29053_, new_n29054_, new_n29055_, new_n29056_, new_n29057_,
    new_n29058_, new_n29059_, new_n29060_, new_n29061_, new_n29062_,
    new_n29063_, new_n29064_, new_n29065_, new_n29066_, new_n29067_,
    new_n29068_, new_n29069_, new_n29070_, new_n29071_, new_n29072_,
    new_n29073_, new_n29074_, new_n29075_, new_n29076_, new_n29077_,
    new_n29078_, new_n29079_, new_n29080_, new_n29081_, new_n29082_,
    new_n29083_, new_n29084_, new_n29085_, new_n29086_, new_n29087_,
    new_n29088_, new_n29089_, new_n29090_, new_n29091_, new_n29092_,
    new_n29093_, new_n29094_, new_n29095_, new_n29096_, new_n29097_,
    new_n29098_, new_n29099_, new_n29100_, new_n29101_, new_n29102_,
    new_n29103_, new_n29104_, new_n29105_, new_n29106_, new_n29107_,
    new_n29108_, new_n29109_, new_n29110_, new_n29111_, new_n29112_,
    new_n29113_, new_n29114_, new_n29115_, new_n29116_, new_n29117_,
    new_n29118_, new_n29119_, new_n29120_, new_n29121_, new_n29122_,
    new_n29123_, new_n29124_, new_n29125_, new_n29126_, new_n29127_,
    new_n29128_, new_n29129_, new_n29130_, new_n29131_, new_n29132_,
    new_n29133_, new_n29134_, new_n29135_, new_n29136_, new_n29137_,
    new_n29138_, new_n29139_, new_n29140_, new_n29141_, new_n29142_,
    new_n29143_, new_n29144_, new_n29145_, new_n29146_, new_n29147_,
    new_n29148_, new_n29149_, new_n29150_, new_n29151_, new_n29152_,
    new_n29153_, new_n29154_, new_n29155_, new_n29156_, new_n29157_,
    new_n29158_, new_n29159_, new_n29160_, new_n29161_, new_n29162_,
    new_n29163_, new_n29164_, new_n29165_, new_n29166_, new_n29167_,
    new_n29168_, new_n29169_, new_n29170_, new_n29171_, new_n29172_,
    new_n29173_, new_n29174_, new_n29175_, new_n29176_, new_n29177_,
    new_n29178_, new_n29179_, new_n29180_, new_n29181_, new_n29182_,
    new_n29183_, new_n29184_, new_n29185_, new_n29186_, new_n29187_,
    new_n29188_, new_n29189_, new_n29190_, new_n29191_, new_n29192_,
    new_n29193_, new_n29194_, new_n29195_, new_n29196_, new_n29197_,
    new_n29198_, new_n29199_, new_n29200_, new_n29201_, new_n29202_,
    new_n29203_, new_n29204_, new_n29205_, new_n29206_, new_n29207_,
    new_n29208_, new_n29209_, new_n29210_, new_n29211_, new_n29212_,
    new_n29213_, new_n29214_, new_n29215_, new_n29216_, new_n29217_,
    new_n29218_, new_n29219_, new_n29220_, new_n29221_, new_n29222_,
    new_n29223_, new_n29224_, new_n29225_, new_n29226_, new_n29227_,
    new_n29228_, new_n29229_, new_n29230_, new_n29231_, new_n29232_,
    new_n29233_, new_n29234_, new_n29235_, new_n29236_, new_n29237_,
    new_n29238_, new_n29239_, new_n29240_, new_n29241_, new_n29242_,
    new_n29243_, new_n29244_, new_n29245_, new_n29246_, new_n29247_,
    new_n29248_, new_n29249_, new_n29250_, new_n29251_, new_n29252_,
    new_n29253_, new_n29254_, new_n29255_, new_n29256_, new_n29257_,
    new_n29258_, new_n29259_, new_n29260_, new_n29261_, new_n29262_,
    new_n29263_, new_n29264_, new_n29265_, new_n29266_, new_n29267_,
    new_n29268_, new_n29269_, new_n29270_, new_n29271_, new_n29272_,
    new_n29273_, new_n29274_, new_n29275_, new_n29276_, new_n29277_,
    new_n29278_, new_n29279_, new_n29280_, new_n29281_, new_n29282_,
    new_n29283_, new_n29284_, new_n29285_, new_n29286_, new_n29287_,
    new_n29288_, new_n29289_, new_n29290_, new_n29291_, new_n29292_,
    new_n29293_, new_n29294_, new_n29295_, new_n29296_, new_n29297_,
    new_n29298_, new_n29299_, new_n29300_, new_n29301_, new_n29302_,
    new_n29303_, new_n29304_, new_n29305_, new_n29306_, new_n29307_,
    new_n29308_, new_n29309_, new_n29310_, new_n29311_, new_n29312_,
    new_n29313_, new_n29314_, new_n29315_, new_n29316_, new_n29317_,
    new_n29318_, new_n29319_, new_n29321_, new_n29322_, new_n29323_,
    new_n29324_, new_n29325_, new_n29327_, new_n29328_, new_n29329_,
    new_n29330_, new_n29331_, new_n29332_, new_n29333_, new_n29334_,
    new_n29335_, new_n29336_, new_n29337_, new_n29338_, new_n29339_,
    new_n29340_, new_n29342_, new_n29343_, new_n29344_, new_n29345_,
    new_n29346_, new_n29347_, new_n29348_, new_n29349_, new_n29350_,
    new_n29351_, new_n29352_, new_n29353_, new_n29354_, new_n29355_,
    new_n29356_, new_n29357_, new_n29358_, new_n29359_, new_n29360_,
    new_n29361_, new_n29362_, new_n29363_, new_n29364_, new_n29365_,
    new_n29366_, new_n29367_, new_n29368_, new_n29369_, new_n29370_,
    new_n29371_, new_n29372_, new_n29373_, new_n29374_, new_n29375_,
    new_n29376_, new_n29377_, new_n29378_, new_n29379_, new_n29380_,
    new_n29381_, new_n29382_, new_n29383_, new_n29384_, new_n29385_,
    new_n29386_, new_n29387_, new_n29388_, new_n29389_, new_n29390_,
    new_n29391_, new_n29392_, new_n29393_, new_n29394_, new_n29395_,
    new_n29396_, new_n29397_, new_n29398_, new_n29399_, new_n29400_,
    new_n29401_, new_n29402_, new_n29403_, new_n29404_, new_n29405_,
    new_n29406_, new_n29407_, new_n29408_, new_n29409_, new_n29410_,
    new_n29411_, new_n29412_, new_n29413_, new_n29414_, new_n29415_,
    new_n29416_, new_n29417_, new_n29418_, new_n29419_, new_n29420_,
    new_n29421_, new_n29422_, new_n29423_, new_n29424_, new_n29425_,
    new_n29426_, new_n29427_, new_n29428_, new_n29430_, new_n29431_,
    new_n29432_, new_n29433_, new_n29434_, new_n29435_, new_n29436_,
    new_n29437_, new_n29438_, new_n29439_, new_n29440_, new_n29441_,
    new_n29442_, new_n29443_, new_n29444_, new_n29445_, new_n29446_,
    new_n29447_, new_n29448_, new_n29449_, new_n29450_, new_n29451_,
    new_n29452_, new_n29453_, new_n29454_, new_n29455_, new_n29456_,
    new_n29457_, new_n29458_, new_n29459_, new_n29460_, new_n29461_,
    new_n29462_, new_n29463_, new_n29464_, new_n29465_, new_n29466_,
    new_n29467_, new_n29468_, new_n29469_, new_n29470_, new_n29471_,
    new_n29472_, new_n29473_, new_n29474_, new_n29475_, new_n29476_,
    new_n29477_, new_n29478_, new_n29479_, new_n29480_, new_n29481_,
    new_n29482_, new_n29483_, new_n29484_, new_n29485_, new_n29486_,
    new_n29487_, new_n29488_, new_n29489_, new_n29490_, new_n29491_,
    new_n29492_, new_n29493_, new_n29494_, new_n29495_, new_n29496_,
    new_n29497_, new_n29498_, new_n29499_, new_n29500_, new_n29501_,
    new_n29502_, new_n29503_, new_n29504_, new_n29505_, new_n29506_,
    new_n29507_, new_n29508_, new_n29509_, new_n29510_, new_n29511_,
    new_n29512_, new_n29513_, new_n29514_, new_n29515_, new_n29516_,
    new_n29517_, new_n29518_, new_n29519_, new_n29520_, new_n29521_,
    new_n29522_, new_n29523_, new_n29524_, new_n29525_, new_n29526_,
    new_n29527_, new_n29528_, new_n29529_, new_n29530_, new_n29531_,
    new_n29532_, new_n29533_, new_n29534_, new_n29535_, new_n29536_,
    new_n29537_, new_n29538_, new_n29539_, new_n29540_, new_n29541_,
    new_n29542_, new_n29543_, new_n29544_, new_n29545_, new_n29546_,
    new_n29547_, new_n29548_, new_n29549_, new_n29550_, new_n29551_,
    new_n29552_, new_n29553_, new_n29554_, new_n29555_, new_n29556_,
    new_n29557_, new_n29558_, new_n29559_, new_n29560_, new_n29561_,
    new_n29562_, new_n29563_, new_n29564_, new_n29565_, new_n29566_,
    new_n29567_, new_n29568_, new_n29569_, new_n29570_, new_n29571_,
    new_n29572_, new_n29573_, new_n29574_, new_n29575_, new_n29576_,
    new_n29577_, new_n29578_, new_n29579_, new_n29580_, new_n29581_,
    new_n29582_, new_n29583_, new_n29584_, new_n29585_, new_n29589_,
    new_n29593_, new_n29594_, new_n29595_, new_n29596_, new_n29597_,
    new_n29598_, new_n29599_, new_n29600_, new_n29601_, new_n29602_,
    new_n29603_, new_n29604_, new_n29605_, new_n29606_, new_n29607_,
    new_n29608_, new_n29609_, new_n29610_, new_n29611_, new_n29612_,
    new_n29613_, new_n29614_, new_n29615_, new_n29616_, new_n29617_,
    new_n29618_, new_n29619_, new_n29620_, new_n29621_, new_n29622_,
    new_n29623_, new_n29624_, new_n29625_, new_n29626_, new_n29627_,
    new_n29628_, new_n29629_, new_n29630_, new_n29631_, new_n29632_,
    new_n29633_, new_n29634_, new_n29635_, new_n29636_, new_n29637_,
    new_n29638_, new_n29639_, new_n29640_, new_n29641_, new_n29642_,
    new_n29643_, new_n29644_, new_n29645_, new_n29646_, new_n29647_,
    new_n29648_, new_n29650_, new_n29651_, new_n29652_, new_n29653_,
    new_n29654_, new_n29655_, new_n29656_, new_n29657_, new_n29658_,
    new_n29659_, new_n29660_, new_n29661_, new_n29662_, new_n29663_,
    new_n29664_, new_n29665_, new_n29666_, new_n29667_, new_n29668_,
    new_n29669_, new_n29670_, new_n29671_, new_n29672_, new_n29673_,
    new_n29674_, new_n29675_, new_n29676_, new_n29677_, new_n29678_,
    new_n29679_, new_n29680_, new_n29681_, new_n29682_, new_n29683_,
    new_n29684_, new_n29685_, new_n29686_, new_n29687_, new_n29688_,
    new_n29689_, new_n29690_, new_n29691_, new_n29692_, new_n29693_,
    new_n29694_, new_n29695_, new_n29696_, new_n29697_, new_n29698_,
    new_n29699_, new_n29700_, new_n29701_, new_n29702_, new_n29703_,
    new_n29704_, new_n29705_, new_n29706_, new_n29707_, new_n29708_,
    new_n29709_, new_n29710_, new_n29711_, new_n29712_, new_n29713_,
    new_n29714_, new_n29715_, new_n29716_, new_n29717_, new_n29718_,
    new_n29719_, new_n29720_, new_n29721_, new_n29722_, new_n29723_,
    new_n29724_, new_n29725_, new_n29726_, new_n29727_, new_n29728_,
    new_n29729_, new_n29730_, new_n29731_, new_n29732_, new_n29733_,
    new_n29734_, new_n29735_, new_n29736_, new_n29737_, new_n29738_,
    new_n29739_, new_n29740_, new_n29741_, new_n29742_, new_n29743_,
    new_n29744_, new_n29745_, new_n29746_, new_n29747_, new_n29748_,
    new_n29749_, new_n29750_, new_n29751_, new_n29752_, new_n29753_,
    new_n29754_, new_n29755_, new_n29756_, new_n29757_, new_n29758_,
    new_n29759_, new_n29760_, new_n29761_, new_n29762_, new_n29763_,
    new_n29764_, new_n29765_, new_n29766_, new_n29767_, new_n29768_,
    new_n29769_, new_n29770_, new_n29771_, new_n29772_, new_n29773_,
    new_n29774_, new_n29775_, new_n29776_, new_n29777_, new_n29778_,
    new_n29779_, new_n29780_, new_n29781_, new_n29782_, new_n29783_,
    new_n29784_, new_n29785_, new_n29786_, new_n29787_, new_n29788_,
    new_n29790_, new_n29791_, new_n29792_, new_n29793_, new_n29794_,
    new_n29795_, new_n29797_, new_n29798_, new_n29799_, new_n29800_,
    new_n29801_, new_n29802_, new_n29803_, new_n29804_, new_n29805_,
    new_n29806_, new_n29807_, new_n29808_, new_n29810_, new_n29811_,
    new_n29812_, new_n29813_, new_n29814_, new_n29815_, new_n29816_,
    new_n29817_, new_n29818_, new_n29819_, new_n29820_, new_n29821_,
    new_n29822_, new_n29823_, new_n29824_, new_n29825_, new_n29826_,
    new_n29827_, new_n29828_, new_n29829_, new_n29830_, new_n29831_,
    new_n29832_, new_n29833_, new_n29834_, new_n29835_, new_n29836_,
    new_n29837_, new_n29838_, new_n29839_, new_n29840_, new_n29841_,
    new_n29842_, new_n29843_, new_n29844_, new_n29845_, new_n29846_,
    new_n29847_, new_n29848_, new_n29849_, new_n29850_, new_n29851_,
    new_n29852_, new_n29853_, new_n29854_, new_n29855_, new_n29856_,
    new_n29857_, new_n29858_, new_n29859_, new_n29860_, new_n29861_,
    new_n29862_, new_n29863_, new_n29864_, new_n29865_, new_n29866_,
    new_n29867_, new_n29868_, new_n29869_, new_n29870_, new_n29871_,
    new_n29872_, new_n29873_, new_n29874_, new_n29875_, new_n29876_,
    new_n29877_, new_n29878_, new_n29879_, new_n29880_, new_n29881_,
    new_n29882_, new_n29883_, new_n29884_, new_n29885_, new_n29886_,
    new_n29887_, new_n29888_, new_n29889_, new_n29890_, new_n29891_,
    new_n29892_, new_n29893_, new_n29894_, new_n29895_, new_n29896_,
    new_n29897_, new_n29898_, new_n29899_, new_n29900_, new_n29901_,
    new_n29902_, new_n29903_, new_n29904_, new_n29905_, new_n29906_,
    new_n29907_, new_n29908_, new_n29909_, new_n29910_, new_n29911_,
    new_n29912_, new_n29913_, new_n29914_, new_n29915_, new_n29916_,
    new_n29917_, new_n29918_, new_n29919_, new_n29920_, new_n29921_,
    new_n29922_, new_n29923_, new_n29924_, new_n29925_, new_n29926_,
    new_n29927_, new_n29928_, new_n29929_, new_n29930_, new_n29931_,
    new_n29932_, new_n29933_, new_n29934_, new_n29935_, new_n29936_,
    new_n29937_, new_n29938_, new_n29939_, new_n29940_, new_n29941_,
    new_n29942_, new_n29943_, new_n29944_, new_n29945_, new_n29946_,
    new_n29947_, new_n29948_, new_n29949_, new_n29950_, new_n29951_,
    new_n29952_, new_n29953_, new_n29954_, new_n29955_, new_n29956_,
    new_n29957_, new_n29958_, new_n29959_, new_n29960_, new_n29961_,
    new_n29962_, new_n29963_, new_n29964_, new_n29965_, new_n29966_,
    new_n29967_, new_n29968_, new_n29969_, new_n29970_, new_n29971_,
    new_n29972_, new_n29973_, new_n29974_, new_n29975_, new_n29976_,
    new_n29977_, new_n29978_, new_n29979_, new_n29980_, new_n29981_,
    new_n29982_, new_n29983_, new_n29984_, new_n29985_, new_n29986_,
    new_n29987_, new_n29988_, new_n29989_, new_n29990_, new_n29991_,
    new_n29992_, new_n29993_, new_n29994_, new_n29995_, new_n29996_,
    new_n29997_, new_n29998_, new_n29999_, new_n30000_, new_n30001_,
    new_n30002_, new_n30003_, new_n30004_, new_n30005_, new_n30006_,
    new_n30007_, new_n30008_, new_n30009_, new_n30010_, new_n30011_,
    new_n30012_, new_n30013_, new_n30014_, new_n30015_, new_n30016_,
    new_n30017_, new_n30018_, new_n30019_, new_n30020_, new_n30021_,
    new_n30022_, new_n30023_, new_n30024_, new_n30025_, new_n30026_,
    new_n30027_, new_n30028_, new_n30029_, new_n30030_, new_n30031_,
    new_n30032_, new_n30033_, new_n30034_, new_n30035_, new_n30036_,
    new_n30037_, new_n30038_, new_n30039_, new_n30040_, new_n30041_,
    new_n30042_, new_n30043_, new_n30044_, new_n30045_, new_n30046_,
    new_n30047_, new_n30048_, new_n30049_, new_n30050_, new_n30051_,
    new_n30052_, new_n30053_, new_n30054_, new_n30055_, new_n30056_,
    new_n30057_, new_n30058_, new_n30059_, new_n30060_, new_n30061_,
    new_n30062_, new_n30063_, new_n30064_, new_n30065_, new_n30066_,
    new_n30067_, new_n30068_, new_n30069_, new_n30070_, new_n30071_,
    new_n30072_, new_n30073_, new_n30074_, new_n30075_, new_n30076_,
    new_n30077_, new_n30078_, new_n30079_, new_n30080_, new_n30081_,
    new_n30082_, new_n30083_, new_n30084_, new_n30085_, new_n30086_,
    new_n30087_, new_n30088_, new_n30089_, new_n30090_, new_n30091_,
    new_n30092_, new_n30093_, new_n30094_, new_n30095_, new_n30096_,
    new_n30097_, new_n30098_, new_n30099_, new_n30100_, new_n30101_,
    new_n30102_, new_n30103_, new_n30104_, new_n30105_, new_n30106_,
    new_n30107_, new_n30108_, new_n30109_, new_n30110_, new_n30111_,
    new_n30112_, new_n30113_, new_n30114_, new_n30115_, new_n30116_,
    new_n30117_, new_n30118_, new_n30119_, new_n30120_, new_n30121_,
    new_n30122_, new_n30123_, new_n30124_, new_n30125_, new_n30126_,
    new_n30127_, new_n30128_, new_n30129_, new_n30130_, new_n30131_,
    new_n30132_, new_n30133_, new_n30134_, new_n30135_, new_n30136_,
    new_n30137_, new_n30138_, new_n30139_, new_n30140_, new_n30141_,
    new_n30142_, new_n30143_, new_n30144_, new_n30145_, new_n30146_,
    new_n30147_, new_n30148_, new_n30149_, new_n30150_, new_n30151_,
    new_n30152_, new_n30153_, new_n30154_, new_n30155_, new_n30156_,
    new_n30157_, new_n30158_, new_n30159_, new_n30160_, new_n30161_,
    new_n30162_, new_n30163_, new_n30164_, new_n30165_, new_n30166_,
    new_n30167_, new_n30168_, new_n30169_, new_n30170_, new_n30171_,
    new_n30172_, new_n30173_, new_n30174_, new_n30175_, new_n30176_,
    new_n30177_, new_n30178_, new_n30179_, new_n30180_, new_n30181_,
    new_n30182_, new_n30183_, new_n30184_, new_n30185_, new_n30186_,
    new_n30187_, new_n30188_, new_n30189_, new_n30190_, new_n30191_,
    new_n30192_, new_n30193_, new_n30194_, new_n30195_, new_n30196_,
    new_n30197_, new_n30198_, new_n30199_, new_n30200_, new_n30201_,
    new_n30202_, new_n30203_, new_n30204_, new_n30205_, new_n30206_,
    new_n30207_, new_n30208_, new_n30209_, new_n30210_, new_n30211_,
    new_n30212_, new_n30213_, new_n30214_, new_n30215_, new_n30216_,
    new_n30217_, new_n30218_, new_n30219_, new_n30220_, new_n30221_,
    new_n30222_, new_n30223_, new_n30224_, new_n30225_, new_n30226_,
    new_n30227_, new_n30228_, new_n30229_, new_n30230_, new_n30231_,
    new_n30232_, new_n30233_, new_n30234_, new_n30235_, new_n30236_,
    new_n30237_, new_n30238_, new_n30239_, new_n30240_, new_n30241_,
    new_n30242_, new_n30243_, new_n30244_, new_n30245_, new_n30246_,
    new_n30247_, new_n30248_, new_n30249_, new_n30250_, new_n30251_,
    new_n30252_, new_n30253_, new_n30254_, new_n30255_, new_n30256_,
    new_n30257_, new_n30258_, new_n30259_, new_n30260_, new_n30261_,
    new_n30262_, new_n30263_, new_n30264_, new_n30265_, new_n30266_,
    new_n30267_, new_n30268_, new_n30269_, new_n30270_, new_n30271_,
    new_n30272_, new_n30273_, new_n30274_, new_n30275_, new_n30276_,
    new_n30277_, new_n30278_, new_n30279_, new_n30280_, new_n30281_,
    new_n30282_, new_n30283_, new_n30284_, new_n30285_, new_n30286_,
    new_n30287_, new_n30288_, new_n30289_, new_n30290_, new_n30291_,
    new_n30292_, new_n30293_, new_n30294_, new_n30295_, new_n30296_,
    new_n30297_, new_n30298_, new_n30299_, new_n30300_, new_n30301_,
    new_n30302_, new_n30303_, new_n30304_, new_n30305_, new_n30306_,
    new_n30307_, new_n30309_, new_n30310_, new_n30311_, new_n30312_,
    new_n30313_, new_n30314_, new_n30315_, new_n30316_, new_n30317_,
    new_n30318_, new_n30319_, new_n30320_, new_n30321_, new_n30322_,
    new_n30323_, new_n30324_, new_n30325_, new_n30326_, new_n30327_,
    new_n30328_, new_n30329_, new_n30330_, new_n30331_, new_n30332_,
    new_n30333_, new_n30334_, new_n30335_, new_n30336_, new_n30337_,
    new_n30338_, new_n30339_, new_n30340_, new_n30341_, new_n30342_,
    new_n30343_, new_n30344_, new_n30345_, new_n30346_, new_n30347_,
    new_n30348_, new_n30349_, new_n30350_, new_n30351_, new_n30352_,
    new_n30353_, new_n30354_, new_n30355_, new_n30356_, new_n30357_,
    new_n30358_, new_n30359_, new_n30360_, new_n30361_, new_n30362_,
    new_n30363_, new_n30364_, new_n30365_, new_n30366_, new_n30367_,
    new_n30368_, new_n30369_, new_n30370_, new_n30371_, new_n30372_,
    new_n30373_, new_n30374_, new_n30375_, new_n30376_, new_n30377_,
    new_n30378_, new_n30379_, new_n30380_, new_n30381_, new_n30383_,
    new_n30384_, new_n30386_, new_n30387_, new_n30388_, new_n30389_,
    new_n30390_, new_n30391_, new_n30392_, new_n30393_, new_n30394_,
    new_n30395_, new_n30396_, new_n30397_, new_n30398_, new_n30399_,
    new_n30400_, new_n30401_, new_n30402_, new_n30403_, new_n30404_,
    new_n30405_, new_n30406_, new_n30407_, new_n30408_, new_n30409_,
    new_n30410_, new_n30411_, new_n30412_, new_n30413_, new_n30414_,
    new_n30415_, new_n30416_, new_n30417_, new_n30418_, new_n30419_,
    new_n30420_, new_n30421_, new_n30422_, new_n30423_, new_n30425_,
    new_n30426_, new_n30427_, new_n30428_, new_n30429_, new_n30430_,
    new_n30431_, new_n30432_, new_n30433_, new_n30434_, new_n30435_,
    new_n30436_, new_n30437_, new_n30438_, new_n30439_, new_n30440_,
    new_n30441_, new_n30442_, new_n30443_, new_n30444_, new_n30446_,
    new_n30447_, new_n30448_, new_n30449_, new_n30450_, new_n30451_,
    new_n30452_, new_n30453_, new_n30455_, new_n30456_, new_n30457_,
    new_n30458_, new_n30459_, new_n30460_, new_n30461_, new_n30462_,
    new_n30463_, new_n30464_, new_n30465_, new_n30466_, new_n30467_,
    new_n30468_, new_n30469_, new_n30470_, new_n30471_, new_n30472_,
    new_n30473_, new_n30474_, new_n30475_, new_n30476_, new_n30477_,
    new_n30478_, new_n30479_, new_n30480_, new_n30481_, new_n30482_,
    new_n30483_, new_n30484_, new_n30485_, new_n30486_, new_n30487_,
    new_n30488_, new_n30489_, new_n30490_, new_n30491_, new_n30492_,
    new_n30493_, new_n30494_, new_n30495_, new_n30496_, new_n30497_,
    new_n30498_, new_n30499_, new_n30500_, new_n30501_, new_n30502_,
    new_n30503_, new_n30504_, new_n30505_, new_n30506_, new_n30507_,
    new_n30508_, new_n30509_, new_n30510_, new_n30511_, new_n30512_,
    new_n30514_, new_n30515_, new_n30516_, new_n30517_, new_n30518_,
    new_n30519_, new_n30520_, new_n30521_, new_n30522_, new_n30523_,
    new_n30524_, new_n30525_, new_n30526_, new_n30527_, new_n30528_,
    new_n30529_, new_n30530_, new_n30531_, new_n30532_, new_n30533_,
    new_n30534_, new_n30535_, new_n30536_, new_n30537_, new_n30538_,
    new_n30539_, new_n30540_, new_n30541_, new_n30542_, new_n30543_,
    new_n30544_, new_n30545_, new_n30546_, new_n30547_, new_n30548_,
    new_n30549_, new_n30550_, new_n30551_, new_n30552_, new_n30553_,
    new_n30554_, new_n30555_, new_n30557_, new_n30558_, new_n30559_,
    new_n30560_, new_n30561_, new_n30562_, new_n30563_, new_n30564_,
    new_n30565_, new_n30566_, new_n30567_, new_n30568_, new_n30569_,
    new_n30570_, new_n30571_, new_n30572_, new_n30573_, new_n30574_,
    new_n30575_, new_n30576_, new_n30577_, new_n30578_, new_n30579_,
    new_n30580_, new_n30581_, new_n30582_, new_n30583_, new_n30584_,
    new_n30585_, new_n30586_, new_n30587_, new_n30588_, new_n30589_,
    new_n30590_, new_n30591_, new_n30592_, new_n30593_, new_n30594_,
    new_n30595_, new_n30596_, new_n30597_, new_n30599_, new_n30600_,
    new_n30601_, new_n30602_, new_n30603_, new_n30604_, new_n30605_,
    new_n30606_, new_n30607_, new_n30608_, new_n30609_, new_n30610_,
    new_n30611_, new_n30612_, new_n30613_, new_n30614_, new_n30615_,
    new_n30616_, new_n30617_, new_n30618_, new_n30619_, new_n30620_,
    new_n30621_, new_n30622_, new_n30623_, new_n30624_, new_n30625_,
    new_n30626_, new_n30627_, new_n30628_, new_n30629_, new_n30630_,
    new_n30631_, new_n30632_, new_n30633_, new_n30634_, new_n30635_,
    new_n30636_, new_n30637_, new_n30638_, new_n30639_, new_n30640_,
    new_n30641_, new_n30642_, new_n30643_, new_n30644_, new_n30645_,
    new_n30646_, new_n30647_, new_n30648_, new_n30649_, new_n30650_,
    new_n30651_, new_n30652_, new_n30653_, new_n30654_, new_n30655_,
    new_n30656_, new_n30657_, new_n30658_, new_n30659_, new_n30660_,
    new_n30661_, new_n30662_, new_n30663_, new_n30664_, new_n30665_,
    new_n30666_, new_n30667_, new_n30668_, new_n30669_, new_n30670_,
    new_n30671_, new_n30672_, new_n30673_, new_n30674_, new_n30675_,
    new_n30676_, new_n30677_, new_n30678_, new_n30679_, new_n30680_,
    new_n30681_, new_n30682_, new_n30683_, new_n30684_, new_n30685_,
    new_n30686_, new_n30687_, new_n30688_, new_n30689_, new_n30690_,
    new_n30691_, new_n30692_, new_n30693_, new_n30694_, new_n30695_,
    new_n30696_, new_n30697_, new_n30698_, new_n30699_, new_n30700_,
    new_n30701_, new_n30702_, new_n30703_, new_n30704_, new_n30705_,
    new_n30706_, new_n30707_, new_n30708_, new_n30709_, new_n30710_,
    new_n30711_, new_n30712_, new_n30713_, new_n30714_, new_n30715_,
    new_n30716_, new_n30717_, new_n30718_, new_n30719_, new_n30720_,
    new_n30721_, new_n30722_, new_n30723_, new_n30724_, new_n30725_,
    new_n30726_, new_n30727_, new_n30728_, new_n30729_, new_n30730_,
    new_n30731_, new_n30732_, new_n30733_, new_n30734_, new_n30735_,
    new_n30736_, new_n30737_, new_n30738_, new_n30739_, new_n30740_,
    new_n30741_, new_n30742_, new_n30743_, new_n30744_, new_n30745_,
    new_n30746_, new_n30747_, new_n30748_, new_n30749_, new_n30750_,
    new_n30751_, new_n30752_, new_n30753_, new_n30754_, new_n30755_,
    new_n30756_, new_n30757_, new_n30758_, new_n30759_, new_n30760_,
    new_n30761_, new_n30762_, new_n30763_, new_n30764_, new_n30765_,
    new_n30766_, new_n30767_, new_n30768_, new_n30769_, new_n30770_,
    new_n30771_, new_n30772_, new_n30773_, new_n30774_, new_n30775_,
    new_n30776_, new_n30777_, new_n30778_, new_n30779_, new_n30780_,
    new_n30781_, new_n30782_, new_n30783_, new_n30784_, new_n30785_,
    new_n30786_, new_n30787_, new_n30788_, new_n30789_, new_n30790_,
    new_n30791_, new_n30792_, new_n30793_, new_n30794_, new_n30795_,
    new_n30796_, new_n30797_, new_n30798_, new_n30799_, new_n30800_,
    new_n30801_, new_n30802_, new_n30803_, new_n30804_, new_n30805_,
    new_n30806_, new_n30807_, new_n30808_, new_n30809_, new_n30810_,
    new_n30811_, new_n30812_, new_n30813_, new_n30814_, new_n30815_,
    new_n30816_, new_n30817_, new_n30818_, new_n30819_, new_n30820_,
    new_n30821_, new_n30822_, new_n30823_, new_n30824_, new_n30825_,
    new_n30826_, new_n30827_, new_n30828_, new_n30829_, new_n30830_,
    new_n30831_, new_n30832_, new_n30833_, new_n30834_, new_n30835_,
    new_n30836_, new_n30837_, new_n30838_, new_n30839_, new_n30840_,
    new_n30841_, new_n30842_, new_n30843_, new_n30844_, new_n30845_,
    new_n30846_, new_n30847_, new_n30848_, new_n30849_, new_n30850_,
    new_n30851_, new_n30852_, new_n30853_, new_n30855_, new_n30856_,
    new_n30857_, new_n30858_, new_n30859_, new_n30860_, new_n30861_,
    new_n30862_, new_n30863_, new_n30864_, new_n30865_, new_n30866_,
    new_n30867_, new_n30868_, new_n30869_, new_n30870_, new_n30871_,
    new_n30872_, new_n30873_, new_n30874_, new_n30875_, new_n30876_,
    new_n30877_, new_n30878_, new_n30879_, new_n30880_, new_n30881_,
    new_n30882_, new_n30883_, new_n30884_, new_n30885_, new_n30886_,
    new_n30887_, new_n30888_, new_n30889_, new_n30890_, new_n30891_,
    new_n30892_, new_n30893_, new_n30894_, new_n30895_, new_n30896_,
    new_n30897_, new_n30898_, new_n30899_, new_n30900_, new_n30901_,
    new_n30902_, new_n30903_, new_n30904_, new_n30905_, new_n30906_,
    new_n30907_, new_n30908_, new_n30909_, new_n30910_, new_n30911_,
    new_n30912_, new_n30913_, new_n30915_, new_n30916_, new_n30917_,
    new_n30918_, new_n30919_, new_n30920_, new_n30921_, new_n30922_,
    new_n30923_, new_n30924_, new_n30925_, new_n30926_, new_n30927_,
    new_n30928_, new_n30929_, new_n30930_, new_n30931_, new_n30932_,
    new_n30933_, new_n30934_, new_n30935_, new_n30936_, new_n30937_,
    new_n30938_, new_n30939_, new_n30940_, new_n30941_, new_n30942_,
    new_n30943_, new_n30944_, new_n30945_, new_n30946_, new_n30947_,
    new_n30948_, new_n30949_, new_n30950_, new_n30951_, new_n30952_,
    new_n30953_, new_n30954_, new_n30955_, new_n30956_, new_n30957_,
    new_n30958_, new_n30959_, new_n30960_, new_n30961_, new_n30962_,
    new_n30963_, new_n30964_, new_n30965_, new_n30966_, new_n30967_,
    new_n30968_, new_n30969_, new_n30970_, new_n30971_, new_n30972_,
    new_n30973_, new_n30974_, new_n30975_, new_n30976_, new_n30977_,
    new_n30978_, new_n30979_, new_n30980_, new_n30981_, new_n30982_,
    new_n30983_, new_n30984_, new_n30985_, new_n30986_, new_n30987_,
    new_n30988_, new_n30989_, new_n30990_, new_n30991_, new_n30992_,
    new_n30993_, new_n30994_, new_n30995_, new_n30996_, new_n30997_,
    new_n30998_, new_n30999_, new_n31000_, new_n31001_, new_n31002_,
    new_n31003_, new_n31004_, new_n31005_, new_n31006_, new_n31007_,
    new_n31008_, new_n31009_, new_n31010_, new_n31011_, new_n31012_,
    new_n31013_, new_n31014_, new_n31015_, new_n31016_, new_n31017_,
    new_n31018_, new_n31019_, new_n31020_, new_n31021_, new_n31022_,
    new_n31023_, new_n31024_, new_n31025_, new_n31026_, new_n31027_,
    new_n31028_, new_n31029_, new_n31030_, new_n31031_, new_n31032_,
    new_n31033_, new_n31034_, new_n31035_, new_n31036_, new_n31037_,
    new_n31038_, new_n31039_, new_n31040_, new_n31041_, new_n31042_,
    new_n31043_, new_n31044_, new_n31045_, new_n31046_, new_n31047_,
    new_n31048_, new_n31049_, new_n31050_, new_n31051_, new_n31052_,
    new_n31053_, new_n31054_, new_n31055_, new_n31056_, new_n31057_,
    new_n31058_, new_n31059_, new_n31060_, new_n31061_, new_n31062_,
    new_n31063_, new_n31064_, new_n31065_, new_n31066_, new_n31067_,
    new_n31068_, new_n31069_, new_n31070_, new_n31071_, new_n31072_,
    new_n31073_, new_n31074_, new_n31075_, new_n31076_, new_n31077_,
    new_n31078_, new_n31079_, new_n31080_, new_n31081_, new_n31082_,
    new_n31083_, new_n31084_, new_n31085_, new_n31086_, new_n31087_,
    new_n31088_, new_n31089_, new_n31090_, new_n31091_, new_n31092_,
    new_n31093_, new_n31094_, new_n31095_, new_n31096_, new_n31097_,
    new_n31098_, new_n31099_, new_n31100_, new_n31101_, new_n31102_,
    new_n31103_, new_n31104_, new_n31105_, new_n31106_, new_n31107_,
    new_n31108_, new_n31109_, new_n31110_, new_n31111_, new_n31112_,
    new_n31113_, new_n31114_, new_n31115_, new_n31116_, new_n31117_,
    new_n31118_, new_n31119_, new_n31120_, new_n31121_, new_n31122_,
    new_n31123_, new_n31124_, new_n31125_, new_n31126_, new_n31127_,
    new_n31128_, new_n31129_, new_n31130_, new_n31131_, new_n31132_,
    new_n31133_, new_n31134_, new_n31135_, new_n31136_, new_n31137_,
    new_n31138_, new_n31139_, new_n31140_, new_n31141_, new_n31142_,
    new_n31143_, new_n31144_, new_n31145_, new_n31146_, new_n31147_,
    new_n31148_, new_n31149_, new_n31150_, new_n31151_, new_n31152_,
    new_n31153_, new_n31154_, new_n31155_, new_n31156_, new_n31157_,
    new_n31158_, new_n31159_, new_n31160_, new_n31161_, new_n31162_,
    new_n31163_, new_n31164_, new_n31165_, new_n31166_, new_n31167_,
    new_n31168_, new_n31169_, new_n31170_, new_n31171_, new_n31172_,
    new_n31173_, new_n31174_, new_n31175_, new_n31176_, new_n31177_,
    new_n31178_, new_n31179_, new_n31180_, new_n31181_, new_n31182_,
    new_n31183_, new_n31184_, new_n31185_, new_n31186_, new_n31187_,
    new_n31188_, new_n31189_, new_n31190_, new_n31191_, new_n31192_,
    new_n31193_, new_n31194_, new_n31195_, new_n31196_, new_n31197_,
    new_n31198_, new_n31199_, new_n31200_, new_n31201_, new_n31203_,
    new_n31204_, new_n31205_, new_n31206_, new_n31207_, new_n31208_,
    new_n31209_, new_n31210_, new_n31211_, new_n31212_, new_n31213_,
    new_n31214_, new_n31215_, new_n31216_, new_n31217_, new_n31218_,
    new_n31219_, new_n31220_, new_n31221_, new_n31222_, new_n31223_,
    new_n31224_, new_n31225_, new_n31226_, new_n31227_, new_n31228_,
    new_n31229_, new_n31230_, new_n31231_, new_n31232_, new_n31233_,
    new_n31234_, new_n31235_, new_n31236_, new_n31237_, new_n31238_,
    new_n31239_, new_n31240_, new_n31241_, new_n31242_, new_n31243_,
    new_n31244_, new_n31245_, new_n31246_, new_n31247_, new_n31248_,
    new_n31249_, new_n31250_, new_n31251_, new_n31252_, new_n31253_,
    new_n31254_, new_n31255_, new_n31256_, new_n31257_, new_n31258_,
    new_n31259_, new_n31260_, new_n31262_, new_n31263_, new_n31264_,
    new_n31265_, new_n31266_, new_n31267_, new_n31268_, new_n31269_,
    new_n31270_, new_n31271_, new_n31272_, new_n31273_, new_n31274_,
    new_n31275_, new_n31276_, new_n31277_, new_n31278_, new_n31279_,
    new_n31280_, new_n31281_, new_n31282_, new_n31283_, new_n31284_,
    new_n31285_, new_n31286_, new_n31287_, new_n31288_, new_n31289_,
    new_n31290_, new_n31291_, new_n31292_, new_n31293_, new_n31294_,
    new_n31295_, new_n31296_, new_n31297_, new_n31298_, new_n31299_,
    new_n31300_, new_n31301_, new_n31302_, new_n31303_, new_n31304_,
    new_n31305_, new_n31306_, new_n31307_, new_n31308_, new_n31309_,
    new_n31310_, new_n31311_, new_n31312_, new_n31313_, new_n31314_,
    new_n31315_, new_n31316_, new_n31317_, new_n31318_, new_n31319_,
    new_n31320_, new_n31321_, new_n31322_, new_n31323_, new_n31324_,
    new_n31325_, new_n31326_, new_n31327_, new_n31328_, new_n31329_,
    new_n31330_, new_n31331_, new_n31332_, new_n31333_, new_n31334_,
    new_n31335_, new_n31336_, new_n31337_, new_n31338_, new_n31339_,
    new_n31340_, new_n31341_, new_n31342_, new_n31343_, new_n31344_,
    new_n31345_, new_n31346_, new_n31347_, new_n31348_, new_n31349_,
    new_n31350_, new_n31351_, new_n31352_, new_n31353_, new_n31354_,
    new_n31355_, new_n31356_, new_n31357_, new_n31358_, new_n31360_,
    new_n31361_, new_n31362_, new_n31363_, new_n31364_, new_n31365_,
    new_n31366_, new_n31368_, new_n31369_, new_n31370_, new_n31371_,
    new_n31372_, new_n31373_, new_n31374_, new_n31375_, new_n31376_,
    new_n31377_, new_n31378_, new_n31379_, new_n31380_, new_n31381_,
    new_n31382_, new_n31383_, new_n31384_, new_n31385_, new_n31386_,
    new_n31387_, new_n31388_, new_n31389_, new_n31390_, new_n31391_,
    new_n31392_, new_n31393_, new_n31394_, new_n31395_, new_n31396_,
    new_n31397_, new_n31398_, new_n31399_, new_n31400_, new_n31401_,
    new_n31402_, new_n31403_, new_n31404_, new_n31405_, new_n31406_,
    new_n31407_, new_n31408_, new_n31409_, new_n31410_, new_n31411_,
    new_n31412_, new_n31413_, new_n31414_, new_n31415_, new_n31416_,
    new_n31417_, new_n31418_, new_n31419_, new_n31420_, new_n31421_,
    new_n31422_, new_n31423_, new_n31424_, new_n31425_, new_n31426_,
    new_n31427_, new_n31428_, new_n31429_, new_n31430_, new_n31431_,
    new_n31432_, new_n31433_, new_n31434_, new_n31435_, new_n31436_,
    new_n31437_, new_n31438_, new_n31439_, new_n31440_, new_n31441_,
    new_n31442_, new_n31443_, new_n31444_, new_n31445_, new_n31446_,
    new_n31447_, new_n31448_, new_n31449_, new_n31450_, new_n31451_,
    new_n31452_, new_n31453_, new_n31454_, new_n31455_, new_n31456_,
    new_n31457_, new_n31458_, new_n31459_, new_n31460_, new_n31461_,
    new_n31462_, new_n31463_, new_n31464_, new_n31465_, new_n31466_,
    new_n31467_, new_n31468_, new_n31469_, new_n31470_, new_n31471_,
    new_n31472_, new_n31473_, new_n31474_, new_n31475_, new_n31476_,
    new_n31477_, new_n31478_, new_n31479_, new_n31480_, new_n31481_,
    new_n31482_, new_n31483_, new_n31484_, new_n31485_, new_n31486_,
    new_n31487_, new_n31488_, new_n31489_, new_n31490_, new_n31491_,
    new_n31492_, new_n31493_, new_n31494_, new_n31495_, new_n31496_,
    new_n31497_, new_n31498_, new_n31499_, new_n31500_, new_n31501_,
    new_n31502_, new_n31503_, new_n31504_, new_n31505_, new_n31506_,
    new_n31507_, new_n31508_, new_n31509_, new_n31510_, new_n31511_,
    new_n31512_, new_n31513_, new_n31514_, new_n31515_, new_n31516_,
    new_n31517_, new_n31518_, new_n31519_, new_n31520_, new_n31521_,
    new_n31522_, new_n31523_, new_n31524_, new_n31525_, new_n31526_,
    new_n31527_, new_n31528_, new_n31529_, new_n31530_, new_n31531_,
    new_n31532_, new_n31533_, new_n31534_, new_n31535_, new_n31536_,
    new_n31537_, new_n31538_, new_n31539_, new_n31540_, new_n31541_,
    new_n31542_, new_n31543_, new_n31544_, new_n31545_, new_n31546_,
    new_n31547_, new_n31548_, new_n31549_, new_n31550_, new_n31551_,
    new_n31552_, new_n31553_, new_n31554_, new_n31555_, new_n31556_,
    new_n31557_, new_n31558_, new_n31559_, new_n31560_, new_n31562_,
    new_n31563_, new_n31564_, new_n31565_, new_n31566_, new_n31567_,
    new_n31568_, new_n31569_, new_n31570_, new_n31571_, new_n31572_,
    new_n31573_, new_n31574_, new_n31575_, new_n31576_, new_n31577_,
    new_n31578_, new_n31579_, new_n31580_, new_n31581_, new_n31582_,
    new_n31583_, new_n31584_, new_n31585_, new_n31586_, new_n31587_,
    new_n31588_, new_n31589_, new_n31590_, new_n31591_, new_n31592_,
    new_n31593_, new_n31594_, new_n31595_, new_n31596_, new_n31597_,
    new_n31598_, new_n31599_, new_n31600_, new_n31601_, new_n31602_,
    new_n31603_, new_n31604_, new_n31605_, new_n31606_, new_n31607_,
    new_n31608_, new_n31609_, new_n31610_, new_n31611_, new_n31612_,
    new_n31613_, new_n31614_, new_n31615_, new_n31616_, new_n31617_,
    new_n31618_, new_n31619_, new_n31620_, new_n31621_, new_n31622_,
    new_n31623_, new_n31624_, new_n31625_, new_n31626_, new_n31627_,
    new_n31628_, new_n31629_, new_n31630_, new_n31631_, new_n31632_,
    new_n31633_, new_n31634_, new_n31635_, new_n31636_, new_n31637_,
    new_n31638_, new_n31639_, new_n31640_, new_n31641_, new_n31642_,
    new_n31643_, new_n31644_, new_n31645_, new_n31646_, new_n31647_,
    new_n31648_, new_n31649_, new_n31650_, new_n31651_, new_n31652_,
    new_n31653_, new_n31654_, new_n31655_, new_n31656_, new_n31657_,
    new_n31658_, new_n31659_, new_n31660_, new_n31661_, new_n31662_,
    new_n31663_, new_n31664_, new_n31665_, new_n31666_, new_n31667_,
    new_n31668_, new_n31669_, new_n31670_, new_n31671_, new_n31672_,
    new_n31673_, new_n31674_, new_n31675_, new_n31676_, new_n31677_,
    new_n31678_, new_n31679_, new_n31680_, new_n31681_, new_n31682_,
    new_n31683_, new_n31684_, new_n31685_, new_n31686_, new_n31687_,
    new_n31688_, new_n31689_, new_n31690_, new_n31691_, new_n31692_,
    new_n31693_, new_n31694_, new_n31695_, new_n31696_, new_n31697_,
    new_n31698_, new_n31699_, new_n31700_, new_n31701_, new_n31702_,
    new_n31703_, new_n31704_, new_n31706_, new_n31708_, new_n31709_,
    new_n31710_, new_n31711_, new_n31712_, new_n31713_, new_n31714_,
    new_n31715_, new_n31716_, new_n31717_, new_n31718_, new_n31719_,
    new_n31720_, new_n31721_, new_n31722_, new_n31723_, new_n31724_,
    new_n31725_, new_n31726_, new_n31727_, new_n31728_, new_n31729_,
    new_n31730_, new_n31731_, new_n31732_, new_n31733_, new_n31734_,
    new_n31735_, new_n31736_, new_n31737_, new_n31738_, new_n31739_,
    new_n31740_, new_n31741_, new_n31742_, new_n31743_, new_n31744_,
    new_n31745_, new_n31746_, new_n31747_, new_n31748_, new_n31749_,
    new_n31750_, new_n31751_, new_n31752_, new_n31753_, new_n31754_,
    new_n31755_, new_n31756_, new_n31757_, new_n31758_, new_n31759_,
    new_n31760_, new_n31761_, new_n31762_, new_n31763_, new_n31764_,
    new_n31765_, new_n31766_, new_n31767_, new_n31768_, new_n31769_,
    new_n31770_, new_n31771_, new_n31772_, new_n31773_, new_n31774_,
    new_n31775_, new_n31776_, new_n31777_, new_n31778_, new_n31779_,
    new_n31780_, new_n31781_, new_n31782_, new_n31783_, new_n31784_,
    new_n31785_, new_n31786_, new_n31787_, new_n31788_, new_n31789_,
    new_n31790_, new_n31791_, new_n31792_, new_n31793_, new_n31794_,
    new_n31795_, new_n31796_, new_n31797_, new_n31798_, new_n31799_,
    new_n31800_, new_n31801_, new_n31802_, new_n31803_, new_n31804_,
    new_n31805_, new_n31806_, new_n31807_, new_n31808_, new_n31809_,
    new_n31810_, new_n31812_, new_n31813_, new_n31814_, new_n31815_,
    new_n31816_, new_n31817_, new_n31818_, new_n31819_, new_n31820_,
    new_n31821_, new_n31822_, new_n31823_, new_n31824_, new_n31825_,
    new_n31826_, new_n31827_, new_n31828_, new_n31829_, new_n31830_,
    new_n31831_, new_n31832_, new_n31833_, new_n31834_, new_n31835_,
    new_n31836_, new_n31838_, new_n31839_, new_n31840_, new_n31841_,
    new_n31842_, new_n31843_, new_n31844_, new_n31845_, new_n31846_,
    new_n31847_, new_n31848_, new_n31849_, new_n31850_, new_n31851_,
    new_n31852_, new_n31853_, new_n31854_, new_n31855_, new_n31856_,
    new_n31857_, new_n31858_, new_n31859_, new_n31860_, new_n31861_,
    new_n31862_, new_n31863_, new_n31864_, new_n31865_, new_n31866_,
    new_n31868_, new_n31869_, new_n31870_, new_n31871_, new_n31872_,
    new_n31873_, new_n31874_, new_n31875_, new_n31876_, new_n31877_,
    new_n31878_, new_n31879_, new_n31880_, new_n31881_, new_n31882_,
    new_n31883_, new_n31884_, new_n31885_, new_n31886_, new_n31887_,
    new_n31888_, new_n31889_, new_n31890_, new_n31891_, new_n31892_,
    new_n31893_, new_n31894_, new_n31895_, new_n31897_, new_n31898_,
    new_n31899_, new_n31900_, new_n31901_, new_n31902_, new_n31903_,
    new_n31904_, new_n31905_, new_n31906_, new_n31907_, new_n31908_,
    new_n31909_, new_n31910_, new_n31911_, new_n31912_, new_n31913_,
    new_n31914_, new_n31915_, new_n31916_, new_n31917_, new_n31918_,
    new_n31919_, new_n31920_, new_n31921_, new_n31922_, new_n31923_,
    new_n31924_, new_n31925_, new_n31926_, new_n31927_, new_n31928_,
    new_n31929_, new_n31930_, new_n31931_, new_n31932_, new_n31933_,
    new_n31934_, new_n31935_, new_n31936_, new_n31937_, new_n31938_,
    new_n31939_, new_n31940_, new_n31941_, new_n31942_, new_n31943_,
    new_n31944_, new_n31945_, new_n31946_, new_n31947_, new_n31948_,
    new_n31949_, new_n31950_, new_n31951_, new_n31952_, new_n31953_,
    new_n31954_, new_n31955_, new_n31956_, new_n31957_, new_n31958_,
    new_n31959_, new_n31960_, new_n31961_, new_n31962_, new_n31963_,
    new_n31965_, new_n31966_, new_n31967_, new_n31968_, new_n31969_,
    new_n31970_, new_n31971_, new_n31972_, new_n31973_, new_n31974_,
    new_n31975_, new_n31976_, new_n31977_, new_n31978_, new_n31979_,
    new_n31980_, new_n31981_, new_n31982_, new_n31983_, new_n31984_,
    new_n31985_, new_n31986_, new_n31987_, new_n31988_, new_n31989_,
    new_n31990_, new_n31991_, new_n31992_, new_n31993_, new_n31994_,
    new_n31995_, new_n31996_, new_n31997_, new_n31998_, new_n31999_,
    new_n32000_, new_n32001_, new_n32002_, new_n32003_, new_n32004_,
    new_n32005_, new_n32006_, new_n32007_, new_n32008_, new_n32009_,
    new_n32010_, new_n32011_, new_n32012_, new_n32013_, new_n32014_,
    new_n32015_, new_n32016_, new_n32017_, new_n32018_, new_n32019_,
    new_n32020_, new_n32021_, new_n32022_, new_n32023_, new_n32024_,
    new_n32025_, new_n32026_, new_n32027_, new_n32028_, new_n32029_,
    new_n32030_, new_n32031_, new_n32032_, new_n32033_, new_n32034_,
    new_n32035_, new_n32036_, new_n32037_, new_n32038_, new_n32039_,
    new_n32040_, new_n32041_, new_n32042_, new_n32043_, new_n32044_,
    new_n32045_, new_n32046_, new_n32047_, new_n32048_, new_n32049_,
    new_n32050_, new_n32051_, new_n32052_, new_n32053_, new_n32054_,
    new_n32055_, new_n32056_, new_n32057_, new_n32058_, new_n32059_,
    new_n32060_, new_n32061_, new_n32062_, new_n32063_, new_n32064_,
    new_n32065_, new_n32066_, new_n32067_, new_n32068_, new_n32069_,
    new_n32070_, new_n32071_, new_n32072_, new_n32073_, new_n32074_,
    new_n32075_, new_n32076_, new_n32077_, new_n32078_, new_n32079_,
    new_n32080_, new_n32081_, new_n32082_, new_n32083_, new_n32084_,
    new_n32085_, new_n32086_, new_n32087_, new_n32088_, new_n32089_,
    new_n32090_, new_n32091_, new_n32092_, new_n32093_, new_n32094_,
    new_n32095_, new_n32096_, new_n32097_, new_n32098_, new_n32099_,
    new_n32100_, new_n32101_, new_n32102_, new_n32103_, new_n32104_,
    new_n32105_, new_n32106_, new_n32107_, new_n32108_, new_n32109_,
    new_n32110_, new_n32111_, new_n32112_, new_n32113_, new_n32114_,
    new_n32115_, new_n32116_, new_n32117_, new_n32118_, new_n32119_,
    new_n32120_, new_n32121_, new_n32122_, new_n32123_, new_n32124_,
    new_n32125_, new_n32126_, new_n32127_, new_n32128_, new_n32129_,
    new_n32130_, new_n32131_, new_n32132_, new_n32133_, new_n32134_,
    new_n32135_, new_n32136_, new_n32137_, new_n32138_, new_n32139_,
    new_n32140_, new_n32141_, new_n32142_, new_n32143_, new_n32144_,
    new_n32145_, new_n32146_, new_n32147_, new_n32148_, new_n32149_,
    new_n32150_, new_n32151_, new_n32152_, new_n32153_, new_n32154_,
    new_n32155_, new_n32156_, new_n32157_, new_n32158_, new_n32159_,
    new_n32160_, new_n32161_, new_n32162_, new_n32163_, new_n32164_,
    new_n32165_, new_n32166_, new_n32167_, new_n32168_, new_n32169_,
    new_n32170_, new_n32171_, new_n32172_, new_n32173_, new_n32174_,
    new_n32175_, new_n32176_, new_n32177_, new_n32178_, new_n32179_,
    new_n32180_, new_n32181_, new_n32182_, new_n32183_, new_n32184_,
    new_n32185_, new_n32186_, new_n32187_, new_n32188_, new_n32189_,
    new_n32190_, new_n32191_, new_n32192_, new_n32193_, new_n32194_,
    new_n32195_, new_n32196_, new_n32197_, new_n32198_, new_n32199_,
    new_n32200_, new_n32201_, new_n32202_, new_n32203_, new_n32204_,
    new_n32205_, new_n32206_, new_n32207_, new_n32208_, new_n32209_,
    new_n32210_, new_n32211_, new_n32212_, new_n32213_, new_n32214_,
    new_n32215_, new_n32216_, new_n32217_, new_n32218_, new_n32219_,
    new_n32220_, new_n32221_, new_n32222_, new_n32223_, new_n32224_,
    new_n32225_, new_n32226_, new_n32227_, new_n32228_, new_n32229_,
    new_n32230_, new_n32231_, new_n32232_, new_n32233_, new_n32234_,
    new_n32235_, new_n32236_, new_n32238_, new_n32239_, new_n32240_,
    new_n32241_, new_n32242_, new_n32243_, new_n32244_, new_n32245_,
    new_n32246_, new_n32247_, new_n32248_, new_n32249_, new_n32250_,
    new_n32251_, new_n32252_, new_n32253_, new_n32254_, new_n32255_,
    new_n32256_, new_n32257_, new_n32258_, new_n32259_, new_n32260_,
    new_n32261_, new_n32262_, new_n32263_, new_n32264_, new_n32265_,
    new_n32266_, new_n32267_, new_n32268_, new_n32269_, new_n32270_,
    new_n32271_, new_n32272_, new_n32273_, new_n32274_, new_n32275_,
    new_n32276_, new_n32277_, new_n32278_, new_n32279_, new_n32280_,
    new_n32281_, new_n32282_, new_n32283_, new_n32284_, new_n32285_,
    new_n32286_, new_n32287_, new_n32288_, new_n32289_, new_n32290_,
    new_n32291_, new_n32292_, new_n32293_, new_n32294_, new_n32295_,
    new_n32296_, new_n32297_, new_n32298_, new_n32299_, new_n32300_,
    new_n32301_, new_n32302_, new_n32303_, new_n32304_, new_n32305_,
    new_n32306_, new_n32307_, new_n32308_, new_n32309_, new_n32310_,
    new_n32311_, new_n32312_, new_n32313_, new_n32314_, new_n32315_,
    new_n32316_, new_n32317_, new_n32318_, new_n32319_, new_n32320_,
    new_n32321_, new_n32322_, new_n32323_, new_n32324_, new_n32325_,
    new_n32326_, new_n32327_, new_n32328_, new_n32329_, new_n32330_,
    new_n32331_, new_n32332_, new_n32333_, new_n32334_, new_n32335_,
    new_n32336_, new_n32337_, new_n32338_, new_n32339_, new_n32340_,
    new_n32341_, new_n32342_, new_n32343_, new_n32344_, new_n32345_,
    new_n32346_, new_n32347_, new_n32348_, new_n32349_, new_n32350_,
    new_n32351_, new_n32352_, new_n32353_, new_n32354_, new_n32355_,
    new_n32356_, new_n32357_, new_n32358_, new_n32359_, new_n32360_,
    new_n32361_, new_n32362_, new_n32363_, new_n32364_, new_n32365_,
    new_n32366_, new_n32367_, new_n32368_, new_n32369_, new_n32370_,
    new_n32371_, new_n32372_, new_n32373_, new_n32374_, new_n32375_,
    new_n32376_, new_n32377_, new_n32378_, new_n32379_, new_n32380_,
    new_n32381_, new_n32382_, new_n32383_, new_n32384_, new_n32385_,
    new_n32386_, new_n32387_, new_n32388_, new_n32389_, new_n32390_,
    new_n32391_, new_n32392_, new_n32393_, new_n32394_, new_n32395_,
    new_n32396_, new_n32397_, new_n32398_, new_n32399_, new_n32400_,
    new_n32401_, new_n32402_, new_n32403_, new_n32404_, new_n32405_,
    new_n32406_, new_n32407_, new_n32408_, new_n32409_, new_n32410_,
    new_n32411_, new_n32412_, new_n32413_, new_n32414_, new_n32415_,
    new_n32416_, new_n32417_, new_n32418_, new_n32419_, new_n32420_,
    new_n32421_, new_n32422_, new_n32423_, new_n32424_, new_n32425_,
    new_n32426_, new_n32427_, new_n32428_, new_n32429_, new_n32430_,
    new_n32431_, new_n32432_, new_n32433_, new_n32434_, new_n32435_,
    new_n32436_, new_n32437_, new_n32438_, new_n32439_, new_n32440_,
    new_n32441_, new_n32442_, new_n32443_, new_n32444_, new_n32445_,
    new_n32446_, new_n32447_, new_n32448_, new_n32449_, new_n32450_,
    new_n32451_, new_n32452_, new_n32453_, new_n32454_, new_n32455_,
    new_n32457_, new_n32458_, new_n32459_, new_n32460_, new_n32461_,
    new_n32462_, new_n32463_, new_n32464_, new_n32465_, new_n32466_,
    new_n32467_, new_n32468_, new_n32469_, new_n32470_, new_n32471_,
    new_n32472_, new_n32473_, new_n32474_, new_n32475_, new_n32476_,
    new_n32477_, new_n32478_, new_n32479_, new_n32480_, new_n32481_,
    new_n32482_, new_n32483_, new_n32484_, new_n32485_, new_n32486_,
    new_n32487_, new_n32488_, new_n32489_, new_n32490_, new_n32491_,
    new_n32492_, new_n32493_, new_n32494_, new_n32495_, new_n32496_,
    new_n32497_, new_n32498_, new_n32499_, new_n32500_, new_n32501_,
    new_n32502_, new_n32503_, new_n32504_, new_n32505_, new_n32506_,
    new_n32507_, new_n32508_, new_n32509_, new_n32510_, new_n32511_,
    new_n32512_, new_n32513_, new_n32514_, new_n32515_, new_n32516_,
    new_n32517_, new_n32518_, new_n32520_, new_n32521_, new_n32522_,
    new_n32524_, new_n32525_, new_n32526_, new_n32528_, new_n32529_,
    new_n32530_, new_n32531_, new_n32532_, new_n32533_, new_n32534_,
    new_n32535_, new_n32536_, new_n32537_, new_n32538_, new_n32539_,
    new_n32540_, new_n32541_, new_n32542_, new_n32543_, new_n32544_,
    new_n32545_, new_n32546_, new_n32547_, new_n32548_, new_n32549_,
    new_n32550_, new_n32551_, new_n32552_, new_n32553_, new_n32554_,
    new_n32555_, new_n32556_, new_n32557_, new_n32558_, new_n32559_,
    new_n32560_, new_n32561_, new_n32562_, new_n32563_, new_n32564_,
    new_n32565_, new_n32566_, new_n32567_, new_n32568_, new_n32569_,
    new_n32570_, new_n32571_, new_n32572_, new_n32573_, new_n32574_,
    new_n32575_, new_n32576_, new_n32577_, new_n32578_, new_n32579_,
    new_n32580_, new_n32581_, new_n32582_, new_n32583_, new_n32584_,
    new_n32585_, new_n32586_, new_n32587_, new_n32588_, new_n32589_,
    new_n32590_, new_n32591_, new_n32592_, new_n32593_, new_n32594_,
    new_n32595_, new_n32596_, new_n32597_, new_n32598_, new_n32599_,
    new_n32600_, new_n32601_, new_n32602_, new_n32603_, new_n32604_,
    new_n32605_, new_n32606_, new_n32607_, new_n32608_, new_n32609_,
    new_n32610_, new_n32611_, new_n32612_, new_n32613_, new_n32614_,
    new_n32615_, new_n32616_, new_n32617_, new_n32618_, new_n32619_,
    new_n32620_, new_n32621_, new_n32622_, new_n32623_, new_n32624_,
    new_n32625_, new_n32626_, new_n32627_, new_n32628_, new_n32629_,
    new_n32630_, new_n32631_, new_n32632_, new_n32633_, new_n32634_,
    new_n32635_, new_n32636_, new_n32637_, new_n32638_, new_n32639_,
    new_n32640_, new_n32641_, new_n32642_, new_n32643_, new_n32644_,
    new_n32645_, new_n32646_, new_n32647_, new_n32648_, new_n32649_,
    new_n32650_, new_n32651_, new_n32652_, new_n32653_, new_n32654_,
    new_n32655_, new_n32656_, new_n32657_, new_n32658_, new_n32659_,
    new_n32660_, new_n32661_, new_n32662_, new_n32663_, new_n32664_,
    new_n32665_, new_n32666_, new_n32667_, new_n32668_, new_n32669_,
    new_n32670_, new_n32671_, new_n32672_, new_n32673_, new_n32674_,
    new_n32675_, new_n32676_, new_n32677_, new_n32678_, new_n32679_,
    new_n32680_, new_n32681_, new_n32682_, new_n32683_, new_n32684_,
    new_n32685_, new_n32686_, new_n32687_, new_n32688_, new_n32689_,
    new_n32690_, new_n32691_, new_n32692_, new_n32693_, new_n32694_,
    new_n32695_, new_n32696_, new_n32697_, new_n32698_, new_n32699_,
    new_n32700_, new_n32701_, new_n32702_, new_n32703_, new_n32704_,
    new_n32705_, new_n32706_, new_n32707_, new_n32708_, new_n32709_,
    new_n32710_, new_n32711_, new_n32712_, new_n32713_, new_n32714_,
    new_n32715_, new_n32716_, new_n32717_, new_n32718_, new_n32719_,
    new_n32720_, new_n32721_, new_n32722_, new_n32723_, new_n32724_,
    new_n32725_, new_n32726_, new_n32727_, new_n32728_, new_n32729_,
    new_n32730_, new_n32731_, new_n32732_, new_n32733_, new_n32734_,
    new_n32735_, new_n32736_, new_n32737_, new_n32738_, new_n32740_,
    new_n32741_, new_n32742_, new_n32743_, new_n32744_, new_n32745_,
    new_n32746_, new_n32747_, new_n32748_, new_n32749_, new_n32750_,
    new_n32751_, new_n32752_, new_n32753_, new_n32754_, new_n32755_,
    new_n32756_, new_n32757_, new_n32758_, new_n32759_, new_n32760_,
    new_n32761_, new_n32762_, new_n32763_, new_n32764_, new_n32765_,
    new_n32766_, new_n32767_, new_n32768_, new_n32769_, new_n32770_,
    new_n32771_, new_n32772_, new_n32773_, new_n32774_, new_n32775_,
    new_n32776_, new_n32777_, new_n32778_, new_n32779_, new_n32780_,
    new_n32781_, new_n32783_, new_n32784_, new_n32785_, new_n32786_,
    new_n32787_, new_n32788_, new_n32789_, new_n32790_, new_n32791_,
    new_n32792_, new_n32793_, new_n32794_, new_n32795_, new_n32796_,
    new_n32797_, new_n32798_, new_n32799_, new_n32800_, new_n32801_,
    new_n32802_, new_n32803_, new_n32804_, new_n32805_, new_n32806_,
    new_n32807_, new_n32809_, new_n32810_, new_n32811_, new_n32812_,
    new_n32813_, new_n32814_, new_n32815_, new_n32816_, new_n32817_,
    new_n32818_, new_n32819_, new_n32820_, new_n32822_, new_n32823_,
    new_n32824_, new_n32825_, new_n32826_, new_n32827_, new_n32828_,
    new_n32829_, new_n32830_, new_n32831_, new_n32832_, new_n32833_,
    new_n32834_, new_n32835_, new_n32836_, new_n32837_, new_n32838_,
    new_n32839_, new_n32840_, new_n32841_, new_n32842_, new_n32843_,
    new_n32844_, new_n32845_, new_n32846_, new_n32848_, new_n32849_,
    new_n32850_, new_n32851_, new_n32852_, new_n32853_, new_n32854_,
    new_n32855_, new_n32856_, new_n32857_, new_n32858_, new_n32859_,
    new_n32860_, new_n32861_, new_n32862_, new_n32863_, new_n32864_,
    new_n32865_, new_n32866_, new_n32867_, new_n32868_, new_n32869_,
    new_n32870_, new_n32871_, new_n32872_, new_n32873_, new_n32874_,
    new_n32875_, new_n32876_, new_n32877_, new_n32878_, new_n32879_,
    new_n32880_, new_n32881_, new_n32882_, new_n32883_, new_n32884_,
    new_n32885_, new_n32886_, new_n32887_, new_n32888_, new_n32889_,
    new_n32890_, new_n32891_, new_n32892_, new_n32893_, new_n32894_,
    new_n32895_, new_n32896_, new_n32897_, new_n32898_, new_n32899_,
    new_n32900_, new_n32901_, new_n32902_, new_n32903_, new_n32905_,
    new_n32906_, new_n32907_, new_n32908_, new_n32909_, new_n32910_,
    new_n32911_, new_n32912_, new_n32913_, new_n32914_, new_n32915_,
    new_n32916_, new_n32917_, new_n32918_, new_n32919_, new_n32920_,
    new_n32921_, new_n32922_, new_n32923_, new_n32924_, new_n32925_,
    new_n32926_, new_n32927_, new_n32928_, new_n32929_, new_n32930_,
    new_n32931_, new_n32932_, new_n32933_, new_n32934_, new_n32935_,
    new_n32936_, new_n32937_, new_n32938_, new_n32939_, new_n32940_,
    new_n32941_, new_n32942_, new_n32943_, new_n32944_, new_n32945_,
    new_n32946_, new_n32947_, new_n32948_, new_n32949_, new_n32950_,
    new_n32951_, new_n32952_, new_n32953_, new_n32954_, new_n32955_,
    new_n32956_, new_n32957_, new_n32958_, new_n32959_, new_n32960_,
    new_n32961_, new_n32962_, new_n32963_, new_n32964_, new_n32965_,
    new_n32966_, new_n32967_, new_n32968_, new_n32969_, new_n32970_,
    new_n32971_, new_n32972_, new_n32973_, new_n32974_, new_n32975_,
    new_n32976_, new_n32977_, new_n32978_, new_n32979_, new_n32980_,
    new_n32981_, new_n32982_, new_n32983_, new_n32984_, new_n32985_,
    new_n32986_, new_n32987_, new_n32988_, new_n32989_, new_n32990_,
    new_n32991_, new_n32992_, new_n32993_, new_n32994_, new_n32995_,
    new_n32996_, new_n32997_, new_n32998_, new_n32999_, new_n33000_,
    new_n33001_, new_n33002_, new_n33003_, new_n33004_, new_n33005_,
    new_n33006_, new_n33007_, new_n33008_, new_n33009_, new_n33010_,
    new_n33011_, new_n33012_, new_n33013_, new_n33014_, new_n33015_,
    new_n33016_, new_n33017_, new_n33018_, new_n33019_, new_n33020_,
    new_n33021_, new_n33022_, new_n33023_, new_n33024_, new_n33025_,
    new_n33026_, new_n33027_, new_n33028_, new_n33029_, new_n33030_,
    new_n33031_, new_n33032_, new_n33033_, new_n33034_, new_n33036_,
    new_n33037_, new_n33038_, new_n33039_, new_n33040_, new_n33041_,
    new_n33042_, new_n33043_, new_n33044_, new_n33045_, new_n33047_,
    new_n33048_, new_n33049_, new_n33050_, new_n33051_, new_n33052_,
    new_n33053_, new_n33054_, new_n33055_, new_n33056_, new_n33057_,
    new_n33058_, new_n33059_, new_n33060_, new_n33061_, new_n33062_,
    new_n33063_, new_n33064_, new_n33065_, new_n33066_, new_n33067_,
    new_n33068_, new_n33069_, new_n33070_, new_n33071_, new_n33072_,
    new_n33073_, new_n33074_, new_n33075_, new_n33076_, new_n33077_,
    new_n33078_, new_n33079_, new_n33080_, new_n33081_, new_n33082_,
    new_n33083_, new_n33084_, new_n33085_, new_n33086_, new_n33087_,
    new_n33088_, new_n33089_, new_n33090_, new_n33091_, new_n33092_,
    new_n33093_, new_n33094_, new_n33095_, new_n33096_, new_n33097_,
    new_n33098_, new_n33099_, new_n33100_, new_n33101_, new_n33102_,
    new_n33103_, new_n33104_, new_n33105_, new_n33106_, new_n33107_,
    new_n33108_, new_n33109_, new_n33110_, new_n33111_, new_n33112_,
    new_n33113_, new_n33114_, new_n33115_, new_n33116_, new_n33117_,
    new_n33118_, new_n33119_, new_n33120_, new_n33121_, new_n33122_,
    new_n33123_, new_n33124_, new_n33125_, new_n33126_, new_n33127_,
    new_n33128_, new_n33129_, new_n33130_, new_n33131_, new_n33132_,
    new_n33133_, new_n33134_, new_n33135_, new_n33136_, new_n33137_,
    new_n33138_, new_n33139_, new_n33140_, new_n33141_, new_n33142_,
    new_n33143_, new_n33144_, new_n33145_, new_n33146_, new_n33147_,
    new_n33148_, new_n33149_, new_n33150_, new_n33151_, new_n33152_,
    new_n33153_, new_n33154_, new_n33155_, new_n33156_, new_n33157_,
    new_n33158_, new_n33159_, new_n33160_, new_n33161_, new_n33162_,
    new_n33163_, new_n33164_, new_n33165_, new_n33166_, new_n33167_,
    new_n33168_, new_n33169_, new_n33170_, new_n33171_, new_n33172_,
    new_n33173_, new_n33174_, new_n33175_, new_n33176_, new_n33177_,
    new_n33178_, new_n33179_, new_n33180_, new_n33181_, new_n33188_,
    new_n33189_, new_n33190_, new_n33191_, new_n33192_, new_n33193_,
    new_n33194_, new_n33195_, new_n33196_, new_n33197_, new_n33198_,
    new_n33199_, new_n33200_, new_n33201_, new_n33202_, new_n33203_,
    new_n33204_, new_n33205_, new_n33206_, new_n33207_, new_n33208_,
    new_n33209_, new_n33210_, new_n33211_, new_n33212_, new_n33213_,
    new_n33214_, new_n33216_, new_n33217_, new_n33218_, new_n33219_,
    new_n33220_, new_n33221_, new_n33222_, new_n33223_, new_n33224_,
    new_n33225_, new_n33226_, new_n33227_, new_n33228_, new_n33229_,
    new_n33230_, new_n33231_, new_n33232_, new_n33233_, new_n33234_,
    new_n33235_, new_n33236_, new_n33237_, new_n33238_, new_n33239_,
    new_n33240_, new_n33241_, new_n33242_, new_n33243_, new_n33244_,
    new_n33245_, new_n33246_, new_n33247_, new_n33248_, new_n33249_,
    new_n33250_, new_n33251_, new_n33252_, new_n33253_, new_n33254_,
    new_n33255_, new_n33256_, new_n33257_, new_n33258_, new_n33259_,
    new_n33260_, new_n33261_, new_n33262_, new_n33263_, new_n33264_,
    new_n33265_, new_n33266_, new_n33267_, new_n33268_, new_n33269_,
    new_n33270_, new_n33271_, new_n33272_, new_n33273_, new_n33274_,
    new_n33275_, new_n33276_, new_n33277_, new_n33278_, new_n33279_,
    new_n33280_, new_n33281_, new_n33282_, new_n33283_, new_n33284_,
    new_n33285_, new_n33286_, new_n33287_, new_n33288_, new_n33289_,
    new_n33290_, new_n33291_, new_n33292_, new_n33293_, new_n33294_,
    new_n33295_, new_n33296_, new_n33297_, new_n33298_, new_n33299_,
    new_n33300_, new_n33301_, new_n33302_, new_n33303_, new_n33304_,
    new_n33305_, new_n33306_, new_n33307_, new_n33308_, new_n33309_,
    new_n33310_, new_n33311_, new_n33312_, new_n33313_, new_n33314_,
    new_n33315_, new_n33316_, new_n33317_, new_n33318_, new_n33319_,
    new_n33320_, new_n33321_, new_n33322_, new_n33323_, new_n33324_,
    new_n33325_, new_n33326_, new_n33327_, new_n33328_, new_n33329_,
    new_n33330_, new_n33331_, new_n33332_, new_n33333_, new_n33334_,
    new_n33335_, new_n33336_, new_n33337_, new_n33338_, new_n33339_,
    new_n33340_, new_n33341_, new_n33342_, new_n33343_, new_n33344_,
    new_n33345_, new_n33346_, new_n33347_, new_n33348_, new_n33349_,
    new_n33350_, new_n33351_, new_n33352_, new_n33353_, new_n33354_,
    new_n33355_, new_n33356_, new_n33357_, new_n33358_, new_n33359_,
    new_n33360_, new_n33361_, new_n33362_, new_n33363_, new_n33364_,
    new_n33365_, new_n33366_, new_n33367_, new_n33368_, new_n33369_,
    new_n33370_, new_n33371_, new_n33372_, new_n33373_, new_n33374_,
    new_n33375_, new_n33376_, new_n33377_, new_n33378_, new_n33379_,
    new_n33380_, new_n33381_, new_n33383_, new_n33384_, new_n33385_,
    new_n33386_, new_n33387_, new_n33388_, new_n33389_, new_n33390_,
    new_n33391_, new_n33392_, new_n33393_, new_n33394_, new_n33395_,
    new_n33397_, new_n33398_, new_n33399_, new_n33400_, new_n33401_,
    new_n33402_, new_n33403_, new_n33404_, new_n33405_, new_n33406_,
    new_n33407_, new_n33408_, new_n33409_, new_n33410_, new_n33411_,
    new_n33412_, new_n33413_, new_n33414_, new_n33415_, new_n33416_,
    new_n33417_, new_n33418_, new_n33419_, new_n33420_, new_n33421_,
    new_n33422_, new_n33423_, new_n33424_, new_n33425_, new_n33426_,
    new_n33427_, new_n33428_, new_n33429_, new_n33430_, new_n33431_,
    new_n33432_, new_n33433_, new_n33434_, new_n33435_, new_n33436_,
    new_n33437_, new_n33438_, new_n33439_, new_n33440_, new_n33441_,
    new_n33442_, new_n33443_, new_n33444_, new_n33445_, new_n33446_,
    new_n33447_, new_n33448_, new_n33449_, new_n33450_, new_n33452_,
    new_n33453_, new_n33454_, new_n33455_, new_n33456_, new_n33457_,
    new_n33458_, new_n33459_, new_n33460_, new_n33461_, new_n33462_,
    new_n33463_, new_n33464_, new_n33465_, new_n33466_, new_n33467_,
    new_n33468_, new_n33469_, new_n33470_, new_n33471_, new_n33472_,
    new_n33473_, new_n33474_, new_n33475_, new_n33476_, new_n33478_,
    new_n33479_, new_n33480_, new_n33481_, new_n33482_, new_n33483_,
    new_n33484_, new_n33485_, new_n33486_, new_n33487_, new_n33488_,
    new_n33489_, new_n33490_, new_n33491_, new_n33492_, new_n33493_,
    new_n33494_, new_n33495_, new_n33496_, new_n33497_, new_n33498_,
    new_n33499_, new_n33500_, new_n33501_, new_n33502_, new_n33503_,
    new_n33504_, new_n33505_, new_n33506_, new_n33507_, new_n33508_,
    new_n33509_, new_n33510_, new_n33511_, new_n33512_, new_n33513_,
    new_n33514_, new_n33515_, new_n33516_, new_n33517_, new_n33518_,
    new_n33519_, new_n33520_, new_n33521_, new_n33522_, new_n33523_,
    new_n33524_, new_n33525_, new_n33526_, new_n33527_, new_n33528_,
    new_n33529_, new_n33530_, new_n33531_, new_n33532_, new_n33533_,
    new_n33534_, new_n33535_, new_n33536_, new_n33537_, new_n33538_,
    new_n33539_, new_n33540_, new_n33541_, new_n33542_, new_n33543_,
    new_n33544_, new_n33545_, new_n33546_, new_n33547_, new_n33548_,
    new_n33549_, new_n33550_, new_n33551_, new_n33552_, new_n33553_,
    new_n33554_, new_n33555_, new_n33556_, new_n33557_, new_n33558_,
    new_n33559_, new_n33560_, new_n33561_, new_n33562_, new_n33563_,
    new_n33564_, new_n33565_, new_n33566_, new_n33567_, new_n33568_,
    new_n33569_, new_n33570_, new_n33571_, new_n33572_, new_n33573_,
    new_n33574_, new_n33575_, new_n33576_, new_n33577_, new_n33578_,
    new_n33579_, new_n33580_, new_n33581_, new_n33582_, new_n33583_,
    new_n33584_, new_n33585_, new_n33586_, new_n33587_, new_n33588_,
    new_n33589_, new_n33590_, new_n33591_, new_n33592_, new_n33593_,
    new_n33594_, new_n33595_, new_n33596_, new_n33598_, new_n33599_,
    new_n33600_, new_n33602_, new_n33603_, new_n33604_, new_n33605_,
    new_n33606_, new_n33607_, new_n33608_, new_n33609_, new_n33610_,
    new_n33611_, new_n33613_, new_n33614_, new_n33615_, new_n33616_,
    new_n33617_, new_n33618_, new_n33619_, new_n33620_, new_n33621_,
    new_n33622_, new_n33623_, new_n33624_, new_n33625_, new_n33626_,
    new_n33627_, new_n33628_, new_n33629_, new_n33630_, new_n33631_,
    new_n33633_, new_n33634_, new_n33635_, new_n33636_, new_n33637_,
    new_n33639_, new_n33640_, new_n33641_, new_n33642_, new_n33643_,
    new_n33644_, new_n33645_, new_n33646_, new_n33649_, new_n33650_,
    new_n33651_, new_n33652_, new_n33653_, new_n33654_, new_n33655_,
    new_n33656_, new_n33657_, new_n33658_, new_n33659_, new_n33660_,
    new_n33661_, new_n33662_, new_n33663_, new_n33664_, new_n33665_,
    new_n33666_, new_n33667_, new_n33668_, new_n33669_, new_n33670_,
    new_n33671_, new_n33672_, new_n33673_, new_n33674_, new_n33675_,
    new_n33676_, new_n33677_, new_n33678_, new_n33679_, new_n33680_,
    new_n33681_, new_n33682_, new_n33683_, new_n33684_, new_n33685_,
    new_n33686_, new_n33687_, new_n33688_, new_n33689_, new_n33690_,
    new_n33691_, new_n33692_, new_n33693_, new_n33694_, new_n33695_,
    new_n33696_, new_n33697_, new_n33698_, new_n33699_, new_n33700_,
    new_n33701_, new_n33702_, new_n33703_, new_n33704_, new_n33705_,
    new_n33706_, new_n33707_, new_n33708_, new_n33709_, new_n33710_,
    new_n33711_, new_n33712_, new_n33713_, new_n33714_, new_n33715_,
    new_n33716_, new_n33717_, new_n33718_, new_n33719_, new_n33720_,
    new_n33721_, new_n33722_, new_n33723_, new_n33724_, new_n33725_,
    new_n33726_, new_n33727_, new_n33728_, new_n33729_, new_n33730_,
    new_n33731_, new_n33732_, new_n33733_, new_n33736_, new_n33737_,
    new_n33738_, new_n33739_, new_n33740_, new_n33741_, new_n33742_,
    new_n33743_, new_n33744_, new_n33745_, new_n33746_, new_n33747_,
    new_n33748_, new_n33749_, new_n33750_, new_n33751_, new_n33752_,
    new_n33753_, new_n33754_, new_n33755_, new_n33756_, new_n33757_,
    new_n33758_, new_n33759_, new_n33760_, new_n33761_, new_n33762_,
    new_n33763_, new_n33764_, new_n33765_, new_n33766_, new_n33767_,
    new_n33768_, new_n33769_, new_n33770_, new_n33771_, new_n33772_,
    new_n33773_, new_n33774_, new_n33775_, new_n33776_, new_n33777_,
    new_n33778_, new_n33779_, new_n33780_, new_n33781_, new_n33782_,
    new_n33783_, new_n33784_, new_n33785_, new_n33786_, new_n33787_,
    new_n33788_, new_n33789_, new_n33790_, new_n33791_, new_n33792_,
    new_n33793_, new_n33794_, new_n33795_, new_n33796_, new_n33800_,
    new_n33801_, new_n33802_, new_n33803_, new_n33804_, new_n33805_,
    new_n33806_, new_n33807_, new_n33808_, new_n33809_, new_n33810_,
    new_n33811_, new_n33812_, new_n33813_, new_n33814_, new_n33815_,
    new_n33816_, new_n33817_, new_n33819_, new_n33820_, new_n33821_,
    new_n33822_, new_n33823_, new_n33824_, new_n33825_, new_n33826_,
    new_n33827_, new_n33828_, new_n33829_, new_n33830_, new_n33831_,
    new_n33832_, new_n33833_, new_n33834_, new_n33835_, new_n33836_,
    new_n33837_, new_n33838_, new_n33839_, new_n33840_, new_n33841_,
    new_n33842_, new_n33843_, new_n33844_, new_n33845_, new_n33846_,
    new_n33847_, new_n33848_, new_n33849_, new_n33850_, new_n33851_,
    new_n33852_, new_n33853_, new_n33854_, new_n33855_, new_n33856_,
    new_n33857_, new_n33858_, new_n33859_, new_n33860_, new_n33861_,
    new_n33862_, new_n33863_, new_n33864_, new_n33865_, new_n33866_,
    new_n33867_, new_n33868_, new_n33869_, new_n33870_, new_n33871_,
    new_n33872_, new_n33873_, new_n33874_, new_n33875_, new_n33876_,
    new_n33877_, new_n33878_, new_n33879_, new_n33880_, new_n33881_,
    new_n33882_, new_n33883_, new_n33884_, new_n33885_, new_n33886_,
    new_n33887_, new_n33888_, new_n33889_, new_n33890_, new_n33891_,
    new_n33892_, new_n33893_, new_n33894_, new_n33895_, new_n33896_,
    new_n33897_, new_n33898_, new_n33899_, new_n33900_, new_n33901_,
    new_n33902_, new_n33903_, new_n33904_, new_n33905_, new_n33906_,
    new_n33907_, new_n33908_, new_n33909_, new_n33910_, new_n33911_,
    new_n33912_, new_n33913_, new_n33914_, new_n33915_, new_n33916_,
    new_n33917_, new_n33918_, new_n33919_, new_n33920_, new_n33921_,
    new_n33922_, new_n33923_, new_n33924_, new_n33925_, new_n33926_,
    new_n33927_, new_n33928_, new_n33929_, new_n33930_, new_n33931_,
    new_n33932_, new_n33933_, new_n33934_, new_n33935_, new_n33936_,
    new_n33937_, new_n33938_, new_n33939_, new_n33940_, new_n33941_,
    new_n33942_, new_n33943_, new_n33944_, new_n33945_, new_n33946_,
    new_n33947_, new_n33948_, new_n33949_, new_n33950_, new_n33951_,
    new_n33952_, new_n33953_, new_n33954_, new_n33955_, new_n33956_,
    new_n33957_, new_n33958_, new_n33959_, new_n33960_, new_n33961_,
    new_n33962_, new_n33963_, new_n33964_, new_n33965_, new_n33966_,
    new_n33967_, new_n33968_, new_n33969_, new_n33970_, new_n33971_,
    new_n33972_, new_n33973_, new_n33974_, new_n33975_, new_n33976_,
    new_n33977_, new_n33978_, new_n33979_, new_n33980_, new_n33981_,
    new_n33982_, new_n33984_, new_n33985_, new_n33986_, new_n33987_,
    new_n33988_, new_n33990_, new_n33991_, new_n33992_, new_n33993_,
    new_n33994_, new_n33996_, new_n33997_, new_n33998_, new_n33999_,
    new_n34000_, new_n34002_, new_n34003_, new_n34004_, new_n34005_,
    new_n34006_, new_n34008_, new_n34009_, new_n34010_, new_n34011_,
    new_n34013_, new_n34014_, new_n34015_, new_n34016_, new_n34017_,
    new_n34018_, new_n34020_, new_n34021_, new_n34022_, new_n34023_,
    new_n34024_, new_n34025_, new_n34027_, new_n34028_, new_n34029_,
    new_n34030_, new_n34031_, new_n34032_, new_n34033_, new_n34034_,
    new_n34035_, new_n34036_, new_n34037_, new_n34038_, new_n34039_,
    new_n34040_, new_n34041_, new_n34042_, new_n34043_, new_n34044_,
    new_n34045_, new_n34046_, new_n34047_, new_n34048_, new_n34049_,
    new_n34050_, new_n34051_, new_n34053_, new_n34054_, new_n34055_,
    new_n34056_, new_n34057_, new_n34058_, new_n34059_, new_n34060_,
    new_n34061_, new_n34062_, new_n34063_, new_n34064_, new_n34065_,
    new_n34066_, new_n34067_, new_n34068_, new_n34069_, new_n34070_,
    new_n34071_, new_n34072_, new_n34073_, new_n34074_, new_n34075_,
    new_n34076_, new_n34077_, new_n34078_, new_n34079_, new_n34080_,
    new_n34081_, new_n34082_, new_n34083_, new_n34084_, new_n34085_,
    new_n34086_, new_n34087_, new_n34088_, new_n34089_, new_n34090_,
    new_n34091_, new_n34092_, new_n34093_, new_n34094_, new_n34095_,
    new_n34096_, new_n34097_, new_n34098_, new_n34099_, new_n34100_,
    new_n34101_, new_n34102_, new_n34103_, new_n34104_, new_n34105_,
    new_n34106_, new_n34107_, new_n34108_, new_n34109_, new_n34110_,
    new_n34111_, new_n34112_, new_n34113_, new_n34114_, new_n34115_,
    new_n34116_, new_n34117_, new_n34118_, new_n34119_, new_n34120_,
    new_n34121_, new_n34122_, new_n34123_, new_n34124_, new_n34125_,
    new_n34126_, new_n34127_, new_n34128_, new_n34129_, new_n34130_,
    new_n34131_, new_n34132_, new_n34133_, new_n34134_, new_n34135_,
    new_n34136_, new_n34137_, new_n34138_, new_n34139_, new_n34140_,
    new_n34141_, new_n34142_, new_n34143_, new_n34144_, new_n34145_,
    new_n34146_, new_n34147_, new_n34148_, new_n34149_, new_n34150_,
    new_n34151_, new_n34152_, new_n34153_, new_n34154_, new_n34155_,
    new_n34156_, new_n34157_, new_n34158_, new_n34159_, new_n34160_,
    new_n34161_, new_n34162_, new_n34163_, new_n34164_, new_n34165_,
    new_n34166_, new_n34167_, new_n34168_, new_n34169_, new_n34170_,
    new_n34171_, new_n34172_, new_n34173_, new_n34174_, new_n34175_,
    new_n34176_, new_n34177_, new_n34178_, new_n34179_, new_n34180_,
    new_n34181_, new_n34182_, new_n34183_, new_n34184_, new_n34185_,
    new_n34186_, new_n34187_, new_n34188_, new_n34189_, new_n34190_,
    new_n34191_, new_n34192_, new_n34193_, new_n34194_, new_n34195_,
    new_n34196_, new_n34197_, new_n34198_, new_n34200_, new_n34201_,
    new_n34202_, new_n34203_, new_n34204_, new_n34205_, new_n34206_,
    new_n34207_, new_n34208_, new_n34209_, new_n34210_, new_n34211_,
    new_n34212_, new_n34213_, new_n34214_, new_n34215_, new_n34216_,
    new_n34217_, new_n34218_, new_n34219_, new_n34220_, new_n34221_,
    new_n34222_, new_n34223_, new_n34224_, new_n34225_, new_n34226_,
    new_n34227_, new_n34228_, new_n34229_, new_n34230_, new_n34231_,
    new_n34232_, new_n34234_, new_n34235_, new_n34236_, new_n34237_,
    new_n34238_, new_n34239_, new_n34240_, new_n34241_, new_n34242_,
    new_n34243_, new_n34244_, new_n34245_, new_n34246_, new_n34247_,
    new_n34248_, new_n34249_, new_n34250_, new_n34251_, new_n34252_,
    new_n34253_, new_n34254_, new_n34255_, new_n34256_, new_n34257_,
    new_n34258_, new_n34259_, new_n34260_, new_n34261_, new_n34262_,
    new_n34264_, new_n34265_, new_n34266_, new_n34267_, new_n34268_,
    new_n34269_, new_n34270_, new_n34271_, new_n34272_, new_n34273_,
    new_n34274_, new_n34275_, new_n34276_, new_n34277_, new_n34278_,
    new_n34279_, new_n34280_, new_n34281_, new_n34282_, new_n34283_,
    new_n34284_, new_n34285_, new_n34286_, new_n34287_, new_n34288_,
    new_n34289_, new_n34290_, new_n34291_, new_n34292_, new_n34293_,
    new_n34294_, new_n34295_, new_n34296_, new_n34297_, new_n34298_,
    new_n34299_, new_n34300_, new_n34301_, new_n34302_, new_n34303_,
    new_n34304_, new_n34305_, new_n34306_, new_n34307_, new_n34308_,
    new_n34309_, new_n34310_, new_n34311_, new_n34312_, new_n34313_,
    new_n34315_, new_n34316_, new_n34317_, new_n34318_, new_n34319_,
    new_n34320_, new_n34321_, new_n34322_, new_n34323_, new_n34324_,
    new_n34325_, new_n34326_, new_n34327_, new_n34328_, new_n34329_,
    new_n34330_, new_n34331_, new_n34332_, new_n34333_, new_n34334_,
    new_n34335_, new_n34336_, new_n34337_, new_n34338_, new_n34339_,
    new_n34340_, new_n34341_, new_n34342_, new_n34343_, new_n34344_,
    new_n34345_, new_n34346_, new_n34347_, new_n34348_, new_n34349_,
    new_n34350_, new_n34351_, new_n34352_, new_n34353_, new_n34354_,
    new_n34355_, new_n34356_, new_n34357_, new_n34358_, new_n34359_,
    new_n34360_, new_n34361_, new_n34362_, new_n34363_, new_n34364_,
    new_n34365_, new_n34366_, new_n34367_, new_n34368_, new_n34369_,
    new_n34370_, new_n34371_, new_n34372_, new_n34373_, new_n34374_,
    new_n34375_, new_n34376_, new_n34377_, new_n34378_, new_n34379_,
    new_n34380_, new_n34381_, new_n34382_, new_n34383_, new_n34384_,
    new_n34385_, new_n34386_, new_n34387_, new_n34388_, new_n34389_,
    new_n34390_, new_n34391_, new_n34392_, new_n34393_, new_n34394_,
    new_n34395_, new_n34396_, new_n34397_, new_n34398_, new_n34399_,
    new_n34400_, new_n34401_, new_n34402_, new_n34403_, new_n34404_,
    new_n34405_, new_n34406_, new_n34407_, new_n34408_, new_n34409_,
    new_n34410_, new_n34411_, new_n34412_, new_n34413_, new_n34414_,
    new_n34415_, new_n34416_, new_n34417_, new_n34418_, new_n34419_,
    new_n34420_, new_n34421_, new_n34422_, new_n34423_, new_n34424_,
    new_n34425_, new_n34426_, new_n34427_, new_n34428_, new_n34429_,
    new_n34430_, new_n34431_, new_n34432_, new_n34433_, new_n34434_,
    new_n34435_, new_n34436_, new_n34437_, new_n34438_, new_n34439_,
    new_n34440_, new_n34441_, new_n34443_, new_n34444_, new_n34445_,
    new_n34446_, new_n34447_, new_n34448_, new_n34449_, new_n34450_,
    new_n34451_, new_n34452_, new_n34453_, new_n34454_, new_n34455_,
    new_n34456_, new_n34458_, new_n34459_, new_n34460_, new_n34461_,
    new_n34462_, new_n34463_, new_n34464_, new_n34465_, new_n34466_,
    new_n34467_, new_n34468_, new_n34469_, new_n34470_, new_n34471_,
    new_n34472_, new_n34473_, new_n34474_, new_n34475_, new_n34476_,
    new_n34477_, new_n34478_, new_n34479_, new_n34480_, new_n34481_,
    new_n34482_, new_n34483_, new_n34484_, new_n34485_, new_n34486_,
    new_n34487_, new_n34488_, new_n34489_, new_n34490_, new_n34491_,
    new_n34492_, new_n34494_, new_n34495_, new_n34496_, new_n34497_,
    new_n34498_, new_n34499_, new_n34500_, new_n34501_, new_n34502_,
    new_n34503_, new_n34504_, new_n34505_, new_n34506_, new_n34507_,
    new_n34508_, new_n34509_, new_n34510_, new_n34511_, new_n34512_,
    new_n34513_, new_n34514_, new_n34515_, new_n34516_, new_n34517_,
    new_n34518_, new_n34519_, new_n34520_, new_n34521_, new_n34522_,
    new_n34523_, new_n34524_, new_n34525_, new_n34526_, new_n34527_,
    new_n34528_, new_n34529_, new_n34530_, new_n34531_, new_n34532_,
    new_n34533_, new_n34534_, new_n34535_, new_n34536_, new_n34537_,
    new_n34538_, new_n34539_, new_n34540_, new_n34541_, new_n34542_,
    new_n34543_, new_n34544_, new_n34545_, new_n34546_, new_n34547_,
    new_n34548_, new_n34549_, new_n34550_, new_n34551_, new_n34552_,
    new_n34553_, new_n34554_, new_n34555_, new_n34556_, new_n34557_,
    new_n34558_, new_n34559_, new_n34560_, new_n34561_, new_n34562_,
    new_n34563_, new_n34564_, new_n34565_, new_n34566_, new_n34567_,
    new_n34568_, new_n34569_, new_n34570_, new_n34571_, new_n34572_,
    new_n34573_, new_n34574_, new_n34575_, new_n34576_, new_n34577_,
    new_n34578_, new_n34579_, new_n34581_, new_n34582_, new_n34583_,
    new_n34584_, new_n34585_, new_n34586_, new_n34587_, new_n34588_,
    new_n34589_, new_n34590_, new_n34591_, new_n34592_, new_n34593_,
    new_n34594_, new_n34595_, new_n34596_, new_n34597_, new_n34598_,
    new_n34599_, new_n34600_, new_n34601_, new_n34602_, new_n34603_,
    new_n34604_, new_n34605_, new_n34606_, new_n34607_, new_n34608_,
    new_n34609_, new_n34610_, new_n34612_, new_n34613_, new_n34614_,
    new_n34615_, new_n34616_, new_n34617_, new_n34618_, new_n34619_,
    new_n34620_, new_n34621_, new_n34626_, new_n34627_, new_n34628_,
    new_n34629_, new_n34630_, new_n34631_, new_n34632_, new_n34633_,
    new_n34634_, new_n34635_, new_n34637_, new_n34638_, new_n34639_,
    new_n34640_, new_n34641_, new_n34642_, new_n34643_, new_n34644_,
    new_n34645_, new_n34646_, new_n34647_, new_n34648_, new_n34649_,
    new_n34650_, new_n34651_, new_n34652_, new_n34653_, new_n34654_,
    new_n34655_, new_n34656_, new_n34657_, new_n34658_, new_n34659_,
    new_n34660_, new_n34661_, new_n34662_, new_n34663_, new_n34664_,
    new_n34665_, new_n34666_, new_n34667_, new_n34668_, new_n34669_,
    new_n34670_, new_n34671_, new_n34672_, new_n34673_, new_n34674_,
    new_n34675_, new_n34676_, new_n34678_, new_n34679_, new_n34680_,
    new_n34681_, new_n34682_, new_n34683_, new_n34684_, new_n34685_,
    new_n34686_, new_n34687_, new_n34688_, new_n34689_, new_n34690_,
    new_n34691_, new_n34692_, new_n34693_, new_n34694_, new_n34695_,
    new_n34696_, new_n34697_, new_n34698_, new_n34699_, new_n34700_,
    new_n34701_, new_n34702_, new_n34703_, new_n34704_, new_n34705_,
    new_n34706_, new_n34709_, new_n34710_, new_n34711_, new_n34712_,
    new_n34713_, new_n34714_, new_n34715_, new_n34716_, new_n34717_,
    new_n34718_, new_n34719_, new_n34720_, new_n34721_, new_n34722_,
    new_n34723_, new_n34724_, new_n34725_, new_n34726_, new_n34727_,
    new_n34728_, new_n34729_, new_n34730_, new_n34731_, new_n34732_,
    new_n34733_, new_n34734_, new_n34735_, new_n34736_, new_n34737_,
    new_n34738_, new_n34739_, new_n34740_, new_n34741_, new_n34742_,
    new_n34743_, new_n34744_, new_n34745_, new_n34747_, new_n34748_,
    new_n34749_, new_n34750_, new_n34751_, new_n34752_, new_n34753_,
    new_n34754_, new_n34755_, new_n34756_, new_n34757_, new_n34758_,
    new_n34759_, new_n34760_, new_n34761_, new_n34762_, new_n34763_,
    new_n34764_, new_n34765_, new_n34766_, new_n34767_, new_n34768_,
    new_n34769_, new_n34770_, new_n34771_, new_n34772_, new_n34773_,
    new_n34774_, new_n34775_, new_n34779_, new_n34780_, new_n34781_,
    new_n34782_, new_n34783_, new_n34785_, new_n34786_, new_n34787_,
    new_n34788_, new_n34789_, new_n34790_, new_n34791_, new_n34792_,
    new_n34793_, new_n34794_, new_n34795_, new_n34796_, new_n34797_,
    new_n34798_, new_n34799_, new_n34800_, new_n34801_, new_n34802_,
    new_n34803_, new_n34804_, new_n34805_, new_n34806_, new_n34807_,
    new_n34808_, new_n34809_, new_n34810_, new_n34811_, new_n34812_,
    new_n34813_, new_n34814_, new_n34815_, new_n34817_, new_n34818_,
    new_n34819_, new_n34820_, new_n34821_, new_n34822_, new_n34823_,
    new_n34824_, new_n34825_, new_n34826_, new_n34827_, new_n34828_,
    new_n34829_, new_n34830_, new_n34831_, new_n34832_, new_n34833_,
    new_n34834_, new_n34835_, new_n34836_, new_n34837_, new_n34838_,
    new_n34839_, new_n34840_, new_n34841_, new_n34842_, new_n34843_,
    new_n34844_, new_n34845_, new_n34846_, new_n34847_, new_n34848_,
    new_n34849_, new_n34850_, new_n34851_, new_n34852_, new_n34853_,
    new_n34854_, new_n34855_, new_n34856_, new_n34857_, new_n34858_,
    new_n34859_, new_n34860_, new_n34861_, new_n34862_, new_n34863_,
    new_n34864_, new_n34865_, new_n34866_, new_n34868_, new_n34869_,
    new_n34870_, new_n34871_, new_n34872_, new_n34873_, new_n34874_,
    new_n34875_, new_n34876_, new_n34877_, new_n34878_, new_n34882_,
    new_n34883_, new_n34884_, new_n34885_, new_n34887_, new_n34888_,
    new_n34889_, new_n34890_, new_n34891_, new_n34892_, new_n34893_,
    new_n34894_, new_n34895_, new_n34896_, new_n34897_, new_n34898_,
    new_n34899_, new_n34900_, new_n34901_, new_n34902_, new_n34903_,
    new_n34904_, new_n34905_, new_n34906_, new_n34907_, new_n34908_,
    new_n34909_, new_n34910_, new_n34911_, new_n34912_, new_n34913_,
    new_n34914_, new_n34915_, new_n34918_, new_n34919_, new_n34920_,
    new_n34921_, new_n34922_, new_n34923_, new_n34924_, new_n34925_,
    new_n34926_, new_n34927_, new_n34928_, new_n34929_, new_n34930_,
    new_n34931_, new_n34932_, new_n34933_, new_n34934_, new_n34935_,
    new_n34936_, new_n34937_, new_n34938_, new_n34939_, new_n34940_,
    new_n34941_, new_n34942_, new_n34943_, new_n34944_, new_n34945_,
    new_n34946_, new_n34947_, new_n34948_, new_n34949_, new_n34950_,
    new_n34951_, new_n34952_, new_n34953_, new_n34954_, new_n34955_,
    new_n34956_, new_n34957_, new_n34958_, new_n34959_, new_n34960_,
    new_n34961_, new_n34962_, new_n34963_, new_n34964_, new_n34965_,
    new_n34966_, new_n34968_, new_n34969_, new_n34970_, new_n34971_,
    new_n34972_, new_n34973_, new_n34974_, new_n34975_, new_n34976_,
    new_n34977_, new_n34978_, new_n34979_, new_n34980_, new_n34981_,
    new_n34982_, new_n34983_, new_n34984_, new_n34985_, new_n34986_,
    new_n34987_, new_n34988_, new_n34989_, new_n34990_, new_n34991_,
    new_n34992_, new_n34993_, new_n34994_, new_n34995_, new_n34996_,
    new_n34997_, new_n34998_, new_n34999_, new_n35000_, new_n35001_,
    new_n35002_, new_n35003_, new_n35004_, new_n35005_, new_n35006_,
    new_n35007_, new_n35008_, new_n35009_, new_n35011_, new_n35012_,
    new_n35013_, new_n35014_, new_n35015_, new_n35016_, new_n35017_,
    new_n35018_, new_n35019_, new_n35020_, new_n35021_, new_n35022_,
    new_n35023_, new_n35024_, new_n35025_, new_n35026_, new_n35027_,
    new_n35028_, new_n35029_, new_n35030_, new_n35031_, new_n35032_,
    new_n35033_, new_n35034_, new_n35035_, new_n35036_, new_n35037_,
    new_n35038_, new_n35039_, new_n35041_, new_n35042_, new_n35043_,
    new_n35044_, new_n35045_, new_n35046_, new_n35047_, new_n35048_,
    new_n35049_, new_n35050_, new_n35051_, new_n35052_, new_n35053_,
    new_n35054_, new_n35055_, new_n35056_, new_n35057_, new_n35058_,
    new_n35059_, new_n35060_, new_n35061_, new_n35062_, new_n35063_,
    new_n35065_, new_n35066_, new_n35067_, new_n35068_, new_n35069_,
    new_n35070_, new_n35071_, new_n35072_, new_n35073_, new_n35074_,
    new_n35075_, new_n35076_, new_n35077_, new_n35078_, new_n35079_,
    new_n35080_, new_n35081_, new_n35082_, new_n35083_, new_n35084_,
    new_n35085_, new_n35088_, new_n35089_, new_n35091_, new_n35092_,
    new_n35093_, new_n35094_, new_n35095_, new_n35096_, new_n35097_,
    new_n35098_, new_n35099_, new_n35100_, new_n35101_, new_n35102_,
    new_n35103_, new_n35104_, new_n35105_, new_n35106_, new_n35107_,
    new_n35108_, new_n35109_, new_n35110_, new_n35111_, new_n35112_,
    new_n35113_, new_n35114_, new_n35115_, new_n35116_, new_n35117_,
    new_n35118_, new_n35119_, new_n35120_, new_n35121_, new_n35122_,
    new_n35123_, new_n35124_, new_n35125_, new_n35126_, new_n35127_,
    new_n35128_, new_n35129_, new_n35131_, new_n35132_, new_n35134_,
    new_n35135_, new_n35136_, new_n35137_, new_n35138_, new_n35139_,
    new_n35140_, new_n35141_, new_n35142_, new_n35143_, new_n35144_,
    new_n35146_, new_n35147_, new_n35148_, new_n35149_, new_n35150_,
    new_n35151_, new_n35152_, new_n35153_, new_n35154_, new_n35155_,
    new_n35156_, new_n35157_, new_n35158_, new_n35161_, new_n35162_,
    new_n35164_, new_n35166_, new_n35167_, new_n35168_, new_n35169_,
    new_n35170_, new_n35171_, new_n35172_, new_n35173_, new_n35175_,
    new_n35176_, new_n35178_, new_n35179_, new_n35181_, new_n35182_,
    new_n35184_, new_n35185_, new_n35187_, new_n35188_, new_n35190_,
    new_n35192_, new_n35194_, new_n35196_, new_n35198_, new_n35199_,
    new_n35200_, new_n35201_, new_n35203_, new_n35204_, new_n35206_,
    new_n35207_, new_n35209_, new_n35210_, new_n35211_, new_n35212_,
    new_n35213_, new_n35214_, new_n35215_, new_n35216_, new_n35217_,
    new_n35218_, new_n35219_, new_n35220_, new_n35221_, new_n35222_,
    new_n35223_, new_n35224_, new_n35226_, new_n35228_, new_n35230_,
    new_n35232_, new_n35234_, new_n35236_, new_n35238_, new_n35240_,
    new_n35241_, new_n35242_, new_n35243_, new_n35244_, new_n35245_,
    new_n35246_, new_n35247_, new_n35248_, new_n35249_, new_n35250_,
    new_n35251_, new_n35252_, new_n35253_, new_n35254_, new_n35255_,
    new_n35256_, new_n35257_, new_n35259_, new_n35260_, new_n35262_,
    new_n35263_, new_n35265_, new_n35266_, new_n35267_, new_n35269_,
    new_n35270_, new_n35271_, new_n35272_, new_n35273_, new_n35274_,
    new_n35275_, new_n35277_, new_n35278_, new_n35279_, new_n35280_,
    new_n35282_, new_n35283_, new_n35285_, new_n35286_, new_n35287_,
    new_n35289_, new_n35290_, new_n35291_, new_n35292_, new_n35294_,
    new_n35296_, new_n35298_, new_n35299_, new_n35301_, new_n35302_,
    new_n35304_, new_n35306_, new_n35307_, new_n35309_, new_n35310_,
    new_n35312_, new_n35313_, new_n35315_, new_n35317_, new_n35319_,
    new_n35320_, new_n35322_, new_n35323_, new_n35324_, new_n35325_,
    new_n35326_, new_n35327_, new_n35328_, new_n35330_, new_n35331_,
    new_n35332_, new_n35333_, new_n35335_, new_n35336_, new_n35337_,
    new_n35338_, new_n35339_, new_n35340_, new_n35341_, new_n35342_,
    new_n35344_, new_n35346_, new_n35348_, new_n35350_, new_n35351_,
    new_n35353_, new_n35354_, new_n35356_, new_n35357_, new_n35359_,
    new_n35364_, new_n35365_, new_n35367_, new_n35369_, new_n35371_,
    new_n35373_, new_n35375_, new_n35377_, new_n35378_, new_n35380_,
    new_n35381_, new_n35383_, new_n35385_, new_n35386_, new_n35388_,
    new_n35389_, new_n35391_, new_n35392_, new_n35394_, new_n35396_,
    new_n35397_, new_n35399_, new_n35401_, new_n35402_, new_n35404_,
    new_n35405_, new_n35407_, new_n35408_, new_n35410_, new_n35411_,
    new_n35413_, new_n35414_, new_n35416_, new_n35418_, new_n35420_,
    new_n35422_, new_n35424_, new_n35425_, new_n35427_, new_n35428_,
    new_n35430_, new_n35432_, new_n35433_, new_n35435_, new_n35437_,
    new_n35439_, new_n35441_, new_n35443_, new_n35444_, new_n35446_,
    new_n35448_, new_n35450_, new_n35451_, new_n35453_, new_n35455_,
    new_n35457_, new_n35458_, new_n35460_, new_n35461_, new_n35463_,
    new_n35465_, new_n35466_, new_n35468_, new_n35469_, new_n35471_,
    new_n35473_, new_n35475_, new_n35477_, new_n35479_, new_n35481_,
    new_n35482_, new_n35484_, new_n35486_, new_n35488_, new_n35490_,
    new_n35492_, new_n35494_, new_n35496_, new_n35498_, new_n35500_,
    new_n35502_, new_n35504_, new_n35506_, new_n35508_, new_n35510_,
    new_n35512_, new_n35514_, new_n35516_, new_n35518_, new_n35520_,
    new_n35522_, new_n35524_, new_n35526_, new_n35528_, new_n35530_,
    new_n35532_, new_n35533_, new_n35535_, new_n35537_, new_n35539_,
    new_n35541_, new_n35543_, new_n35545_, new_n35547_, new_n35549_,
    new_n35551_, new_n35553_, new_n35555_, new_n35557_, new_n35559_,
    new_n35561_, new_n35563_, new_n35565_, new_n35567_, new_n35569_,
    new_n35571_, new_n35573_, new_n35575_, new_n35577_, new_n35579_,
    new_n35581_, new_n35583_, new_n35584_, new_n35586_, new_n35588_,
    new_n35590_, new_n35592_, new_n35594_, new_n35596_, new_n35598_,
    new_n35600_, new_n35601_, new_n35603_, new_n35605_, new_n35607_,
    new_n35609_, new_n35611_, new_n35613_, new_n35615_, new_n35617_,
    new_n35619_, new_n35621_, new_n35622_, new_n35623_, new_n35624_,
    new_n35625_, new_n35626_, new_n35627_, new_n35628_, new_n35629_,
    new_n35630_, new_n35631_, new_n35632_, new_n35633_, new_n35634_,
    new_n35635_, new_n35636_, new_n35637_, new_n35638_, new_n35639_,
    new_n35640_, new_n35641_, new_n35642_, new_n35644_, new_n35646_,
    new_n35648_, new_n35650_, new_n35652_, new_n35654_, new_n35656_,
    new_n35658_, new_n35659_, new_n35660_, new_n35661_, new_n35662_,
    new_n35663_, new_n35664_, new_n35665_, new_n35666_, new_n35667_,
    new_n35668_, new_n35669_, new_n35670_, new_n35671_, new_n35672_,
    new_n35673_, new_n35674_, new_n35675_, new_n35676_, new_n35678_,
    new_n35679_, new_n35680_, new_n35681_, new_n35682_, new_n35683_,
    new_n35684_, new_n35685_, new_n35686_, new_n35687_, new_n35688_,
    new_n35689_, new_n35690_, new_n35691_, new_n35692_, new_n35694_,
    new_n35695_, new_n35696_, new_n35697_, new_n35698_, new_n35699_,
    new_n35700_, new_n35701_, new_n35702_, new_n35703_, new_n35704_,
    new_n35705_, new_n35706_, new_n35708_, new_n35709_, new_n35710_,
    new_n35711_, new_n35712_, new_n35713_, new_n35714_, new_n35715_,
    new_n35717_, new_n35719_, new_n35720_, new_n35721_, new_n35722_,
    new_n35723_, new_n35724_, new_n35725_, new_n35726_, new_n35727_,
    new_n35728_, new_n35729_, new_n35731_, new_n35732_, new_n35733_,
    new_n35734_, new_n35735_, new_n35736_, new_n35737_, new_n35738_,
    new_n35739_, new_n35740_, new_n35741_, new_n35743_, new_n35744_,
    new_n35745_, new_n35746_, new_n35747_, new_n35748_, new_n35749_,
    new_n35750_, new_n35751_, new_n35752_, new_n35753_, new_n35755_,
    new_n35756_, new_n35757_, new_n35758_, new_n35759_, new_n35760_,
    new_n35761_, new_n35762_, new_n35763_, new_n35764_, new_n35765_,
    new_n35767_, new_n35768_, new_n35769_, new_n35770_, new_n35771_,
    new_n35772_, new_n35774_, new_n35775_, new_n35776_, new_n35777_,
    new_n35778_, new_n35779_, new_n35781_, new_n35782_, new_n35783_,
    new_n35784_, new_n35785_, new_n35786_, new_n35788_, new_n35789_,
    new_n35790_, new_n35791_, new_n35792_, new_n35793_, new_n35797_,
    new_n35798_, new_n35800_, new_n35801_, new_n35803_, new_n35804_,
    new_n35806_, new_n35808_, new_n35809_, new_n35811_, new_n35812_,
    new_n35814_, new_n35815_, new_n35817_, new_n35819_, new_n35820_,
    new_n35822_, new_n35824_, new_n35826_, new_n35828_, new_n35829_,
    new_n35831_, new_n35832_, new_n35833_, new_n35835_, new_n35837_,
    new_n35838_, new_n35840_, new_n35841_, new_n35843_, new_n35844_,
    new_n35846_, new_n35848_, new_n35850_, new_n35852_, new_n35854_,
    new_n35856_, new_n35857_, new_n35859_, new_n35860_, new_n35861_,
    new_n35862_, new_n35863_, new_n35864_, new_n35866_, new_n35867_,
    new_n35869_, new_n35870_, new_n35872_, new_n35873_, new_n35875_,
    new_n35876_, new_n35878_, new_n35879_, new_n35881_, new_n35882_,
    new_n35883_, new_n35884_, new_n35885_, new_n35886_, new_n35887_,
    new_n35889_, new_n35890_, new_n35892_, new_n35893_, new_n35895_,
    new_n35896_, new_n35898_, new_n35899_, new_n35901_, new_n35902_,
    new_n35904_, new_n35905_, new_n35907_, new_n35908_, new_n35910_,
    new_n35912_, new_n35914_, new_n35916_, new_n35918_, new_n35919_,
    new_n35921_, new_n35922_, new_n35924_, new_n35926_, new_n35928_,
    new_n35930_, new_n35932_, new_n35934_, new_n35936_, new_n35937_,
    new_n35939_, new_n35940_, new_n35942_, new_n35943_, new_n35945_,
    new_n35947_, new_n35948_, new_n35950_, new_n35951_, new_n35953_,
    new_n35954_, new_n35956_, new_n35957_, new_n35959_, new_n35961_,
    new_n35963_, new_n35965_, new_n35967_, new_n35969_, new_n35971_,
    new_n35973_, new_n35975_, new_n35977_, new_n35979_, new_n35980_,
    new_n35982_, new_n35984_, new_n35985_, new_n35987_, new_n35988_,
    new_n35990_, new_n35991_, new_n35993_, new_n35994_, new_n35996_,
    new_n35997_, new_n35999_, new_n36000_, new_n36002_, new_n36004_,
    new_n36005_, new_n36007_, new_n36008_, new_n36010_, new_n36011_,
    new_n36013_, new_n36015_, new_n36017_, new_n36018_, new_n36020_,
    new_n36022_, new_n36024_, new_n36025_, new_n36027_, new_n36028_,
    new_n36029_, new_n36030_, new_n36031_, new_n36032_, new_n36033_,
    new_n36034_, new_n36035_, new_n36036_, new_n36037_, new_n36038_,
    new_n36039_, new_n36040_, new_n36041_, new_n36042_, new_n36043_,
    new_n36044_, new_n36045_, new_n36046_, new_n36047_, new_n36048_,
    new_n36049_, new_n36050_, new_n36051_, new_n36052_, new_n36053_,
    new_n36054_, new_n36055_, new_n36056_, new_n36057_, new_n36058_,
    new_n36059_, new_n36060_, new_n36061_, new_n36062_, new_n36063_,
    new_n36064_, new_n36065_, new_n36066_, new_n36067_, new_n36068_,
    new_n36069_, new_n36070_, new_n36071_, new_n36072_, new_n36073_,
    new_n36074_, new_n36075_, new_n36076_, new_n36077_, new_n36078_,
    new_n36079_, new_n36080_, new_n36081_, new_n36082_, new_n36083_,
    new_n36084_, new_n36085_, new_n36086_, new_n36087_, new_n36088_,
    new_n36089_, new_n36090_, new_n36091_, new_n36092_, new_n36093_,
    new_n36094_, new_n36095_, new_n36097_, new_n36098_, new_n36100_,
    new_n36102_, new_n36104_, new_n36106_, new_n36108_, new_n36110_,
    new_n36112_, new_n36114_, new_n36116_, new_n36117_, new_n36119_,
    new_n36121_, new_n36122_, new_n36124_, new_n36125_, new_n36127_,
    new_n36129_, new_n36131_, new_n36133_, new_n36135_, new_n36137_,
    new_n36138_, new_n36140_, new_n36141_, new_n36142_, new_n36143_,
    new_n36145_, new_n36146_, new_n36147_, new_n36148_, new_n36149_,
    new_n36151_, new_n36152_, new_n36154_, new_n36155_, new_n36157_,
    new_n36158_, new_n36160_, new_n36161_, new_n36162_, new_n36163_,
    new_n36164_, new_n36165_, new_n36166_, new_n36167_, new_n36168_,
    new_n36169_, new_n36170_, new_n36171_, new_n36172_, new_n36173_,
    new_n36174_, new_n36175_, new_n36176_, new_n36177_, new_n36178_,
    new_n36179_, new_n36180_, new_n36181_, new_n36182_, new_n36183_,
    new_n36184_, new_n36185_, new_n36186_, new_n36187_, new_n36188_,
    new_n36189_, new_n36190_, new_n36191_, new_n36192_, new_n36193_,
    new_n36194_, new_n36195_, new_n36196_, new_n36197_, new_n36198_,
    new_n36199_, new_n36200_, new_n36201_, new_n36202_, new_n36203_,
    new_n36204_, new_n36205_, new_n36206_, new_n36207_, new_n36208_,
    new_n36209_, new_n36210_, new_n36211_, new_n36212_, new_n36213_,
    new_n36214_, new_n36215_, new_n36216_, new_n36217_, new_n36218_,
    new_n36219_, new_n36220_, new_n36221_, new_n36222_, new_n36223_,
    new_n36224_, new_n36225_, new_n36226_, new_n36227_, new_n36228_,
    new_n36229_, new_n36230_, new_n36231_, new_n36232_, new_n36233_,
    new_n36234_, new_n36235_, new_n36236_, new_n36237_, new_n36238_,
    new_n36239_, new_n36240_, new_n36241_, new_n36242_, new_n36243_,
    new_n36244_, new_n36245_, new_n36246_, new_n36247_, new_n36248_,
    new_n36249_, new_n36250_, new_n36251_, new_n36252_, new_n36253_,
    new_n36254_, new_n36255_, new_n36256_, new_n36257_, new_n36258_,
    new_n36259_, new_n36260_, new_n36261_, new_n36262_, new_n36263_,
    new_n36264_, new_n36265_, new_n36266_, new_n36267_, new_n36268_,
    new_n36269_, new_n36270_, new_n36271_, new_n36272_, new_n36273_,
    new_n36274_, new_n36275_, new_n36276_, new_n36277_, new_n36278_,
    new_n36279_, new_n36280_, new_n36281_, new_n36282_, new_n36283_,
    new_n36284_, new_n36285_, new_n36286_, new_n36287_, new_n36288_,
    new_n36289_, new_n36290_, new_n36291_, new_n36292_, new_n36293_,
    new_n36294_, new_n36295_, new_n36296_, new_n36297_, new_n36298_,
    new_n36299_, new_n36300_, new_n36301_, new_n36302_, new_n36303_,
    new_n36304_, new_n36305_, new_n36306_, new_n36307_, new_n36308_,
    new_n36309_, new_n36310_, new_n36311_, new_n36312_, new_n36313_,
    new_n36314_, new_n36315_, new_n36316_, new_n36317_, new_n36318_,
    new_n36319_, new_n36320_, new_n36321_, new_n36322_, new_n36323_,
    new_n36324_, new_n36325_, new_n36326_, new_n36327_, new_n36328_,
    new_n36329_, new_n36330_, new_n36331_, new_n36332_, new_n36333_,
    new_n36334_, new_n36335_, new_n36336_, new_n36337_, new_n36338_,
    new_n36339_, new_n36340_, new_n36341_, new_n36342_, new_n36343_,
    new_n36344_, new_n36345_, new_n36346_, new_n36347_, new_n36348_,
    new_n36349_, new_n36350_, new_n36351_, new_n36352_, new_n36353_,
    new_n36354_, new_n36355_, new_n36356_, new_n36357_, new_n36358_,
    new_n36359_, new_n36360_, new_n36361_, new_n36362_, new_n36363_,
    new_n36364_, new_n36365_, new_n36366_, new_n36367_, new_n36368_,
    new_n36369_, new_n36370_, new_n36371_, new_n36372_, new_n36373_,
    new_n36374_, new_n36375_, new_n36376_, new_n36377_, new_n36378_,
    new_n36379_, new_n36380_, new_n36381_, new_n36382_, new_n36383_,
    new_n36384_, new_n36385_, new_n36386_, new_n36387_, new_n36388_,
    new_n36389_, new_n36390_, new_n36391_, new_n36392_, new_n36393_,
    new_n36394_, new_n36395_, new_n36396_, new_n36397_, new_n36398_,
    new_n36399_, new_n36400_, new_n36401_, new_n36402_, new_n36403_,
    new_n36404_, new_n36405_, new_n36406_, new_n36407_, new_n36408_,
    new_n36409_, new_n36410_, new_n36411_, new_n36412_, new_n36413_,
    new_n36414_, new_n36415_, new_n36416_, new_n36417_, new_n36418_,
    new_n36419_, new_n36420_, new_n36421_, new_n36422_, new_n36423_,
    new_n36424_, new_n36425_, new_n36426_, new_n36427_, new_n36428_,
    new_n36429_, new_n36430_, new_n36431_, new_n36432_, new_n36433_,
    new_n36434_, new_n36435_, new_n36436_, new_n36437_, new_n36438_,
    new_n36439_, new_n36440_, new_n36441_, new_n36442_, new_n36443_,
    new_n36444_, new_n36445_, new_n36446_, new_n36447_, new_n36448_,
    new_n36449_, new_n36450_, new_n36451_, new_n36452_, new_n36453_,
    new_n36454_, new_n36455_, new_n36456_, new_n36457_, new_n36458_,
    new_n36459_, new_n36460_, new_n36461_, new_n36462_, new_n36463_,
    new_n36464_, new_n36465_, new_n36466_, new_n36467_, new_n36468_,
    new_n36469_, new_n36470_, new_n36471_, new_n36472_, new_n36473_,
    new_n36474_, new_n36475_, new_n36476_, new_n36477_, new_n36478_,
    new_n36479_, new_n36480_, new_n36481_, new_n36482_, new_n36483_,
    new_n36484_, new_n36485_, new_n36486_, new_n36487_, new_n36488_,
    new_n36489_, new_n36490_, new_n36491_, new_n36492_, new_n36493_,
    new_n36494_, new_n36495_, new_n36496_, new_n36497_, new_n36498_,
    new_n36499_, new_n36500_, new_n36501_, new_n36502_, new_n36503_,
    new_n36504_, new_n36505_, new_n36506_, new_n36507_, new_n36508_,
    new_n36509_, new_n36510_, new_n36511_, new_n36512_, new_n36513_,
    new_n36514_, new_n36515_, new_n36516_, new_n36517_, new_n36518_,
    new_n36519_, new_n36520_, new_n36521_, new_n36522_, new_n36523_,
    new_n36524_, new_n36525_, new_n36526_, new_n36527_, new_n36528_,
    new_n36529_, new_n36530_, new_n36531_, new_n36532_, new_n36533_,
    new_n36534_, new_n36535_, new_n36536_, new_n36537_, new_n36538_,
    new_n36539_, new_n36540_, new_n36541_, new_n36542_, new_n36543_,
    new_n36544_, new_n36545_, new_n36546_, new_n36547_, new_n36548_,
    new_n36549_, new_n36550_, new_n36551_, new_n36552_, new_n36553_,
    new_n36554_, new_n36555_, new_n36556_, new_n36557_, new_n36558_,
    new_n36559_, new_n36560_, new_n36561_, new_n36562_, new_n36563_,
    new_n36564_, new_n36565_, new_n36566_, new_n36567_, new_n36568_,
    new_n36569_, new_n36570_, new_n36571_, new_n36572_, new_n36573_,
    new_n36574_, new_n36575_, new_n36576_, new_n36577_, new_n36578_,
    new_n36579_, new_n36580_, new_n36581_, new_n36582_, new_n36583_,
    new_n36584_, new_n36585_, new_n36586_, new_n36587_, new_n36588_,
    new_n36589_, new_n36590_, new_n36591_, new_n36592_, new_n36593_,
    new_n36594_, new_n36595_, new_n36596_, new_n36597_, new_n36598_,
    new_n36599_, new_n36600_, new_n36601_, new_n36602_, new_n36603_,
    new_n36604_, new_n36605_, new_n36606_, new_n36607_, new_n36608_,
    new_n36609_, new_n36610_, new_n36611_, new_n36612_, new_n36613_,
    new_n36614_, new_n36615_, new_n36616_, new_n36617_, new_n36618_,
    new_n36619_, new_n36620_, new_n36621_, new_n36622_, new_n36623_,
    new_n36624_, new_n36625_, new_n36626_, new_n36627_, new_n36628_,
    new_n36629_, new_n36630_, new_n36631_, new_n36632_, new_n36633_,
    new_n36634_, new_n36635_, new_n36636_, new_n36637_, new_n36638_,
    new_n36639_, new_n36640_, new_n36641_, new_n36642_, new_n36643_,
    new_n36644_, new_n36645_, new_n36646_, new_n36647_, new_n36648_,
    new_n36649_, new_n36650_, new_n36651_, new_n36652_, new_n36653_,
    new_n36654_, new_n36655_, new_n36656_, new_n36657_, new_n36658_,
    new_n36659_, new_n36660_, new_n36661_, new_n36662_, new_n36663_,
    new_n36664_, new_n36665_, new_n36666_, new_n36667_, new_n36668_,
    new_n36669_, new_n36670_, new_n36671_, new_n36672_, new_n36673_,
    new_n36674_, new_n36675_, new_n36676_, new_n36677_, new_n36678_,
    new_n36679_, new_n36680_, new_n36681_, new_n36682_, new_n36683_,
    new_n36684_, new_n36685_, new_n36686_, new_n36687_, new_n36688_,
    new_n36689_, new_n36690_, new_n36691_, new_n36692_, new_n36693_,
    new_n36694_, new_n36695_, new_n36696_, new_n36697_, new_n36698_,
    new_n36699_, new_n36700_, new_n36701_, new_n36702_, new_n36703_,
    new_n36704_, new_n36705_, new_n36706_, new_n36707_, new_n36708_,
    new_n36709_, new_n36710_, new_n36711_, new_n36712_, new_n36713_,
    new_n36714_, new_n36715_, new_n36716_, new_n36717_, new_n36718_,
    new_n36719_, new_n36720_, new_n36721_, new_n36722_, new_n36723_,
    new_n36724_, new_n36725_, new_n36726_, new_n36727_, new_n36728_,
    new_n36729_, new_n36730_, new_n36731_, new_n36732_, new_n36733_,
    new_n36734_, new_n36735_, new_n36736_, new_n36737_, new_n36738_,
    new_n36739_, new_n36740_, new_n36741_, new_n36742_, new_n36743_,
    new_n36744_, new_n36745_, new_n36746_, new_n36747_, new_n36748_,
    new_n36749_, new_n36750_, new_n36751_, new_n36752_, new_n36753_,
    new_n36754_, new_n36755_, new_n36756_, new_n36757_, new_n36758_,
    new_n36759_, new_n36760_, new_n36761_, new_n36762_, new_n36763_,
    new_n36764_, new_n36765_, new_n36766_, new_n36767_, new_n36768_,
    new_n36769_, new_n36770_, new_n36771_, new_n36772_, new_n36773_,
    new_n36774_, new_n36775_, new_n36776_, new_n36777_, new_n36778_,
    new_n36779_, new_n36780_, new_n36781_, new_n36782_, new_n36783_,
    new_n36784_, new_n36785_, new_n36787_, new_n36788_, new_n36789_,
    new_n36790_, new_n36791_, new_n36792_, new_n36793_, new_n36794_,
    new_n36795_, new_n36796_, new_n36797_, new_n36798_, new_n36799_,
    new_n36800_, new_n36801_, new_n36802_, new_n36803_, new_n36805_,
    new_n36806_, new_n36807_, new_n36808_, new_n36809_, new_n36810_,
    new_n36811_, new_n36812_, new_n36813_, new_n36814_, new_n36815_,
    new_n36816_, new_n36817_, new_n36818_, new_n36819_, new_n36820_,
    new_n36821_, new_n36822_, new_n36823_, new_n36824_, new_n36825_,
    new_n36826_, new_n36827_, new_n36828_, new_n36829_, new_n36830_,
    new_n36831_, new_n36832_, new_n36833_, new_n36834_, new_n36835_,
    new_n36836_, new_n36837_, new_n36838_, new_n36839_, new_n36840_,
    new_n36841_, new_n36842_, new_n36843_, new_n36844_, new_n36845_,
    new_n36846_, new_n36847_, new_n36848_, new_n36849_, new_n36850_,
    new_n36851_, new_n36852_, new_n36853_, new_n36854_, new_n36855_,
    new_n36856_, new_n36857_, new_n36858_, new_n36859_, new_n36860_,
    new_n36861_, new_n36862_, new_n36863_, new_n36864_, new_n36865_,
    new_n36866_, new_n36867_, new_n36868_, new_n36869_, new_n36870_,
    new_n36871_, new_n36872_, new_n36873_, new_n36874_, new_n36875_,
    new_n36876_, new_n36877_, new_n36878_, new_n36879_, new_n36880_,
    new_n36881_, new_n36882_, new_n36883_, new_n36884_, new_n36885_,
    new_n36886_, new_n36887_, new_n36888_, new_n36889_, new_n36890_,
    new_n36891_, new_n36892_, new_n36893_, new_n36894_, new_n36897_,
    new_n36898_, new_n36899_, new_n36901_, new_n36902_, new_n36903_,
    new_n36904_, new_n36905_, new_n36907_, new_n36908_, new_n36910_,
    new_n36911_, new_n36912_, new_n36913_, new_n36914_, new_n36916_,
    new_n36917_, new_n36919_, new_n36920_, new_n36922_, new_n36923_,
    new_n36924_, new_n36926_, new_n36927_, new_n36928_, new_n36929_,
    new_n36931_, new_n36932_, new_n36933_, new_n36934_, new_n36935_,
    new_n36936_, new_n36937_, new_n36938_, new_n36940_, new_n36941_,
    new_n36942_, new_n36943_, new_n36944_, new_n36945_, new_n36947_,
    new_n36948_, new_n36950_, new_n36951_, new_n36952_, new_n36953_,
    new_n36954_, new_n36957_, new_n36958_, new_n36959_, new_n36960_,
    new_n36962_, new_n36963_, new_n36964_, new_n36966_, new_n36967_,
    new_n36968_, new_n36970_, new_n36971_, new_n36972_, new_n36973_,
    new_n36975_, new_n36976_, new_n36977_, new_n36978_, new_n36980_,
    new_n36981_, new_n36982_, new_n36984_, new_n36985_, new_n36986_,
    new_n36987_, new_n36989_, new_n36990_, new_n36991_, new_n36993_,
    new_n36994_, new_n36995_, new_n36996_, new_n36997_, new_n36999_,
    new_n37000_, new_n37002_, new_n37003_, new_n37004_, new_n37005_,
    new_n37007_, new_n37008_, new_n37009_, new_n37011_, new_n37012_,
    new_n37013_, new_n37015_, new_n37016_, new_n37017_, new_n37018_,
    new_n37020_, new_n37021_, new_n37022_, new_n37024_, new_n37025_,
    new_n37026_, new_n37028_, new_n37029_, new_n37030_, new_n37032_,
    new_n37033_, new_n37034_, new_n37035_, new_n37036_, new_n37038_,
    new_n37039_, new_n37040_, new_n37041_, new_n37042_, new_n37044_,
    new_n37045_, new_n37046_, new_n37048_, new_n37049_, new_n37050_,
    new_n37052_, new_n37053_, new_n37055_, new_n37056_, new_n37057_,
    new_n37059_, new_n37060_, new_n37062_, new_n37063_, new_n37064_,
    new_n37066_, new_n37067_, new_n37068_, new_n37070_, new_n37071_,
    new_n37072_, new_n37074_, new_n37075_, new_n37076_, new_n37078_,
    new_n37079_, new_n37081_, new_n37082_, new_n37083_, new_n37085_,
    new_n37086_, new_n37087_, new_n37088_, new_n37090_, new_n37091_,
    new_n37093_, new_n37094_, new_n37096_, new_n37097_, new_n37099_,
    new_n37100_, new_n37101_, new_n37102_, new_n37104_, new_n37105_,
    new_n37107_, new_n37108_, new_n37109_, new_n37111_, new_n37112_,
    new_n37114_, new_n37115_, new_n37116_, new_n37118_, new_n37119_,
    new_n37120_, new_n37121_, new_n37123_, new_n37124_, new_n37125_,
    new_n37127_, new_n37128_, new_n37130_, new_n37131_, new_n37133_,
    new_n37134_, new_n37135_, new_n37136_, new_n37138_, new_n37139_,
    new_n37140_, new_n37142_, new_n37143_, new_n37144_, new_n37145_,
    new_n37147_, new_n37148_, new_n37149_, new_n37150_, new_n37152_,
    new_n37153_, new_n37154_, new_n37155_, new_n37157_, new_n37158_,
    new_n37159_, new_n37161_, new_n37162_, new_n37163_, new_n37164_,
    new_n37166_, new_n37167_, new_n37168_, new_n37170_, new_n37171_,
    new_n37172_, new_n37174_, new_n37175_, new_n37176_, new_n37178_,
    new_n37179_, new_n37180_, new_n37181_, new_n37182_, new_n37183_,
    new_n37184_, new_n37185_, new_n37187_, new_n37188_, new_n37190_,
    new_n37191_, new_n37192_, new_n37194_, new_n37195_, new_n37196_,
    new_n37198_, new_n37199_, new_n37200_, new_n37201_, new_n37202_,
    new_n37203_, new_n37204_, new_n37205_, new_n37206_, new_n37207_,
    new_n37208_, new_n37209_, new_n37210_, new_n37211_, new_n37212_,
    new_n37213_, new_n37214_, new_n37215_, new_n37216_, new_n37217_,
    new_n37218_, new_n37219_, new_n37220_, new_n37221_, new_n37222_,
    new_n37223_, new_n37224_, new_n37225_, new_n37226_, new_n37227_,
    new_n37228_, new_n37229_, new_n37230_, new_n37231_, new_n37232_,
    new_n37234_, new_n37235_, new_n37236_, new_n37237_, new_n37238_,
    new_n37239_, new_n37240_, new_n37241_, new_n37242_, new_n37243_,
    new_n37244_, new_n37245_, new_n37246_, new_n37247_, new_n37248_,
    new_n37249_, new_n37250_, new_n37251_, new_n37252_, new_n37253_,
    new_n37254_, new_n37255_, new_n37256_, new_n37257_, new_n37259_,
    new_n37260_, new_n37262_, new_n37263_, new_n37264_, new_n37265_,
    new_n37266_, new_n37267_, new_n37268_, new_n37269_, new_n37270_,
    new_n37271_, new_n37272_, new_n37273_, new_n37274_, new_n37275_,
    new_n37276_, new_n37277_, new_n37278_, new_n37279_, new_n37280_,
    new_n37281_, new_n37282_, new_n37283_, new_n37285_, new_n37286_,
    new_n37287_, new_n37288_, new_n37289_, new_n37290_, new_n37291_,
    new_n37292_, new_n37293_, new_n37294_, new_n37295_, new_n37296_,
    new_n37297_, new_n37298_, new_n37299_, new_n37300_, new_n37301_,
    new_n37302_, new_n37303_, new_n37305_, new_n37306_, new_n37307_,
    new_n37308_, new_n37309_, new_n37310_, new_n37311_, new_n37312_,
    new_n37313_, new_n37314_, new_n37315_, new_n37316_, new_n37317_,
    new_n37318_, new_n37319_, new_n37320_, new_n37321_, new_n37323_,
    new_n37324_, new_n37325_, new_n37327_, new_n37328_, new_n37329_,
    new_n37330_, new_n37331_, new_n37332_, new_n37333_, new_n37334_,
    new_n37335_, new_n37336_, new_n37337_, new_n37338_, new_n37339_,
    new_n37340_, new_n37341_, new_n37342_, new_n37343_, new_n37344_,
    new_n37345_, new_n37347_, new_n37348_, new_n37349_, new_n37350_,
    new_n37351_, new_n37352_, new_n37353_, new_n37354_, new_n37355_,
    new_n37356_, new_n37357_, new_n37358_, new_n37359_, new_n37360_,
    new_n37361_, new_n37362_, new_n37363_, new_n37364_, new_n37365_,
    new_n37367_, new_n37368_, new_n37369_, new_n37370_, new_n37371_,
    new_n37372_, new_n37373_, new_n37374_, new_n37375_, new_n37376_,
    new_n37377_, new_n37378_, new_n37379_, new_n37380_, new_n37381_,
    new_n37382_, new_n37383_, new_n37385_, new_n37386_, new_n37387_,
    new_n37388_, new_n37389_, new_n37390_, new_n37391_, new_n37392_,
    new_n37393_, new_n37394_, new_n37395_, new_n37396_, new_n37397_,
    new_n37398_, new_n37399_, new_n37400_, new_n37401_, new_n37403_,
    new_n37404_, new_n37405_, new_n37406_, new_n37407_, new_n37408_,
    new_n37409_, new_n37410_, new_n37411_, new_n37412_, new_n37413_,
    new_n37414_, new_n37415_, new_n37416_, new_n37417_, new_n37418_,
    new_n37419_, new_n37420_, new_n37421_, new_n37422_, new_n37423_,
    new_n37424_, new_n37426_, new_n37427_, new_n37428_, new_n37429_,
    new_n37430_, new_n37431_, new_n37432_, new_n37433_, new_n37434_,
    new_n37438_, new_n37439_, new_n37440_, new_n37441_, new_n37442_,
    new_n37443_, new_n37445_, new_n37446_, new_n37447_, new_n37448_,
    new_n37449_, new_n37450_, new_n37451_, new_n37452_, new_n37453_,
    new_n37454_, new_n37455_, new_n37456_, new_n37457_, new_n37458_,
    new_n37459_, new_n37460_, new_n37461_, new_n37462_, new_n37464_,
    new_n37465_, new_n37466_, new_n37467_, new_n37468_, new_n37469_,
    new_n37470_, new_n37471_, new_n37472_, new_n37473_, new_n37474_,
    new_n37475_, new_n37476_, new_n37477_, new_n37478_, new_n37479_,
    new_n37480_, new_n37481_, new_n37482_, new_n37484_, new_n37485_,
    new_n37486_, new_n37487_, new_n37488_, new_n37489_, new_n37490_,
    new_n37491_, new_n37492_, new_n37493_, new_n37494_, new_n37495_,
    new_n37496_, new_n37497_, new_n37498_, new_n37499_, new_n37500_,
    new_n37502_, new_n37503_, new_n37504_, new_n37505_, new_n37506_,
    new_n37507_, new_n37508_, new_n37509_, new_n37510_, new_n37511_,
    new_n37512_, new_n37513_, new_n37514_, new_n37515_, new_n37516_,
    new_n37517_, new_n37518_, new_n37519_, new_n37520_, new_n37522_,
    new_n37523_, new_n37524_, new_n37526_, new_n37527_, new_n37529_,
    new_n37530_, new_n37531_, new_n37532_, new_n37533_, new_n37534_,
    new_n37535_, new_n37536_, new_n37537_, new_n37538_, new_n37539_,
    new_n37540_, new_n37541_, new_n37542_, new_n37543_, new_n37544_,
    new_n37545_, new_n37547_, new_n37548_, new_n37550_, new_n37551_,
    new_n37553_, new_n37554_, new_n37555_, new_n37556_, new_n37557_,
    new_n37558_, new_n37559_, new_n37560_, new_n37561_, new_n37562_,
    new_n37563_, new_n37564_, new_n37565_, new_n37566_, new_n37567_,
    new_n37568_, new_n37569_, new_n37570_, new_n37571_, new_n37572_,
    new_n37573_, new_n37574_, new_n37575_, new_n37576_, new_n37577_,
    new_n37578_, new_n37579_, new_n37580_, new_n37582_, new_n37583_,
    new_n37585_, new_n37586_, new_n37588_, new_n37589_, new_n37591_,
    new_n37592_, new_n37593_, new_n37594_, new_n37595_, new_n37596_,
    new_n37597_, new_n37598_, new_n37599_, new_n37600_, new_n37601_,
    new_n37602_, new_n37603_, new_n37604_, new_n37605_, new_n37606_,
    new_n37607_, new_n37608_, new_n37610_, new_n37611_, new_n37613_,
    new_n37614_, new_n37616_, new_n37617_, new_n37618_, new_n37619_,
    new_n37620_, new_n37621_, new_n37622_, new_n37623_, new_n37624_,
    new_n37625_, new_n37626_, new_n37627_, new_n37628_, new_n37629_,
    new_n37630_, new_n37631_, new_n37632_, new_n37633_, new_n37634_,
    new_n37635_, new_n37637_, new_n37638_, new_n37639_, new_n37641_,
    new_n37642_, new_n37643_, new_n37645_, new_n37646_, new_n37648_,
    new_n37649_, new_n37651_, new_n37652_, new_n37653_, new_n37655_,
    new_n37656_, new_n37658_, new_n37659_, new_n37661_, new_n37662_,
    new_n37664_, new_n37665_, new_n37667_, new_n37668_, new_n37670_,
    new_n37671_, new_n37673_, new_n37674_, new_n37676_, new_n37677_,
    new_n37679_, new_n37680_, new_n37682_, new_n37683_, new_n37684_,
    new_n37685_, new_n37686_, new_n37692_, new_n37693_, new_n37694_,
    new_n37695_, new_n37696_, new_n37697_, new_n37698_, new_n37699_,
    new_n37700_, new_n37701_, new_n37702_, new_n37703_, new_n37705_,
    new_n37706_, new_n37707_, new_n37708_, new_n37709_, new_n37710_,
    new_n37711_, new_n37712_, new_n37713_, new_n37714_, new_n37715_,
    new_n37716_, new_n37717_, new_n37718_, new_n37719_, new_n37720_,
    new_n37721_, new_n37722_, new_n37723_, new_n37724_, new_n37725_,
    new_n37726_, new_n37727_, new_n37728_, new_n37730_, new_n37731_,
    new_n37733_, new_n37734_, new_n37736_, new_n37737_, new_n37738_,
    new_n37739_, new_n37740_, new_n37746_, new_n37747_, new_n37748_,
    new_n37749_, new_n37750_, new_n37751_, new_n37752_, new_n37753_,
    new_n37754_, new_n37756_, new_n37757_, new_n37758_, new_n37759_,
    new_n37760_, new_n37761_, new_n37762_, new_n37763_, new_n37764_,
    new_n37765_, new_n37766_, new_n37767_, new_n37768_, new_n37769_,
    new_n37770_, new_n37771_, new_n37772_, new_n37773_, new_n37774_,
    new_n37775_, new_n37776_, new_n37778_, new_n37779_, new_n37780_,
    new_n37781_, new_n37782_, new_n37788_, new_n37789_, new_n37790_,
    new_n37791_, new_n37792_, new_n37793_, new_n37794_, new_n37795_,
    new_n37796_, new_n37798_, new_n37799_, new_n37800_, new_n37801_,
    new_n37802_, new_n37803_, new_n37804_, new_n37805_, new_n37806_,
    new_n37807_, new_n37808_, new_n37809_, new_n37810_, new_n37811_,
    new_n37812_, new_n37813_, new_n37814_, new_n37815_, new_n37816_,
    new_n37817_, new_n37818_, new_n37819_, new_n37821_, new_n37822_,
    new_n37824_, new_n37825_, new_n37826_, new_n37827_, new_n37828_,
    new_n37829_, new_n37830_, new_n37831_, new_n37832_, new_n37833_,
    new_n37834_, new_n37835_, new_n37836_, new_n37837_, new_n37838_,
    new_n37839_, new_n37840_, new_n37841_, new_n37842_, new_n37843_,
    new_n37845_, new_n37846_, new_n37847_, new_n37848_, new_n37849_,
    new_n37850_, new_n37851_, new_n37852_, new_n37853_, new_n37854_,
    new_n37855_, new_n37856_, new_n37857_, new_n37858_, new_n37859_,
    new_n37860_, new_n37861_, new_n37862_, new_n37863_, new_n37864_,
    new_n37865_, new_n37867_, new_n37868_, new_n37869_, new_n37870_,
    new_n37871_, new_n37872_, new_n37873_, new_n37874_, new_n37875_,
    new_n37876_, new_n37877_, new_n37878_, new_n37879_, new_n37880_,
    new_n37881_, new_n37882_, new_n37883_, new_n37884_, new_n37885_,
    new_n37886_, new_n37888_, new_n37889_, new_n37890_, new_n37891_,
    new_n37892_, new_n37893_, new_n37894_, new_n37895_, new_n37896_,
    new_n37897_, new_n37898_, new_n37899_, new_n37900_, new_n37901_,
    new_n37902_, new_n37903_, new_n37904_, new_n37905_, new_n37907_,
    new_n37908_, new_n37909_, new_n37910_, new_n37911_, new_n37912_,
    new_n37913_, new_n37914_, new_n37915_, new_n37916_, new_n37917_,
    new_n37918_, new_n37919_, new_n37920_, new_n37921_, new_n37922_,
    new_n37923_, new_n37924_, new_n37925_, new_n37926_, new_n37927_,
    new_n37929_, new_n37930_, new_n37931_, new_n37932_, new_n37933_,
    new_n37934_, new_n37935_, new_n37936_, new_n37937_, new_n37938_,
    new_n37939_, new_n37940_, new_n37941_, new_n37942_, new_n37943_,
    new_n37944_, new_n37945_, new_n37946_, new_n37947_, new_n37948_,
    new_n37949_, new_n37950_, new_n37951_, new_n37952_, new_n37953_,
    new_n37954_, new_n37955_, new_n37956_, new_n37957_, new_n37958_,
    new_n37959_, new_n37960_, new_n37961_, new_n37962_, new_n37963_,
    new_n37964_, new_n37965_, new_n37966_, new_n37967_, new_n37968_,
    new_n37969_, new_n37970_, new_n37971_, new_n37972_, new_n37973_,
    new_n37974_, new_n37975_, new_n37976_, new_n37977_, new_n37978_,
    new_n37979_, new_n37980_, new_n37981_, new_n37982_, new_n37983_,
    new_n37985_, new_n37986_, new_n37987_, new_n37988_, new_n37989_,
    new_n37990_, new_n37991_, new_n37992_, new_n37993_, new_n37994_,
    new_n37995_, new_n37996_, new_n37997_, new_n37998_, new_n38003_,
    new_n38004_, new_n38005_, new_n38006_, new_n38007_, new_n38008_,
    new_n38010_, new_n38011_, new_n38013_, new_n38014_, new_n38016_,
    new_n38017_, new_n38019_, new_n38020_, new_n38022_, new_n38023_,
    new_n38025_, new_n38026_, new_n38027_, new_n38029_, new_n38030_,
    new_n38032_, new_n38033_, new_n38035_, new_n38036_, new_n38037_,
    new_n38038_, new_n38039_, new_n38040_, new_n38041_, new_n38042_,
    new_n38043_, new_n38044_, new_n38045_, new_n38046_, new_n38047_,
    new_n38048_, new_n38049_, new_n38050_, new_n38051_, new_n38053_,
    new_n38054_, new_n38056_, new_n38057_, new_n38058_, new_n38059_,
    new_n38060_, new_n38061_, new_n38062_, new_n38063_, new_n38064_,
    new_n38065_, new_n38066_, new_n38067_, new_n38068_, new_n38069_,
    new_n38070_, new_n38071_, new_n38072_, new_n38073_, new_n38074_,
    new_n38075_, new_n38077_, new_n38078_, new_n38080_, new_n38081_,
    new_n38083_, new_n38084_, new_n38086_, new_n38087_, new_n38089_,
    new_n38090_, new_n38092_, new_n38093_, new_n38095_, new_n38096_,
    new_n38098_, new_n38099_, new_n38101_, new_n38102_, new_n38104_,
    new_n38105_, new_n38107_, new_n38108_, new_n38110_, new_n38111_,
    new_n38113_, new_n38114_, new_n38116_, new_n38117_, new_n38118_,
    new_n38119_, new_n38120_, new_n38121_, new_n38122_, new_n38123_,
    new_n38124_, new_n38126_, new_n38127_, new_n38129_, new_n38130_,
    new_n38132_, new_n38133_, new_n38135_, new_n38136_, new_n38138_,
    new_n38139_, new_n38141_, new_n38142_, new_n38144_, new_n38145_,
    new_n38147_, new_n38148_, new_n38150_, new_n38151_, new_n38153_,
    new_n38154_, new_n38156_, new_n38157_, new_n38159_, new_n38161_,
    new_n38162_, new_n38164_, new_n38165_, new_n38167_, new_n38168_,
    new_n38170_, new_n38171_, new_n38173_, new_n38174_, new_n38176_,
    new_n38178_, new_n38179_, new_n38180_, new_n38181_, new_n38182_,
    new_n38183_, new_n38184_, new_n38185_, new_n38186_, new_n38187_,
    new_n38188_, new_n38189_, new_n38190_, new_n38191_, new_n38192_,
    new_n38193_, new_n38194_, new_n38195_, new_n38196_, new_n38198_,
    new_n38199_, new_n38201_, new_n38202_, new_n38204_, new_n38205_,
    new_n38207_, new_n38208_, new_n38209_, new_n38210_, new_n38211_,
    new_n38212_, new_n38213_, new_n38214_, new_n38215_, new_n38216_,
    new_n38217_, new_n38219_, new_n38220_, new_n38222_, new_n38223_,
    new_n38224_, new_n38226_, new_n38227_, new_n38228_, new_n38230_,
    new_n38231_, new_n38233_, new_n38234_, new_n38235_, new_n38236_,
    new_n38238_, new_n38239_, new_n38241_, new_n38242_, new_n38243_,
    new_n38244_, new_n38245_, new_n38246_, new_n38247_, new_n38248_,
    new_n38250_, new_n38251_, new_n38252_, new_n38254_, new_n38255_,
    new_n38257_, new_n38258_, new_n38259_, new_n38260_, new_n38264_,
    new_n38266_, new_n38268_, new_n38270_, new_n38271_, new_n38273_,
    new_n38275_, new_n38277_, new_n38279_, new_n38281_, new_n38283_,
    new_n38285_, new_n38286_, new_n38288_, new_n38290_, new_n38291_,
    new_n38292_, new_n38294_, new_n38296_, new_n38297_, new_n38299_,
    new_n38300_, new_n38302_, new_n38304_, new_n38306_, new_n38309_,
    new_n38311_, new_n38313_, new_n38314_, new_n38316_, new_n38318_,
    new_n38319_, new_n38321_, new_n38323_, new_n38325_, new_n38327_,
    new_n38329_, new_n38331_, new_n38333_, new_n38335_, new_n38339_,
    new_n38340_, new_n38342_, new_n38345_, new_n38346_, new_n38348_,
    new_n38349_, new_n38350_, new_n38351_, new_n38352_, new_n38353_,
    new_n38354_, new_n38355_, new_n38356_, new_n38357_, new_n38358_,
    new_n38359_, new_n38360_, new_n38361_, new_n38363_, new_n38364_,
    new_n38365_, new_n38366_, new_n38367_, new_n38368_, new_n38369_,
    new_n38370_, new_n38371_, new_n38372_, new_n38373_, new_n38374_,
    new_n38376_, new_n38377_, new_n38378_, new_n38379_, new_n38380_,
    new_n38381_, new_n38382_, new_n38383_, new_n38384_, new_n38385_,
    new_n38386_, new_n38387_, new_n38389_, new_n38390_, new_n38391_,
    new_n38392_, new_n38393_, new_n38394_, new_n38395_, new_n38396_,
    new_n38397_, new_n38398_, new_n38399_, new_n38400_, new_n38402_,
    new_n38406_, new_n38407_, new_n38409_, new_n38412_, new_n38414_,
    new_n38416_, new_n38418_, new_n38420_, new_n38422_, new_n38424_,
    new_n38426_, new_n38428_, new_n38430_, new_n38432_, new_n38434_,
    new_n38436_, new_n38438_, new_n38440_, new_n38442_, new_n38444_,
    new_n38446_, new_n38448_, new_n38450_, new_n38452_, new_n38454_,
    new_n38456_, new_n38458_, new_n38460_, new_n38461_, new_n38462_,
    new_n38463_, new_n38464_, new_n38465_, new_n38467_, new_n38469_,
    new_n38471_, new_n38473_, new_n38475_, new_n38477_, new_n38479_,
    new_n38481_, new_n38482_, new_n38483_, new_n38484_, new_n38486_,
    new_n38488_, new_n38490_, new_n38492_, new_n38494_, new_n38496_,
    new_n38497_, new_n38498_, new_n38499_, new_n38501_, new_n38503_,
    new_n38504_, new_n38505_, new_n38506_, new_n38508_, new_n38509_,
    new_n38510_, new_n38511_, new_n38513_, new_n38514_, new_n38515_,
    new_n38516_, new_n38518_, new_n38520_, new_n38523_, new_n38526_,
    new_n38529_, new_n38532_, new_n38535_, new_n38538_, new_n38541_,
    new_n38544_, new_n38547_, new_n38550_, new_n38554_, new_n38557_,
    new_n38560_, new_n38563_, new_n38566_, new_n38569_, new_n38572_,
    new_n38575_, new_n38578_, new_n38581_, new_n38584_, new_n38586_,
    new_n38587_, new_n38588_, new_n38589_, new_n38590_, new_n38591_,
    new_n38592_, new_n38593_, new_n38596_, new_n38599_, new_n38602_,
    new_n38605_, new_n38608_, new_n38611_, new_n38613_, new_n38616_,
    new_n38619_, new_n38622_, new_n38625_, new_n38628_, new_n38630_,
    new_n38632_, new_n38634_, new_n38636_, new_n38639_, new_n38641_,
    new_n38643_, new_n38645_, new_n38647_, new_n38649_, new_n38651_,
    new_n38653_, new_n38655_, new_n38657_, new_n38659_, new_n38661_,
    new_n38663_, new_n38665_, new_n38667_, new_n38669_, new_n38671_,
    new_n38673_, new_n38675_, new_n38677_, new_n38682_;
  INV_X1     g00000(.I(pi0095), .ZN(new_n2436_));
  INV_X1     g00001(.I(pi0072), .ZN(new_n2437_));
  NAND4_X1   g00002(.A1(pi0061), .A2(pi0076), .A3(pi0085), .A4(pi0106), .ZN(new_n2438_));
  NAND3_X1   g00003(.A1(pi0048), .A2(pi0049), .A3(pi0089), .ZN(new_n2439_));
  NOR2_X1    g00004(.A1(new_n2438_), .A2(new_n2439_), .ZN(new_n2440_));
  NAND3_X1   g00005(.A1(pi0036), .A2(pi0068), .A3(pi0084), .ZN(new_n2441_));
  NAND2_X1   g00006(.A1(pi0045), .A2(pi0104), .ZN(new_n2442_));
  NOR4_X1    g00007(.A1(new_n2441_), .A2(pi0082), .A3(new_n2442_), .A4(pi0111), .ZN(new_n2443_));
  NOR2_X1    g00008(.A1(pi0067), .A2(pi0069), .ZN(new_n2444_));
  NOR2_X1    g00009(.A1(pi0066), .A2(pi0073), .ZN(new_n2445_));
  NOR2_X1    g00010(.A1(pi0083), .A2(pi0103), .ZN(new_n2446_));
  AND3_X2    g00011(.A1(new_n2444_), .A2(new_n2445_), .A3(new_n2446_), .Z(new_n2447_));
  OR2_X2     g00012(.A1(pi0063), .A2(pi0107), .Z(new_n2448_));
  INV_X1     g00013(.I(pi0065), .ZN(new_n2449_));
  INV_X1     g00014(.I(pi0071), .ZN(new_n2450_));
  NAND3_X1   g00015(.A1(new_n2449_), .A2(new_n2450_), .A3(pi0064), .ZN(new_n2451_));
  NOR2_X1    g00016(.A1(new_n2451_), .A2(new_n2448_), .ZN(new_n2452_));
  NAND4_X1   g00017(.A1(new_n2447_), .A2(new_n2452_), .A3(new_n2443_), .A4(new_n2440_), .ZN(new_n2453_));
  INV_X1     g00018(.I(pi0102), .ZN(new_n2454_));
  OR3_X2     g00019(.A1(pi0077), .A2(pi0088), .A3(pi0098), .Z(new_n2455_));
  NOR2_X1    g00020(.A1(new_n2455_), .A2(pi0050), .ZN(new_n2456_));
  NAND2_X1   g00021(.A1(new_n2456_), .A2(new_n2454_), .ZN(new_n2457_));
  NOR3_X1    g00022(.A1(new_n2453_), .A2(pi0081), .A3(new_n2457_), .ZN(new_n2458_));
  INV_X1     g00023(.I(new_n2458_), .ZN(new_n2459_));
  OR3_X2     g00024(.A1(pi0053), .A2(pi0060), .A3(pi0086), .Z(new_n2460_));
  INV_X1     g00025(.I(pi0097), .ZN(new_n2461_));
  INV_X1     g00026(.I(pi0108), .ZN(new_n2462_));
  NAND4_X1   g00027(.A1(new_n2461_), .A2(new_n2462_), .A3(pi0046), .A4(pi0094), .ZN(new_n2463_));
  NOR2_X1    g00028(.A1(new_n2463_), .A2(new_n2460_), .ZN(new_n2464_));
  INV_X1     g00029(.I(new_n2464_), .ZN(new_n2465_));
  NOR2_X1    g00030(.A1(new_n2459_), .A2(new_n2465_), .ZN(new_n2466_));
  INV_X1     g00031(.I(new_n2466_), .ZN(new_n2467_));
  NOR2_X1    g00032(.A1(pi0058), .A2(pi0091), .ZN(new_n2468_));
  NAND4_X1   g00033(.A1(new_n2468_), .A2(pi0047), .A3(pi0109), .A4(pi0110), .ZN(new_n2469_));
  NOR2_X1    g00034(.A1(new_n2467_), .A2(new_n2469_), .ZN(new_n2470_));
  INV_X1     g00035(.I(new_n2470_), .ZN(new_n2471_));
  NOR2_X1    g00036(.A1(pi0070), .A2(pi0096), .ZN(new_n2472_));
  INV_X1     g00037(.I(new_n2472_), .ZN(new_n2473_));
  NOR2_X1    g00038(.A1(pi0035), .A2(pi0051), .ZN(new_n2474_));
  INV_X1     g00039(.I(new_n2474_), .ZN(new_n2475_));
  NOR2_X1    g00040(.A1(new_n2473_), .A2(new_n2475_), .ZN(new_n2476_));
  INV_X1     g00041(.I(new_n2476_), .ZN(new_n2477_));
  NOR2_X1    g00042(.A1(pi0090), .A2(pi0093), .ZN(new_n2478_));
  INV_X1     g00043(.I(new_n2478_), .ZN(new_n2479_));
  NOR2_X1    g00044(.A1(new_n2477_), .A2(new_n2479_), .ZN(new_n2480_));
  INV_X1     g00045(.I(new_n2480_), .ZN(new_n2481_));
  NOR2_X1    g00046(.A1(new_n2471_), .A2(new_n2481_), .ZN(new_n2482_));
  NOR2_X1    g00047(.A1(new_n2482_), .A2(new_n2437_), .ZN(new_n2483_));
  NOR2_X1    g00048(.A1(new_n2483_), .A2(pi0040), .ZN(new_n2484_));
  INV_X1     g00049(.I(new_n2484_), .ZN(new_n2485_));
  INV_X1     g00050(.I(pi0040), .ZN(new_n2486_));
  NOR2_X1    g00051(.A1(pi0058), .A2(pi0090), .ZN(new_n2487_));
  NOR2_X1    g00052(.A1(pi0109), .A2(pi0110), .ZN(new_n2488_));
  INV_X1     g00053(.I(new_n2488_), .ZN(new_n2489_));
  OR2_X2     g00054(.A1(pi0047), .A2(pi0091), .Z(new_n2490_));
  NOR4_X1    g00055(.A1(new_n2463_), .A2(new_n2460_), .A3(new_n2489_), .A4(new_n2490_), .ZN(new_n2491_));
  INV_X1     g00056(.I(pi0081), .ZN(new_n2492_));
  NOR4_X1    g00057(.A1(new_n2455_), .A2(pi0050), .A3(new_n2492_), .A4(pi0102), .ZN(new_n2493_));
  NAND2_X1   g00058(.A1(new_n2491_), .A2(new_n2493_), .ZN(new_n2494_));
  NOR2_X1    g00059(.A1(new_n2494_), .A2(new_n2453_), .ZN(new_n2495_));
  NOR2_X1    g00060(.A1(pi0035), .A2(pi0093), .ZN(new_n2496_));
  NOR2_X1    g00061(.A1(pi0072), .A2(pi0096), .ZN(new_n2497_));
  NOR2_X1    g00062(.A1(pi0051), .A2(pi0070), .ZN(new_n2498_));
  NAND2_X1   g00063(.A1(new_n2497_), .A2(new_n2498_), .ZN(new_n2499_));
  INV_X1     g00064(.I(new_n2499_), .ZN(new_n2500_));
  NAND4_X1   g00065(.A1(new_n2495_), .A2(new_n2487_), .A3(new_n2496_), .A4(new_n2500_), .ZN(new_n2501_));
  NOR2_X1    g00066(.A1(new_n2501_), .A2(new_n2486_), .ZN(new_n2502_));
  NOR2_X1    g00067(.A1(new_n2502_), .A2(pi0032), .ZN(new_n2503_));
  INV_X1     g00068(.I(new_n2503_), .ZN(new_n2504_));
  NOR2_X1    g00069(.A1(new_n2485_), .A2(new_n2504_), .ZN(new_n2505_));
  NOR2_X1    g00070(.A1(new_n2505_), .A2(pi0072), .ZN(new_n2506_));
  NAND2_X1   g00071(.A1(new_n2495_), .A2(new_n2487_), .ZN(new_n2507_));
  INV_X1     g00072(.I(new_n2507_), .ZN(new_n2508_));
  INV_X1     g00073(.I(pi0093), .ZN(new_n2509_));
  NOR2_X1    g00074(.A1(pi0047), .A2(pi0110), .ZN(new_n2510_));
  NAND2_X1   g00075(.A1(new_n2510_), .A2(pi0109), .ZN(new_n2511_));
  INV_X1     g00076(.I(new_n2510_), .ZN(new_n2512_));
  NOR2_X1    g00077(.A1(pi0088), .A2(pi0098), .ZN(new_n2513_));
  NOR2_X1    g00078(.A1(new_n2453_), .A2(new_n2492_), .ZN(new_n2514_));
  NAND3_X1   g00079(.A1(new_n2514_), .A2(pi0102), .A3(new_n2513_), .ZN(new_n2515_));
  NOR2_X1    g00080(.A1(pi0086), .A2(pi0094), .ZN(new_n2516_));
  INV_X1     g00081(.I(pi0050), .ZN(new_n2517_));
  INV_X1     g00082(.I(pi0053), .ZN(new_n2518_));
  INV_X1     g00083(.I(pi0060), .ZN(new_n2519_));
  NAND3_X1   g00084(.A1(new_n2517_), .A2(new_n2518_), .A3(new_n2519_), .ZN(new_n2520_));
  NOR2_X1    g00085(.A1(new_n2520_), .A2(pi0077), .ZN(new_n2521_));
  NAND2_X1   g00086(.A1(new_n2521_), .A2(new_n2516_), .ZN(new_n2522_));
  NOR2_X1    g00087(.A1(new_n2515_), .A2(new_n2522_), .ZN(new_n2523_));
  NOR2_X1    g00088(.A1(new_n2523_), .A2(new_n2461_), .ZN(new_n2524_));
  AOI21_X1   g00089(.A1(new_n2523_), .A2(new_n2461_), .B(new_n2462_), .ZN(new_n2525_));
  NOR2_X1    g00090(.A1(new_n2525_), .A2(pi0046), .ZN(new_n2526_));
  INV_X1     g00091(.I(new_n2526_), .ZN(new_n2527_));
  NOR2_X1    g00092(.A1(new_n2527_), .A2(new_n2462_), .ZN(new_n2528_));
  INV_X1     g00093(.I(new_n2528_), .ZN(new_n2529_));
  INV_X1     g00094(.I(pi0094), .ZN(new_n2530_));
  AND4_X2    g00095(.A1(pi0061), .A2(pi0076), .A3(pi0085), .A4(pi0106), .Z(new_n2531_));
  AND3_X2    g00096(.A1(pi0048), .A2(pi0049), .A3(pi0089), .Z(new_n2532_));
  NAND2_X1   g00097(.A1(new_n2531_), .A2(new_n2532_), .ZN(new_n2533_));
  NOR2_X1    g00098(.A1(pi0082), .A2(pi0111), .ZN(new_n2534_));
  AND3_X2    g00099(.A1(pi0036), .A2(pi0068), .A3(pi0084), .Z(new_n2535_));
  AND2_X2    g00100(.A1(pi0045), .A2(pi0104), .Z(new_n2536_));
  NAND3_X1   g00101(.A1(new_n2535_), .A2(new_n2536_), .A3(new_n2534_), .ZN(new_n2537_));
  NAND3_X1   g00102(.A1(new_n2444_), .A2(new_n2445_), .A3(new_n2446_), .ZN(new_n2538_));
  NOR2_X1    g00103(.A1(pi0063), .A2(pi0107), .ZN(new_n2539_));
  NOR2_X1    g00104(.A1(pi0065), .A2(pi0071), .ZN(new_n2540_));
  NAND3_X1   g00105(.A1(new_n2539_), .A2(new_n2540_), .A3(pi0064), .ZN(new_n2541_));
  NOR4_X1    g00106(.A1(new_n2533_), .A2(new_n2537_), .A3(new_n2538_), .A4(new_n2541_), .ZN(new_n2542_));
  NOR2_X1    g00107(.A1(pi0081), .A2(pi0102), .ZN(new_n2543_));
  NAND2_X1   g00108(.A1(new_n2542_), .A2(new_n2543_), .ZN(new_n2544_));
  NOR2_X1    g00109(.A1(new_n2544_), .A2(new_n2455_), .ZN(new_n2545_));
  INV_X1     g00110(.I(new_n2545_), .ZN(new_n2546_));
  NOR2_X1    g00111(.A1(new_n2546_), .A2(new_n2520_), .ZN(new_n2547_));
  INV_X1     g00112(.I(new_n2547_), .ZN(new_n2548_));
  NOR3_X1    g00113(.A1(new_n2548_), .A2(pi0086), .A3(new_n2530_), .ZN(new_n2549_));
  NOR2_X1    g00114(.A1(new_n2549_), .A2(pi0097), .ZN(new_n2550_));
  INV_X1     g00115(.I(new_n2550_), .ZN(new_n2551_));
  AOI21_X1   g00116(.A1(new_n2546_), .A2(pi0050), .B(pi0060), .ZN(new_n2552_));
  INV_X1     g00117(.I(pi0077), .ZN(new_n2553_));
  NOR2_X1    g00118(.A1(new_n2515_), .A2(new_n2553_), .ZN(new_n2554_));
  NOR2_X1    g00119(.A1(new_n2554_), .A2(pi0050), .ZN(new_n2555_));
  INV_X1     g00120(.I(new_n2555_), .ZN(new_n2556_));
  INV_X1     g00121(.I(new_n2544_), .ZN(new_n2557_));
  INV_X1     g00122(.I(pi0098), .ZN(new_n2558_));
  AOI21_X1   g00123(.A1(pi0077), .A2(pi0098), .B(pi0088), .ZN(new_n2559_));
  AOI21_X1   g00124(.A1(new_n2553_), .A2(new_n2558_), .B(new_n2559_), .ZN(new_n2560_));
  NAND2_X1   g00125(.A1(new_n2557_), .A2(new_n2560_), .ZN(new_n2561_));
  INV_X1     g00126(.I(new_n2543_), .ZN(new_n2562_));
  NOR2_X1    g00127(.A1(new_n2492_), .A2(new_n2454_), .ZN(new_n2563_));
  OAI21_X1   g00128(.A1(new_n2453_), .A2(new_n2563_), .B(new_n2562_), .ZN(new_n2564_));
  INV_X1     g00129(.I(pi0107), .ZN(new_n2565_));
  NOR2_X1    g00130(.A1(new_n2533_), .A2(new_n2537_), .ZN(new_n2566_));
  INV_X1     g00131(.I(new_n2566_), .ZN(new_n2567_));
  NOR2_X1    g00132(.A1(new_n2567_), .A2(new_n2538_), .ZN(new_n2568_));
  INV_X1     g00133(.I(new_n2568_), .ZN(new_n2569_));
  AOI21_X1   g00134(.A1(new_n2569_), .A2(pi0071), .B(pi0065), .ZN(new_n2570_));
  INV_X1     g00135(.I(pi0066), .ZN(new_n2571_));
  INV_X1     g00136(.I(pi0045), .ZN(new_n2572_));
  NOR2_X1    g00137(.A1(new_n2438_), .A2(pi0048), .ZN(new_n2573_));
  INV_X1     g00138(.I(pi0049), .ZN(new_n2574_));
  INV_X1     g00139(.I(pi0085), .ZN(new_n2575_));
  INV_X1     g00140(.I(pi0106), .ZN(new_n2576_));
  NOR4_X1    g00141(.A1(new_n2575_), .A2(new_n2576_), .A3(pi0061), .A4(pi0076), .ZN(new_n2577_));
  NOR2_X1    g00142(.A1(new_n2577_), .A2(pi0048), .ZN(new_n2578_));
  NOR2_X1    g00143(.A1(new_n2573_), .A2(pi0089), .ZN(new_n2579_));
  NOR4_X1    g00144(.A1(new_n2579_), .A2(new_n2574_), .A3(new_n2531_), .A4(new_n2578_), .ZN(new_n2580_));
  AOI21_X1   g00145(.A1(pi0089), .A2(new_n2573_), .B(new_n2580_), .ZN(new_n2581_));
  XOR2_X1    g00146(.A1(new_n2581_), .A2(new_n2572_), .Z(new_n2582_));
  NOR2_X1    g00147(.A1(new_n2533_), .A2(pi0045), .ZN(new_n2583_));
  XOR2_X1    g00148(.A1(new_n2582_), .A2(new_n2583_), .Z(new_n2584_));
  INV_X1     g00149(.I(pi0104), .ZN(new_n2585_));
  AOI21_X1   g00150(.A1(pi0045), .A2(new_n2585_), .B(new_n2533_), .ZN(new_n2586_));
  NAND2_X1   g00151(.A1(new_n2584_), .A2(new_n2586_), .ZN(new_n2587_));
  NOR2_X1    g00152(.A1(new_n2587_), .A2(new_n2571_), .ZN(new_n2588_));
  NOR3_X1    g00153(.A1(new_n2533_), .A2(pi0045), .A3(pi0104), .ZN(new_n2589_));
  INV_X1     g00154(.I(pi0073), .ZN(new_n2590_));
  NOR2_X1    g00155(.A1(new_n2571_), .A2(new_n2590_), .ZN(new_n2591_));
  INV_X1     g00156(.I(new_n2591_), .ZN(new_n2592_));
  XOR2_X1    g00157(.A1(new_n2587_), .A2(new_n2592_), .Z(new_n2593_));
  NAND2_X1   g00158(.A1(new_n2593_), .A2(new_n2589_), .ZN(new_n2594_));
  NOR2_X1    g00159(.A1(pi0068), .A2(pi0111), .ZN(new_n2595_));
  OAI21_X1   g00160(.A1(new_n2594_), .A2(new_n2588_), .B(new_n2595_), .ZN(new_n2596_));
  AOI21_X1   g00161(.A1(new_n2588_), .A2(new_n2594_), .B(new_n2596_), .ZN(new_n2597_));
  INV_X1     g00162(.I(pi0084), .ZN(new_n2598_));
  NOR3_X1    g00163(.A1(new_n2598_), .A2(pi0068), .A3(pi0111), .ZN(new_n2599_));
  XOR2_X1    g00164(.A1(new_n2597_), .A2(new_n2599_), .Z(new_n2600_));
  INV_X1     g00165(.I(new_n2445_), .ZN(new_n2601_));
  INV_X1     g00166(.I(new_n2589_), .ZN(new_n2602_));
  NOR3_X1    g00167(.A1(new_n2602_), .A2(pi0084), .A3(new_n2601_), .ZN(new_n2603_));
  NAND3_X1   g00168(.A1(new_n2603_), .A2(pi0082), .A3(new_n2595_), .ZN(new_n2604_));
  INV_X1     g00169(.I(pi0036), .ZN(new_n2605_));
  INV_X1     g00170(.I(pi0067), .ZN(new_n2606_));
  NAND2_X1   g00171(.A1(new_n2605_), .A2(new_n2606_), .ZN(new_n2607_));
  NAND2_X1   g00172(.A1(new_n2604_), .A2(new_n2607_), .ZN(new_n2608_));
  NOR2_X1    g00173(.A1(new_n2602_), .A2(new_n2601_), .ZN(new_n2609_));
  INV_X1     g00174(.I(new_n2534_), .ZN(new_n2610_));
  INV_X1     g00175(.I(pi0068), .ZN(new_n2611_));
  NAND2_X1   g00176(.A1(pi0082), .A2(pi0111), .ZN(new_n2612_));
  NAND2_X1   g00177(.A1(new_n2612_), .A2(new_n2611_), .ZN(new_n2613_));
  AND3_X2    g00178(.A1(new_n2603_), .A2(new_n2610_), .A3(new_n2613_), .Z(new_n2614_));
  NAND4_X1   g00179(.A1(new_n2600_), .A2(new_n2608_), .A3(new_n2609_), .A4(new_n2614_), .ZN(new_n2615_));
  NAND2_X1   g00180(.A1(new_n2603_), .A2(new_n2611_), .ZN(new_n2616_));
  INV_X1     g00181(.I(new_n2616_), .ZN(new_n2617_));
  AOI21_X1   g00182(.A1(new_n2617_), .A2(new_n2534_), .B(new_n2605_), .ZN(new_n2618_));
  NOR2_X1    g00183(.A1(new_n2567_), .A2(new_n2601_), .ZN(new_n2619_));
  INV_X1     g00184(.I(new_n2619_), .ZN(new_n2620_));
  AOI21_X1   g00185(.A1(pi0067), .A2(new_n2620_), .B(new_n2618_), .ZN(new_n2621_));
  NAND2_X1   g00186(.A1(new_n2615_), .A2(new_n2621_), .ZN(new_n2622_));
  INV_X1     g00187(.I(pi0069), .ZN(new_n2623_));
  INV_X1     g00188(.I(new_n2444_), .ZN(new_n2624_));
  NOR2_X1    g00189(.A1(new_n2620_), .A2(new_n2624_), .ZN(new_n2625_));
  INV_X1     g00190(.I(new_n2625_), .ZN(new_n2626_));
  AOI21_X1   g00191(.A1(new_n2626_), .A2(pi0083), .B(pi0103), .ZN(new_n2627_));
  INV_X1     g00192(.I(new_n2627_), .ZN(new_n2628_));
  OAI21_X1   g00193(.A1(new_n2628_), .A2(new_n2623_), .B(new_n2620_), .ZN(new_n2629_));
  INV_X1     g00194(.I(pi0083), .ZN(new_n2630_));
  NAND2_X1   g00195(.A1(new_n2623_), .A2(new_n2630_), .ZN(new_n2631_));
  INV_X1     g00196(.I(pi0103), .ZN(new_n2632_));
  NOR2_X1    g00197(.A1(new_n2620_), .A2(new_n2606_), .ZN(new_n2633_));
  INV_X1     g00198(.I(new_n2633_), .ZN(new_n2634_));
  NOR3_X1    g00199(.A1(new_n2634_), .A2(new_n2632_), .A3(new_n2631_), .ZN(new_n2635_));
  INV_X1     g00200(.I(new_n2635_), .ZN(new_n2636_));
  AOI21_X1   g00201(.A1(new_n2636_), .A2(new_n2450_), .B(new_n2631_), .ZN(new_n2637_));
  NAND4_X1   g00202(.A1(new_n2622_), .A2(pi0067), .A3(new_n2629_), .A4(new_n2637_), .ZN(new_n2638_));
  NAND2_X1   g00203(.A1(new_n2638_), .A2(new_n2570_), .ZN(new_n2639_));
  INV_X1     g00204(.I(new_n2540_), .ZN(new_n2640_));
  NOR2_X1    g00205(.A1(new_n2569_), .A2(new_n2640_), .ZN(new_n2641_));
  INV_X1     g00206(.I(new_n2641_), .ZN(new_n2642_));
  AOI21_X1   g00207(.A1(new_n2642_), .A2(pi0107), .B(pi0063), .ZN(new_n2643_));
  INV_X1     g00208(.I(pi0064), .ZN(new_n2644_));
  AOI21_X1   g00209(.A1(new_n2641_), .A2(new_n2539_), .B(new_n2644_), .ZN(new_n2645_));
  AND3_X2    g00210(.A1(new_n2639_), .A2(new_n2565_), .A3(new_n2643_), .Z(new_n2647_));
  NAND2_X1   g00211(.A1(new_n2639_), .A2(new_n2565_), .ZN(new_n2648_));
  NAND2_X1   g00212(.A1(new_n2643_), .A2(pi0064), .ZN(new_n2649_));
  NAND2_X1   g00213(.A1(new_n2648_), .A2(new_n2649_), .ZN(new_n2650_));
  INV_X1     g00214(.I(new_n2645_), .ZN(new_n2651_));
  NAND3_X1   g00215(.A1(new_n2568_), .A2(pi0065), .A3(new_n2450_), .ZN(new_n2652_));
  NOR3_X1    g00216(.A1(new_n2651_), .A2(new_n2543_), .A3(new_n2652_), .ZN(new_n2653_));
  NAND2_X1   g00217(.A1(new_n2650_), .A2(new_n2653_), .ZN(new_n2654_));
  OAI21_X1   g00218(.A1(new_n2654_), .A2(new_n2647_), .B(new_n2564_), .ZN(new_n2655_));
  AOI21_X1   g00219(.A1(new_n2655_), .A2(new_n2513_), .B(new_n2561_), .ZN(new_n2656_));
  OAI21_X1   g00220(.A1(new_n2656_), .A2(new_n2556_), .B(new_n2552_), .ZN(new_n2657_));
  AOI21_X1   g00221(.A1(new_n2548_), .A2(pi0086), .B(pi0094), .ZN(new_n2658_));
  NAND2_X1   g00222(.A1(new_n2658_), .A2(pi0086), .ZN(new_n2659_));
  AOI21_X1   g00223(.A1(new_n2657_), .A2(new_n2659_), .B(new_n2518_), .ZN(new_n2660_));
  OAI21_X1   g00224(.A1(new_n2660_), .A2(new_n2551_), .B(new_n2529_), .ZN(new_n2661_));
  AOI21_X1   g00225(.A1(new_n2661_), .A2(new_n2524_), .B(new_n2512_), .ZN(new_n2662_));
  XNOR2_X1   g00226(.A1(new_n2662_), .A2(new_n2511_), .ZN(new_n2663_));
  INV_X1     g00227(.I(pi0109), .ZN(new_n2664_));
  INV_X1     g00228(.I(pi0110), .ZN(new_n2665_));
  AOI21_X1   g00229(.A1(new_n2466_), .A2(new_n2664_), .B(new_n2665_), .ZN(new_n2666_));
  NOR3_X1    g00230(.A1(pi0053), .A2(pi0060), .A3(pi0086), .ZN(new_n2667_));
  NOR2_X1    g00231(.A1(pi0097), .A2(pi0108), .ZN(new_n2668_));
  INV_X1     g00232(.I(pi0046), .ZN(new_n2669_));
  NOR2_X1    g00233(.A1(new_n2669_), .A2(new_n2530_), .ZN(new_n2670_));
  NAND4_X1   g00234(.A1(new_n2670_), .A2(new_n2667_), .A3(new_n2668_), .A4(new_n2488_), .ZN(new_n2671_));
  INV_X1     g00235(.I(new_n2671_), .ZN(new_n2672_));
  INV_X1     g00236(.I(pi0047), .ZN(new_n2673_));
  INV_X1     g00237(.I(pi0091), .ZN(new_n2674_));
  NOR2_X1    g00238(.A1(new_n2673_), .A2(new_n2674_), .ZN(new_n2675_));
  OAI21_X1   g00239(.A1(new_n2458_), .A2(new_n2675_), .B(new_n2672_), .ZN(new_n2676_));
  NOR2_X1    g00240(.A1(new_n2666_), .A2(new_n2676_), .ZN(new_n2677_));
  INV_X1     g00241(.I(new_n2487_), .ZN(new_n2678_));
  INV_X1     g00242(.I(pi0090), .ZN(new_n2679_));
  NOR2_X1    g00243(.A1(new_n2470_), .A2(new_n2679_), .ZN(new_n2680_));
  NOR2_X1    g00244(.A1(new_n2671_), .A2(pi0047), .ZN(new_n2681_));
  INV_X1     g00245(.I(new_n2681_), .ZN(new_n2682_));
  NOR2_X1    g00246(.A1(new_n2459_), .A2(new_n2682_), .ZN(new_n2683_));
  INV_X1     g00247(.I(new_n2683_), .ZN(new_n2684_));
  NOR2_X1    g00248(.A1(new_n2684_), .A2(new_n2674_), .ZN(new_n2685_));
  INV_X1     g00249(.I(pi0058), .ZN(new_n2686_));
  NOR2_X1    g00250(.A1(new_n2495_), .A2(new_n2686_), .ZN(new_n2687_));
  NOR4_X1    g00251(.A1(new_n2680_), .A2(new_n2678_), .A3(new_n2685_), .A4(new_n2687_), .ZN(new_n2688_));
  NOR2_X1    g00252(.A1(new_n2688_), .A2(new_n2677_), .ZN(new_n2689_));
  NOR2_X1    g00253(.A1(new_n2689_), .A2(new_n2467_), .ZN(new_n2690_));
  AOI21_X1   g00254(.A1(new_n2663_), .A2(new_n2690_), .B(new_n2509_), .ZN(new_n2691_));
  INV_X1     g00255(.I(pi0035), .ZN(new_n2692_));
  NOR2_X1    g00256(.A1(new_n2692_), .A2(new_n2509_), .ZN(new_n2693_));
  XOR2_X1    g00257(.A1(new_n2691_), .A2(new_n2693_), .Z(new_n2694_));
  INV_X1     g00258(.I(pi0225), .ZN(new_n2695_));
  NOR2_X1    g00259(.A1(new_n2507_), .A2(pi0093), .ZN(new_n2696_));
  INV_X1     g00260(.I(new_n2696_), .ZN(new_n2697_));
  NOR2_X1    g00261(.A1(pi0035), .A2(pi0070), .ZN(new_n2698_));
  AOI21_X1   g00262(.A1(new_n2697_), .A2(new_n2698_), .B(new_n2695_), .ZN(new_n2699_));
  INV_X1     g00263(.I(new_n2699_), .ZN(new_n2700_));
  NOR2_X1    g00264(.A1(new_n2700_), .A2(pi0051), .ZN(new_n2701_));
  INV_X1     g00265(.I(pi0051), .ZN(new_n2702_));
  NOR3_X1    g00266(.A1(pi0077), .A2(pi0088), .A3(pi0098), .ZN(new_n2703_));
  NAND4_X1   g00267(.A1(new_n2703_), .A2(new_n2517_), .A3(pi0081), .A4(new_n2454_), .ZN(new_n2704_));
  NOR3_X1    g00268(.A1(new_n2671_), .A2(new_n2490_), .A3(new_n2704_), .ZN(new_n2705_));
  NAND2_X1   g00269(.A1(new_n2542_), .A2(new_n2705_), .ZN(new_n2706_));
  INV_X1     g00270(.I(pi0070), .ZN(new_n2707_));
  INV_X1     g00271(.I(new_n2496_), .ZN(new_n2708_));
  NOR3_X1    g00272(.A1(new_n2678_), .A2(new_n2708_), .A3(new_n2707_), .ZN(new_n2709_));
  INV_X1     g00273(.I(new_n2709_), .ZN(new_n2710_));
  NOR2_X1    g00274(.A1(new_n2706_), .A2(new_n2710_), .ZN(new_n2711_));
  NOR2_X1    g00275(.A1(new_n2711_), .A2(new_n2702_), .ZN(new_n2712_));
  NOR2_X1    g00276(.A1(new_n2712_), .A2(pi0096), .ZN(new_n2713_));
  INV_X1     g00277(.I(new_n2713_), .ZN(new_n2714_));
  NOR2_X1    g00278(.A1(new_n2507_), .A2(new_n2708_), .ZN(new_n2715_));
  NOR2_X1    g00279(.A1(new_n2715_), .A2(new_n2707_), .ZN(new_n2716_));
  INV_X1     g00280(.I(new_n2716_), .ZN(new_n2717_));
  NAND2_X1   g00281(.A1(new_n2717_), .A2(new_n2714_), .ZN(new_n2718_));
  NAND4_X1   g00282(.A1(new_n2694_), .A2(new_n2508_), .A3(new_n2701_), .A4(new_n2718_), .ZN(new_n2719_));
  NOR2_X1    g00283(.A1(new_n2719_), .A2(new_n2506_), .ZN(new_n2720_));
  INV_X1     g00284(.I(pi0829), .ZN(new_n2721_));
  INV_X1     g00285(.I(pi0950), .ZN(new_n2722_));
  NAND2_X1   g00286(.A1(pi1092), .A2(pi1093), .ZN(new_n2723_));
  NOR3_X1    g00287(.A1(new_n2723_), .A2(new_n2721_), .A3(new_n2722_), .ZN(new_n2724_));
  INV_X1     g00288(.I(new_n2724_), .ZN(new_n2725_));
  INV_X1     g00289(.I(pi1091), .ZN(new_n2726_));
  INV_X1     g00290(.I(pi0957), .ZN(new_n2727_));
  NOR2_X1    g00291(.A1(new_n2727_), .A2(pi0833), .ZN(new_n2728_));
  NOR2_X1    g00292(.A1(new_n2728_), .A2(new_n2726_), .ZN(new_n2729_));
  INV_X1     g00293(.I(new_n2729_), .ZN(new_n2730_));
  NOR2_X1    g00294(.A1(new_n2730_), .A2(new_n2725_), .ZN(new_n2731_));
  INV_X1     g00295(.I(pi0841), .ZN(new_n2732_));
  INV_X1     g00296(.I(new_n2482_), .ZN(new_n2733_));
  NOR2_X1    g00297(.A1(pi0040), .A2(pi0072), .ZN(new_n2734_));
  INV_X1     g00298(.I(new_n2734_), .ZN(new_n2735_));
  NOR2_X1    g00299(.A1(new_n2733_), .A2(new_n2735_), .ZN(new_n2736_));
  NAND2_X1   g00300(.A1(new_n2736_), .A2(pi0032), .ZN(new_n2737_));
  AOI21_X1   g00301(.A1(new_n2737_), .A2(new_n2732_), .B(new_n2695_), .ZN(new_n2738_));
  INV_X1     g00302(.I(new_n2738_), .ZN(new_n2739_));
  AOI21_X1   g00303(.A1(new_n2528_), .A2(pi0097), .B(new_n2512_), .ZN(new_n2740_));
  XNOR2_X1   g00304(.A1(new_n2740_), .A2(new_n2511_), .ZN(new_n2741_));
  AOI21_X1   g00305(.A1(new_n2741_), .A2(new_n2690_), .B(new_n2509_), .ZN(new_n2742_));
  XOR2_X1    g00306(.A1(new_n2742_), .A2(new_n2693_), .Z(new_n2743_));
  NAND4_X1   g00307(.A1(new_n2743_), .A2(new_n2508_), .A3(new_n2701_), .A4(new_n2718_), .ZN(new_n2744_));
  INV_X1     g00308(.I(new_n2731_), .ZN(new_n2745_));
  NOR3_X1    g00309(.A1(new_n2485_), .A2(new_n2504_), .A3(new_n2745_), .ZN(new_n2746_));
  NOR2_X1    g00310(.A1(new_n2746_), .A2(pi0072), .ZN(new_n2747_));
  OAI21_X1   g00311(.A1(new_n2744_), .A2(new_n2747_), .B(new_n2739_), .ZN(new_n2748_));
  NAND3_X1   g00312(.A1(new_n2720_), .A2(new_n2731_), .A3(new_n2748_), .ZN(new_n2749_));
  INV_X1     g00313(.I(new_n2501_), .ZN(new_n2750_));
  NOR2_X1    g00314(.A1(pi0032), .A2(pi0040), .ZN(new_n2751_));
  AOI21_X1   g00315(.A1(new_n2750_), .A2(new_n2751_), .B(new_n2436_), .ZN(new_n2752_));
  NOR2_X1    g00316(.A1(new_n2436_), .A2(pi0479), .ZN(new_n2753_));
  NOR2_X1    g00317(.A1(new_n2752_), .A2(new_n2753_), .ZN(new_n2754_));
  INV_X1     g00318(.I(pi0096), .ZN(new_n2755_));
  NAND2_X1   g00319(.A1(new_n2702_), .A2(new_n2755_), .ZN(new_n2756_));
  NOR2_X1    g00320(.A1(new_n2716_), .A2(new_n2756_), .ZN(new_n2757_));
  INV_X1     g00321(.I(new_n2757_), .ZN(new_n2758_));
  NOR2_X1    g00322(.A1(new_n2734_), .A2(pi0032), .ZN(new_n2759_));
  AOI21_X1   g00323(.A1(new_n2758_), .A2(new_n2759_), .B(new_n2700_), .ZN(new_n2760_));
  INV_X1     g00324(.I(new_n2760_), .ZN(new_n2761_));
  NOR2_X1    g00325(.A1(pi0095), .A2(pi0137), .ZN(new_n2762_));
  AOI21_X1   g00326(.A1(new_n2739_), .A2(new_n2762_), .B(new_n2761_), .ZN(new_n2763_));
  AND2_X2    g00327(.A1(new_n2763_), .A2(pi0210), .Z(new_n2764_));
  OAI21_X1   g00328(.A1(new_n2764_), .A2(pi0137), .B(new_n2754_), .ZN(new_n2765_));
  AOI21_X1   g00329(.A1(new_n2749_), .A2(new_n2436_), .B(new_n2765_), .ZN(new_n2766_));
  NOR2_X1    g00330(.A1(pi0146), .A2(pi0210), .ZN(new_n2767_));
  INV_X1     g00331(.I(pi0234), .ZN(new_n2768_));
  NOR2_X1    g00332(.A1(new_n2768_), .A2(pi0332), .ZN(new_n2769_));
  AOI21_X1   g00333(.A1(new_n2720_), .A2(pi0032), .B(new_n2736_), .ZN(new_n2770_));
  NOR2_X1    g00334(.A1(new_n2754_), .A2(pi0137), .ZN(new_n2771_));
  NOR4_X1    g00335(.A1(new_n2770_), .A2(new_n2436_), .A3(new_n2695_), .A4(new_n2771_), .ZN(new_n2772_));
  INV_X1     g00336(.I(new_n2736_), .ZN(new_n2773_));
  NAND2_X1   g00337(.A1(pi0032), .A2(pi0095), .ZN(new_n2774_));
  AOI21_X1   g00338(.A1(new_n2773_), .A2(new_n2774_), .B(new_n2695_), .ZN(new_n2775_));
  INV_X1     g00339(.I(pi0137), .ZN(new_n2776_));
  INV_X1     g00340(.I(pi0210), .ZN(new_n2777_));
  NAND2_X1   g00341(.A1(new_n2776_), .A2(new_n2777_), .ZN(new_n2778_));
  OAI21_X1   g00342(.A1(new_n2775_), .A2(new_n2778_), .B(new_n2760_), .ZN(new_n2779_));
  OAI21_X1   g00343(.A1(new_n2772_), .A2(new_n2779_), .B(new_n2769_), .ZN(new_n2780_));
  INV_X1     g00344(.I(new_n2754_), .ZN(new_n2781_));
  NOR2_X1    g00345(.A1(new_n2781_), .A2(new_n2436_), .ZN(new_n2782_));
  NOR2_X1    g00346(.A1(new_n2720_), .A2(new_n2782_), .ZN(new_n2783_));
  OAI21_X1   g00347(.A1(new_n2783_), .A2(new_n2739_), .B(new_n2776_), .ZN(new_n2784_));
  NOR2_X1    g00348(.A1(pi0152), .A2(pi0161), .ZN(new_n2785_));
  INV_X1     g00349(.I(new_n2785_), .ZN(new_n2786_));
  NOR2_X1    g00350(.A1(new_n2786_), .A2(pi0166), .ZN(new_n2787_));
  INV_X1     g00351(.I(new_n2787_), .ZN(new_n2788_));
  NOR2_X1    g00352(.A1(new_n2763_), .A2(new_n2788_), .ZN(new_n2789_));
  NAND2_X1   g00353(.A1(new_n2784_), .A2(new_n2789_), .ZN(new_n2790_));
  AOI21_X1   g00354(.A1(new_n2780_), .A2(new_n2767_), .B(new_n2790_), .ZN(new_n2791_));
  OAI21_X1   g00355(.A1(new_n2791_), .A2(pi0146), .B(new_n2766_), .ZN(new_n2792_));
  INV_X1     g00356(.I(new_n2752_), .ZN(new_n2793_));
  INV_X1     g00357(.I(pi0032), .ZN(new_n2794_));
  NOR2_X1    g00358(.A1(new_n2475_), .A2(pi0070), .ZN(new_n2795_));
  INV_X1     g00359(.I(new_n2795_), .ZN(new_n2796_));
  NOR2_X1    g00360(.A1(new_n2678_), .A2(pi0093), .ZN(new_n2797_));
  INV_X1     g00361(.I(new_n2797_), .ZN(new_n2798_));
  NOR2_X1    g00362(.A1(new_n2798_), .A2(new_n2674_), .ZN(new_n2799_));
  INV_X1     g00363(.I(new_n2799_), .ZN(new_n2800_));
  NOR2_X1    g00364(.A1(new_n2800_), .A2(new_n2796_), .ZN(new_n2801_));
  INV_X1     g00365(.I(new_n2801_), .ZN(new_n2802_));
  NOR2_X1    g00366(.A1(new_n2684_), .A2(new_n2802_), .ZN(new_n2803_));
  INV_X1     g00367(.I(new_n2803_), .ZN(new_n2804_));
  NOR2_X1    g00368(.A1(new_n2804_), .A2(new_n2755_), .ZN(new_n2805_));
  NOR2_X1    g00369(.A1(new_n2805_), .A2(pi0072), .ZN(new_n2806_));
  NOR2_X1    g00370(.A1(new_n2505_), .A2(new_n2806_), .ZN(new_n2807_));
  NOR2_X1    g00371(.A1(new_n2719_), .A2(new_n2807_), .ZN(new_n2808_));
  INV_X1     g00372(.I(new_n2808_), .ZN(new_n2809_));
  OAI21_X1   g00373(.A1(new_n2809_), .A2(new_n2794_), .B(new_n2773_), .ZN(new_n2810_));
  NAND2_X1   g00374(.A1(new_n2810_), .A2(pi0225), .ZN(new_n2811_));
  NAND2_X1   g00375(.A1(new_n2811_), .A2(new_n2436_), .ZN(new_n2812_));
  NAND3_X1   g00376(.A1(new_n2812_), .A2(new_n2776_), .A3(new_n2793_), .ZN(new_n2813_));
  NOR2_X1    g00377(.A1(pi0234), .A2(pi0332), .ZN(new_n2814_));
  NOR2_X1    g00378(.A1(new_n2814_), .A2(pi0210), .ZN(new_n2815_));
  INV_X1     g00379(.I(new_n2751_), .ZN(new_n2816_));
  INV_X1     g00380(.I(new_n2805_), .ZN(new_n2817_));
  NOR3_X1    g00381(.A1(new_n2817_), .A2(pi0072), .A3(new_n2816_), .ZN(new_n2818_));
  NOR2_X1    g00382(.A1(new_n2818_), .A2(new_n2761_), .ZN(new_n2819_));
  INV_X1     g00383(.I(new_n2753_), .ZN(new_n2820_));
  NOR2_X1    g00384(.A1(new_n2820_), .A2(new_n2816_), .ZN(new_n2821_));
  NAND2_X1   g00385(.A1(new_n2750_), .A2(new_n2821_), .ZN(new_n2822_));
  NOR2_X1    g00386(.A1(new_n2822_), .A2(new_n2776_), .ZN(new_n2823_));
  OAI21_X1   g00387(.A1(new_n2775_), .A2(new_n2823_), .B(new_n2819_), .ZN(new_n2824_));
  AOI21_X1   g00388(.A1(new_n2813_), .A2(new_n2815_), .B(new_n2824_), .ZN(new_n2825_));
  NAND2_X1   g00389(.A1(new_n2739_), .A2(new_n2436_), .ZN(new_n2826_));
  INV_X1     g00390(.I(new_n2822_), .ZN(new_n2827_));
  NOR2_X1    g00391(.A1(new_n2827_), .A2(new_n2776_), .ZN(new_n2828_));
  OAI21_X1   g00392(.A1(new_n2826_), .A2(new_n2819_), .B(new_n2828_), .ZN(new_n2829_));
  NOR2_X1    g00393(.A1(new_n2746_), .A2(new_n2806_), .ZN(new_n2830_));
  OAI21_X1   g00394(.A1(new_n2744_), .A2(new_n2830_), .B(new_n2739_), .ZN(new_n2831_));
  OAI21_X1   g00395(.A1(new_n2793_), .A2(new_n2776_), .B(new_n2436_), .ZN(new_n2832_));
  NAND4_X1   g00396(.A1(new_n2808_), .A2(new_n2731_), .A3(new_n2831_), .A4(new_n2832_), .ZN(new_n2833_));
  NAND2_X1   g00397(.A1(new_n2833_), .A2(new_n2829_), .ZN(new_n2834_));
  NAND2_X1   g00398(.A1(new_n2834_), .A2(new_n2777_), .ZN(new_n2835_));
  AND2_X2    g00399(.A1(new_n2825_), .A2(new_n2835_), .Z(new_n2836_));
  INV_X1     g00400(.I(pi0153), .ZN(new_n2837_));
  NOR2_X1    g00401(.A1(new_n2788_), .A2(new_n2837_), .ZN(new_n2838_));
  INV_X1     g00402(.I(new_n2838_), .ZN(new_n2839_));
  OAI21_X1   g00403(.A1(new_n2836_), .A2(new_n2839_), .B(new_n2780_), .ZN(new_n2840_));
  NAND3_X1   g00404(.A1(new_n2840_), .A2(pi0228), .A3(new_n2766_), .ZN(new_n2841_));
  INV_X1     g00405(.I(new_n2767_), .ZN(new_n2842_));
  NOR2_X1    g00406(.A1(new_n2793_), .A2(new_n2436_), .ZN(new_n2843_));
  NOR2_X1    g00407(.A1(new_n2808_), .A2(new_n2843_), .ZN(new_n2844_));
  OAI21_X1   g00408(.A1(new_n2844_), .A2(new_n2739_), .B(new_n2776_), .ZN(new_n2845_));
  AOI21_X1   g00409(.A1(new_n2845_), .A2(new_n2829_), .B(new_n2842_), .ZN(new_n2846_));
  INV_X1     g00410(.I(pi0146), .ZN(new_n2847_));
  NOR2_X1    g00411(.A1(new_n2835_), .A2(new_n2847_), .ZN(new_n2848_));
  OAI21_X1   g00412(.A1(new_n2825_), .A2(new_n2846_), .B(new_n2848_), .ZN(new_n2849_));
  AOI21_X1   g00413(.A1(new_n2841_), .A2(new_n2792_), .B(new_n2849_), .ZN(new_n2850_));
  AOI21_X1   g00414(.A1(new_n2736_), .A2(pi0225), .B(new_n2794_), .ZN(new_n2851_));
  INV_X1     g00415(.I(new_n2851_), .ZN(new_n2852_));
  INV_X1     g00416(.I(new_n2715_), .ZN(new_n2853_));
  NOR4_X1    g00417(.A1(new_n2853_), .A2(new_n2486_), .A3(new_n2702_), .A4(new_n2437_), .ZN(new_n2854_));
  INV_X1     g00418(.I(new_n2854_), .ZN(new_n2855_));
  NOR2_X1    g00419(.A1(new_n2817_), .A2(new_n2855_), .ZN(new_n2856_));
  INV_X1     g00420(.I(new_n2856_), .ZN(new_n2857_));
  NOR2_X1    g00421(.A1(new_n2714_), .A2(new_n2702_), .ZN(new_n2858_));
  AOI21_X1   g00422(.A1(new_n2458_), .A2(pi0060), .B(pi0053), .ZN(new_n2859_));
  NOR2_X1    g00423(.A1(new_n2459_), .A2(pi0060), .ZN(new_n2860_));
  NOR2_X1    g00424(.A1(new_n2860_), .A2(new_n2518_), .ZN(new_n2861_));
  AOI21_X1   g00425(.A1(new_n2530_), .A2(new_n2461_), .B(pi0086), .ZN(new_n2862_));
  OR2_X2     g00426(.A1(new_n2861_), .A2(new_n2862_), .Z(new_n2863_));
  AOI21_X1   g00427(.A1(new_n2657_), .A2(new_n2859_), .B(new_n2863_), .ZN(new_n2864_));
  OAI21_X1   g00428(.A1(new_n2864_), .A2(new_n2528_), .B(new_n2524_), .ZN(new_n2865_));
  INV_X1     g00429(.I(new_n2677_), .ZN(new_n2866_));
  NOR2_X1    g00430(.A1(new_n2680_), .A2(pi0093), .ZN(new_n2867_));
  INV_X1     g00431(.I(new_n2685_), .ZN(new_n2868_));
  NOR2_X1    g00432(.A1(new_n2706_), .A2(new_n2686_), .ZN(new_n2869_));
  NAND3_X1   g00433(.A1(new_n2868_), .A2(new_n2487_), .A3(new_n2869_), .ZN(new_n2870_));
  OAI21_X1   g00434(.A1(new_n2867_), .A2(new_n2870_), .B(new_n2866_), .ZN(new_n2871_));
  INV_X1     g00435(.I(new_n2871_), .ZN(new_n2872_));
  INV_X1     g00436(.I(new_n2668_), .ZN(new_n2873_));
  INV_X1     g00437(.I(new_n2523_), .ZN(new_n2874_));
  NOR3_X1    g00438(.A1(new_n2874_), .A2(new_n2669_), .A3(new_n2873_), .ZN(new_n2875_));
  NOR2_X1    g00439(.A1(new_n2875_), .A2(pi0109), .ZN(new_n2876_));
  NOR2_X1    g00440(.A1(new_n2466_), .A2(new_n2664_), .ZN(new_n2877_));
  AOI21_X1   g00441(.A1(new_n2510_), .A2(new_n2877_), .B(new_n2876_), .ZN(new_n2878_));
  NOR2_X1    g00442(.A1(new_n2507_), .A2(new_n2509_), .ZN(new_n2879_));
  INV_X1     g00443(.I(new_n2879_), .ZN(new_n2880_));
  NAND2_X1   g00444(.A1(new_n2880_), .A2(new_n2692_), .ZN(new_n2881_));
  AOI21_X1   g00445(.A1(new_n2696_), .A2(pi0225), .B(new_n2692_), .ZN(new_n2882_));
  INV_X1     g00446(.I(new_n2882_), .ZN(new_n2883_));
  NOR2_X1    g00447(.A1(new_n2883_), .A2(new_n2881_), .ZN(new_n2884_));
  NOR4_X1    g00448(.A1(new_n2865_), .A2(new_n2872_), .A3(new_n2878_), .A4(new_n2884_), .ZN(new_n2885_));
  OAI21_X1   g00449(.A1(new_n2885_), .A2(new_n2858_), .B(pi0070), .ZN(new_n2886_));
  NOR2_X1    g00450(.A1(new_n2886_), .A2(new_n2506_), .ZN(new_n2887_));
  NAND2_X1   g00451(.A1(new_n2887_), .A2(new_n2857_), .ZN(new_n2888_));
  AOI21_X1   g00452(.A1(new_n2888_), .A2(new_n2852_), .B(pi0095), .ZN(new_n2889_));
  INV_X1     g00453(.I(pi0479), .ZN(new_n2890_));
  OAI21_X1   g00454(.A1(new_n2793_), .A2(new_n2890_), .B(pi0137), .ZN(new_n2891_));
  NAND2_X1   g00455(.A1(new_n2852_), .A2(pi0095), .ZN(new_n2892_));
  AOI21_X1   g00456(.A1(new_n2804_), .A2(pi0096), .B(new_n2735_), .ZN(new_n2893_));
  NAND2_X1   g00457(.A1(new_n2697_), .A2(pi0035), .ZN(new_n2894_));
  NAND2_X1   g00458(.A1(new_n2701_), .A2(new_n2894_), .ZN(new_n2895_));
  INV_X1     g00459(.I(new_n2859_), .ZN(new_n2896_));
  INV_X1     g00460(.I(new_n2516_), .ZN(new_n2897_));
  NOR2_X1    g00461(.A1(new_n2861_), .A2(new_n2897_), .ZN(new_n2898_));
  INV_X1     g00462(.I(new_n2898_), .ZN(new_n2899_));
  NOR3_X1    g00463(.A1(pi0046), .A2(pi0109), .A3(pi0110), .ZN(new_n2900_));
  NAND3_X1   g00464(.A1(new_n2675_), .A2(new_n2668_), .A3(new_n2900_), .ZN(new_n2901_));
  NOR2_X1    g00465(.A1(new_n2901_), .A2(pi0058), .ZN(new_n2902_));
  INV_X1     g00466(.I(new_n2902_), .ZN(new_n2903_));
  NOR4_X1    g00467(.A1(new_n2899_), .A2(new_n2479_), .A3(new_n2896_), .A4(new_n2903_), .ZN(new_n2904_));
  INV_X1     g00468(.I(new_n2904_), .ZN(new_n2905_));
  AOI21_X1   g00469(.A1(new_n2692_), .A2(new_n2905_), .B(new_n2895_), .ZN(new_n2906_));
  NOR2_X1    g00470(.A1(new_n2906_), .A2(pi0096), .ZN(new_n2907_));
  INV_X1     g00471(.I(new_n2907_), .ZN(new_n2908_));
  NAND2_X1   g00472(.A1(new_n2908_), .A2(new_n2893_), .ZN(new_n2909_));
  NAND4_X1   g00473(.A1(new_n2909_), .A2(new_n2794_), .A3(pi0095), .A4(pi0479), .ZN(new_n2910_));
  XNOR2_X1   g00474(.A1(new_n2910_), .A2(new_n2892_), .ZN(new_n2911_));
  INV_X1     g00475(.I(new_n2911_), .ZN(new_n2912_));
  OAI22_X1   g00476(.A1(new_n2889_), .A2(new_n2891_), .B1(pi0137), .B2(new_n2912_), .ZN(new_n2913_));
  NAND2_X1   g00477(.A1(new_n2913_), .A2(pi0210), .ZN(new_n2914_));
  NOR2_X1    g00478(.A1(new_n2697_), .A2(new_n2732_), .ZN(new_n2915_));
  INV_X1     g00479(.I(new_n2915_), .ZN(new_n2916_));
  NOR3_X1    g00480(.A1(new_n2916_), .A2(pi0051), .A3(pi0072), .ZN(new_n2917_));
  NOR4_X1    g00481(.A1(new_n2473_), .A2(new_n2692_), .A3(new_n2486_), .A4(new_n2695_), .ZN(new_n2918_));
  NAND2_X1   g00482(.A1(new_n2917_), .A2(new_n2918_), .ZN(new_n2919_));
  NAND2_X1   g00483(.A1(new_n2919_), .A2(pi0032), .ZN(new_n2920_));
  AOI21_X1   g00484(.A1(new_n2888_), .A2(new_n2920_), .B(pi0095), .ZN(new_n2921_));
  NAND2_X1   g00485(.A1(new_n2921_), .A2(pi0137), .ZN(new_n2922_));
  AOI21_X1   g00486(.A1(new_n2922_), .A2(new_n2890_), .B(new_n2793_), .ZN(new_n2923_));
  NOR2_X1    g00487(.A1(new_n2923_), .A2(new_n2730_), .ZN(new_n2924_));
  NAND2_X1   g00488(.A1(new_n2920_), .A2(pi0095), .ZN(new_n2925_));
  XNOR2_X1   g00489(.A1(new_n2910_), .A2(new_n2925_), .ZN(new_n2926_));
  INV_X1     g00490(.I(new_n2926_), .ZN(new_n2927_));
  AOI21_X1   g00491(.A1(new_n2776_), .A2(new_n2926_), .B(new_n2923_), .ZN(new_n2928_));
  NOR3_X1    g00492(.A1(new_n2524_), .A2(pi0108), .A3(pi0110), .ZN(new_n2929_));
  INV_X1     g00493(.I(new_n2929_), .ZN(new_n2930_));
  NOR4_X1    g00494(.A1(new_n2669_), .A2(new_n2673_), .A3(new_n2674_), .A4(new_n2664_), .ZN(new_n2931_));
  AOI21_X1   g00495(.A1(new_n2797_), .A2(new_n2931_), .B(pi0035), .ZN(new_n2932_));
  OAI21_X1   g00496(.A1(new_n2899_), .A2(new_n2859_), .B(new_n2461_), .ZN(new_n2933_));
  AOI21_X1   g00497(.A1(new_n2930_), .A2(new_n2932_), .B(new_n2933_), .ZN(new_n2934_));
  OAI21_X1   g00498(.A1(new_n2934_), .A2(new_n2895_), .B(new_n2755_), .ZN(new_n2935_));
  AOI21_X1   g00499(.A1(new_n2919_), .A2(pi0032), .B(new_n2893_), .ZN(new_n2936_));
  OAI21_X1   g00500(.A1(new_n2935_), .A2(new_n2936_), .B(new_n2724_), .ZN(new_n2937_));
  NAND2_X1   g00501(.A1(new_n2724_), .A2(pi0095), .ZN(new_n2938_));
  XOR2_X1    g00502(.A1(new_n2937_), .A2(new_n2938_), .Z(new_n2939_));
  NAND2_X1   g00503(.A1(new_n2939_), .A2(pi0479), .ZN(new_n2940_));
  NAND2_X1   g00504(.A1(new_n2940_), .A2(new_n2776_), .ZN(new_n2941_));
  NAND4_X1   g00505(.A1(new_n2928_), .A2(new_n2731_), .A3(new_n2927_), .A4(new_n2941_), .ZN(new_n2942_));
  XOR2_X1    g00506(.A1(new_n2942_), .A2(new_n2924_), .Z(new_n2943_));
  NAND2_X1   g00507(.A1(new_n2943_), .A2(new_n2777_), .ZN(new_n2944_));
  NAND2_X1   g00508(.A1(new_n2944_), .A2(new_n2914_), .ZN(new_n2945_));
  INV_X1     g00509(.I(new_n2928_), .ZN(new_n2946_));
  NOR2_X1    g00510(.A1(new_n2913_), .A2(new_n2777_), .ZN(new_n2947_));
  NAND2_X1   g00511(.A1(pi0146), .A2(pi0210), .ZN(new_n2948_));
  XOR2_X1    g00512(.A1(new_n2947_), .A2(new_n2948_), .Z(new_n2949_));
  NOR2_X1    g00513(.A1(new_n2949_), .A2(new_n2946_), .ZN(new_n2950_));
  OAI21_X1   g00514(.A1(new_n2950_), .A2(new_n2769_), .B(pi0146), .ZN(new_n2951_));
  INV_X1     g00515(.I(new_n2951_), .ZN(new_n2952_));
  AOI21_X1   g00516(.A1(new_n2945_), .A2(new_n2952_), .B(new_n2788_), .ZN(new_n2953_));
  NAND3_X1   g00517(.A1(new_n2945_), .A2(pi0234), .A3(pi0332), .ZN(new_n2954_));
  INV_X1     g00518(.I(pi0332), .ZN(new_n2955_));
  NAND4_X1   g00519(.A1(new_n2944_), .A2(pi0234), .A3(new_n2955_), .A4(new_n2914_), .ZN(new_n2956_));
  NAND2_X1   g00520(.A1(new_n2954_), .A2(new_n2956_), .ZN(new_n2957_));
  INV_X1     g00521(.I(new_n2497_), .ZN(new_n2958_));
  NOR2_X1    g00522(.A1(new_n2958_), .A2(pi0040), .ZN(new_n2959_));
  NAND2_X1   g00523(.A1(new_n2906_), .A2(new_n2959_), .ZN(new_n2960_));
  NAND2_X1   g00524(.A1(new_n2960_), .A2(new_n2794_), .ZN(new_n2961_));
  AOI21_X1   g00525(.A1(new_n2961_), .A2(new_n2762_), .B(new_n2852_), .ZN(new_n2962_));
  OAI21_X1   g00526(.A1(new_n2887_), .A2(new_n2782_), .B(new_n2851_), .ZN(new_n2963_));
  AOI21_X1   g00527(.A1(new_n2963_), .A2(pi0137), .B(new_n2962_), .ZN(new_n2964_));
  INV_X1     g00528(.I(new_n2964_), .ZN(new_n2965_));
  INV_X1     g00529(.I(new_n2920_), .ZN(new_n2966_));
  NOR2_X1    g00530(.A1(new_n2966_), .A2(pi0095), .ZN(new_n2967_));
  INV_X1     g00531(.I(new_n2967_), .ZN(new_n2968_));
  AOI21_X1   g00532(.A1(new_n2794_), .A2(new_n2960_), .B(new_n2968_), .ZN(new_n2969_));
  NOR2_X1    g00533(.A1(new_n2969_), .A2(pi0137), .ZN(new_n2970_));
  OAI21_X1   g00534(.A1(new_n2887_), .A2(new_n2966_), .B(new_n2436_), .ZN(new_n2971_));
  AOI21_X1   g00535(.A1(new_n2971_), .A2(new_n2754_), .B(new_n2776_), .ZN(new_n2972_));
  NOR2_X1    g00536(.A1(new_n2972_), .A2(new_n2970_), .ZN(new_n2973_));
  NOR2_X1    g00537(.A1(new_n2973_), .A2(new_n2777_), .ZN(new_n2974_));
  XOR2_X1    g00538(.A1(new_n2974_), .A2(new_n2948_), .Z(new_n2975_));
  NOR2_X1    g00539(.A1(new_n2975_), .A2(new_n2965_), .ZN(new_n2976_));
  NOR2_X1    g00540(.A1(new_n2976_), .A2(new_n2814_), .ZN(new_n2977_));
  INV_X1     g00541(.I(new_n2972_), .ZN(new_n2978_));
  INV_X1     g00542(.I(pi1092), .ZN(new_n2979_));
  NOR2_X1    g00543(.A1(new_n2722_), .A2(new_n2979_), .ZN(new_n2980_));
  INV_X1     g00544(.I(new_n2980_), .ZN(new_n2981_));
  NOR2_X1    g00545(.A1(new_n2981_), .A2(new_n2721_), .ZN(new_n2982_));
  INV_X1     g00546(.I(new_n2728_), .ZN(new_n2983_));
  INV_X1     g00547(.I(pi1093), .ZN(new_n2984_));
  NOR2_X1    g00548(.A1(new_n2726_), .A2(new_n2984_), .ZN(new_n2985_));
  INV_X1     g00549(.I(new_n2985_), .ZN(new_n2986_));
  NOR2_X1    g00550(.A1(new_n2986_), .A2(new_n2983_), .ZN(new_n2987_));
  NAND4_X1   g00551(.A1(new_n2934_), .A2(new_n2731_), .A3(new_n2982_), .A4(new_n2987_), .ZN(new_n2988_));
  INV_X1     g00552(.I(new_n2959_), .ZN(new_n2989_));
  NAND3_X1   g00553(.A1(new_n2895_), .A2(new_n2794_), .A3(new_n2989_), .ZN(new_n2990_));
  NAND2_X1   g00554(.A1(new_n2990_), .A2(new_n2904_), .ZN(new_n2991_));
  AOI21_X1   g00555(.A1(new_n2988_), .A2(new_n2692_), .B(new_n2991_), .ZN(new_n2992_));
  OAI21_X1   g00556(.A1(new_n2992_), .A2(new_n2968_), .B(new_n2776_), .ZN(new_n2993_));
  NAND2_X1   g00557(.A1(new_n2978_), .A2(new_n2993_), .ZN(new_n2994_));
  NOR2_X1    g00558(.A1(new_n2994_), .A2(pi0210), .ZN(new_n2995_));
  NOR2_X1    g00559(.A1(new_n2965_), .A2(new_n2777_), .ZN(new_n2996_));
  NOR2_X1    g00560(.A1(new_n2788_), .A2(new_n2847_), .ZN(new_n2997_));
  OAI21_X1   g00561(.A1(new_n2995_), .A2(new_n2996_), .B(new_n2997_), .ZN(new_n2998_));
  NOR2_X1    g00562(.A1(new_n2977_), .A2(new_n2998_), .ZN(new_n2999_));
  NAND2_X1   g00563(.A1(new_n2957_), .A2(new_n2999_), .ZN(new_n3000_));
  NAND2_X1   g00564(.A1(new_n3000_), .A2(new_n2953_), .ZN(new_n3001_));
  INV_X1     g00565(.I(new_n3001_), .ZN(new_n3002_));
  OAI21_X1   g00566(.A1(new_n3000_), .A2(new_n2953_), .B(pi0228), .ZN(new_n3003_));
  INV_X1     g00567(.I(pi0105), .ZN(new_n3004_));
  INV_X1     g00568(.I(pi0228), .ZN(new_n3005_));
  NOR2_X1    g00569(.A1(new_n3004_), .A2(new_n3005_), .ZN(new_n3006_));
  OAI21_X1   g00570(.A1(new_n3002_), .A2(new_n3003_), .B(new_n3006_), .ZN(new_n3007_));
  INV_X1     g00571(.I(new_n3003_), .ZN(new_n3008_));
  INV_X1     g00572(.I(new_n3006_), .ZN(new_n3009_));
  NAND3_X1   g00573(.A1(new_n3008_), .A2(new_n3001_), .A3(new_n3009_), .ZN(new_n3010_));
  INV_X1     g00574(.I(pi0216), .ZN(new_n3011_));
  NOR2_X1    g00575(.A1(new_n2837_), .A2(pi0332), .ZN(new_n3012_));
  INV_X1     g00576(.I(new_n3012_), .ZN(new_n3013_));
  NOR2_X1    g00577(.A1(new_n3013_), .A2(new_n3011_), .ZN(new_n3014_));
  INV_X1     g00578(.I(new_n3014_), .ZN(new_n3015_));
  AOI21_X1   g00579(.A1(new_n3010_), .A2(new_n3007_), .B(new_n3015_), .ZN(new_n3016_));
  NOR2_X1    g00580(.A1(pi0210), .A2(pi0234), .ZN(new_n3017_));
  NOR4_X1    g00581(.A1(new_n2911_), .A2(pi0137), .A3(new_n2752_), .A4(new_n3017_), .ZN(new_n3018_));
  OR3_X2     g00582(.A1(new_n2865_), .A2(new_n2664_), .A3(new_n2512_), .Z(new_n3019_));
  NAND3_X1   g00583(.A1(new_n2865_), .A2(new_n2664_), .A3(new_n2510_), .ZN(new_n3020_));
  NOR2_X1    g00584(.A1(new_n2872_), .A2(new_n2467_), .ZN(new_n3021_));
  INV_X1     g00585(.I(new_n3021_), .ZN(new_n3022_));
  AOI21_X1   g00586(.A1(new_n3019_), .A2(new_n3020_), .B(new_n3022_), .ZN(new_n3023_));
  NOR2_X1    g00587(.A1(new_n3023_), .A2(new_n2881_), .ZN(new_n3024_));
  NOR2_X1    g00588(.A1(new_n3024_), .A2(new_n2882_), .ZN(new_n3025_));
  NOR2_X1    g00589(.A1(new_n3025_), .A2(new_n2858_), .ZN(new_n3026_));
  NOR3_X1    g00590(.A1(new_n3026_), .A2(new_n2707_), .A3(new_n2506_), .ZN(new_n3027_));
  NOR2_X1    g00591(.A1(new_n3027_), .A2(new_n2782_), .ZN(new_n3028_));
  NAND2_X1   g00592(.A1(new_n2993_), .A2(new_n3017_), .ZN(new_n3029_));
  NOR2_X1    g00593(.A1(new_n2787_), .A2(pi0146), .ZN(new_n3030_));
  NAND2_X1   g00594(.A1(new_n3030_), .A2(new_n3017_), .ZN(new_n3031_));
  XNOR2_X1   g00595(.A1(new_n3029_), .A2(new_n3031_), .ZN(new_n3032_));
  NOR2_X1    g00596(.A1(new_n2962_), .A2(pi0210), .ZN(new_n3033_));
  NAND3_X1   g00597(.A1(new_n2970_), .A2(pi0137), .A3(new_n2851_), .ZN(new_n3034_));
  NOR4_X1    g00598(.A1(new_n3028_), .A2(new_n3032_), .A3(new_n3033_), .A4(new_n3034_), .ZN(new_n3035_));
  NOR3_X1    g00599(.A1(new_n3028_), .A2(new_n2768_), .A3(new_n2920_), .ZN(new_n3036_));
  OAI21_X1   g00600(.A1(new_n3035_), .A2(pi0137), .B(new_n3036_), .ZN(new_n3037_));
  NAND2_X1   g00601(.A1(new_n2926_), .A2(new_n2793_), .ZN(new_n3038_));
  NOR3_X1    g00602(.A1(new_n3030_), .A2(new_n2725_), .A3(new_n2730_), .ZN(new_n3039_));
  AOI21_X1   g00603(.A1(new_n3038_), .A2(new_n3039_), .B(new_n2776_), .ZN(new_n3040_));
  INV_X1     g00604(.I(new_n2843_), .ZN(new_n3041_));
  NAND2_X1   g00605(.A1(new_n3027_), .A2(new_n2857_), .ZN(new_n3042_));
  NAND2_X1   g00606(.A1(new_n3042_), .A2(new_n3041_), .ZN(new_n3043_));
  INV_X1     g00607(.I(new_n3030_), .ZN(new_n3044_));
  NAND3_X1   g00608(.A1(new_n3044_), .A2(pi0137), .A3(new_n2729_), .ZN(new_n3045_));
  NOR4_X1    g00609(.A1(new_n2940_), .A2(new_n2752_), .A3(new_n2920_), .A4(new_n3045_), .ZN(new_n3046_));
  NAND2_X1   g00610(.A1(new_n3043_), .A2(new_n3046_), .ZN(new_n3047_));
  XOR2_X1    g00611(.A1(new_n3047_), .A2(new_n3040_), .Z(new_n3048_));
  NAND2_X1   g00612(.A1(new_n3048_), .A2(new_n3037_), .ZN(new_n3049_));
  AND3_X2    g00613(.A1(new_n3049_), .A2(pi0210), .A3(new_n3012_), .Z(new_n3050_));
  NAND3_X1   g00614(.A1(new_n2793_), .A2(pi0095), .A3(pi0137), .ZN(new_n3051_));
  AOI21_X1   g00615(.A1(new_n3042_), .A2(new_n3051_), .B(new_n2852_), .ZN(new_n3052_));
  OAI21_X1   g00616(.A1(new_n3050_), .A2(new_n3018_), .B(new_n3052_), .ZN(new_n3053_));
  INV_X1     g00617(.I(new_n3053_), .ZN(new_n3054_));
  OAI21_X1   g00618(.A1(new_n3016_), .A2(new_n2850_), .B(new_n3054_), .ZN(new_n3055_));
  NAND2_X1   g00619(.A1(new_n3055_), .A2(pi0221), .ZN(new_n3056_));
  INV_X1     g00620(.I(pi1144), .ZN(new_n3057_));
  INV_X1     g00621(.I(pi0833), .ZN(new_n3058_));
  NOR2_X1    g00622(.A1(new_n3058_), .A2(pi0216), .ZN(new_n3059_));
  NAND3_X1   g00623(.A1(new_n3059_), .A2(pi0332), .A3(pi0929), .ZN(new_n3060_));
  INV_X1     g00624(.I(pi0929), .ZN(new_n3061_));
  NAND3_X1   g00625(.A1(new_n3059_), .A2(new_n2955_), .A3(new_n3061_), .ZN(new_n3062_));
  AOI21_X1   g00626(.A1(new_n3060_), .A2(new_n3062_), .B(new_n3057_), .ZN(new_n3063_));
  INV_X1     g00627(.I(new_n3063_), .ZN(new_n3064_));
  AOI21_X1   g00628(.A1(pi0265), .A2(new_n2955_), .B(new_n3011_), .ZN(new_n3065_));
  NAND2_X1   g00629(.A1(new_n3065_), .A2(pi0221), .ZN(new_n3066_));
  NOR2_X1    g00630(.A1(new_n3064_), .A2(new_n3066_), .ZN(new_n3067_));
  NAND2_X1   g00631(.A1(new_n3056_), .A2(new_n3067_), .ZN(new_n3068_));
  INV_X1     g00632(.I(new_n3067_), .ZN(new_n3069_));
  NAND3_X1   g00633(.A1(new_n3055_), .A2(pi0221), .A3(new_n3069_), .ZN(new_n3070_));
  NOR2_X1    g00634(.A1(new_n2768_), .A2(new_n2955_), .ZN(new_n3071_));
  INV_X1     g00635(.I(pi0198), .ZN(new_n3072_));
  AND2_X2    g00636(.A1(new_n2913_), .A2(pi0198), .Z(new_n3073_));
  AOI21_X1   g00637(.A1(new_n2943_), .A2(new_n3072_), .B(new_n3073_), .ZN(new_n3074_));
  NAND2_X1   g00638(.A1(new_n3074_), .A2(pi0234), .ZN(new_n3075_));
  XNOR2_X1   g00639(.A1(new_n3075_), .A2(new_n3071_), .ZN(new_n3076_));
  NAND2_X1   g00640(.A1(new_n2964_), .A2(pi0198), .ZN(new_n3077_));
  OAI21_X1   g00641(.A1(new_n2994_), .A2(pi0198), .B(new_n3077_), .ZN(new_n3078_));
  NOR3_X1    g00642(.A1(pi0144), .A2(pi0174), .A3(pi0189), .ZN(new_n3079_));
  INV_X1     g00643(.I(new_n3079_), .ZN(new_n3080_));
  NAND2_X1   g00644(.A1(pi0142), .A2(pi0198), .ZN(new_n3081_));
  NOR2_X1    g00645(.A1(new_n2913_), .A2(new_n3072_), .ZN(new_n3082_));
  XOR2_X1    g00646(.A1(new_n3082_), .A2(new_n3081_), .Z(new_n3083_));
  OAI22_X1   g00647(.A1(new_n3083_), .A2(new_n2946_), .B1(new_n2768_), .B2(pi0332), .ZN(new_n3084_));
  INV_X1     g00648(.I(new_n2814_), .ZN(new_n3085_));
  NOR2_X1    g00649(.A1(new_n2973_), .A2(new_n3072_), .ZN(new_n3086_));
  XOR2_X1    g00650(.A1(new_n3086_), .A2(new_n3081_), .Z(new_n3087_));
  OAI21_X1   g00651(.A1(new_n3087_), .A2(new_n2965_), .B(new_n3085_), .ZN(new_n3088_));
  INV_X1     g00652(.I(pi0142), .ZN(new_n3089_));
  INV_X1     g00653(.I(pi0223), .ZN(new_n3090_));
  NOR2_X1    g00654(.A1(pi0222), .A2(pi0224), .ZN(new_n3091_));
  INV_X1     g00655(.I(new_n3091_), .ZN(new_n3092_));
  NOR4_X1    g00656(.A1(new_n3080_), .A2(new_n3089_), .A3(new_n3092_), .A4(new_n3090_), .ZN(new_n3093_));
  NAND4_X1   g00657(.A1(new_n3084_), .A2(new_n3088_), .A3(new_n3078_), .A4(new_n3093_), .ZN(new_n3094_));
  OAI22_X1   g00658(.A1(new_n3074_), .A2(new_n3094_), .B1(pi0223), .B2(new_n3080_), .ZN(new_n3095_));
  NAND3_X1   g00659(.A1(new_n3076_), .A2(new_n3078_), .A3(new_n3095_), .ZN(new_n3096_));
  NOR2_X1    g00660(.A1(pi0039), .A2(pi0299), .ZN(new_n3097_));
  INV_X1     g00661(.I(pi0299), .ZN(new_n3098_));
  INV_X1     g00662(.I(pi0222), .ZN(new_n3099_));
  INV_X1     g00663(.I(pi0224), .ZN(new_n3100_));
  NOR2_X1    g00664(.A1(new_n3099_), .A2(new_n3100_), .ZN(new_n3101_));
  OAI21_X1   g00665(.A1(new_n3101_), .A2(pi0265), .B(pi0332), .ZN(new_n3102_));
  NOR2_X1    g00666(.A1(new_n3058_), .A2(pi0224), .ZN(new_n3103_));
  NOR2_X1    g00667(.A1(new_n3103_), .A2(pi0929), .ZN(new_n3104_));
  NOR2_X1    g00668(.A1(pi0332), .A2(pi1144), .ZN(new_n3105_));
  NAND2_X1   g00669(.A1(new_n3105_), .A2(pi0332), .ZN(new_n3106_));
  AOI21_X1   g00670(.A1(new_n3102_), .A2(new_n3104_), .B(new_n3106_), .ZN(new_n3107_));
  NOR2_X1    g00671(.A1(new_n3103_), .A2(new_n3099_), .ZN(new_n3108_));
  NOR2_X1    g00672(.A1(new_n3108_), .A2(pi0223), .ZN(new_n3109_));
  AOI21_X1   g00673(.A1(pi0223), .A2(new_n3109_), .B(new_n3107_), .ZN(new_n3110_));
  INV_X1     g00674(.I(pi0215), .ZN(new_n3111_));
  NOR2_X1    g00675(.A1(new_n3105_), .A2(new_n3111_), .ZN(new_n3112_));
  OR3_X2     g00676(.A1(new_n3110_), .A2(new_n3098_), .A3(new_n3112_), .Z(new_n3113_));
  AOI21_X1   g00677(.A1(new_n3096_), .A2(new_n3097_), .B(new_n3113_), .ZN(new_n3114_));
  INV_X1     g00678(.I(pi0054), .ZN(new_n3115_));
  NAND2_X1   g00679(.A1(new_n3110_), .A2(pi0299), .ZN(new_n3116_));
  NOR2_X1    g00680(.A1(new_n2820_), .A2(new_n2768_), .ZN(new_n3117_));
  NOR2_X1    g00681(.A1(new_n3117_), .A2(pi0332), .ZN(new_n3118_));
  INV_X1     g00682(.I(new_n3118_), .ZN(new_n3119_));
  NAND2_X1   g00683(.A1(new_n3105_), .A2(pi0215), .ZN(new_n3120_));
  INV_X1     g00684(.I(pi0221), .ZN(new_n3121_));
  AOI21_X1   g00685(.A1(new_n3009_), .A2(new_n3012_), .B(pi0216), .ZN(new_n3122_));
  NAND2_X1   g00686(.A1(new_n3118_), .A2(new_n3006_), .ZN(new_n3123_));
  AOI21_X1   g00687(.A1(new_n3123_), .A2(new_n3122_), .B(new_n3121_), .ZN(new_n3124_));
  XOR2_X1    g00688(.A1(new_n3124_), .A2(new_n3067_), .Z(new_n3125_));
  NAND2_X1   g00689(.A1(new_n3125_), .A2(new_n3111_), .ZN(new_n3126_));
  NAND2_X1   g00690(.A1(new_n3126_), .A2(new_n3120_), .ZN(new_n3127_));
  NOR2_X1    g00691(.A1(new_n3092_), .A2(pi0223), .ZN(new_n3128_));
  NAND4_X1   g00692(.A1(new_n3127_), .A2(pi0299), .A3(new_n3119_), .A4(new_n3128_), .ZN(new_n3129_));
  XNOR2_X1   g00693(.A1(new_n3129_), .A2(new_n3116_), .ZN(new_n3130_));
  INV_X1     g00694(.I(new_n3130_), .ZN(new_n3131_));
  NOR2_X1    g00695(.A1(pi0038), .A2(pi0100), .ZN(new_n3132_));
  INV_X1     g00696(.I(new_n3132_), .ZN(new_n3133_));
  NOR2_X1    g00697(.A1(new_n3133_), .A2(pi0039), .ZN(new_n3134_));
  NOR2_X1    g00698(.A1(new_n3130_), .A2(new_n3134_), .ZN(new_n3135_));
  INV_X1     g00699(.I(new_n3128_), .ZN(new_n3136_));
  NOR2_X1    g00700(.A1(new_n2816_), .A2(pi0095), .ZN(new_n3137_));
  INV_X1     g00701(.I(new_n3137_), .ZN(new_n3138_));
  NOR2_X1    g00702(.A1(new_n2501_), .A2(new_n3138_), .ZN(new_n3139_));
  INV_X1     g00703(.I(new_n3139_), .ZN(new_n3140_));
  NAND2_X1   g00704(.A1(new_n3140_), .A2(pi0234), .ZN(new_n3141_));
  NOR2_X1    g00705(.A1(pi0032), .A2(pi0095), .ZN(new_n3142_));
  NAND4_X1   g00706(.A1(new_n2734_), .A2(new_n3142_), .A3(new_n2702_), .A4(new_n2755_), .ZN(new_n3143_));
  INV_X1     g00707(.I(new_n3143_), .ZN(new_n3144_));
  NAND4_X1   g00708(.A1(new_n2542_), .A2(new_n2705_), .A3(new_n2709_), .A4(new_n3144_), .ZN(new_n3145_));
  NOR3_X1    g00709(.A1(new_n3145_), .A2(new_n2768_), .A3(new_n2820_), .ZN(new_n3146_));
  XOR2_X1    g00710(.A1(new_n3141_), .A2(new_n3146_), .Z(new_n3147_));
  AOI21_X1   g00711(.A1(new_n3147_), .A2(pi0137), .B(new_n3119_), .ZN(new_n3148_));
  INV_X1     g00712(.I(new_n3148_), .ZN(new_n3149_));
  NOR2_X1    g00713(.A1(new_n3110_), .A2(new_n3098_), .ZN(new_n3150_));
  INV_X1     g00714(.I(new_n3150_), .ZN(new_n3151_));
  AOI21_X1   g00715(.A1(new_n3136_), .A2(new_n3151_), .B(new_n3149_), .ZN(new_n3152_));
  INV_X1     g00716(.I(new_n3152_), .ZN(new_n3153_));
  OAI21_X1   g00717(.A1(new_n3063_), .A2(new_n3121_), .B(pi0215), .ZN(new_n3154_));
  NOR4_X1    g00718(.A1(new_n3140_), .A2(new_n2776_), .A3(new_n2837_), .A4(new_n2955_), .ZN(new_n3155_));
  INV_X1     g00719(.I(new_n3155_), .ZN(new_n3156_));
  NAND2_X1   g00720(.A1(new_n3156_), .A2(pi0228), .ZN(new_n3157_));
  NAND2_X1   g00721(.A1(new_n3012_), .A2(new_n3004_), .ZN(new_n3158_));
  OAI21_X1   g00722(.A1(new_n3149_), .A2(new_n3004_), .B(new_n3158_), .ZN(new_n3159_));
  NOR4_X1    g00723(.A1(new_n2494_), .A2(new_n2453_), .A3(new_n2710_), .A4(new_n3143_), .ZN(new_n3160_));
  NAND2_X1   g00724(.A1(new_n3160_), .A2(pi0137), .ZN(new_n3161_));
  NAND4_X1   g00725(.A1(new_n3159_), .A2(pi0228), .A3(new_n3012_), .A4(new_n3161_), .ZN(new_n3162_));
  XOR2_X1    g00726(.A1(new_n3162_), .A2(new_n3157_), .Z(new_n3163_));
  AOI21_X1   g00727(.A1(new_n3066_), .A2(new_n3011_), .B(new_n3120_), .ZN(new_n3164_));
  NAND2_X1   g00728(.A1(new_n3163_), .A2(new_n3164_), .ZN(new_n3165_));
  XNOR2_X1   g00729(.A1(new_n3165_), .A2(new_n3154_), .ZN(new_n3166_));
  NAND2_X1   g00730(.A1(new_n3166_), .A2(pi0299), .ZN(new_n3167_));
  NAND2_X1   g00731(.A1(new_n3167_), .A2(new_n3153_), .ZN(new_n3168_));
  AOI21_X1   g00732(.A1(new_n3168_), .A2(new_n3134_), .B(new_n3135_), .ZN(new_n3169_));
  NAND2_X1   g00733(.A1(new_n3169_), .A2(pi0092), .ZN(new_n3170_));
  NOR2_X1    g00734(.A1(pi0075), .A2(pi0087), .ZN(new_n3171_));
  NAND2_X1   g00735(.A1(new_n3171_), .A2(pi0092), .ZN(new_n3172_));
  XOR2_X1    g00736(.A1(new_n3170_), .A2(new_n3172_), .Z(new_n3173_));
  NAND2_X1   g00737(.A1(new_n3173_), .A2(new_n3131_), .ZN(new_n3174_));
  INV_X1     g00738(.I(pi0074), .ZN(new_n3175_));
  INV_X1     g00739(.I(new_n3127_), .ZN(new_n3176_));
  INV_X1     g00740(.I(new_n3122_), .ZN(new_n3177_));
  NAND2_X1   g00741(.A1(pi0215), .A2(pi0221), .ZN(new_n3178_));
  NOR3_X1    g00742(.A1(new_n3149_), .A2(new_n3177_), .A3(new_n3178_), .ZN(new_n3179_));
  INV_X1     g00743(.I(new_n3179_), .ZN(new_n3180_));
  NAND2_X1   g00744(.A1(new_n3152_), .A2(pi0299), .ZN(new_n3181_));
  AOI21_X1   g00745(.A1(new_n3181_), .A2(new_n3176_), .B(new_n3180_), .ZN(new_n3182_));
  INV_X1     g00746(.I(pi0039), .ZN(new_n3183_));
  NOR2_X1    g00747(.A1(pi0087), .A2(pi0100), .ZN(new_n3184_));
  INV_X1     g00748(.I(new_n3184_), .ZN(new_n3185_));
  NOR2_X1    g00749(.A1(new_n3185_), .A2(pi0038), .ZN(new_n3186_));
  INV_X1     g00750(.I(new_n3186_), .ZN(new_n3187_));
  NOR2_X1    g00751(.A1(pi0075), .A2(pi0092), .ZN(new_n3188_));
  INV_X1     g00752(.I(new_n3188_), .ZN(new_n3189_));
  NOR3_X1    g00753(.A1(new_n3187_), .A2(new_n3189_), .A3(new_n3183_), .ZN(new_n3190_));
  NOR2_X1    g00754(.A1(pi0039), .A2(pi0087), .ZN(new_n3191_));
  INV_X1     g00755(.I(new_n3191_), .ZN(new_n3192_));
  NOR2_X1    g00756(.A1(new_n3133_), .A2(new_n3192_), .ZN(new_n3193_));
  INV_X1     g00757(.I(new_n3193_), .ZN(new_n3194_));
  NOR2_X1    g00758(.A1(new_n3194_), .A2(new_n3189_), .ZN(new_n3195_));
  INV_X1     g00759(.I(new_n3195_), .ZN(new_n3196_));
  AOI22_X1   g00760(.A1(new_n3182_), .A2(new_n3190_), .B1(new_n3131_), .B2(new_n3196_), .ZN(new_n3197_));
  NAND2_X1   g00761(.A1(new_n3131_), .A2(new_n3175_), .ZN(new_n3198_));
  NOR4_X1    g00762(.A1(new_n3197_), .A2(pi0054), .A3(new_n3175_), .A4(new_n3198_), .ZN(new_n3199_));
  AOI21_X1   g00763(.A1(new_n3174_), .A2(new_n3115_), .B(new_n3199_), .ZN(new_n3200_));
  INV_X1     g00764(.I(pi0062), .ZN(new_n3201_));
  NOR2_X1    g00765(.A1(pi0054), .A2(pi0074), .ZN(new_n3202_));
  INV_X1     g00766(.I(new_n3202_), .ZN(new_n3203_));
  INV_X1     g00767(.I(new_n3171_), .ZN(new_n3204_));
  NOR2_X1    g00768(.A1(new_n3204_), .A2(pi0092), .ZN(new_n3205_));
  INV_X1     g00769(.I(new_n3205_), .ZN(new_n3206_));
  NOR2_X1    g00770(.A1(new_n3206_), .A2(new_n3203_), .ZN(new_n3207_));
  INV_X1     g00771(.I(new_n3207_), .ZN(new_n3208_));
  NOR2_X1    g00772(.A1(new_n3208_), .A2(pi0055), .ZN(new_n3209_));
  INV_X1     g00773(.I(new_n3209_), .ZN(new_n3210_));
  NOR2_X1    g00774(.A1(pi0038), .A2(pi0039), .ZN(new_n3211_));
  INV_X1     g00775(.I(new_n3211_), .ZN(new_n3212_));
  NOR2_X1    g00776(.A1(new_n3212_), .A2(pi0100), .ZN(new_n3213_));
  INV_X1     g00777(.I(new_n3213_), .ZN(new_n3214_));
  NOR2_X1    g00778(.A1(new_n3210_), .A2(new_n3214_), .ZN(new_n3215_));
  NAND2_X1   g00779(.A1(new_n3166_), .A2(new_n3215_), .ZN(new_n3216_));
  OAI21_X1   g00780(.A1(new_n3127_), .A2(new_n3215_), .B(new_n3216_), .ZN(new_n3217_));
  NOR2_X1    g00781(.A1(new_n3217_), .A2(new_n3201_), .ZN(new_n3218_));
  INV_X1     g00782(.I(pi0056), .ZN(new_n3219_));
  NOR2_X1    g00783(.A1(new_n3219_), .A2(new_n3201_), .ZN(new_n3220_));
  INV_X1     g00784(.I(new_n3220_), .ZN(new_n3221_));
  XOR2_X1    g00785(.A1(new_n3218_), .A2(new_n3221_), .Z(new_n3222_));
  NOR2_X1    g00786(.A1(new_n3222_), .A2(new_n3176_), .ZN(new_n3223_));
  INV_X1     g00787(.I(new_n3215_), .ZN(new_n3224_));
  NOR2_X1    g00788(.A1(pi0056), .A2(pi0062), .ZN(new_n3225_));
  INV_X1     g00789(.I(new_n3225_), .ZN(new_n3226_));
  NOR3_X1    g00790(.A1(new_n3180_), .A2(new_n3224_), .A3(new_n3226_), .ZN(new_n3227_));
  AOI21_X1   g00791(.A1(pi0057), .A2(new_n3127_), .B(new_n3227_), .ZN(new_n3228_));
  INV_X1     g00792(.I(pi0059), .ZN(new_n3229_));
  NOR2_X1    g00793(.A1(pi0057), .A2(pi0059), .ZN(new_n3230_));
  AOI21_X1   g00794(.A1(new_n3176_), .A2(new_n3230_), .B(new_n3229_), .ZN(new_n3231_));
  NAND2_X1   g00795(.A1(new_n3227_), .A2(new_n3231_), .ZN(new_n3232_));
  OAI22_X1   g00796(.A1(new_n3223_), .A2(pi0059), .B1(new_n3228_), .B2(new_n3232_), .ZN(new_n3233_));
  AND2_X2    g00797(.A1(new_n3169_), .A2(pi0087), .Z(new_n3234_));
  INV_X1     g00798(.I(pi0075), .ZN(new_n3235_));
  INV_X1     g00799(.I(new_n3147_), .ZN(new_n3236_));
  AOI21_X1   g00800(.A1(pi0095), .A2(pi0234), .B(pi0137), .ZN(new_n3237_));
  NAND2_X1   g00801(.A1(new_n3236_), .A2(new_n3237_), .ZN(new_n3238_));
  NOR2_X1    g00802(.A1(new_n3004_), .A2(new_n3005_), .ZN(new_n3239_));
  OAI21_X1   g00803(.A1(pi0332), .A2(new_n3239_), .B(new_n3030_), .ZN(new_n3240_));
  AOI21_X1   g00804(.A1(new_n3238_), .A2(new_n2777_), .B(new_n3240_), .ZN(new_n3241_));
  AOI21_X1   g00805(.A1(new_n3177_), .A2(new_n3066_), .B(new_n3120_), .ZN(new_n3242_));
  NAND2_X1   g00806(.A1(new_n3241_), .A2(new_n3242_), .ZN(new_n3243_));
  XNOR2_X1   g00807(.A1(new_n3243_), .A2(new_n3154_), .ZN(new_n3244_));
  OAI21_X1   g00808(.A1(new_n3147_), .A2(new_n2776_), .B(new_n3089_), .ZN(new_n3245_));
  NAND2_X1   g00809(.A1(new_n3080_), .A2(new_n3090_), .ZN(new_n3246_));
  NAND4_X1   g00810(.A1(new_n3245_), .A2(pi0198), .A3(new_n3118_), .A4(new_n3246_), .ZN(new_n3247_));
  OAI21_X1   g00811(.A1(new_n3145_), .A2(new_n3085_), .B(new_n3072_), .ZN(new_n3248_));
  AOI22_X1   g00812(.A1(new_n3248_), .A2(pi0137), .B1(new_n3090_), .B2(new_n3079_), .ZN(new_n3249_));
  AND3_X2    g00813(.A1(new_n2769_), .A2(pi0198), .A3(new_n2762_), .Z(new_n3250_));
  AOI21_X1   g00814(.A1(new_n3151_), .A2(new_n3092_), .B(new_n2820_), .ZN(new_n3251_));
  OAI21_X1   g00815(.A1(new_n3139_), .A2(new_n3250_), .B(new_n3251_), .ZN(new_n3252_));
  AOI21_X1   g00816(.A1(new_n3247_), .A2(new_n3249_), .B(new_n3252_), .ZN(new_n3253_));
  OAI21_X1   g00817(.A1(new_n3253_), .A2(new_n3193_), .B(pi0299), .ZN(new_n3254_));
  OAI21_X1   g00818(.A1(new_n3244_), .A2(new_n3254_), .B(new_n3235_), .ZN(new_n3255_));
  NAND4_X1   g00819(.A1(new_n3255_), .A2(pi0092), .A3(new_n3131_), .A4(new_n3193_), .ZN(new_n3256_));
  OAI21_X1   g00820(.A1(new_n3234_), .A2(pi0075), .B(new_n3256_), .ZN(new_n3257_));
  INV_X1     g00821(.I(pi0055), .ZN(new_n3258_));
  INV_X1     g00822(.I(pi0038), .ZN(new_n3259_));
  NAND2_X1   g00823(.A1(new_n3168_), .A2(pi0039), .ZN(new_n3260_));
  NOR2_X1    g00824(.A1(new_n3182_), .A2(new_n3259_), .ZN(new_n3261_));
  NOR2_X1    g00825(.A1(new_n3259_), .A2(new_n3183_), .ZN(new_n3262_));
  XOR2_X1    g00826(.A1(new_n3261_), .A2(new_n3262_), .Z(new_n3263_));
  NAND2_X1   g00827(.A1(new_n3263_), .A2(new_n3131_), .ZN(new_n3264_));
  NOR2_X1    g00828(.A1(pi0087), .A2(pi0100), .ZN(new_n3278_));
  AOI22_X1   g00829(.A1(new_n3260_), .A2(new_n3259_), .B1(new_n3264_), .B2(new_n3278_), .ZN(new_n3279_));
  OAI21_X1   g00830(.A1(new_n3236_), .A2(new_n3239_), .B(pi0332), .ZN(new_n3280_));
  NOR2_X1    g00831(.A1(new_n3065_), .A2(pi0216), .ZN(new_n3281_));
  NAND2_X1   g00832(.A1(new_n3280_), .A2(new_n3281_), .ZN(new_n3282_));
  NOR3_X1    g00833(.A1(new_n3160_), .A2(pi0228), .A3(new_n3013_), .ZN(new_n3283_));
  AOI21_X1   g00834(.A1(new_n3282_), .A2(new_n3283_), .B(new_n3121_), .ZN(new_n3284_));
  XOR2_X1    g00835(.A1(new_n3284_), .A2(new_n3178_), .Z(new_n3285_));
  INV_X1     g00836(.I(new_n3112_), .ZN(new_n3286_));
  NOR2_X1    g00837(.A1(new_n3189_), .A2(new_n3203_), .ZN(new_n3287_));
  INV_X1     g00838(.I(new_n3287_), .ZN(new_n3288_));
  NOR2_X1    g00839(.A1(new_n3288_), .A2(new_n3185_), .ZN(new_n3289_));
  INV_X1     g00840(.I(new_n3289_), .ZN(new_n3290_));
  NOR2_X1    g00841(.A1(new_n3290_), .A2(new_n3212_), .ZN(new_n3291_));
  INV_X1     g00842(.I(new_n3291_), .ZN(new_n3292_));
  NAND2_X1   g00843(.A1(new_n3127_), .A2(new_n3292_), .ZN(new_n3293_));
  NOR2_X1    g00844(.A1(new_n3258_), .A2(new_n3219_), .ZN(new_n3294_));
  AOI22_X1   g00845(.A1(new_n3293_), .A2(new_n3294_), .B1(new_n3286_), .B2(new_n3291_), .ZN(new_n3295_));
  NOR4_X1    g00846(.A1(new_n3285_), .A2(pi0062), .A3(new_n3064_), .A4(new_n3295_), .ZN(new_n3296_));
  OAI21_X1   g00847(.A1(new_n3217_), .A2(new_n3219_), .B(new_n3296_), .ZN(new_n3297_));
  AOI21_X1   g00848(.A1(new_n3297_), .A2(new_n3258_), .B(new_n3279_), .ZN(new_n3298_));
  NAND3_X1   g00849(.A1(new_n3233_), .A2(new_n3257_), .A3(new_n3298_), .ZN(new_n3299_));
  NOR2_X1    g00850(.A1(new_n3299_), .A2(new_n3200_), .ZN(new_n3300_));
  OAI21_X1   g00851(.A1(new_n3114_), .A2(pi0215), .B(new_n3300_), .ZN(new_n3301_));
  AOI21_X1   g00852(.A1(new_n3068_), .A2(new_n3070_), .B(new_n3301_), .ZN(po0153));
  INV_X1     g00853(.I(pi0092), .ZN(new_n3303_));
  NAND2_X1   g00854(.A1(new_n2734_), .A2(new_n3142_), .ZN(new_n3304_));
  NOR2_X1    g00855(.A1(new_n2817_), .A2(new_n3304_), .ZN(new_n3305_));
  NOR2_X1    g00856(.A1(new_n3305_), .A2(new_n2753_), .ZN(new_n3306_));
  NOR2_X1    g00857(.A1(new_n3306_), .A2(new_n2752_), .ZN(new_n3307_));
  INV_X1     g00858(.I(new_n3307_), .ZN(new_n3308_));
  NOR2_X1    g00859(.A1(new_n3306_), .A2(new_n3004_), .ZN(new_n3309_));
  NAND2_X1   g00860(.A1(new_n3309_), .A2(pi0228), .ZN(new_n3310_));
  OAI21_X1   g00861(.A1(pi0228), .A2(new_n3308_), .B(new_n3310_), .ZN(new_n3311_));
  NOR2_X1    g00862(.A1(pi0216), .A2(pi0221), .ZN(new_n3312_));
  INV_X1     g00863(.I(new_n3312_), .ZN(new_n3313_));
  NOR2_X1    g00864(.A1(new_n3313_), .A2(pi0215), .ZN(new_n3314_));
  NOR2_X1    g00865(.A1(new_n3306_), .A2(new_n3005_), .ZN(new_n3315_));
  INV_X1     g00866(.I(new_n3315_), .ZN(new_n3316_));
  NOR3_X1    g00867(.A1(new_n3023_), .A2(pi0070), .A3(new_n2881_), .ZN(new_n3317_));
  NAND2_X1   g00868(.A1(new_n2717_), .A2(new_n2894_), .ZN(new_n3318_));
  OAI21_X1   g00869(.A1(new_n3317_), .A2(new_n3318_), .B(new_n2702_), .ZN(new_n3319_));
  NAND4_X1   g00870(.A1(new_n3319_), .A2(pi0072), .A3(new_n2713_), .A4(new_n2751_), .ZN(new_n3320_));
  NAND2_X1   g00871(.A1(new_n3319_), .A2(new_n2713_), .ZN(new_n3321_));
  NAND3_X1   g00872(.A1(new_n3321_), .A2(new_n2437_), .A3(new_n2751_), .ZN(new_n3322_));
  INV_X1     g00873(.I(new_n2782_), .ZN(new_n3323_));
  NOR2_X1    g00874(.A1(new_n2750_), .A2(new_n2486_), .ZN(new_n3324_));
  NOR2_X1    g00875(.A1(new_n2736_), .A2(new_n2794_), .ZN(new_n3325_));
  NOR2_X1    g00876(.A1(new_n3325_), .A2(new_n3324_), .ZN(new_n3326_));
  INV_X1     g00877(.I(new_n3326_), .ZN(new_n3327_));
  AOI21_X1   g00878(.A1(new_n3327_), .A2(new_n3323_), .B(new_n2733_), .ZN(new_n3328_));
  INV_X1     g00879(.I(new_n3328_), .ZN(new_n3329_));
  AOI21_X1   g00880(.A1(new_n3322_), .A2(new_n3320_), .B(new_n3329_), .ZN(new_n3330_));
  NAND3_X1   g00881(.A1(new_n3330_), .A2(new_n3006_), .A3(new_n3316_), .ZN(new_n3331_));
  AOI21_X1   g00882(.A1(new_n3330_), .A2(new_n3006_), .B(new_n3316_), .ZN(new_n3332_));
  INV_X1     g00883(.I(new_n3332_), .ZN(new_n3333_));
  NAND2_X1   g00884(.A1(new_n3333_), .A2(new_n3331_), .ZN(new_n3334_));
  NAND3_X1   g00885(.A1(new_n3334_), .A2(pi0154), .A3(new_n3314_), .ZN(new_n3335_));
  INV_X1     g00886(.I(pi0154), .ZN(new_n3336_));
  INV_X1     g00887(.I(new_n3331_), .ZN(new_n3337_));
  NOR2_X1    g00888(.A1(new_n3337_), .A2(new_n3332_), .ZN(new_n3338_));
  NAND3_X1   g00889(.A1(new_n3338_), .A2(new_n3336_), .A3(new_n3314_), .ZN(new_n3339_));
  NAND2_X1   g00890(.A1(new_n3335_), .A2(new_n3339_), .ZN(new_n3340_));
  AOI21_X1   g00891(.A1(new_n3340_), .A2(new_n3311_), .B(new_n3098_), .ZN(new_n3341_));
  INV_X1     g00892(.I(pi0939), .ZN(new_n3342_));
  NAND2_X1   g00893(.A1(new_n3342_), .A2(pi0222), .ZN(new_n3343_));
  NAND2_X1   g00894(.A1(new_n3103_), .A2(pi0222), .ZN(new_n3344_));
  XOR2_X1    g00895(.A1(new_n3344_), .A2(new_n3343_), .Z(new_n3345_));
  NAND2_X1   g00896(.A1(new_n3345_), .A2(pi1146), .ZN(new_n3346_));
  NAND2_X1   g00897(.A1(new_n3346_), .A2(pi0223), .ZN(new_n3347_));
  NOR2_X1    g00898(.A1(new_n3306_), .A2(new_n3100_), .ZN(new_n3348_));
  XOR2_X1    g00899(.A1(new_n3348_), .A2(new_n3101_), .Z(new_n3349_));
  INV_X1     g00900(.I(pi1146), .ZN(new_n3350_));
  NOR2_X1    g00901(.A1(new_n3090_), .A2(new_n3350_), .ZN(new_n3351_));
  NAND3_X1   g00902(.A1(new_n3349_), .A2(pi0276), .A3(new_n3351_), .ZN(new_n3352_));
  XOR2_X1    g00903(.A1(new_n3352_), .A2(new_n3347_), .Z(new_n3353_));
  NOR2_X1    g00904(.A1(new_n3121_), .A2(pi0939), .ZN(new_n3354_));
  INV_X1     g00905(.I(new_n3059_), .ZN(new_n3355_));
  NOR2_X1    g00906(.A1(new_n3355_), .A2(new_n3121_), .ZN(new_n3356_));
  XNOR2_X1   g00907(.A1(new_n3356_), .A2(new_n3354_), .ZN(new_n3357_));
  NOR2_X1    g00908(.A1(new_n3357_), .A2(new_n3350_), .ZN(new_n3358_));
  INV_X1     g00909(.I(new_n3358_), .ZN(new_n3359_));
  NOR2_X1    g00910(.A1(pi0216), .A2(pi0276), .ZN(new_n3360_));
  NOR2_X1    g00911(.A1(new_n3121_), .A2(pi0215), .ZN(new_n3361_));
  INV_X1     g00912(.I(new_n3361_), .ZN(new_n3362_));
  AOI21_X1   g00913(.A1(new_n3359_), .A2(new_n3360_), .B(new_n3362_), .ZN(new_n3363_));
  AOI21_X1   g00914(.A1(pi0215), .A2(new_n3350_), .B(new_n3363_), .ZN(new_n3364_));
  INV_X1     g00915(.I(new_n3364_), .ZN(new_n3365_));
  NAND3_X1   g00916(.A1(new_n3353_), .A2(pi0299), .A3(new_n3365_), .ZN(new_n3366_));
  XNOR2_X1   g00917(.A1(new_n3341_), .A2(new_n3366_), .ZN(new_n3367_));
  INV_X1     g00918(.I(new_n3314_), .ZN(new_n3368_));
  NOR2_X1    g00919(.A1(new_n3009_), .A2(new_n2820_), .ZN(new_n3369_));
  INV_X1     g00920(.I(new_n3369_), .ZN(new_n3370_));
  OAI21_X1   g00921(.A1(new_n3368_), .A2(new_n3370_), .B(new_n3365_), .ZN(new_n3371_));
  NOR2_X1    g00922(.A1(new_n3006_), .A2(new_n3011_), .ZN(new_n3372_));
  NOR2_X1    g00923(.A1(new_n3011_), .A2(new_n3121_), .ZN(new_n3373_));
  XOR2_X1    g00924(.A1(new_n3372_), .A2(new_n3373_), .Z(new_n3374_));
  AOI21_X1   g00925(.A1(new_n3374_), .A2(pi0276), .B(new_n3111_), .ZN(new_n3375_));
  NOR2_X1    g00926(.A1(new_n3111_), .A2(new_n3350_), .ZN(new_n3376_));
  NAND2_X1   g00927(.A1(new_n3358_), .A2(new_n3376_), .ZN(new_n3377_));
  XOR2_X1    g00928(.A1(new_n3377_), .A2(new_n3375_), .Z(new_n3378_));
  NOR3_X1    g00929(.A1(new_n3378_), .A2(pi0154), .A3(pi0215), .ZN(new_n3379_));
  NAND2_X1   g00930(.A1(new_n3371_), .A2(new_n3379_), .ZN(new_n3380_));
  NOR2_X1    g00931(.A1(pi0223), .A2(pi0299), .ZN(new_n3381_));
  INV_X1     g00932(.I(new_n3381_), .ZN(new_n3382_));
  NOR2_X1    g00933(.A1(new_n3092_), .A2(new_n3382_), .ZN(new_n3383_));
  INV_X1     g00934(.I(new_n3383_), .ZN(new_n3384_));
  NOR2_X1    g00935(.A1(new_n3384_), .A2(new_n2820_), .ZN(new_n3385_));
  NOR2_X1    g00936(.A1(new_n3100_), .A2(pi0222), .ZN(new_n3386_));
  NAND2_X1   g00937(.A1(new_n3386_), .A2(pi0276), .ZN(new_n3387_));
  AOI21_X1   g00938(.A1(new_n3346_), .A2(new_n3090_), .B(new_n3387_), .ZN(new_n3388_));
  OAI21_X1   g00939(.A1(new_n3385_), .A2(new_n3351_), .B(pi0299), .ZN(new_n3389_));
  NOR2_X1    g00940(.A1(new_n3380_), .A2(new_n3389_), .ZN(new_n3390_));
  AOI21_X1   g00941(.A1(pi0146), .A2(pi0252), .B(new_n3145_), .ZN(new_n3391_));
  INV_X1     g00942(.I(new_n3391_), .ZN(new_n3392_));
  NOR2_X1    g00943(.A1(new_n3145_), .A2(pi0252), .ZN(new_n3393_));
  NOR2_X1    g00944(.A1(pi0161), .A2(pi0166), .ZN(new_n3394_));
  NAND3_X1   g00945(.A1(new_n3393_), .A2(pi0152), .A3(new_n3394_), .ZN(new_n3395_));
  INV_X1     g00946(.I(new_n3393_), .ZN(new_n3396_));
  NAND2_X1   g00947(.A1(new_n3394_), .A2(pi0152), .ZN(new_n3397_));
  NAND3_X1   g00948(.A1(new_n3396_), .A2(new_n3394_), .A3(new_n3397_), .ZN(new_n3398_));
  AOI21_X1   g00949(.A1(new_n3398_), .A2(new_n3395_), .B(new_n3392_), .ZN(new_n3399_));
  AOI21_X1   g00950(.A1(pi0152), .A2(new_n3392_), .B(new_n3399_), .ZN(new_n3400_));
  NOR2_X1    g00951(.A1(new_n3358_), .A2(new_n3376_), .ZN(new_n3401_));
  INV_X1     g00952(.I(new_n3401_), .ZN(new_n3402_));
  NAND3_X1   g00953(.A1(new_n3259_), .A2(new_n3011_), .A3(new_n3005_), .ZN(new_n3403_));
  NAND2_X1   g00954(.A1(pi0039), .A2(pi0154), .ZN(new_n3404_));
  NOR4_X1    g00955(.A1(new_n3402_), .A2(new_n3098_), .A3(new_n3403_), .A4(new_n3404_), .ZN(new_n3405_));
  NAND2_X1   g00956(.A1(new_n3400_), .A2(new_n3405_), .ZN(new_n3406_));
  NAND2_X1   g00957(.A1(new_n3406_), .A2(pi0100), .ZN(new_n3407_));
  NAND2_X1   g00958(.A1(new_n3390_), .A2(pi0100), .ZN(new_n3408_));
  XOR2_X1    g00959(.A1(new_n3408_), .A2(new_n3407_), .Z(new_n3409_));
  INV_X1     g00960(.I(new_n3380_), .ZN(new_n3410_));
  NOR2_X1    g00961(.A1(new_n3145_), .A2(pi0228), .ZN(new_n3411_));
  INV_X1     g00962(.I(new_n3411_), .ZN(new_n3412_));
  NOR3_X1    g00963(.A1(new_n3402_), .A2(new_n3412_), .A3(pi0216), .ZN(new_n3413_));
  INV_X1     g00964(.I(new_n3413_), .ZN(new_n3414_));
  AOI21_X1   g00965(.A1(new_n3371_), .A2(pi0154), .B(new_n3414_), .ZN(new_n3415_));
  OAI21_X1   g00966(.A1(new_n3410_), .A2(new_n3415_), .B(pi0299), .ZN(new_n3416_));
  NAND2_X1   g00967(.A1(new_n3132_), .A2(pi0039), .ZN(new_n3417_));
  NAND2_X1   g00968(.A1(new_n3416_), .A2(new_n3417_), .ZN(new_n3418_));
  NAND4_X1   g00969(.A1(new_n3409_), .A2(pi0038), .A3(new_n3390_), .A4(new_n3418_), .ZN(new_n3419_));
  NAND2_X1   g00970(.A1(new_n3419_), .A2(new_n3183_), .ZN(new_n3420_));
  OAI21_X1   g00971(.A1(new_n3390_), .A2(pi0087), .B(new_n3134_), .ZN(new_n3421_));
  OAI21_X1   g00972(.A1(new_n3421_), .A2(new_n3416_), .B(new_n3235_), .ZN(new_n3422_));
  NAND4_X1   g00973(.A1(new_n3367_), .A2(pi0087), .A3(new_n3420_), .A4(new_n3422_), .ZN(new_n3423_));
  NAND2_X1   g00974(.A1(new_n3390_), .A2(pi0075), .ZN(new_n3424_));
  AOI21_X1   g00975(.A1(new_n3423_), .A2(new_n3303_), .B(new_n3424_), .ZN(new_n3425_));
  INV_X1     g00976(.I(new_n3230_), .ZN(new_n3426_));
  NOR2_X1    g00977(.A1(new_n3410_), .A2(new_n3415_), .ZN(new_n3427_));
  NOR2_X1    g00978(.A1(new_n3292_), .A2(pi0055), .ZN(new_n3428_));
  NAND3_X1   g00979(.A1(new_n3427_), .A2(new_n3410_), .A3(new_n3428_), .ZN(new_n3429_));
  NOR2_X1    g00980(.A1(new_n3210_), .A2(pi0056), .ZN(new_n3430_));
  INV_X1     g00981(.I(new_n3430_), .ZN(new_n3431_));
  NOR2_X1    g00982(.A1(new_n3431_), .A2(new_n3214_), .ZN(new_n3432_));
  AOI21_X1   g00983(.A1(new_n3432_), .A2(pi0056), .B(new_n3201_), .ZN(new_n3433_));
  AOI21_X1   g00984(.A1(new_n3429_), .A2(new_n3433_), .B(new_n3426_), .ZN(new_n3434_));
  NAND3_X1   g00985(.A1(new_n3410_), .A2(pi0056), .A3(new_n3215_), .ZN(new_n3435_));
  NAND2_X1   g00986(.A1(new_n3435_), .A2(new_n3201_), .ZN(new_n3436_));
  NOR2_X1    g00987(.A1(new_n3214_), .A2(new_n3204_), .ZN(new_n3437_));
  OAI21_X1   g00988(.A1(new_n3390_), .A2(pi0092), .B(new_n3437_), .ZN(new_n3438_));
  NOR2_X1    g00989(.A1(new_n3438_), .A2(new_n3416_), .ZN(new_n3439_));
  AOI21_X1   g00990(.A1(new_n3380_), .A2(new_n3258_), .B(new_n3292_), .ZN(new_n3440_));
  AOI21_X1   g00991(.A1(new_n3440_), .A2(new_n3415_), .B(pi0056), .ZN(new_n3441_));
  NAND2_X1   g00992(.A1(new_n3390_), .A2(new_n3203_), .ZN(new_n3442_));
  NOR2_X1    g00993(.A1(new_n3378_), .A2(pi0154), .ZN(new_n3443_));
  NOR2_X1    g00994(.A1(new_n3364_), .A2(new_n3336_), .ZN(new_n3444_));
  NOR2_X1    g00995(.A1(new_n3443_), .A2(new_n3444_), .ZN(new_n3445_));
  INV_X1     g00996(.I(new_n3445_), .ZN(new_n3446_));
  NAND2_X1   g00997(.A1(new_n3446_), .A2(new_n3426_), .ZN(new_n3447_));
  NOR2_X1    g00998(.A1(pi0055), .A2(pi0239), .ZN(new_n3448_));
  NAND4_X1   g00999(.A1(new_n3442_), .A2(new_n3202_), .A3(new_n3447_), .A4(new_n3448_), .ZN(new_n3449_));
  NOR3_X1    g01000(.A1(new_n3449_), .A2(new_n3439_), .A3(new_n3441_), .ZN(new_n3450_));
  OAI21_X1   g01001(.A1(new_n3434_), .A2(new_n3436_), .B(new_n3450_), .ZN(new_n3451_));
  OAI21_X1   g01002(.A1(new_n3388_), .A2(pi0299), .B(new_n3351_), .ZN(new_n3452_));
  INV_X1     g01003(.I(new_n3452_), .ZN(new_n3453_));
  AOI21_X1   g01004(.A1(new_n3445_), .A2(pi0299), .B(new_n3453_), .ZN(new_n3454_));
  INV_X1     g01005(.I(pi0087), .ZN(new_n3455_));
  NOR3_X1    g01006(.A1(new_n2482_), .A2(new_n2437_), .A3(new_n2816_), .ZN(new_n3456_));
  OAI22_X1   g01007(.A1(new_n3326_), .A2(new_n2843_), .B1(new_n2806_), .B2(new_n3456_), .ZN(new_n3457_));
  INV_X1     g01008(.I(new_n3457_), .ZN(new_n3458_));
  NAND3_X1   g01009(.A1(new_n3319_), .A2(new_n2713_), .A3(new_n3458_), .ZN(new_n3459_));
  NAND2_X1   g01010(.A1(new_n3160_), .A2(pi0039), .ZN(new_n3460_));
  OAI21_X1   g01011(.A1(new_n3459_), .A2(pi0039), .B(new_n3460_), .ZN(new_n3461_));
  INV_X1     g01012(.I(pi0100), .ZN(new_n3462_));
  INV_X1     g01013(.I(new_n3454_), .ZN(new_n3463_));
  OAI21_X1   g01014(.A1(new_n3463_), .A2(new_n3259_), .B(new_n3462_), .ZN(new_n3464_));
  NAND2_X1   g01015(.A1(new_n3453_), .A2(pi0154), .ZN(new_n3465_));
  AOI21_X1   g01016(.A1(new_n3465_), .A2(new_n3098_), .B(new_n3364_), .ZN(new_n3466_));
  NOR2_X1    g01017(.A1(new_n3466_), .A2(pi0038), .ZN(new_n3467_));
  NAND2_X1   g01018(.A1(new_n3378_), .A2(pi0299), .ZN(new_n3468_));
  NAND2_X1   g01019(.A1(new_n3468_), .A2(new_n3465_), .ZN(new_n3469_));
  NAND4_X1   g01020(.A1(new_n3469_), .A2(pi0216), .A3(pi0228), .A4(new_n3401_), .ZN(new_n3470_));
  AOI21_X1   g01021(.A1(new_n3464_), .A2(new_n3467_), .B(new_n3470_), .ZN(new_n3471_));
  AOI21_X1   g01022(.A1(new_n3461_), .A2(new_n3471_), .B(new_n3455_), .ZN(new_n3472_));
  NAND2_X1   g01023(.A1(new_n3469_), .A2(new_n3413_), .ZN(new_n3473_));
  INV_X1     g01024(.I(new_n3134_), .ZN(new_n3474_));
  NOR2_X1    g01025(.A1(new_n3466_), .A2(new_n3474_), .ZN(new_n3475_));
  NAND2_X1   g01026(.A1(new_n3473_), .A2(new_n3475_), .ZN(new_n3476_));
  NOR2_X1    g01027(.A1(new_n3455_), .A2(new_n3462_), .ZN(new_n3477_));
  NAND2_X1   g01028(.A1(new_n3463_), .A2(new_n3477_), .ZN(new_n3478_));
  AOI21_X1   g01029(.A1(new_n3474_), .A2(new_n3454_), .B(new_n3478_), .ZN(new_n3479_));
  NAND3_X1   g01030(.A1(new_n3479_), .A2(new_n3406_), .A3(new_n3476_), .ZN(new_n3480_));
  OAI21_X1   g01031(.A1(new_n3472_), .A2(new_n3480_), .B(pi0075), .ZN(new_n3481_));
  AOI21_X1   g01032(.A1(new_n3472_), .A2(new_n3480_), .B(new_n3481_), .ZN(new_n3482_));
  NAND2_X1   g01033(.A1(pi0075), .A2(pi0092), .ZN(new_n3483_));
  XNOR2_X1   g01034(.A1(new_n3482_), .A2(new_n3483_), .ZN(new_n3484_));
  OAI21_X1   g01035(.A1(new_n3454_), .A2(pi0055), .B(new_n3203_), .ZN(new_n3485_));
  AOI21_X1   g01036(.A1(new_n3484_), .A2(new_n3454_), .B(new_n3485_), .ZN(new_n3486_));
  NAND3_X1   g01037(.A1(new_n3445_), .A2(new_n3413_), .A3(new_n3428_), .ZN(new_n3487_));
  AOI21_X1   g01038(.A1(new_n3487_), .A2(new_n3336_), .B(new_n3364_), .ZN(new_n3488_));
  INV_X1     g01039(.I(new_n3488_), .ZN(new_n3489_));
  NAND2_X1   g01040(.A1(new_n3446_), .A2(new_n3215_), .ZN(new_n3490_));
  AOI21_X1   g01041(.A1(new_n3489_), .A2(new_n3219_), .B(new_n3490_), .ZN(new_n3491_));
  NAND2_X1   g01042(.A1(new_n3414_), .A2(new_n3292_), .ZN(new_n3492_));
  NAND2_X1   g01043(.A1(new_n3258_), .A2(new_n3219_), .ZN(new_n3493_));
  AOI21_X1   g01044(.A1(new_n3492_), .A2(new_n3444_), .B(new_n3493_), .ZN(new_n3494_));
  INV_X1     g01045(.I(new_n3437_), .ZN(new_n3495_));
  AOI21_X1   g01046(.A1(new_n3454_), .A2(new_n3495_), .B(pi0092), .ZN(new_n3496_));
  NAND2_X1   g01047(.A1(new_n3446_), .A2(new_n3171_), .ZN(new_n3497_));
  NOR4_X1    g01048(.A1(new_n3496_), .A2(new_n3476_), .A3(new_n3494_), .A4(new_n3497_), .ZN(new_n3498_));
  OAI21_X1   g01049(.A1(new_n3491_), .A2(pi0062), .B(new_n3498_), .ZN(new_n3499_));
  OAI21_X1   g01050(.A1(new_n3489_), .A2(new_n3201_), .B(new_n3445_), .ZN(new_n3500_));
  NAND2_X1   g01051(.A1(new_n3230_), .A2(pi0239), .ZN(new_n3501_));
  AOI21_X1   g01052(.A1(new_n3500_), .A2(new_n3432_), .B(new_n3501_), .ZN(new_n3502_));
  OAI21_X1   g01053(.A1(new_n3486_), .A2(new_n3499_), .B(new_n3502_), .ZN(new_n3503_));
  OAI21_X1   g01054(.A1(new_n3425_), .A2(new_n3451_), .B(new_n3503_), .ZN(po0154));
  INV_X1     g01055(.I(pi0274), .ZN(new_n3505_));
  INV_X1     g01056(.I(pi0927), .ZN(new_n3506_));
  NAND2_X1   g01057(.A1(new_n3506_), .A2(pi0222), .ZN(new_n3507_));
  XOR2_X1    g01058(.A1(new_n3344_), .A2(new_n3507_), .Z(new_n3508_));
  NAND2_X1   g01059(.A1(new_n3508_), .A2(pi1145), .ZN(new_n3509_));
  NAND3_X1   g01060(.A1(new_n3509_), .A2(new_n3100_), .A3(new_n3505_), .ZN(new_n3510_));
  AOI21_X1   g01061(.A1(new_n3510_), .A2(pi0222), .B(new_n3090_), .ZN(new_n3511_));
  NOR2_X1    g01062(.A1(new_n3090_), .A2(new_n3098_), .ZN(new_n3512_));
  XOR2_X1    g01063(.A1(new_n3511_), .A2(new_n3512_), .Z(new_n3513_));
  NAND2_X1   g01064(.A1(new_n3513_), .A2(pi1145), .ZN(new_n3514_));
  INV_X1     g01065(.I(new_n3514_), .ZN(new_n3515_));
  NOR2_X1    g01066(.A1(new_n3515_), .A2(new_n3385_), .ZN(new_n3516_));
  INV_X1     g01067(.I(new_n3516_), .ZN(new_n3517_));
  INV_X1     g01068(.I(pi1145), .ZN(new_n3518_));
  NOR2_X1    g01069(.A1(new_n3121_), .A2(pi0927), .ZN(new_n3519_));
  XNOR2_X1   g01070(.A1(new_n3356_), .A2(new_n3519_), .ZN(new_n3520_));
  NOR2_X1    g01071(.A1(new_n3520_), .A2(new_n3518_), .ZN(new_n3521_));
  INV_X1     g01072(.I(new_n3521_), .ZN(new_n3522_));
  NAND2_X1   g01073(.A1(new_n3522_), .A2(pi0215), .ZN(new_n3523_));
  NOR2_X1    g01074(.A1(new_n3009_), .A2(new_n2753_), .ZN(new_n3524_));
  AOI21_X1   g01075(.A1(pi0151), .A2(new_n3009_), .B(new_n3524_), .ZN(new_n3525_));
  NOR2_X1    g01076(.A1(new_n3525_), .A2(new_n3011_), .ZN(new_n3526_));
  OAI21_X1   g01077(.A1(new_n3411_), .A2(new_n3526_), .B(pi0151), .ZN(new_n3527_));
  NOR2_X1    g01078(.A1(new_n3011_), .A2(new_n3505_), .ZN(new_n3528_));
  NOR2_X1    g01079(.A1(new_n3528_), .A2(pi0221), .ZN(new_n3529_));
  NOR2_X1    g01080(.A1(new_n3111_), .A2(new_n3518_), .ZN(new_n3530_));
  NAND3_X1   g01081(.A1(new_n3527_), .A2(new_n3529_), .A3(new_n3530_), .ZN(new_n3531_));
  XNOR2_X1   g01082(.A1(new_n3531_), .A2(new_n3523_), .ZN(new_n3532_));
  AND2_X2    g01083(.A1(new_n3532_), .A2(pi0299), .Z(new_n3533_));
  OAI21_X1   g01084(.A1(new_n3517_), .A2(new_n3533_), .B(new_n3134_), .ZN(new_n3534_));
  NOR2_X1    g01085(.A1(pi0215), .A2(pi0221), .ZN(new_n3535_));
  INV_X1     g01086(.I(new_n3535_), .ZN(new_n3536_));
  NOR2_X1    g01087(.A1(new_n3370_), .A2(new_n3536_), .ZN(new_n3537_));
  INV_X1     g01088(.I(pi0151), .ZN(new_n3538_));
  AOI21_X1   g01089(.A1(new_n3529_), .A2(pi0216), .B(new_n3006_), .ZN(new_n3539_));
  OAI21_X1   g01090(.A1(new_n3539_), .A2(new_n3538_), .B(pi0215), .ZN(new_n3540_));
  INV_X1     g01091(.I(new_n3530_), .ZN(new_n3541_));
  NOR2_X1    g01092(.A1(new_n3522_), .A2(new_n3541_), .ZN(new_n3542_));
  AND2_X2    g01093(.A1(new_n3542_), .A2(new_n3540_), .Z(new_n3543_));
  NOR2_X1    g01094(.A1(new_n3542_), .A2(new_n3540_), .ZN(new_n3544_));
  NOR2_X1    g01095(.A1(new_n3543_), .A2(new_n3544_), .ZN(new_n3545_));
  INV_X1     g01096(.I(new_n3545_), .ZN(new_n3546_));
  NAND2_X1   g01097(.A1(new_n3546_), .A2(new_n3537_), .ZN(new_n3547_));
  AOI21_X1   g01098(.A1(new_n3547_), .A2(new_n3505_), .B(new_n3011_), .ZN(new_n3548_));
  INV_X1     g01099(.I(new_n3548_), .ZN(new_n3549_));
  AOI21_X1   g01100(.A1(new_n3549_), .A2(pi0299), .B(new_n3517_), .ZN(new_n3550_));
  OAI21_X1   g01101(.A1(new_n3550_), .A2(new_n3134_), .B(new_n3534_), .ZN(new_n3551_));
  INV_X1     g01102(.I(new_n3529_), .ZN(new_n3552_));
  NAND3_X1   g01103(.A1(new_n3334_), .A2(pi0151), .A3(pi0216), .ZN(new_n3553_));
  NAND4_X1   g01104(.A1(new_n3333_), .A2(pi0151), .A3(new_n3331_), .A4(new_n3011_), .ZN(new_n3554_));
  NAND2_X1   g01105(.A1(new_n3553_), .A2(new_n3554_), .ZN(new_n3555_));
  AOI21_X1   g01106(.A1(new_n3555_), .A2(new_n3311_), .B(new_n3552_), .ZN(new_n3556_));
  NOR4_X1    g01107(.A1(new_n3556_), .A2(new_n3111_), .A3(new_n3098_), .A4(new_n3521_), .ZN(new_n3557_));
  NOR3_X1    g01108(.A1(new_n3338_), .A2(new_n3538_), .A3(new_n3011_), .ZN(new_n3558_));
  INV_X1     g01109(.I(new_n3554_), .ZN(new_n3559_));
  OAI21_X1   g01110(.A1(new_n3558_), .A2(new_n3559_), .B(new_n3311_), .ZN(new_n3560_));
  AOI21_X1   g01111(.A1(new_n3560_), .A2(new_n3529_), .B(new_n3521_), .ZN(new_n3561_));
  NOR3_X1    g01112(.A1(new_n3561_), .A2(pi0215), .A3(new_n3098_), .ZN(new_n3562_));
  OAI21_X1   g01113(.A1(new_n3562_), .A2(new_n3557_), .B(pi1145), .ZN(new_n3563_));
  NOR2_X1    g01114(.A1(new_n3259_), .A2(pi0039), .ZN(new_n3564_));
  INV_X1     g01115(.I(new_n3512_), .ZN(new_n3565_));
  NAND2_X1   g01116(.A1(new_n3349_), .A2(pi0274), .ZN(new_n3566_));
  AOI21_X1   g01117(.A1(new_n3566_), .A2(new_n3509_), .B(new_n3090_), .ZN(new_n3567_));
  XOR2_X1    g01118(.A1(new_n3567_), .A2(new_n3565_), .Z(new_n3568_));
  NOR2_X1    g01119(.A1(new_n3568_), .A2(new_n3518_), .ZN(new_n3569_));
  INV_X1     g01120(.I(new_n3569_), .ZN(new_n3570_));
  AOI21_X1   g01121(.A1(new_n3563_), .A2(new_n3564_), .B(new_n3570_), .ZN(new_n3571_));
  INV_X1     g01122(.I(new_n3550_), .ZN(new_n3572_));
  NOR2_X1    g01123(.A1(new_n3572_), .A2(new_n3259_), .ZN(new_n3573_));
  OAI21_X1   g01124(.A1(new_n3571_), .A2(pi0100), .B(new_n3573_), .ZN(new_n3574_));
  AND2_X2    g01125(.A1(new_n3400_), .A2(new_n3005_), .Z(new_n3575_));
  NOR2_X1    g01126(.A1(new_n3575_), .A2(new_n3524_), .ZN(new_n3576_));
  INV_X1     g01127(.I(new_n3576_), .ZN(new_n3577_));
  OAI21_X1   g01128(.A1(new_n3527_), .A2(new_n3552_), .B(new_n3577_), .ZN(new_n3578_));
  NAND4_X1   g01129(.A1(new_n3578_), .A2(pi0151), .A3(pi0215), .A4(pi1145), .ZN(new_n3579_));
  XNOR2_X1   g01130(.A1(new_n3579_), .A2(new_n3523_), .ZN(new_n3580_));
  OAI21_X1   g01131(.A1(new_n3516_), .A2(new_n3211_), .B(pi0299), .ZN(new_n3581_));
  AOI21_X1   g01132(.A1(new_n3550_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n3582_));
  OAI21_X1   g01133(.A1(new_n3580_), .A2(new_n3581_), .B(new_n3582_), .ZN(new_n3583_));
  NAND4_X1   g01134(.A1(new_n3574_), .A2(pi0075), .A3(pi0087), .A4(new_n3583_), .ZN(new_n3584_));
  NAND2_X1   g01135(.A1(new_n3574_), .A2(new_n3583_), .ZN(new_n3585_));
  NAND3_X1   g01136(.A1(new_n3585_), .A2(new_n3235_), .A3(pi0087), .ZN(new_n3586_));
  NAND2_X1   g01137(.A1(new_n3586_), .A2(new_n3584_), .ZN(new_n3587_));
  AOI21_X1   g01138(.A1(new_n3587_), .A2(new_n3551_), .B(pi0092), .ZN(new_n3588_));
  NAND2_X1   g01139(.A1(new_n3550_), .A2(pi0075), .ZN(new_n3589_));
  NOR2_X1    g01140(.A1(new_n3551_), .A2(new_n3303_), .ZN(new_n3590_));
  XOR2_X1    g01141(.A1(new_n3590_), .A2(new_n3172_), .Z(new_n3591_));
  NOR2_X1    g01142(.A1(new_n3591_), .A2(new_n3572_), .ZN(new_n3592_));
  NAND2_X1   g01143(.A1(new_n3532_), .A2(pi0062), .ZN(new_n3593_));
  NAND2_X1   g01144(.A1(new_n3432_), .A2(pi0062), .ZN(new_n3594_));
  XOR2_X1    g01145(.A1(new_n3593_), .A2(new_n3594_), .Z(new_n3595_));
  NAND2_X1   g01146(.A1(new_n3230_), .A2(pi0235), .ZN(new_n3596_));
  AOI21_X1   g01147(.A1(new_n3595_), .A2(new_n3548_), .B(new_n3596_), .ZN(new_n3597_));
  NAND2_X1   g01148(.A1(new_n3532_), .A2(pi0056), .ZN(new_n3598_));
  NOR2_X1    g01149(.A1(new_n3224_), .A2(new_n3219_), .ZN(new_n3599_));
  XOR2_X1    g01150(.A1(new_n3598_), .A2(new_n3599_), .Z(new_n3600_));
  OAI21_X1   g01151(.A1(new_n3549_), .A2(new_n3600_), .B(new_n3201_), .ZN(new_n3601_));
  NOR2_X1    g01152(.A1(new_n3601_), .A2(new_n3597_), .ZN(new_n3602_));
  NAND2_X1   g01153(.A1(new_n3532_), .A2(pi0055), .ZN(new_n3603_));
  NOR2_X1    g01154(.A1(new_n3292_), .A2(new_n3258_), .ZN(new_n3604_));
  INV_X1     g01155(.I(new_n3604_), .ZN(new_n3605_));
  XOR2_X1    g01156(.A1(new_n3603_), .A2(new_n3605_), .Z(new_n3606_));
  AOI21_X1   g01157(.A1(new_n3606_), .A2(new_n3548_), .B(pi0056), .ZN(new_n3607_));
  NAND2_X1   g01158(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n3608_));
  NOR4_X1    g01159(.A1(new_n3592_), .A2(new_n3602_), .A3(new_n3607_), .A4(new_n3608_), .ZN(new_n3609_));
  OAI21_X1   g01160(.A1(new_n3588_), .A2(new_n3589_), .B(new_n3609_), .ZN(new_n3610_));
  INV_X1     g01161(.I(pi0235), .ZN(new_n3611_));
  INV_X1     g01162(.I(new_n3537_), .ZN(new_n3612_));
  NAND2_X1   g01163(.A1(new_n3612_), .A2(new_n3611_), .ZN(new_n3613_));
  AOI21_X1   g01164(.A1(new_n3613_), .A2(new_n3528_), .B(new_n3230_), .ZN(new_n3614_));
  NAND2_X1   g01165(.A1(new_n3546_), .A2(new_n3614_), .ZN(new_n3615_));
  NOR2_X1    g01166(.A1(new_n3546_), .A2(new_n3098_), .ZN(new_n3616_));
  NOR2_X1    g01167(.A1(new_n3462_), .A2(pi0039), .ZN(new_n3617_));
  NAND3_X1   g01168(.A1(new_n3461_), .A2(pi0100), .A3(new_n3400_), .ZN(new_n3618_));
  XNOR2_X1   g01169(.A1(new_n3618_), .A2(new_n3617_), .ZN(new_n3619_));
  INV_X1     g01170(.I(new_n3616_), .ZN(new_n3620_));
  NAND2_X1   g01171(.A1(new_n3522_), .A2(new_n3541_), .ZN(new_n3621_));
  NAND3_X1   g01172(.A1(new_n3620_), .A2(new_n3403_), .A3(new_n3621_), .ZN(new_n3622_));
  AOI21_X1   g01173(.A1(new_n3619_), .A2(new_n3622_), .B(new_n3455_), .ZN(new_n3623_));
  NAND2_X1   g01174(.A1(new_n3514_), .A2(new_n3214_), .ZN(new_n3624_));
  NOR3_X1    g01175(.A1(new_n3621_), .A2(new_n3412_), .A3(pi0216), .ZN(new_n3625_));
  NAND3_X1   g01176(.A1(new_n3616_), .A2(new_n3624_), .A3(new_n3625_), .ZN(new_n3626_));
  NOR2_X1    g01177(.A1(new_n3616_), .A2(new_n3515_), .ZN(new_n3627_));
  NAND2_X1   g01178(.A1(new_n3627_), .A2(new_n3474_), .ZN(new_n3628_));
  NAND4_X1   g01179(.A1(new_n3628_), .A2(pi0087), .A3(new_n3515_), .A4(new_n3626_), .ZN(new_n3629_));
  OAI21_X1   g01180(.A1(new_n3623_), .A2(new_n3629_), .B(pi0075), .ZN(new_n3630_));
  AOI21_X1   g01181(.A1(new_n3623_), .A2(new_n3629_), .B(new_n3630_), .ZN(new_n3631_));
  XOR2_X1    g01182(.A1(new_n3631_), .A2(new_n3483_), .Z(new_n3632_));
  NOR3_X1    g01183(.A1(new_n3632_), .A2(new_n3515_), .A3(new_n3616_), .ZN(new_n3633_));
  OAI21_X1   g01184(.A1(new_n3627_), .A2(pi0055), .B(new_n3203_), .ZN(new_n3634_));
  NAND2_X1   g01185(.A1(new_n3625_), .A2(new_n3215_), .ZN(new_n3635_));
  AOI21_X1   g01186(.A1(new_n3221_), .A2(new_n3635_), .B(new_n3545_), .ZN(new_n3636_));
  NAND2_X1   g01187(.A1(new_n3545_), .A2(new_n3258_), .ZN(new_n3637_));
  AND3_X2    g01188(.A1(new_n3637_), .A2(new_n3291_), .A3(new_n3625_), .Z(new_n3638_));
  NOR3_X1    g01189(.A1(new_n3638_), .A2(pi0056), .A3(new_n3636_), .ZN(new_n3639_));
  OAI21_X1   g01190(.A1(new_n3546_), .A2(pi0062), .B(pi0056), .ZN(new_n3640_));
  NOR3_X1    g01191(.A1(new_n3204_), .A2(new_n3426_), .A3(pi0235), .ZN(new_n3641_));
  OAI21_X1   g01192(.A1(new_n3640_), .A2(new_n3635_), .B(new_n3641_), .ZN(new_n3642_));
  AOI21_X1   g01193(.A1(new_n3627_), .A2(new_n3495_), .B(pi0092), .ZN(new_n3643_));
  NOR4_X1    g01194(.A1(new_n3639_), .A2(new_n3643_), .A3(new_n3626_), .A4(new_n3642_), .ZN(new_n3644_));
  OAI21_X1   g01195(.A1(new_n3633_), .A2(new_n3634_), .B(new_n3644_), .ZN(new_n3645_));
  AOI21_X1   g01196(.A1(new_n3610_), .A2(new_n3615_), .B(new_n3645_), .ZN(po0155));
  NAND2_X1   g01197(.A1(new_n2820_), .A2(pi0284), .ZN(new_n3647_));
  AOI21_X1   g01198(.A1(pi0224), .A2(pi0264), .B(pi0222), .ZN(new_n3648_));
  INV_X1     g01199(.I(new_n3648_), .ZN(new_n3649_));
  INV_X1     g01200(.I(pi1143), .ZN(new_n3650_));
  NAND3_X1   g01201(.A1(new_n3103_), .A2(pi0222), .A3(pi0944), .ZN(new_n3651_));
  INV_X1     g01202(.I(pi0944), .ZN(new_n3652_));
  NAND3_X1   g01203(.A1(new_n3344_), .A2(pi0222), .A3(new_n3652_), .ZN(new_n3653_));
  AOI21_X1   g01204(.A1(new_n3653_), .A2(new_n3651_), .B(new_n3650_), .ZN(new_n3654_));
  INV_X1     g01205(.I(new_n3654_), .ZN(new_n3655_));
  OAI21_X1   g01206(.A1(new_n3655_), .A2(new_n3649_), .B(new_n3647_), .ZN(new_n3656_));
  AOI21_X1   g01207(.A1(new_n3656_), .A2(pi0224), .B(new_n3090_), .ZN(new_n3657_));
  XOR2_X1    g01208(.A1(new_n3657_), .A2(new_n3512_), .Z(new_n3658_));
  NAND2_X1   g01209(.A1(new_n3658_), .A2(pi1143), .ZN(new_n3659_));
  NOR2_X1    g01210(.A1(new_n3136_), .A2(new_n2820_), .ZN(new_n3660_));
  NOR2_X1    g01211(.A1(new_n3659_), .A2(new_n3660_), .ZN(new_n3661_));
  NAND3_X1   g01212(.A1(new_n3059_), .A2(pi0221), .A3(pi0944), .ZN(new_n3662_));
  NAND3_X1   g01213(.A1(new_n3355_), .A2(pi0221), .A3(new_n3652_), .ZN(new_n3663_));
  AOI21_X1   g01214(.A1(new_n3663_), .A2(new_n3662_), .B(new_n3650_), .ZN(new_n3664_));
  NOR2_X1    g01215(.A1(new_n3664_), .A2(new_n3111_), .ZN(new_n3665_));
  INV_X1     g01216(.I(new_n3665_), .ZN(new_n3666_));
  NOR2_X1    g01217(.A1(new_n3111_), .A2(new_n3650_), .ZN(new_n3667_));
  INV_X1     g01218(.I(new_n3667_), .ZN(new_n3668_));
  INV_X1     g01219(.I(pi0264), .ZN(new_n3669_));
  OAI21_X1   g01220(.A1(new_n3011_), .A2(new_n3669_), .B(new_n3121_), .ZN(new_n3670_));
  NAND2_X1   g01221(.A1(new_n3647_), .A2(pi0228), .ZN(new_n3671_));
  XOR2_X1    g01222(.A1(new_n3671_), .A2(new_n3009_), .Z(new_n3672_));
  NAND2_X1   g01223(.A1(new_n3672_), .A2(pi0146), .ZN(new_n3673_));
  INV_X1     g01224(.I(new_n3673_), .ZN(new_n3674_));
  NOR2_X1    g01225(.A1(new_n3674_), .A2(new_n3369_), .ZN(new_n3675_));
  NAND2_X1   g01226(.A1(new_n2847_), .A2(new_n3005_), .ZN(new_n3676_));
  AOI21_X1   g01227(.A1(new_n3675_), .A2(new_n3676_), .B(pi0216), .ZN(new_n3677_));
  NOR3_X1    g01228(.A1(new_n3677_), .A2(new_n3668_), .A3(new_n3670_), .ZN(new_n3678_));
  XOR2_X1    g01229(.A1(new_n3678_), .A2(new_n3666_), .Z(new_n3679_));
  AOI21_X1   g01230(.A1(new_n3679_), .A2(pi0299), .B(new_n3661_), .ZN(new_n3680_));
  NAND3_X1   g01231(.A1(new_n3160_), .A2(pi0228), .A3(pi0284), .ZN(new_n3681_));
  INV_X1     g01232(.I(pi0284), .ZN(new_n3682_));
  NAND3_X1   g01233(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n3682_), .ZN(new_n3683_));
  AOI21_X1   g01234(.A1(new_n3681_), .A2(new_n3683_), .B(new_n2847_), .ZN(new_n3684_));
  INV_X1     g01235(.I(new_n3684_), .ZN(new_n3685_));
  NOR2_X1    g01236(.A1(new_n3670_), .A2(new_n3011_), .ZN(new_n3686_));
  OAI21_X1   g01237(.A1(new_n3675_), .A2(new_n3686_), .B(new_n3667_), .ZN(new_n3687_));
  NOR2_X1    g01238(.A1(new_n3687_), .A2(new_n3685_), .ZN(new_n3688_));
  XOR2_X1    g01239(.A1(new_n3688_), .A2(new_n3666_), .Z(new_n3689_));
  INV_X1     g01240(.I(new_n3689_), .ZN(new_n3690_));
  OAI22_X1   g01241(.A1(new_n3690_), .A2(new_n3098_), .B1(new_n3659_), .B2(new_n3660_), .ZN(new_n3691_));
  NOR2_X1    g01242(.A1(new_n3680_), .A2(new_n3134_), .ZN(new_n3692_));
  AOI21_X1   g01243(.A1(new_n3134_), .A2(new_n3691_), .B(new_n3692_), .ZN(new_n3693_));
  NOR2_X1    g01244(.A1(new_n3235_), .A2(new_n3455_), .ZN(new_n3694_));
  NOR2_X1    g01245(.A1(new_n3111_), .A2(new_n3098_), .ZN(new_n3695_));
  INV_X1     g01246(.I(new_n3459_), .ZN(new_n3696_));
  NAND3_X1   g01247(.A1(new_n3308_), .A2(new_n2847_), .A3(pi0284), .ZN(new_n3697_));
  NAND2_X1   g01248(.A1(new_n2847_), .A2(pi0284), .ZN(new_n3698_));
  NAND4_X1   g01249(.A1(new_n3696_), .A2(pi0146), .A3(new_n3308_), .A4(new_n3698_), .ZN(new_n3699_));
  AOI21_X1   g01250(.A1(new_n3699_), .A2(new_n3697_), .B(new_n3005_), .ZN(new_n3700_));
  OAI21_X1   g01251(.A1(new_n3700_), .A2(pi0146), .B(new_n3330_), .ZN(new_n3701_));
  INV_X1     g01252(.I(new_n3306_), .ZN(new_n3702_));
  NAND2_X1   g01253(.A1(new_n3702_), .A2(new_n3006_), .ZN(new_n3703_));
  INV_X1     g01254(.I(new_n3664_), .ZN(new_n3704_));
  OAI21_X1   g01255(.A1(new_n3704_), .A2(new_n3670_), .B(new_n3011_), .ZN(new_n3705_));
  AND3_X2    g01256(.A1(new_n3703_), .A2(new_n3673_), .A3(new_n3705_), .Z(new_n3706_));
  AOI21_X1   g01257(.A1(new_n3701_), .A2(new_n3706_), .B(new_n3098_), .ZN(new_n3707_));
  XOR2_X1    g01258(.A1(new_n3707_), .A2(new_n3695_), .Z(new_n3708_));
  AOI21_X1   g01259(.A1(pi0223), .A2(pi1143), .B(pi0299), .ZN(new_n3709_));
  NOR2_X1    g01260(.A1(new_n3649_), .A2(new_n3100_), .ZN(new_n3710_));
  OAI21_X1   g01261(.A1(new_n3306_), .A2(new_n3710_), .B(pi0284), .ZN(new_n3711_));
  AND3_X2    g01262(.A1(new_n3711_), .A2(pi0223), .A3(new_n3655_), .Z(new_n3712_));
  OAI21_X1   g01263(.A1(new_n3712_), .A2(new_n3648_), .B(new_n3306_), .ZN(new_n3713_));
  AOI21_X1   g01264(.A1(new_n3713_), .A2(new_n3709_), .B(pi0039), .ZN(new_n3714_));
  AOI21_X1   g01265(.A1(new_n3708_), .A2(pi1143), .B(new_n3714_), .ZN(new_n3715_));
  NAND3_X1   g01266(.A1(new_n3711_), .A2(new_n3655_), .A3(new_n3709_), .ZN(new_n3716_));
  OAI21_X1   g01267(.A1(new_n3715_), .A2(new_n3716_), .B(new_n3259_), .ZN(new_n3717_));
  NOR2_X1    g01268(.A1(new_n3691_), .A2(new_n3183_), .ZN(new_n3718_));
  AOI21_X1   g01269(.A1(new_n3717_), .A2(new_n3718_), .B(pi0100), .ZN(new_n3719_));
  NAND2_X1   g01270(.A1(new_n3680_), .A2(pi0038), .ZN(new_n3720_));
  INV_X1     g01271(.I(pi0252), .ZN(new_n3721_));
  NOR2_X1    g01272(.A1(new_n2788_), .A2(new_n3721_), .ZN(new_n3722_));
  OAI21_X1   g01273(.A1(new_n3160_), .A2(pi0284), .B(new_n3722_), .ZN(new_n3723_));
  NAND2_X1   g01274(.A1(new_n3723_), .A2(new_n3005_), .ZN(new_n3724_));
  NAND3_X1   g01275(.A1(new_n3724_), .A2(pi0146), .A3(new_n3393_), .ZN(new_n3725_));
  NOR2_X1    g01276(.A1(new_n3687_), .A2(new_n3725_), .ZN(new_n3726_));
  XOR2_X1    g01277(.A1(new_n3726_), .A2(new_n3666_), .Z(new_n3727_));
  OAI21_X1   g01278(.A1(new_n3661_), .A2(new_n3211_), .B(pi0299), .ZN(new_n3728_));
  NOR2_X1    g01279(.A1(new_n3727_), .A2(new_n3728_), .ZN(new_n3729_));
  INV_X1     g01280(.I(new_n3680_), .ZN(new_n3730_));
  OAI21_X1   g01281(.A1(new_n3730_), .A2(new_n3211_), .B(pi0100), .ZN(new_n3731_));
  OAI22_X1   g01282(.A1(new_n3719_), .A2(new_n3720_), .B1(new_n3729_), .B2(new_n3731_), .ZN(new_n3732_));
  NAND2_X1   g01283(.A1(new_n3732_), .A2(pi0087), .ZN(new_n3733_));
  XOR2_X1    g01284(.A1(new_n3733_), .A2(new_n3694_), .Z(new_n3734_));
  OAI21_X1   g01285(.A1(new_n3734_), .A2(new_n3693_), .B(new_n3303_), .ZN(new_n3735_));
  NAND3_X1   g01286(.A1(new_n3735_), .A2(pi0075), .A3(new_n3680_), .ZN(new_n3736_));
  NAND2_X1   g01287(.A1(new_n3693_), .A2(pi0092), .ZN(new_n3737_));
  XNOR2_X1   g01288(.A1(new_n3737_), .A2(new_n3172_), .ZN(new_n3738_));
  NOR2_X1    g01289(.A1(new_n3738_), .A2(new_n3730_), .ZN(new_n3739_));
  INV_X1     g01290(.I(new_n3679_), .ZN(new_n3740_));
  NAND2_X1   g01291(.A1(new_n3689_), .A2(pi0062), .ZN(new_n3741_));
  XOR2_X1    g01292(.A1(new_n3741_), .A2(new_n3594_), .Z(new_n3742_));
  INV_X1     g01293(.I(pi0238), .ZN(new_n3743_));
  NAND2_X1   g01294(.A1(new_n3230_), .A2(new_n3743_), .ZN(new_n3744_));
  AOI21_X1   g01295(.A1(new_n3742_), .A2(new_n3740_), .B(new_n3744_), .ZN(new_n3745_));
  NAND2_X1   g01296(.A1(new_n3689_), .A2(pi0056), .ZN(new_n3746_));
  XOR2_X1    g01297(.A1(new_n3746_), .A2(new_n3599_), .Z(new_n3747_));
  OAI21_X1   g01298(.A1(new_n3747_), .A2(new_n3679_), .B(new_n3201_), .ZN(new_n3748_));
  NOR2_X1    g01299(.A1(new_n3745_), .A2(new_n3748_), .ZN(new_n3749_));
  NAND2_X1   g01300(.A1(new_n3689_), .A2(pi0055), .ZN(new_n3750_));
  XOR2_X1    g01301(.A1(new_n3750_), .A2(new_n3605_), .Z(new_n3751_));
  AOI21_X1   g01302(.A1(new_n3751_), .A2(new_n3740_), .B(pi0056), .ZN(new_n3752_));
  NAND2_X1   g01303(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n3753_));
  NOR4_X1    g01304(.A1(new_n3739_), .A2(new_n3749_), .A3(new_n3752_), .A4(new_n3753_), .ZN(new_n3754_));
  NOR2_X1    g01305(.A1(new_n3740_), .A2(new_n3230_), .ZN(new_n3755_));
  AOI21_X1   g01306(.A1(pi0216), .A2(pi0264), .B(new_n3612_), .ZN(new_n3756_));
  NAND2_X1   g01307(.A1(new_n3756_), .A2(pi0238), .ZN(new_n3757_));
  NOR2_X1    g01308(.A1(new_n3679_), .A2(new_n3756_), .ZN(new_n3758_));
  OAI21_X1   g01309(.A1(new_n3758_), .A2(new_n3098_), .B(new_n3659_), .ZN(new_n3759_));
  NOR2_X1    g01310(.A1(new_n3673_), .A2(new_n3668_), .ZN(new_n3760_));
  OAI21_X1   g01311(.A1(new_n3684_), .A2(new_n3686_), .B(new_n3760_), .ZN(new_n3761_));
  XOR2_X1    g01312(.A1(new_n3761_), .A2(new_n3665_), .Z(new_n3762_));
  NAND2_X1   g01313(.A1(new_n3762_), .A2(pi0299), .ZN(new_n3763_));
  NAND2_X1   g01314(.A1(new_n3763_), .A2(new_n3659_), .ZN(new_n3764_));
  INV_X1     g01315(.I(new_n3759_), .ZN(new_n3765_));
  NOR2_X1    g01316(.A1(new_n3765_), .A2(new_n3134_), .ZN(new_n3766_));
  AOI21_X1   g01317(.A1(new_n3134_), .A2(new_n3764_), .B(new_n3766_), .ZN(new_n3767_));
  INV_X1     g01318(.I(new_n3767_), .ZN(new_n3768_));
  NOR2_X1    g01319(.A1(pi0146), .A2(pi0284), .ZN(new_n3769_));
  NAND2_X1   g01320(.A1(new_n3696_), .A2(new_n3674_), .ZN(new_n3770_));
  OAI21_X1   g01321(.A1(new_n3770_), .A2(new_n3769_), .B(new_n3310_), .ZN(new_n3771_));
  AOI21_X1   g01322(.A1(new_n3771_), .A2(new_n3705_), .B(new_n3098_), .ZN(new_n3772_));
  XOR2_X1    g01323(.A1(new_n3772_), .A2(new_n3695_), .Z(new_n3773_));
  NAND2_X1   g01324(.A1(new_n3764_), .A2(pi0039), .ZN(new_n3774_));
  NOR2_X1    g01325(.A1(pi0038), .A2(pi0100), .ZN(new_n3775_));
  AOI21_X1   g01326(.A1(new_n3774_), .A2(new_n3775_), .B(new_n3714_), .ZN(new_n3776_));
  NOR2_X1    g01327(.A1(new_n3776_), .A2(new_n3650_), .ZN(new_n3777_));
  INV_X1     g01328(.I(new_n3686_), .ZN(new_n3778_));
  NAND2_X1   g01329(.A1(new_n3725_), .A2(new_n3778_), .ZN(new_n3779_));
  NAND2_X1   g01330(.A1(new_n3779_), .A2(new_n3760_), .ZN(new_n3780_));
  XOR2_X1    g01331(.A1(new_n3780_), .A2(new_n3666_), .Z(new_n3781_));
  AOI21_X1   g01332(.A1(new_n3659_), .A2(new_n3212_), .B(new_n3098_), .ZN(new_n3782_));
  NAND2_X1   g01333(.A1(new_n3781_), .A2(new_n3782_), .ZN(new_n3783_));
  AOI21_X1   g01334(.A1(new_n3765_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n3784_));
  AOI22_X1   g01335(.A1(new_n3773_), .A2(new_n3777_), .B1(new_n3783_), .B2(new_n3784_), .ZN(new_n3785_));
  NOR2_X1    g01336(.A1(new_n3785_), .A2(new_n3455_), .ZN(new_n3786_));
  XOR2_X1    g01337(.A1(new_n3786_), .A2(new_n3694_), .Z(new_n3787_));
  AOI21_X1   g01338(.A1(new_n3787_), .A2(new_n3768_), .B(pi0092), .ZN(new_n3788_));
  NOR3_X1    g01339(.A1(new_n3788_), .A2(new_n3235_), .A3(new_n3759_), .ZN(new_n3789_));
  NAND2_X1   g01340(.A1(new_n3767_), .A2(pi0092), .ZN(new_n3790_));
  XOR2_X1    g01341(.A1(new_n3790_), .A2(new_n3172_), .Z(new_n3791_));
  NAND2_X1   g01342(.A1(new_n3791_), .A2(new_n3765_), .ZN(new_n3792_));
  NAND2_X1   g01343(.A1(new_n3762_), .A2(pi0062), .ZN(new_n3793_));
  XOR2_X1    g01344(.A1(new_n3793_), .A2(new_n3594_), .Z(new_n3794_));
  NAND2_X1   g01345(.A1(new_n3794_), .A2(new_n3758_), .ZN(new_n3795_));
  NAND3_X1   g01346(.A1(new_n3795_), .A2(pi0238), .A3(new_n3230_), .ZN(new_n3796_));
  INV_X1     g01347(.I(new_n3599_), .ZN(new_n3797_));
  NAND2_X1   g01348(.A1(new_n3762_), .A2(pi0056), .ZN(new_n3798_));
  XOR2_X1    g01349(.A1(new_n3798_), .A2(new_n3797_), .Z(new_n3799_));
  AOI21_X1   g01350(.A1(new_n3799_), .A2(new_n3758_), .B(pi0062), .ZN(new_n3800_));
  NAND2_X1   g01351(.A1(new_n3796_), .A2(new_n3800_), .ZN(new_n3801_));
  NAND2_X1   g01352(.A1(new_n3762_), .A2(pi0055), .ZN(new_n3802_));
  XOR2_X1    g01353(.A1(new_n3802_), .A2(new_n3605_), .Z(new_n3803_));
  NAND2_X1   g01354(.A1(new_n3803_), .A2(new_n3758_), .ZN(new_n3804_));
  NAND2_X1   g01355(.A1(new_n3804_), .A2(new_n3219_), .ZN(new_n3805_));
  NOR2_X1    g01356(.A1(new_n3203_), .A2(pi0055), .ZN(new_n3806_));
  NAND4_X1   g01357(.A1(new_n3792_), .A2(new_n3801_), .A3(new_n3805_), .A4(new_n3806_), .ZN(new_n3807_));
  OAI22_X1   g01358(.A1(new_n3789_), .A2(new_n3807_), .B1(new_n3755_), .B2(new_n3757_), .ZN(new_n3808_));
  AOI21_X1   g01359(.A1(new_n3736_), .A2(new_n3754_), .B(new_n3808_), .ZN(po0156));
  INV_X1     g01360(.I(pi0249), .ZN(new_n3810_));
  INV_X1     g01361(.I(pi0262), .ZN(new_n3811_));
  NOR2_X1    g01362(.A1(new_n2753_), .A2(new_n3811_), .ZN(new_n3812_));
  AOI21_X1   g01363(.A1(pi0224), .A2(pi0277), .B(pi0222), .ZN(new_n3813_));
  INV_X1     g01364(.I(pi1142), .ZN(new_n3814_));
  NAND3_X1   g01365(.A1(new_n3103_), .A2(pi0222), .A3(pi0932), .ZN(new_n3815_));
  INV_X1     g01366(.I(pi0932), .ZN(new_n3816_));
  NAND3_X1   g01367(.A1(new_n3344_), .A2(pi0222), .A3(new_n3816_), .ZN(new_n3817_));
  AOI21_X1   g01368(.A1(new_n3817_), .A2(new_n3815_), .B(new_n3814_), .ZN(new_n3818_));
  AOI21_X1   g01369(.A1(new_n3818_), .A2(new_n3813_), .B(new_n3812_), .ZN(new_n3819_));
  OAI21_X1   g01370(.A1(new_n3819_), .A2(new_n3100_), .B(pi0223), .ZN(new_n3820_));
  XOR2_X1    g01371(.A1(new_n3820_), .A2(new_n3565_), .Z(new_n3821_));
  NAND2_X1   g01372(.A1(new_n3821_), .A2(pi1142), .ZN(new_n3822_));
  NAND3_X1   g01373(.A1(new_n3059_), .A2(pi0221), .A3(pi0932), .ZN(new_n3823_));
  NAND3_X1   g01374(.A1(new_n3355_), .A2(pi0221), .A3(new_n3816_), .ZN(new_n3824_));
  AOI21_X1   g01375(.A1(new_n3824_), .A2(new_n3823_), .B(new_n3814_), .ZN(new_n3825_));
  NOR2_X1    g01376(.A1(new_n3825_), .A2(new_n3111_), .ZN(new_n3826_));
  INV_X1     g01377(.I(pi0172), .ZN(new_n3827_));
  NAND3_X1   g01378(.A1(new_n3160_), .A2(pi0228), .A3(pi0262), .ZN(new_n3828_));
  NAND3_X1   g01379(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n3811_), .ZN(new_n3829_));
  AOI21_X1   g01380(.A1(new_n3828_), .A2(new_n3829_), .B(new_n3827_), .ZN(new_n3830_));
  AOI21_X1   g01381(.A1(pi0216), .A2(pi0277), .B(pi0221), .ZN(new_n3831_));
  INV_X1     g01382(.I(new_n3831_), .ZN(new_n3832_));
  NOR2_X1    g01383(.A1(new_n3832_), .A2(new_n3011_), .ZN(new_n3833_));
  NAND3_X1   g01384(.A1(new_n3812_), .A2(pi0105), .A3(pi0228), .ZN(new_n3834_));
  OR3_X2     g01385(.A1(new_n3812_), .A2(pi0105), .A3(new_n3005_), .Z(new_n3835_));
  AOI21_X1   g01386(.A1(new_n3835_), .A2(new_n3834_), .B(new_n3827_), .ZN(new_n3836_));
  INV_X1     g01387(.I(new_n3836_), .ZN(new_n3837_));
  NOR2_X1    g01388(.A1(new_n3111_), .A2(new_n3814_), .ZN(new_n3838_));
  INV_X1     g01389(.I(new_n3838_), .ZN(new_n3839_));
  NOR2_X1    g01390(.A1(new_n3837_), .A2(new_n3839_), .ZN(new_n3840_));
  OAI21_X1   g01391(.A1(new_n3830_), .A2(new_n3833_), .B(new_n3840_), .ZN(new_n3841_));
  XOR2_X1    g01392(.A1(new_n3841_), .A2(new_n3826_), .Z(new_n3842_));
  NAND2_X1   g01393(.A1(new_n3842_), .A2(pi0299), .ZN(new_n3843_));
  NAND2_X1   g01394(.A1(new_n3843_), .A2(new_n3822_), .ZN(new_n3844_));
  INV_X1     g01395(.I(new_n3822_), .ZN(new_n3845_));
  INV_X1     g01396(.I(new_n3826_), .ZN(new_n3846_));
  NAND2_X1   g01397(.A1(new_n3005_), .A2(pi0172), .ZN(new_n3847_));
  AOI21_X1   g01398(.A1(new_n3837_), .A2(new_n3847_), .B(pi0216), .ZN(new_n3848_));
  NOR3_X1    g01399(.A1(new_n3848_), .A2(new_n3832_), .A3(new_n3839_), .ZN(new_n3849_));
  XOR2_X1    g01400(.A1(new_n3849_), .A2(new_n3846_), .Z(new_n3850_));
  AOI21_X1   g01401(.A1(pi0299), .A2(new_n3850_), .B(new_n3845_), .ZN(new_n3851_));
  NOR2_X1    g01402(.A1(new_n3851_), .A2(new_n3134_), .ZN(new_n3852_));
  AOI21_X1   g01403(.A1(new_n3844_), .A2(new_n3134_), .B(new_n3852_), .ZN(new_n3853_));
  INV_X1     g01404(.I(new_n3853_), .ZN(new_n3854_));
  INV_X1     g01405(.I(new_n3695_), .ZN(new_n3855_));
  INV_X1     g01406(.I(new_n3825_), .ZN(new_n3856_));
  NAND3_X1   g01407(.A1(new_n3696_), .A2(pi0172), .A3(pi0262), .ZN(new_n3857_));
  NAND3_X1   g01408(.A1(new_n3459_), .A2(pi0172), .A3(new_n3811_), .ZN(new_n3858_));
  NAND2_X1   g01409(.A1(new_n3857_), .A2(new_n3858_), .ZN(new_n3859_));
  NOR2_X1    g01410(.A1(new_n3308_), .A2(new_n3827_), .ZN(new_n3860_));
  AOI21_X1   g01411(.A1(new_n3859_), .A2(new_n3860_), .B(pi0262), .ZN(new_n3861_));
  INV_X1     g01412(.I(new_n3330_), .ZN(new_n3862_));
  AOI21_X1   g01413(.A1(new_n3004_), .A2(pi0172), .B(new_n3005_), .ZN(new_n3863_));
  NOR3_X1    g01414(.A1(new_n3812_), .A2(pi0105), .A3(new_n3863_), .ZN(new_n3864_));
  NOR3_X1    g01415(.A1(new_n2817_), .A2(new_n3304_), .A3(new_n3864_), .ZN(new_n3865_));
  NOR2_X1    g01416(.A1(new_n3865_), .A2(pi0216), .ZN(new_n3866_));
  OR3_X2     g01417(.A1(new_n3862_), .A2(new_n3005_), .A3(new_n3866_), .Z(new_n3867_));
  OAI21_X1   g01418(.A1(new_n3867_), .A2(new_n3861_), .B(new_n3831_), .ZN(new_n3868_));
  AOI21_X1   g01419(.A1(new_n3868_), .A2(new_n3856_), .B(new_n3098_), .ZN(new_n3869_));
  XOR2_X1    g01420(.A1(new_n3869_), .A2(new_n3855_), .Z(new_n3870_));
  AOI21_X1   g01421(.A1(pi0223), .A2(pi1142), .B(pi0299), .ZN(new_n3871_));
  NAND2_X1   g01422(.A1(new_n3813_), .A2(pi0224), .ZN(new_n3872_));
  AOI21_X1   g01423(.A1(new_n3702_), .A2(new_n3872_), .B(new_n3811_), .ZN(new_n3873_));
  NOR3_X1    g01424(.A1(new_n3873_), .A2(new_n3090_), .A3(new_n3818_), .ZN(new_n3874_));
  OAI21_X1   g01425(.A1(new_n3874_), .A2(new_n3813_), .B(new_n3306_), .ZN(new_n3875_));
  AOI21_X1   g01426(.A1(new_n3875_), .A2(new_n3871_), .B(pi0039), .ZN(new_n3876_));
  NOR2_X1    g01427(.A1(pi0038), .A2(pi0100), .ZN(new_n3877_));
  INV_X1     g01428(.I(new_n3877_), .ZN(new_n3878_));
  AOI21_X1   g01429(.A1(new_n3844_), .A2(pi0039), .B(new_n3878_), .ZN(new_n3879_));
  OAI21_X1   g01430(.A1(new_n3876_), .A2(new_n3879_), .B(pi1142), .ZN(new_n3880_));
  NOR2_X1    g01431(.A1(new_n3870_), .A2(new_n3880_), .ZN(new_n3881_));
  NAND3_X1   g01432(.A1(new_n3400_), .A2(pi0228), .A3(pi0262), .ZN(new_n3882_));
  NAND3_X1   g01433(.A1(new_n3400_), .A2(new_n3005_), .A3(new_n3811_), .ZN(new_n3883_));
  AOI21_X1   g01434(.A1(new_n3882_), .A2(new_n3883_), .B(new_n3827_), .ZN(new_n3884_));
  OAI21_X1   g01435(.A1(new_n3884_), .A2(new_n3833_), .B(new_n3840_), .ZN(new_n3885_));
  XOR2_X1    g01436(.A1(new_n3885_), .A2(new_n3846_), .Z(new_n3886_));
  AOI21_X1   g01437(.A1(new_n3822_), .A2(new_n3212_), .B(new_n3098_), .ZN(new_n3887_));
  INV_X1     g01438(.I(new_n3851_), .ZN(new_n3888_));
  OAI21_X1   g01439(.A1(new_n3888_), .A2(new_n3211_), .B(pi0100), .ZN(new_n3889_));
  AOI21_X1   g01440(.A1(new_n3886_), .A2(new_n3887_), .B(new_n3889_), .ZN(new_n3890_));
  NOR4_X1    g01441(.A1(new_n3881_), .A2(new_n3235_), .A3(new_n3455_), .A4(new_n3890_), .ZN(new_n3891_));
  OAI21_X1   g01442(.A1(new_n3881_), .A2(new_n3890_), .B(pi0087), .ZN(new_n3892_));
  NOR2_X1    g01443(.A1(new_n3892_), .A2(new_n3694_), .ZN(new_n3893_));
  OAI21_X1   g01444(.A1(new_n3893_), .A2(new_n3891_), .B(new_n3854_), .ZN(new_n3894_));
  NAND2_X1   g01445(.A1(new_n3851_), .A2(pi0075), .ZN(new_n3895_));
  AOI21_X1   g01446(.A1(new_n3894_), .A2(new_n3303_), .B(new_n3895_), .ZN(new_n3896_));
  NAND2_X1   g01447(.A1(new_n3853_), .A2(pi0092), .ZN(new_n3897_));
  XNOR2_X1   g01448(.A1(new_n3897_), .A2(new_n3172_), .ZN(new_n3898_));
  INV_X1     g01449(.I(new_n3850_), .ZN(new_n3899_));
  NAND2_X1   g01450(.A1(new_n3842_), .A2(pi0055), .ZN(new_n3900_));
  XOR2_X1    g01451(.A1(new_n3900_), .A2(new_n3605_), .Z(new_n3901_));
  NAND2_X1   g01452(.A1(new_n3901_), .A2(new_n3899_), .ZN(new_n3902_));
  NAND2_X1   g01453(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n3903_));
  AOI21_X1   g01454(.A1(new_n3902_), .A2(new_n3219_), .B(new_n3903_), .ZN(new_n3904_));
  OAI21_X1   g01455(.A1(new_n3898_), .A2(new_n3888_), .B(new_n3904_), .ZN(new_n3905_));
  NAND2_X1   g01456(.A1(new_n3842_), .A2(pi0056), .ZN(new_n3906_));
  XOR2_X1    g01457(.A1(new_n3906_), .A2(new_n3797_), .Z(new_n3907_));
  AOI21_X1   g01458(.A1(new_n3907_), .A2(new_n3899_), .B(pi0062), .ZN(new_n3908_));
  OAI21_X1   g01459(.A1(new_n3896_), .A2(new_n3905_), .B(new_n3908_), .ZN(new_n3909_));
  NAND2_X1   g01460(.A1(new_n3842_), .A2(pi0062), .ZN(new_n3910_));
  XOR2_X1    g01461(.A1(new_n3910_), .A2(new_n3594_), .Z(new_n3911_));
  NAND2_X1   g01462(.A1(new_n3911_), .A2(new_n3899_), .ZN(new_n3912_));
  NOR2_X1    g01463(.A1(new_n3370_), .A2(new_n3368_), .ZN(new_n3913_));
  NOR2_X1    g01464(.A1(new_n3899_), .A2(new_n3913_), .ZN(new_n3914_));
  NAND4_X1   g01465(.A1(new_n3909_), .A2(new_n3810_), .A3(new_n3230_), .A4(new_n3912_), .ZN(new_n3915_));
  NOR2_X1    g01466(.A1(new_n3822_), .A2(new_n3660_), .ZN(new_n3916_));
  INV_X1     g01467(.I(new_n3833_), .ZN(new_n3917_));
  NAND2_X1   g01468(.A1(new_n3837_), .A2(new_n3370_), .ZN(new_n3918_));
  AOI21_X1   g01469(.A1(new_n3918_), .A2(new_n3917_), .B(new_n3839_), .ZN(new_n3919_));
  NAND2_X1   g01470(.A1(new_n3919_), .A2(new_n3830_), .ZN(new_n3920_));
  XOR2_X1    g01471(.A1(new_n3920_), .A2(new_n3826_), .Z(new_n3921_));
  AOI21_X1   g01472(.A1(new_n3921_), .A2(pi0299), .B(new_n3916_), .ZN(new_n3922_));
  NOR2_X1    g01473(.A1(new_n3922_), .A2(new_n3474_), .ZN(new_n3923_));
  AOI21_X1   g01474(.A1(new_n3914_), .A2(pi0299), .B(new_n3916_), .ZN(new_n3924_));
  INV_X1     g01475(.I(new_n3924_), .ZN(new_n3925_));
  AOI21_X1   g01476(.A1(new_n3925_), .A2(new_n3474_), .B(new_n3923_), .ZN(new_n3926_));
  NAND2_X1   g01477(.A1(new_n3811_), .A2(pi0172), .ZN(new_n3927_));
  NAND4_X1   g01478(.A1(new_n3330_), .A2(pi0262), .A3(new_n3308_), .A4(new_n3927_), .ZN(new_n3928_));
  NAND3_X1   g01479(.A1(new_n3308_), .A2(pi0172), .A3(new_n3811_), .ZN(new_n3929_));
  NAND3_X1   g01480(.A1(new_n3928_), .A2(new_n3005_), .A3(new_n3929_), .ZN(new_n3930_));
  INV_X1     g01481(.I(new_n3309_), .ZN(new_n3931_));
  AOI21_X1   g01482(.A1(new_n3931_), .A2(new_n3865_), .B(pi0216), .ZN(new_n3932_));
  NOR2_X1    g01483(.A1(new_n3856_), .A2(new_n3832_), .ZN(new_n3933_));
  OAI21_X1   g01484(.A1(new_n3932_), .A2(new_n3933_), .B(pi0262), .ZN(new_n3934_));
  NOR2_X1    g01485(.A1(new_n3459_), .A2(new_n3934_), .ZN(new_n3935_));
  NAND4_X1   g01486(.A1(new_n3930_), .A2(pi0215), .A3(pi0299), .A4(new_n3935_), .ZN(new_n3936_));
  NAND2_X1   g01487(.A1(new_n3930_), .A2(new_n3935_), .ZN(new_n3937_));
  NAND3_X1   g01488(.A1(new_n3937_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n3938_));
  AOI21_X1   g01489(.A1(new_n3938_), .A2(new_n3936_), .B(new_n3814_), .ZN(new_n3939_));
  INV_X1     g01490(.I(new_n3871_), .ZN(new_n3940_));
  NOR3_X1    g01491(.A1(new_n3873_), .A2(new_n3818_), .A3(new_n3940_), .ZN(new_n3941_));
  OAI21_X1   g01492(.A1(new_n3939_), .A2(new_n3876_), .B(new_n3941_), .ZN(new_n3942_));
  NAND2_X1   g01493(.A1(new_n3922_), .A2(pi0039), .ZN(new_n3943_));
  AOI21_X1   g01494(.A1(new_n3942_), .A2(new_n3259_), .B(new_n3943_), .ZN(new_n3944_));
  NOR2_X1    g01495(.A1(new_n3925_), .A2(new_n3259_), .ZN(new_n3945_));
  OAI21_X1   g01496(.A1(new_n3944_), .A2(pi0100), .B(new_n3945_), .ZN(new_n3946_));
  NAND2_X1   g01497(.A1(new_n3884_), .A2(new_n3919_), .ZN(new_n3947_));
  XOR2_X1    g01498(.A1(new_n3947_), .A2(new_n3826_), .Z(new_n3948_));
  OAI21_X1   g01499(.A1(new_n3916_), .A2(new_n3211_), .B(pi0299), .ZN(new_n3949_));
  AOI21_X1   g01500(.A1(new_n3924_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n3950_));
  OAI21_X1   g01501(.A1(new_n3948_), .A2(new_n3949_), .B(new_n3950_), .ZN(new_n3951_));
  NAND4_X1   g01502(.A1(new_n3946_), .A2(pi0075), .A3(pi0087), .A4(new_n3951_), .ZN(new_n3952_));
  INV_X1     g01503(.I(new_n3694_), .ZN(new_n3953_));
  NAND2_X1   g01504(.A1(new_n3946_), .A2(new_n3951_), .ZN(new_n3954_));
  NAND3_X1   g01505(.A1(new_n3954_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n3955_));
  AOI21_X1   g01506(.A1(new_n3955_), .A2(new_n3952_), .B(new_n3926_), .ZN(new_n3956_));
  NOR2_X1    g01507(.A1(new_n3925_), .A2(new_n3235_), .ZN(new_n3957_));
  OAI21_X1   g01508(.A1(new_n3956_), .A2(pi0092), .B(new_n3957_), .ZN(new_n3958_));
  NAND2_X1   g01509(.A1(new_n3926_), .A2(pi0092), .ZN(new_n3959_));
  XOR2_X1    g01510(.A1(new_n3959_), .A2(new_n3172_), .Z(new_n3960_));
  INV_X1     g01511(.I(new_n3914_), .ZN(new_n3961_));
  NAND2_X1   g01512(.A1(new_n3921_), .A2(pi0055), .ZN(new_n3962_));
  XOR2_X1    g01513(.A1(new_n3962_), .A2(new_n3604_), .Z(new_n3963_));
  OAI21_X1   g01514(.A1(new_n3963_), .A2(new_n3961_), .B(new_n3219_), .ZN(new_n3964_));
  NOR2_X1    g01515(.A1(new_n3203_), .A2(pi0055), .ZN(new_n3965_));
  NAND2_X1   g01516(.A1(new_n3964_), .A2(new_n3965_), .ZN(new_n3966_));
  AOI21_X1   g01517(.A1(new_n3960_), .A2(new_n3924_), .B(new_n3966_), .ZN(new_n3967_));
  NAND2_X1   g01518(.A1(new_n3921_), .A2(pi0056), .ZN(new_n3968_));
  XOR2_X1    g01519(.A1(new_n3968_), .A2(new_n3599_), .Z(new_n3969_));
  OAI21_X1   g01520(.A1(new_n3969_), .A2(new_n3961_), .B(new_n3201_), .ZN(new_n3970_));
  AOI21_X1   g01521(.A1(new_n3958_), .A2(new_n3967_), .B(new_n3970_), .ZN(new_n3971_));
  INV_X1     g01522(.I(new_n3594_), .ZN(new_n3972_));
  NAND2_X1   g01523(.A1(new_n3921_), .A2(pi0062), .ZN(new_n3973_));
  XOR2_X1    g01524(.A1(new_n3973_), .A2(new_n3972_), .Z(new_n3974_));
  NOR2_X1    g01525(.A1(new_n3426_), .A2(new_n3810_), .ZN(new_n3975_));
  OAI21_X1   g01526(.A1(new_n3974_), .A2(new_n3961_), .B(new_n3975_), .ZN(new_n3976_));
  OAI21_X1   g01527(.A1(new_n3971_), .A2(new_n3976_), .B(new_n3915_), .ZN(po0157));
  NAND2_X1   g01528(.A1(new_n2820_), .A2(pi0861), .ZN(new_n3978_));
  AOI21_X1   g01529(.A1(pi0224), .A2(pi0270), .B(pi0222), .ZN(new_n3979_));
  INV_X1     g01530(.I(pi1141), .ZN(new_n3980_));
  NAND3_X1   g01531(.A1(new_n3103_), .A2(pi0222), .A3(pi0935), .ZN(new_n3981_));
  INV_X1     g01532(.I(pi0935), .ZN(new_n3982_));
  NAND3_X1   g01533(.A1(new_n3344_), .A2(pi0222), .A3(new_n3982_), .ZN(new_n3983_));
  AOI21_X1   g01534(.A1(new_n3983_), .A2(new_n3981_), .B(new_n3980_), .ZN(new_n3984_));
  AOI21_X1   g01535(.A1(new_n3984_), .A2(new_n3979_), .B(pi0224), .ZN(new_n3985_));
  OAI21_X1   g01536(.A1(new_n3985_), .A2(new_n3978_), .B(pi0223), .ZN(new_n3986_));
  XOR2_X1    g01537(.A1(new_n3986_), .A2(new_n3565_), .Z(new_n3987_));
  NAND2_X1   g01538(.A1(new_n3987_), .A2(pi1141), .ZN(new_n3988_));
  INV_X1     g01539(.I(pi0171), .ZN(new_n3989_));
  NAND3_X1   g01540(.A1(new_n3160_), .A2(pi0228), .A3(pi0861), .ZN(new_n3990_));
  INV_X1     g01541(.I(pi0861), .ZN(new_n3991_));
  NAND3_X1   g01542(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n3991_), .ZN(new_n3992_));
  AOI21_X1   g01543(.A1(new_n3990_), .A2(new_n3992_), .B(new_n3989_), .ZN(new_n3993_));
  NAND4_X1   g01544(.A1(new_n2820_), .A2(pi0105), .A3(pi0228), .A4(pi0861), .ZN(new_n3994_));
  NAND3_X1   g01545(.A1(new_n3978_), .A2(new_n3004_), .A3(pi0228), .ZN(new_n3995_));
  AOI21_X1   g01546(.A1(new_n3995_), .A2(new_n3994_), .B(new_n3989_), .ZN(new_n3996_));
  NOR2_X1    g01547(.A1(new_n3996_), .A2(pi0216), .ZN(new_n3997_));
  INV_X1     g01548(.I(new_n3997_), .ZN(new_n3998_));
  NOR2_X1    g01549(.A1(new_n3121_), .A2(pi0935), .ZN(new_n3999_));
  XOR2_X1    g01550(.A1(new_n3356_), .A2(new_n3999_), .Z(new_n4000_));
  AOI21_X1   g01551(.A1(pi0216), .A2(pi0270), .B(pi0221), .ZN(new_n4001_));
  NAND3_X1   g01552(.A1(new_n4000_), .A2(pi1141), .A3(new_n4001_), .ZN(new_n4002_));
  NAND2_X1   g01553(.A1(new_n3998_), .A2(new_n4002_), .ZN(new_n4003_));
  NAND3_X1   g01554(.A1(new_n4003_), .A2(new_n3993_), .A3(new_n3111_), .ZN(new_n4004_));
  OAI21_X1   g01555(.A1(new_n3111_), .A2(pi1141), .B(new_n4004_), .ZN(new_n4005_));
  OAI21_X1   g01556(.A1(new_n4005_), .A2(new_n3098_), .B(new_n3988_), .ZN(new_n4006_));
  INV_X1     g01557(.I(new_n3988_), .ZN(new_n4007_));
  NAND2_X1   g01558(.A1(new_n4000_), .A2(pi1141), .ZN(new_n4008_));
  NAND2_X1   g01559(.A1(new_n4008_), .A2(pi0215), .ZN(new_n4009_));
  NAND2_X1   g01560(.A1(new_n3997_), .A2(new_n4001_), .ZN(new_n4010_));
  NAND2_X1   g01561(.A1(new_n4010_), .A2(new_n3005_), .ZN(new_n4011_));
  NAND4_X1   g01562(.A1(new_n4011_), .A2(pi0171), .A3(pi0215), .A4(pi1141), .ZN(new_n4012_));
  XNOR2_X1   g01563(.A1(new_n4012_), .A2(new_n4009_), .ZN(new_n4013_));
  AOI21_X1   g01564(.A1(new_n4013_), .A2(pi0299), .B(new_n4007_), .ZN(new_n4014_));
  NOR2_X1    g01565(.A1(new_n4014_), .A2(new_n3134_), .ZN(new_n4015_));
  AOI21_X1   g01566(.A1(new_n3134_), .A2(new_n4006_), .B(new_n4015_), .ZN(new_n4016_));
  NAND2_X1   g01567(.A1(new_n3307_), .A2(pi0861), .ZN(new_n4017_));
  AOI21_X1   g01568(.A1(new_n3459_), .A2(new_n3989_), .B(new_n4017_), .ZN(new_n4018_));
  NAND3_X1   g01569(.A1(new_n3330_), .A2(pi0171), .A3(pi0861), .ZN(new_n4019_));
  NAND3_X1   g01570(.A1(new_n3862_), .A2(new_n3989_), .A3(pi0861), .ZN(new_n4020_));
  AOI21_X1   g01571(.A1(new_n4020_), .A2(new_n4019_), .B(new_n3308_), .ZN(new_n4021_));
  NAND2_X1   g01572(.A1(new_n3931_), .A2(new_n3996_), .ZN(new_n4022_));
  NAND2_X1   g01573(.A1(new_n4022_), .A2(new_n3011_), .ZN(new_n4023_));
  AOI21_X1   g01574(.A1(new_n4023_), .A2(new_n4002_), .B(pi0228), .ZN(new_n4024_));
  OAI21_X1   g01575(.A1(new_n4021_), .A2(new_n4018_), .B(new_n4024_), .ZN(new_n4025_));
  OR3_X2     g01576(.A1(new_n4025_), .A2(new_n3111_), .A3(new_n3098_), .Z(new_n4026_));
  NAND3_X1   g01577(.A1(new_n4025_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n4027_));
  AOI21_X1   g01578(.A1(new_n4026_), .A2(new_n4027_), .B(new_n3980_), .ZN(new_n4028_));
  AOI21_X1   g01579(.A1(pi0223), .A2(pi1141), .B(pi0299), .ZN(new_n4029_));
  AOI21_X1   g01580(.A1(new_n3979_), .A2(pi0224), .B(pi0861), .ZN(new_n4030_));
  NOR2_X1    g01581(.A1(new_n3702_), .A2(new_n4030_), .ZN(new_n4031_));
  NOR3_X1    g01582(.A1(new_n4031_), .A2(new_n3090_), .A3(new_n3984_), .ZN(new_n4032_));
  OAI21_X1   g01583(.A1(new_n4032_), .A2(new_n3979_), .B(new_n3306_), .ZN(new_n4033_));
  AOI21_X1   g01584(.A1(new_n4033_), .A2(new_n4029_), .B(pi0039), .ZN(new_n4034_));
  INV_X1     g01585(.I(new_n4029_), .ZN(new_n4035_));
  NOR3_X1    g01586(.A1(new_n4031_), .A2(new_n3984_), .A3(new_n4035_), .ZN(new_n4036_));
  OAI21_X1   g01587(.A1(new_n4028_), .A2(new_n4034_), .B(new_n4036_), .ZN(new_n4037_));
  OR2_X2     g01588(.A1(new_n4006_), .A2(new_n3183_), .Z(new_n4038_));
  AOI21_X1   g01589(.A1(new_n4037_), .A2(new_n3259_), .B(new_n4038_), .ZN(new_n4039_));
  INV_X1     g01590(.I(new_n4014_), .ZN(new_n4040_));
  NOR2_X1    g01591(.A1(new_n4040_), .A2(new_n3259_), .ZN(new_n4041_));
  OAI21_X1   g01592(.A1(new_n4039_), .A2(pi0100), .B(new_n4041_), .ZN(new_n4042_));
  NAND3_X1   g01593(.A1(new_n3400_), .A2(pi0228), .A3(pi0861), .ZN(new_n4043_));
  NAND3_X1   g01594(.A1(new_n3400_), .A2(new_n3005_), .A3(new_n3991_), .ZN(new_n4044_));
  AOI21_X1   g01595(.A1(new_n4043_), .A2(new_n4044_), .B(new_n3989_), .ZN(new_n4045_));
  AOI21_X1   g01596(.A1(new_n4045_), .A2(new_n4003_), .B(new_n3098_), .ZN(new_n4046_));
  XOR2_X1    g01597(.A1(new_n4046_), .A2(new_n3855_), .Z(new_n4047_));
  NOR2_X1    g01598(.A1(new_n4047_), .A2(new_n3980_), .ZN(new_n4048_));
  NAND2_X1   g01599(.A1(new_n3988_), .A2(new_n3211_), .ZN(new_n4049_));
  AOI21_X1   g01600(.A1(new_n4014_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4050_));
  OAI21_X1   g01601(.A1(new_n4048_), .A2(new_n4049_), .B(new_n4050_), .ZN(new_n4051_));
  NAND4_X1   g01602(.A1(new_n4042_), .A2(pi0075), .A3(pi0087), .A4(new_n4051_), .ZN(new_n4052_));
  NAND2_X1   g01603(.A1(new_n4042_), .A2(new_n4051_), .ZN(new_n4053_));
  NAND3_X1   g01604(.A1(new_n4053_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4054_));
  AOI21_X1   g01605(.A1(new_n4054_), .A2(new_n4052_), .B(new_n4016_), .ZN(new_n4055_));
  NOR2_X1    g01606(.A1(new_n4040_), .A2(new_n3235_), .ZN(new_n4056_));
  OAI21_X1   g01607(.A1(new_n4055_), .A2(pi0092), .B(new_n4056_), .ZN(new_n4057_));
  NAND2_X1   g01608(.A1(new_n4016_), .A2(pi0092), .ZN(new_n4058_));
  XNOR2_X1   g01609(.A1(new_n4058_), .A2(new_n3172_), .ZN(new_n4059_));
  NOR2_X1    g01610(.A1(new_n4059_), .A2(new_n4040_), .ZN(new_n4060_));
  INV_X1     g01611(.I(new_n4013_), .ZN(new_n4061_));
  NOR2_X1    g01612(.A1(new_n4005_), .A2(new_n3201_), .ZN(new_n4062_));
  XOR2_X1    g01613(.A1(new_n4062_), .A2(new_n3972_), .Z(new_n4063_));
  INV_X1     g01614(.I(pi0241), .ZN(new_n4064_));
  NAND2_X1   g01615(.A1(new_n3230_), .A2(new_n4064_), .ZN(new_n4065_));
  AOI21_X1   g01616(.A1(new_n4063_), .A2(new_n4061_), .B(new_n4065_), .ZN(new_n4066_));
  NOR2_X1    g01617(.A1(new_n4005_), .A2(new_n3219_), .ZN(new_n4067_));
  XOR2_X1    g01618(.A1(new_n4067_), .A2(new_n3797_), .Z(new_n4068_));
  OAI21_X1   g01619(.A1(new_n4068_), .A2(new_n4013_), .B(new_n3201_), .ZN(new_n4069_));
  NOR2_X1    g01620(.A1(new_n4066_), .A2(new_n4069_), .ZN(new_n4070_));
  NOR2_X1    g01621(.A1(new_n4005_), .A2(new_n3258_), .ZN(new_n4071_));
  XOR2_X1    g01622(.A1(new_n4071_), .A2(new_n3604_), .Z(new_n4072_));
  AOI21_X1   g01623(.A1(new_n4072_), .A2(new_n4061_), .B(pi0056), .ZN(new_n4073_));
  NAND2_X1   g01624(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n4074_));
  NOR4_X1    g01625(.A1(new_n4060_), .A2(new_n4070_), .A3(new_n4073_), .A4(new_n4074_), .ZN(new_n4075_));
  NOR2_X1    g01626(.A1(new_n4061_), .A2(new_n3230_), .ZN(new_n4076_));
  AOI21_X1   g01627(.A1(pi0216), .A2(pi0270), .B(new_n3612_), .ZN(new_n4077_));
  NAND2_X1   g01628(.A1(new_n4077_), .A2(pi0241), .ZN(new_n4078_));
  NOR2_X1    g01629(.A1(new_n4007_), .A2(new_n3385_), .ZN(new_n4079_));
  NOR2_X1    g01630(.A1(new_n3997_), .A2(new_n4001_), .ZN(new_n4080_));
  INV_X1     g01631(.I(new_n4080_), .ZN(new_n4081_));
  NOR3_X1    g01632(.A1(new_n3370_), .A2(new_n3111_), .A3(new_n3980_), .ZN(new_n4082_));
  OAI21_X1   g01633(.A1(new_n4081_), .A2(new_n3993_), .B(new_n4082_), .ZN(new_n4083_));
  XNOR2_X1   g01634(.A1(new_n4083_), .A2(new_n4009_), .ZN(new_n4084_));
  NAND2_X1   g01635(.A1(new_n4084_), .A2(pi0299), .ZN(new_n4085_));
  NAND2_X1   g01636(.A1(new_n4085_), .A2(new_n4079_), .ZN(new_n4086_));
  NOR2_X1    g01637(.A1(new_n4013_), .A2(new_n4077_), .ZN(new_n4087_));
  OAI21_X1   g01638(.A1(new_n4087_), .A2(new_n3098_), .B(new_n4079_), .ZN(new_n4088_));
  INV_X1     g01639(.I(new_n4088_), .ZN(new_n4089_));
  NOR2_X1    g01640(.A1(new_n4089_), .A2(new_n3134_), .ZN(new_n4090_));
  AOI21_X1   g01641(.A1(new_n4086_), .A2(new_n3134_), .B(new_n4090_), .ZN(new_n4091_));
  INV_X1     g01642(.I(new_n4091_), .ZN(new_n4092_));
  NAND3_X1   g01643(.A1(new_n3696_), .A2(pi0171), .A3(pi0861), .ZN(new_n4093_));
  NAND3_X1   g01644(.A1(new_n3459_), .A2(pi0171), .A3(new_n3991_), .ZN(new_n4094_));
  NAND2_X1   g01645(.A1(new_n3307_), .A2(pi0171), .ZN(new_n4095_));
  AOI21_X1   g01646(.A1(new_n4093_), .A2(new_n4094_), .B(new_n4095_), .ZN(new_n4096_));
  NAND2_X1   g01647(.A1(pi0228), .A2(pi0861), .ZN(new_n4097_));
  AOI21_X1   g01648(.A1(new_n3703_), .A2(new_n3998_), .B(new_n4097_), .ZN(new_n4098_));
  OAI21_X1   g01649(.A1(new_n4096_), .A2(new_n3330_), .B(new_n4098_), .ZN(new_n4099_));
  NAND2_X1   g01650(.A1(new_n4099_), .A2(new_n4001_), .ZN(new_n4100_));
  AOI21_X1   g01651(.A1(new_n4100_), .A2(new_n4008_), .B(new_n3098_), .ZN(new_n4101_));
  XOR2_X1    g01652(.A1(new_n4101_), .A2(new_n3855_), .Z(new_n4102_));
  NOR2_X1    g01653(.A1(pi0038), .A2(pi0100), .ZN(new_n4103_));
  INV_X1     g01654(.I(new_n4103_), .ZN(new_n4104_));
  AOI21_X1   g01655(.A1(new_n4086_), .A2(pi0039), .B(new_n4104_), .ZN(new_n4105_));
  OAI21_X1   g01656(.A1(new_n4034_), .A2(new_n4105_), .B(pi1141), .ZN(new_n4106_));
  NOR2_X1    g01657(.A1(new_n4102_), .A2(new_n4106_), .ZN(new_n4107_));
  OAI21_X1   g01658(.A1(new_n4045_), .A2(new_n4081_), .B(new_n4082_), .ZN(new_n4108_));
  XOR2_X1    g01659(.A1(new_n4108_), .A2(new_n4009_), .Z(new_n4109_));
  NOR2_X1    g01660(.A1(new_n4079_), .A2(new_n3211_), .ZN(new_n4110_));
  NOR2_X1    g01661(.A1(new_n4110_), .A2(new_n3098_), .ZN(new_n4111_));
  OAI21_X1   g01662(.A1(new_n4088_), .A2(new_n3211_), .B(pi0100), .ZN(new_n4112_));
  AOI21_X1   g01663(.A1(new_n4109_), .A2(new_n4111_), .B(new_n4112_), .ZN(new_n4113_));
  NOR4_X1    g01664(.A1(new_n4107_), .A2(new_n3235_), .A3(new_n3455_), .A4(new_n4113_), .ZN(new_n4114_));
  OAI21_X1   g01665(.A1(new_n4107_), .A2(new_n4113_), .B(pi0087), .ZN(new_n4115_));
  NOR2_X1    g01666(.A1(new_n4115_), .A2(new_n3694_), .ZN(new_n4116_));
  OAI21_X1   g01667(.A1(new_n4116_), .A2(new_n4114_), .B(new_n4092_), .ZN(new_n4117_));
  NAND2_X1   g01668(.A1(new_n4089_), .A2(pi0075), .ZN(new_n4118_));
  AOI21_X1   g01669(.A1(new_n4117_), .A2(new_n3303_), .B(new_n4118_), .ZN(new_n4119_));
  NAND2_X1   g01670(.A1(new_n4091_), .A2(pi0092), .ZN(new_n4120_));
  XOR2_X1    g01671(.A1(new_n4120_), .A2(new_n3172_), .Z(new_n4121_));
  NAND2_X1   g01672(.A1(new_n4121_), .A2(new_n4089_), .ZN(new_n4122_));
  NAND2_X1   g01673(.A1(new_n4084_), .A2(pi0062), .ZN(new_n4123_));
  XOR2_X1    g01674(.A1(new_n4123_), .A2(new_n3594_), .Z(new_n4124_));
  NAND2_X1   g01675(.A1(new_n4124_), .A2(new_n4087_), .ZN(new_n4125_));
  NAND3_X1   g01676(.A1(new_n4125_), .A2(pi0241), .A3(new_n3230_), .ZN(new_n4126_));
  NAND2_X1   g01677(.A1(new_n4084_), .A2(pi0056), .ZN(new_n4127_));
  XOR2_X1    g01678(.A1(new_n4127_), .A2(new_n3797_), .Z(new_n4128_));
  AOI21_X1   g01679(.A1(new_n4128_), .A2(new_n4087_), .B(pi0062), .ZN(new_n4129_));
  NAND2_X1   g01680(.A1(new_n4126_), .A2(new_n4129_), .ZN(new_n4130_));
  NAND2_X1   g01681(.A1(new_n4084_), .A2(pi0055), .ZN(new_n4131_));
  XOR2_X1    g01682(.A1(new_n4131_), .A2(new_n3605_), .Z(new_n4132_));
  NAND2_X1   g01683(.A1(new_n4132_), .A2(new_n4087_), .ZN(new_n4133_));
  NAND2_X1   g01684(.A1(new_n4133_), .A2(new_n3219_), .ZN(new_n4134_));
  NOR2_X1    g01685(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4135_));
  NAND4_X1   g01686(.A1(new_n4122_), .A2(new_n4130_), .A3(new_n4134_), .A4(new_n4135_), .ZN(new_n4136_));
  OAI22_X1   g01687(.A1(new_n4119_), .A2(new_n4136_), .B1(new_n4076_), .B2(new_n4078_), .ZN(new_n4137_));
  AOI21_X1   g01688(.A1(new_n4057_), .A2(new_n4075_), .B(new_n4137_), .ZN(po0158));
  NAND2_X1   g01689(.A1(new_n2820_), .A2(pi0869), .ZN(new_n4139_));
  AOI21_X1   g01690(.A1(pi0224), .A2(pi0282), .B(pi0222), .ZN(new_n4140_));
  INV_X1     g01691(.I(pi1140), .ZN(new_n4141_));
  NAND3_X1   g01692(.A1(new_n3103_), .A2(pi0222), .A3(pi0921), .ZN(new_n4142_));
  INV_X1     g01693(.I(pi0921), .ZN(new_n4143_));
  NAND3_X1   g01694(.A1(new_n3344_), .A2(pi0222), .A3(new_n4143_), .ZN(new_n4144_));
  AOI21_X1   g01695(.A1(new_n4144_), .A2(new_n4142_), .B(new_n4141_), .ZN(new_n4145_));
  AOI21_X1   g01696(.A1(new_n4145_), .A2(new_n4140_), .B(pi0224), .ZN(new_n4146_));
  OAI21_X1   g01697(.A1(new_n4146_), .A2(new_n4139_), .B(pi0223), .ZN(new_n4147_));
  XOR2_X1    g01698(.A1(new_n4147_), .A2(new_n3565_), .Z(new_n4148_));
  NAND2_X1   g01699(.A1(new_n4148_), .A2(pi1140), .ZN(new_n4149_));
  INV_X1     g01700(.I(pi0170), .ZN(new_n4150_));
  NAND3_X1   g01701(.A1(new_n3160_), .A2(pi0228), .A3(pi0869), .ZN(new_n4151_));
  INV_X1     g01702(.I(pi0869), .ZN(new_n4152_));
  NAND3_X1   g01703(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n4152_), .ZN(new_n4153_));
  AOI21_X1   g01704(.A1(new_n4151_), .A2(new_n4153_), .B(new_n4150_), .ZN(new_n4154_));
  NAND4_X1   g01705(.A1(new_n2820_), .A2(pi0105), .A3(pi0228), .A4(pi0869), .ZN(new_n4155_));
  NAND3_X1   g01706(.A1(new_n4139_), .A2(new_n3004_), .A3(pi0228), .ZN(new_n4156_));
  AOI21_X1   g01707(.A1(new_n4156_), .A2(new_n4155_), .B(new_n4150_), .ZN(new_n4157_));
  NOR2_X1    g01708(.A1(new_n4157_), .A2(pi0216), .ZN(new_n4158_));
  INV_X1     g01709(.I(new_n4158_), .ZN(new_n4159_));
  NOR2_X1    g01710(.A1(new_n3121_), .A2(pi0921), .ZN(new_n4160_));
  XOR2_X1    g01711(.A1(new_n3356_), .A2(new_n4160_), .Z(new_n4161_));
  AOI21_X1   g01712(.A1(pi0216), .A2(pi0282), .B(pi0221), .ZN(new_n4162_));
  NAND3_X1   g01713(.A1(new_n4161_), .A2(pi1140), .A3(new_n4162_), .ZN(new_n4163_));
  NAND2_X1   g01714(.A1(new_n4159_), .A2(new_n4163_), .ZN(new_n4164_));
  NAND3_X1   g01715(.A1(new_n4164_), .A2(new_n4154_), .A3(new_n3111_), .ZN(new_n4165_));
  OAI21_X1   g01716(.A1(new_n3111_), .A2(pi1140), .B(new_n4165_), .ZN(new_n4166_));
  OAI21_X1   g01717(.A1(new_n4166_), .A2(new_n3098_), .B(new_n4149_), .ZN(new_n4167_));
  INV_X1     g01718(.I(new_n4149_), .ZN(new_n4168_));
  NAND2_X1   g01719(.A1(new_n4161_), .A2(pi1140), .ZN(new_n4169_));
  NAND2_X1   g01720(.A1(new_n4169_), .A2(pi0215), .ZN(new_n4170_));
  NAND2_X1   g01721(.A1(new_n4158_), .A2(new_n4162_), .ZN(new_n4171_));
  NAND2_X1   g01722(.A1(new_n4171_), .A2(new_n3005_), .ZN(new_n4172_));
  NAND4_X1   g01723(.A1(new_n4172_), .A2(pi0170), .A3(pi0215), .A4(pi1140), .ZN(new_n4173_));
  XNOR2_X1   g01724(.A1(new_n4173_), .A2(new_n4170_), .ZN(new_n4174_));
  AOI21_X1   g01725(.A1(new_n4174_), .A2(pi0299), .B(new_n4168_), .ZN(new_n4175_));
  NOR2_X1    g01726(.A1(new_n4175_), .A2(new_n3134_), .ZN(new_n4176_));
  AOI21_X1   g01727(.A1(new_n3134_), .A2(new_n4167_), .B(new_n4176_), .ZN(new_n4177_));
  NAND2_X1   g01728(.A1(new_n3307_), .A2(pi0869), .ZN(new_n4178_));
  AOI21_X1   g01729(.A1(new_n3459_), .A2(new_n4150_), .B(new_n4178_), .ZN(new_n4179_));
  NAND3_X1   g01730(.A1(new_n3330_), .A2(pi0170), .A3(pi0869), .ZN(new_n4180_));
  NAND3_X1   g01731(.A1(new_n3862_), .A2(new_n4150_), .A3(pi0869), .ZN(new_n4181_));
  AOI21_X1   g01732(.A1(new_n4181_), .A2(new_n4180_), .B(new_n3308_), .ZN(new_n4182_));
  NAND2_X1   g01733(.A1(new_n3931_), .A2(new_n4157_), .ZN(new_n4183_));
  NAND2_X1   g01734(.A1(new_n4183_), .A2(new_n3011_), .ZN(new_n4184_));
  AOI21_X1   g01735(.A1(new_n4184_), .A2(new_n4163_), .B(pi0228), .ZN(new_n4185_));
  OAI21_X1   g01736(.A1(new_n4182_), .A2(new_n4179_), .B(new_n4185_), .ZN(new_n4186_));
  OR3_X2     g01737(.A1(new_n4186_), .A2(new_n3111_), .A3(new_n3098_), .Z(new_n4187_));
  NAND3_X1   g01738(.A1(new_n4186_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n4188_));
  AOI21_X1   g01739(.A1(new_n4187_), .A2(new_n4188_), .B(new_n4141_), .ZN(new_n4189_));
  AOI21_X1   g01740(.A1(pi0223), .A2(pi1140), .B(pi0299), .ZN(new_n4190_));
  AOI21_X1   g01741(.A1(new_n4140_), .A2(pi0224), .B(pi0869), .ZN(new_n4191_));
  NOR2_X1    g01742(.A1(new_n3702_), .A2(new_n4191_), .ZN(new_n4192_));
  NOR3_X1    g01743(.A1(new_n4192_), .A2(new_n3090_), .A3(new_n4145_), .ZN(new_n4193_));
  OAI21_X1   g01744(.A1(new_n4193_), .A2(new_n4140_), .B(new_n3306_), .ZN(new_n4194_));
  AOI21_X1   g01745(.A1(new_n4194_), .A2(new_n4190_), .B(pi0039), .ZN(new_n4195_));
  INV_X1     g01746(.I(new_n4190_), .ZN(new_n4196_));
  NOR3_X1    g01747(.A1(new_n4192_), .A2(new_n4145_), .A3(new_n4196_), .ZN(new_n4197_));
  OAI21_X1   g01748(.A1(new_n4189_), .A2(new_n4195_), .B(new_n4197_), .ZN(new_n4198_));
  OR2_X2     g01749(.A1(new_n4167_), .A2(new_n3183_), .Z(new_n4199_));
  AOI21_X1   g01750(.A1(new_n4198_), .A2(new_n3259_), .B(new_n4199_), .ZN(new_n4200_));
  INV_X1     g01751(.I(new_n4175_), .ZN(new_n4201_));
  NOR2_X1    g01752(.A1(new_n4201_), .A2(new_n3259_), .ZN(new_n4202_));
  OAI21_X1   g01753(.A1(new_n4200_), .A2(pi0100), .B(new_n4202_), .ZN(new_n4203_));
  NAND3_X1   g01754(.A1(new_n3400_), .A2(pi0228), .A3(pi0869), .ZN(new_n4204_));
  NAND3_X1   g01755(.A1(new_n3400_), .A2(new_n3005_), .A3(new_n4152_), .ZN(new_n4205_));
  AOI21_X1   g01756(.A1(new_n4204_), .A2(new_n4205_), .B(new_n4150_), .ZN(new_n4206_));
  AOI21_X1   g01757(.A1(new_n4206_), .A2(new_n4164_), .B(new_n3098_), .ZN(new_n4207_));
  XOR2_X1    g01758(.A1(new_n4207_), .A2(new_n3855_), .Z(new_n4208_));
  NOR2_X1    g01759(.A1(new_n4208_), .A2(new_n4141_), .ZN(new_n4209_));
  NAND2_X1   g01760(.A1(new_n4149_), .A2(new_n3211_), .ZN(new_n4210_));
  AOI21_X1   g01761(.A1(new_n4175_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4211_));
  OAI21_X1   g01762(.A1(new_n4209_), .A2(new_n4210_), .B(new_n4211_), .ZN(new_n4212_));
  NAND4_X1   g01763(.A1(new_n4203_), .A2(pi0075), .A3(pi0087), .A4(new_n4212_), .ZN(new_n4213_));
  NAND2_X1   g01764(.A1(new_n4203_), .A2(new_n4212_), .ZN(new_n4214_));
  NAND3_X1   g01765(.A1(new_n4214_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4215_));
  AOI21_X1   g01766(.A1(new_n4215_), .A2(new_n4213_), .B(new_n4177_), .ZN(new_n4216_));
  NOR2_X1    g01767(.A1(new_n4201_), .A2(new_n3235_), .ZN(new_n4217_));
  OAI21_X1   g01768(.A1(new_n4216_), .A2(pi0092), .B(new_n4217_), .ZN(new_n4218_));
  NAND2_X1   g01769(.A1(new_n4177_), .A2(pi0092), .ZN(new_n4219_));
  XNOR2_X1   g01770(.A1(new_n4219_), .A2(new_n3172_), .ZN(new_n4220_));
  NOR2_X1    g01771(.A1(new_n4220_), .A2(new_n4201_), .ZN(new_n4221_));
  INV_X1     g01772(.I(new_n4174_), .ZN(new_n4222_));
  NOR2_X1    g01773(.A1(new_n4166_), .A2(new_n3201_), .ZN(new_n4223_));
  XOR2_X1    g01774(.A1(new_n4223_), .A2(new_n3972_), .Z(new_n4224_));
  INV_X1     g01775(.I(pi0248), .ZN(new_n4225_));
  NAND2_X1   g01776(.A1(new_n3230_), .A2(new_n4225_), .ZN(new_n4226_));
  AOI21_X1   g01777(.A1(new_n4224_), .A2(new_n4222_), .B(new_n4226_), .ZN(new_n4227_));
  NOR2_X1    g01778(.A1(new_n4166_), .A2(new_n3219_), .ZN(new_n4228_));
  XOR2_X1    g01779(.A1(new_n4228_), .A2(new_n3797_), .Z(new_n4229_));
  OAI21_X1   g01780(.A1(new_n4229_), .A2(new_n4174_), .B(new_n3201_), .ZN(new_n4230_));
  NOR2_X1    g01781(.A1(new_n4227_), .A2(new_n4230_), .ZN(new_n4231_));
  NOR2_X1    g01782(.A1(new_n4166_), .A2(new_n3258_), .ZN(new_n4232_));
  XOR2_X1    g01783(.A1(new_n4232_), .A2(new_n3604_), .Z(new_n4233_));
  AOI21_X1   g01784(.A1(new_n4233_), .A2(new_n4222_), .B(pi0056), .ZN(new_n4234_));
  NAND2_X1   g01785(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n4235_));
  NOR4_X1    g01786(.A1(new_n4221_), .A2(new_n4231_), .A3(new_n4234_), .A4(new_n4235_), .ZN(new_n4236_));
  NOR2_X1    g01787(.A1(new_n4222_), .A2(new_n3230_), .ZN(new_n4237_));
  AOI21_X1   g01788(.A1(pi0216), .A2(pi0282), .B(new_n3612_), .ZN(new_n4238_));
  NAND2_X1   g01789(.A1(new_n4238_), .A2(pi0248), .ZN(new_n4239_));
  NOR2_X1    g01790(.A1(new_n4168_), .A2(new_n3385_), .ZN(new_n4240_));
  NOR2_X1    g01791(.A1(new_n4158_), .A2(new_n4162_), .ZN(new_n4241_));
  INV_X1     g01792(.I(new_n4241_), .ZN(new_n4242_));
  NOR3_X1    g01793(.A1(new_n3370_), .A2(new_n3111_), .A3(new_n4141_), .ZN(new_n4243_));
  OAI21_X1   g01794(.A1(new_n4242_), .A2(new_n4154_), .B(new_n4243_), .ZN(new_n4244_));
  XNOR2_X1   g01795(.A1(new_n4244_), .A2(new_n4170_), .ZN(new_n4245_));
  NAND2_X1   g01796(.A1(new_n4245_), .A2(pi0299), .ZN(new_n4246_));
  NAND2_X1   g01797(.A1(new_n4246_), .A2(new_n4240_), .ZN(new_n4247_));
  NOR2_X1    g01798(.A1(new_n4174_), .A2(new_n4238_), .ZN(new_n4248_));
  OAI21_X1   g01799(.A1(new_n4248_), .A2(new_n3098_), .B(new_n4240_), .ZN(new_n4249_));
  INV_X1     g01800(.I(new_n4249_), .ZN(new_n4250_));
  NOR2_X1    g01801(.A1(new_n4250_), .A2(new_n3134_), .ZN(new_n4251_));
  AOI21_X1   g01802(.A1(new_n4247_), .A2(new_n3134_), .B(new_n4251_), .ZN(new_n4252_));
  INV_X1     g01803(.I(new_n4252_), .ZN(new_n4253_));
  NAND3_X1   g01804(.A1(new_n3696_), .A2(pi0170), .A3(pi0869), .ZN(new_n4254_));
  NAND3_X1   g01805(.A1(new_n3459_), .A2(pi0170), .A3(new_n4152_), .ZN(new_n4255_));
  NAND2_X1   g01806(.A1(new_n3307_), .A2(pi0170), .ZN(new_n4256_));
  AOI21_X1   g01807(.A1(new_n4254_), .A2(new_n4255_), .B(new_n4256_), .ZN(new_n4257_));
  NAND2_X1   g01808(.A1(pi0228), .A2(pi0869), .ZN(new_n4258_));
  AOI21_X1   g01809(.A1(new_n3703_), .A2(new_n4159_), .B(new_n4258_), .ZN(new_n4259_));
  OAI21_X1   g01810(.A1(new_n4257_), .A2(new_n3330_), .B(new_n4259_), .ZN(new_n4260_));
  NAND2_X1   g01811(.A1(new_n4260_), .A2(new_n4162_), .ZN(new_n4261_));
  AOI21_X1   g01812(.A1(new_n4261_), .A2(new_n4169_), .B(new_n3098_), .ZN(new_n4262_));
  XOR2_X1    g01813(.A1(new_n4262_), .A2(new_n3855_), .Z(new_n4263_));
  NOR2_X1    g01814(.A1(pi0038), .A2(pi0100), .ZN(new_n4264_));
  INV_X1     g01815(.I(new_n4264_), .ZN(new_n4265_));
  AOI21_X1   g01816(.A1(new_n4247_), .A2(pi0039), .B(new_n4265_), .ZN(new_n4266_));
  OAI21_X1   g01817(.A1(new_n4195_), .A2(new_n4266_), .B(pi1140), .ZN(new_n4267_));
  NOR2_X1    g01818(.A1(new_n4263_), .A2(new_n4267_), .ZN(new_n4268_));
  OAI21_X1   g01819(.A1(new_n4206_), .A2(new_n4242_), .B(new_n4243_), .ZN(new_n4269_));
  XOR2_X1    g01820(.A1(new_n4269_), .A2(new_n4170_), .Z(new_n4270_));
  NOR2_X1    g01821(.A1(new_n4240_), .A2(new_n3211_), .ZN(new_n4271_));
  NOR2_X1    g01822(.A1(new_n4271_), .A2(new_n3098_), .ZN(new_n4272_));
  OAI21_X1   g01823(.A1(new_n4249_), .A2(new_n3211_), .B(pi0100), .ZN(new_n4273_));
  AOI21_X1   g01824(.A1(new_n4270_), .A2(new_n4272_), .B(new_n4273_), .ZN(new_n4274_));
  NOR4_X1    g01825(.A1(new_n4268_), .A2(new_n3235_), .A3(new_n3455_), .A4(new_n4274_), .ZN(new_n4275_));
  OAI21_X1   g01826(.A1(new_n4268_), .A2(new_n4274_), .B(pi0087), .ZN(new_n4276_));
  NOR2_X1    g01827(.A1(new_n4276_), .A2(new_n3694_), .ZN(new_n4277_));
  OAI21_X1   g01828(.A1(new_n4277_), .A2(new_n4275_), .B(new_n4253_), .ZN(new_n4278_));
  NAND2_X1   g01829(.A1(new_n4250_), .A2(pi0075), .ZN(new_n4279_));
  AOI21_X1   g01830(.A1(new_n4278_), .A2(new_n3303_), .B(new_n4279_), .ZN(new_n4280_));
  NAND2_X1   g01831(.A1(new_n4252_), .A2(pi0092), .ZN(new_n4281_));
  XOR2_X1    g01832(.A1(new_n4281_), .A2(new_n3172_), .Z(new_n4282_));
  NAND2_X1   g01833(.A1(new_n4282_), .A2(new_n4250_), .ZN(new_n4283_));
  NAND2_X1   g01834(.A1(new_n4245_), .A2(pi0062), .ZN(new_n4284_));
  XOR2_X1    g01835(.A1(new_n4284_), .A2(new_n3594_), .Z(new_n4285_));
  NAND2_X1   g01836(.A1(new_n4285_), .A2(new_n4248_), .ZN(new_n4286_));
  NAND3_X1   g01837(.A1(new_n4286_), .A2(pi0248), .A3(new_n3230_), .ZN(new_n4287_));
  NAND2_X1   g01838(.A1(new_n4245_), .A2(pi0056), .ZN(new_n4288_));
  XOR2_X1    g01839(.A1(new_n4288_), .A2(new_n3797_), .Z(new_n4289_));
  AOI21_X1   g01840(.A1(new_n4289_), .A2(new_n4248_), .B(pi0062), .ZN(new_n4290_));
  NAND2_X1   g01841(.A1(new_n4287_), .A2(new_n4290_), .ZN(new_n4291_));
  NAND2_X1   g01842(.A1(new_n4245_), .A2(pi0055), .ZN(new_n4292_));
  XOR2_X1    g01843(.A1(new_n4292_), .A2(new_n3605_), .Z(new_n4293_));
  NAND2_X1   g01844(.A1(new_n4293_), .A2(new_n4248_), .ZN(new_n4294_));
  NAND2_X1   g01845(.A1(new_n4294_), .A2(new_n3219_), .ZN(new_n4295_));
  NOR2_X1    g01846(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4296_));
  NAND4_X1   g01847(.A1(new_n4283_), .A2(new_n4291_), .A3(new_n4295_), .A4(new_n4296_), .ZN(new_n4297_));
  OAI22_X1   g01848(.A1(new_n4280_), .A2(new_n4297_), .B1(new_n4237_), .B2(new_n4239_), .ZN(new_n4298_));
  AOI21_X1   g01849(.A1(new_n4218_), .A2(new_n4236_), .B(new_n4298_), .ZN(po0159));
  INV_X1     g01850(.I(pi1139), .ZN(new_n4300_));
  NAND3_X1   g01851(.A1(new_n3103_), .A2(pi0222), .A3(pi0920), .ZN(new_n4301_));
  INV_X1     g01852(.I(pi0920), .ZN(new_n4302_));
  NAND3_X1   g01853(.A1(new_n3344_), .A2(pi0222), .A3(new_n4302_), .ZN(new_n4303_));
  AOI21_X1   g01854(.A1(new_n4303_), .A2(new_n4301_), .B(new_n4300_), .ZN(new_n4304_));
  NOR2_X1    g01855(.A1(new_n3090_), .A2(new_n4300_), .ZN(new_n4305_));
  OAI21_X1   g01856(.A1(new_n4304_), .A2(pi0224), .B(new_n4305_), .ZN(new_n4306_));
  INV_X1     g01857(.I(new_n4306_), .ZN(new_n4307_));
  AOI21_X1   g01858(.A1(new_n4304_), .A2(pi0222), .B(pi0281), .ZN(new_n4308_));
  NAND2_X1   g01859(.A1(new_n3090_), .A2(pi0224), .ZN(new_n4309_));
  OAI22_X1   g01860(.A1(new_n4308_), .A2(new_n4309_), .B1(new_n3090_), .B2(pi1139), .ZN(new_n4310_));
  NOR2_X1    g01861(.A1(new_n4310_), .A2(pi0299), .ZN(new_n4311_));
  INV_X1     g01862(.I(new_n4311_), .ZN(new_n4312_));
  NOR3_X1    g01863(.A1(new_n4312_), .A2(new_n2820_), .A3(new_n3384_), .ZN(new_n4313_));
  OAI21_X1   g01864(.A1(new_n4313_), .A2(new_n4307_), .B(pi0862), .ZN(new_n4314_));
  NOR2_X1    g01865(.A1(new_n3411_), .A2(new_n3524_), .ZN(new_n4315_));
  INV_X1     g01866(.I(new_n4315_), .ZN(new_n4316_));
  INV_X1     g01867(.I(pi0862), .ZN(new_n4317_));
  NOR3_X1    g01868(.A1(new_n3011_), .A2(new_n3058_), .A3(new_n4302_), .ZN(new_n4318_));
  NOR3_X1    g01869(.A1(new_n3058_), .A2(pi0216), .A3(pi0920), .ZN(new_n4319_));
  OAI21_X1   g01870(.A1(new_n4318_), .A2(new_n4319_), .B(pi1139), .ZN(new_n4320_));
  NAND2_X1   g01871(.A1(new_n4320_), .A2(pi0221), .ZN(new_n4321_));
  AOI21_X1   g01872(.A1(pi0216), .A2(new_n4300_), .B(new_n4321_), .ZN(new_n4322_));
  AOI21_X1   g01873(.A1(pi0216), .A2(pi0281), .B(pi0221), .ZN(new_n4323_));
  AOI22_X1   g01874(.A1(new_n4322_), .A2(new_n4323_), .B1(new_n3011_), .B2(new_n4317_), .ZN(new_n4324_));
  NOR2_X1    g01875(.A1(new_n4316_), .A2(new_n4324_), .ZN(new_n4325_));
  INV_X1     g01876(.I(new_n4325_), .ZN(new_n4326_));
  NOR2_X1    g01877(.A1(new_n3111_), .A2(new_n4300_), .ZN(new_n4327_));
  INV_X1     g01878(.I(new_n4327_), .ZN(new_n4328_));
  INV_X1     g01879(.I(pi0148), .ZN(new_n4329_));
  NOR2_X1    g01880(.A1(new_n4329_), .A2(pi0215), .ZN(new_n4330_));
  INV_X1     g01881(.I(new_n4330_), .ZN(new_n4331_));
  NAND2_X1   g01882(.A1(new_n4328_), .A2(new_n4331_), .ZN(new_n4332_));
  NOR2_X1    g01883(.A1(new_n4325_), .A2(new_n4332_), .ZN(new_n4333_));
  NAND2_X1   g01884(.A1(new_n4321_), .A2(new_n3011_), .ZN(new_n4334_));
  NOR3_X1    g01885(.A1(new_n4333_), .A2(new_n4316_), .A3(new_n4334_), .ZN(new_n4335_));
  INV_X1     g01886(.I(new_n4335_), .ZN(new_n4336_));
  NOR2_X1    g01887(.A1(pi0148), .A2(pi0215), .ZN(new_n4337_));
  AOI21_X1   g01888(.A1(new_n4334_), .A2(new_n4337_), .B(new_n3009_), .ZN(new_n4338_));
  AOI21_X1   g01889(.A1(new_n4326_), .A2(new_n4338_), .B(new_n4336_), .ZN(new_n4339_));
  NOR2_X1    g01890(.A1(new_n4339_), .A2(new_n3098_), .ZN(new_n4340_));
  NOR2_X1    g01891(.A1(new_n4340_), .A2(new_n4314_), .ZN(new_n4341_));
  INV_X1     g01892(.I(new_n4341_), .ZN(new_n4342_));
  INV_X1     g01893(.I(new_n4338_), .ZN(new_n4343_));
  NOR2_X1    g01894(.A1(pi0216), .A2(pi0862), .ZN(new_n4344_));
  NOR3_X1    g01895(.A1(new_n3006_), .A2(new_n4344_), .A3(new_n4323_), .ZN(new_n4345_));
  OAI22_X1   g01896(.A1(new_n4343_), .A2(new_n4328_), .B1(new_n2820_), .B2(new_n4345_), .ZN(new_n4346_));
  NAND2_X1   g01897(.A1(new_n4346_), .A2(new_n4322_), .ZN(new_n4347_));
  INV_X1     g01898(.I(new_n4347_), .ZN(new_n4348_));
  NOR2_X1    g01899(.A1(new_n4348_), .A2(new_n3098_), .ZN(new_n4349_));
  NOR2_X1    g01900(.A1(new_n4314_), .A2(new_n4349_), .ZN(new_n4350_));
  NOR2_X1    g01901(.A1(new_n4350_), .A2(new_n3134_), .ZN(new_n4351_));
  AOI21_X1   g01902(.A1(new_n4342_), .A2(new_n3134_), .B(new_n4351_), .ZN(new_n4352_));
  INV_X1     g01903(.I(new_n4337_), .ZN(new_n4353_));
  NOR2_X1    g01904(.A1(new_n3338_), .A2(new_n4324_), .ZN(new_n4354_));
  NOR2_X1    g01905(.A1(new_n4354_), .A2(new_n4353_), .ZN(new_n4355_));
  NOR3_X1    g01906(.A1(new_n3306_), .A2(new_n4307_), .A3(new_n4311_), .ZN(new_n4356_));
  NAND2_X1   g01907(.A1(pi0299), .A2(pi0862), .ZN(new_n4357_));
  OAI22_X1   g01908(.A1(new_n4355_), .A2(new_n4327_), .B1(new_n4356_), .B2(new_n4357_), .ZN(new_n4358_));
  NOR2_X1    g01909(.A1(new_n3696_), .A2(pi0228), .ZN(new_n4359_));
  OAI21_X1   g01910(.A1(new_n3005_), .A2(pi0105), .B(pi0862), .ZN(new_n4360_));
  NOR2_X1    g01911(.A1(new_n4359_), .A2(new_n4360_), .ZN(new_n4361_));
  NOR2_X1    g01912(.A1(new_n3011_), .A2(new_n4317_), .ZN(new_n4362_));
  XOR2_X1    g01913(.A1(new_n4361_), .A2(new_n4362_), .Z(new_n4363_));
  NAND2_X1   g01914(.A1(new_n4363_), .A2(new_n3311_), .ZN(new_n4364_));
  AOI21_X1   g01915(.A1(new_n4322_), .A2(new_n4330_), .B(new_n4323_), .ZN(new_n4365_));
  NOR2_X1    g01916(.A1(new_n4364_), .A2(new_n4365_), .ZN(new_n4366_));
  NAND4_X1   g01917(.A1(new_n4358_), .A2(pi0038), .A3(pi0039), .A4(new_n4366_), .ZN(new_n4367_));
  INV_X1     g01918(.I(new_n3262_), .ZN(new_n4368_));
  NAND2_X1   g01919(.A1(new_n4358_), .A2(new_n4366_), .ZN(new_n4369_));
  NAND3_X1   g01920(.A1(new_n4369_), .A2(pi0039), .A3(new_n4368_), .ZN(new_n4370_));
  AOI21_X1   g01921(.A1(new_n4370_), .A2(new_n4367_), .B(new_n4342_), .ZN(new_n4371_));
  INV_X1     g01922(.I(new_n4350_), .ZN(new_n4372_));
  NOR2_X1    g01923(.A1(new_n4372_), .A2(new_n3259_), .ZN(new_n4373_));
  OAI21_X1   g01924(.A1(new_n4371_), .A2(pi0100), .B(new_n4373_), .ZN(new_n4374_));
  AOI21_X1   g01925(.A1(new_n3576_), .A2(new_n4323_), .B(new_n4326_), .ZN(new_n4375_));
  NOR2_X1    g01926(.A1(new_n4375_), .A2(new_n4353_), .ZN(new_n4376_));
  AND4_X2    g01927(.A1(pi0216), .A2(new_n3575_), .A3(new_n3006_), .A4(new_n4322_), .Z(new_n4377_));
  NAND2_X1   g01928(.A1(new_n4325_), .A2(pi0299), .ZN(new_n4378_));
  AOI21_X1   g01929(.A1(new_n4314_), .A2(new_n3212_), .B(new_n4378_), .ZN(new_n4379_));
  OAI21_X1   g01930(.A1(new_n4377_), .A2(new_n4332_), .B(new_n4379_), .ZN(new_n4380_));
  AOI21_X1   g01931(.A1(new_n4350_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4381_));
  OAI21_X1   g01932(.A1(new_n4380_), .A2(new_n4376_), .B(new_n4381_), .ZN(new_n4382_));
  NAND4_X1   g01933(.A1(new_n4374_), .A2(pi0075), .A3(pi0087), .A4(new_n4382_), .ZN(new_n4383_));
  NAND2_X1   g01934(.A1(new_n4374_), .A2(new_n4382_), .ZN(new_n4384_));
  NAND3_X1   g01935(.A1(new_n4384_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4385_));
  AOI21_X1   g01936(.A1(new_n4385_), .A2(new_n4383_), .B(new_n4352_), .ZN(new_n4386_));
  NOR2_X1    g01937(.A1(new_n4372_), .A2(new_n3235_), .ZN(new_n4387_));
  OAI21_X1   g01938(.A1(new_n4386_), .A2(pi0092), .B(new_n4387_), .ZN(new_n4388_));
  NAND2_X1   g01939(.A1(new_n4352_), .A2(pi0092), .ZN(new_n4389_));
  XOR2_X1    g01940(.A1(new_n4389_), .A2(new_n3172_), .Z(new_n4390_));
  NOR2_X1    g01941(.A1(new_n4339_), .A2(new_n3258_), .ZN(new_n4391_));
  XOR2_X1    g01942(.A1(new_n4391_), .A2(new_n3605_), .Z(new_n4392_));
  OAI21_X1   g01943(.A1(new_n4392_), .A2(new_n4347_), .B(new_n3219_), .ZN(new_n4393_));
  NOR2_X1    g01944(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4394_));
  NAND2_X1   g01945(.A1(new_n4393_), .A2(new_n4394_), .ZN(new_n4395_));
  AOI21_X1   g01946(.A1(new_n4390_), .A2(new_n4350_), .B(new_n4395_), .ZN(new_n4396_));
  NOR2_X1    g01947(.A1(new_n4339_), .A2(new_n3219_), .ZN(new_n4397_));
  XOR2_X1    g01948(.A1(new_n4397_), .A2(new_n3797_), .Z(new_n4398_));
  OAI21_X1   g01949(.A1(new_n4398_), .A2(new_n4347_), .B(new_n3201_), .ZN(new_n4399_));
  AOI21_X1   g01950(.A1(new_n4388_), .A2(new_n4396_), .B(new_n4399_), .ZN(new_n4400_));
  NOR2_X1    g01951(.A1(new_n4339_), .A2(new_n3201_), .ZN(new_n4401_));
  XOR2_X1    g01952(.A1(new_n4401_), .A2(new_n3594_), .Z(new_n4402_));
  NOR2_X1    g01953(.A1(new_n4348_), .A2(new_n3913_), .ZN(new_n4403_));
  NOR2_X1    g01954(.A1(new_n3426_), .A2(pi0247), .ZN(new_n4404_));
  OAI21_X1   g01955(.A1(new_n4402_), .A2(new_n4347_), .B(new_n4404_), .ZN(new_n4405_));
  OAI21_X1   g01956(.A1(new_n4312_), .A2(new_n4306_), .B(new_n4317_), .ZN(new_n4406_));
  NAND2_X1   g01957(.A1(new_n4406_), .A2(new_n2753_), .ZN(new_n4407_));
  AOI21_X1   g01958(.A1(new_n3370_), .A2(pi0862), .B(pi0216), .ZN(new_n4408_));
  OAI21_X1   g01959(.A1(new_n3411_), .A2(new_n3006_), .B(new_n4408_), .ZN(new_n4409_));
  AOI21_X1   g01960(.A1(new_n4409_), .A2(new_n4323_), .B(new_n4322_), .ZN(new_n4410_));
  OAI21_X1   g01961(.A1(new_n4353_), .A2(new_n4410_), .B(new_n4335_), .ZN(new_n4411_));
  NAND2_X1   g01962(.A1(new_n4411_), .A2(pi0299), .ZN(new_n4412_));
  NAND2_X1   g01963(.A1(new_n4412_), .A2(new_n4407_), .ZN(new_n4413_));
  INV_X1     g01964(.I(new_n4403_), .ZN(new_n4414_));
  OAI21_X1   g01965(.A1(new_n4414_), .A2(new_n3098_), .B(new_n4407_), .ZN(new_n4415_));
  INV_X1     g01966(.I(new_n4415_), .ZN(new_n4416_));
  NOR2_X1    g01967(.A1(new_n4416_), .A2(new_n3134_), .ZN(new_n4417_));
  AOI21_X1   g01968(.A1(new_n3134_), .A2(new_n4413_), .B(new_n4417_), .ZN(new_n4418_));
  OAI21_X1   g01969(.A1(new_n3338_), .A2(new_n4324_), .B(new_n4331_), .ZN(new_n4419_));
  AOI21_X1   g01970(.A1(new_n4322_), .A2(new_n4337_), .B(new_n4323_), .ZN(new_n4420_));
  NAND4_X1   g01971(.A1(new_n4321_), .A2(new_n3011_), .A3(pi0299), .A4(new_n4327_), .ZN(new_n4421_));
  NOR4_X1    g01972(.A1(new_n4364_), .A2(new_n3338_), .A3(new_n4420_), .A4(new_n4421_), .ZN(new_n4422_));
  AOI21_X1   g01973(.A1(new_n4422_), .A2(new_n4419_), .B(pi0039), .ZN(new_n4423_));
  AOI21_X1   g01974(.A1(new_n4310_), .A2(new_n4307_), .B(pi0862), .ZN(new_n4424_));
  OR3_X2     g01975(.A1(new_n3702_), .A2(new_n3098_), .A3(new_n4424_), .Z(new_n4425_));
  OAI21_X1   g01976(.A1(new_n4423_), .A2(new_n4425_), .B(new_n3259_), .ZN(new_n4426_));
  NOR2_X1    g01977(.A1(new_n4413_), .A2(new_n3183_), .ZN(new_n4427_));
  AOI21_X1   g01978(.A1(new_n4426_), .A2(new_n4427_), .B(pi0100), .ZN(new_n4428_));
  NAND2_X1   g01979(.A1(new_n4416_), .A2(pi0038), .ZN(new_n4429_));
  OR2_X2     g01980(.A1(new_n4375_), .A2(new_n4330_), .Z(new_n4430_));
  NOR2_X1    g01981(.A1(new_n3577_), .A2(new_n4334_), .ZN(new_n4431_));
  NAND2_X1   g01982(.A1(new_n4430_), .A2(new_n4431_), .ZN(new_n4432_));
  OR3_X2     g01983(.A1(new_n4410_), .A2(new_n3006_), .A3(new_n4323_), .Z(new_n4433_));
  NAND2_X1   g01984(.A1(new_n4407_), .A2(new_n3212_), .ZN(new_n4434_));
  NOR2_X1    g01985(.A1(new_n4353_), .A2(new_n3098_), .ZN(new_n4435_));
  NAND4_X1   g01986(.A1(new_n3575_), .A2(new_n4433_), .A3(new_n4434_), .A4(new_n4435_), .ZN(new_n4436_));
  AOI21_X1   g01987(.A1(new_n4432_), .A2(new_n4328_), .B(new_n4436_), .ZN(new_n4437_));
  OAI21_X1   g01988(.A1(new_n4415_), .A2(new_n3211_), .B(pi0100), .ZN(new_n4438_));
  OAI22_X1   g01989(.A1(new_n4428_), .A2(new_n4429_), .B1(new_n4437_), .B2(new_n4438_), .ZN(new_n4439_));
  OR3_X2     g01990(.A1(new_n4439_), .A2(new_n3235_), .A3(new_n3455_), .Z(new_n4440_));
  NAND3_X1   g01991(.A1(new_n4439_), .A2(new_n3235_), .A3(pi0087), .ZN(new_n4441_));
  AOI21_X1   g01992(.A1(new_n4440_), .A2(new_n4441_), .B(new_n4418_), .ZN(new_n4442_));
  NOR2_X1    g01993(.A1(new_n4415_), .A2(new_n3235_), .ZN(new_n4443_));
  OAI21_X1   g01994(.A1(new_n4442_), .A2(pi0092), .B(new_n4443_), .ZN(new_n4444_));
  NAND2_X1   g01995(.A1(new_n4418_), .A2(pi0092), .ZN(new_n4445_));
  XOR2_X1    g01996(.A1(new_n4445_), .A2(new_n3172_), .Z(new_n4446_));
  NAND2_X1   g01997(.A1(new_n4411_), .A2(pi0055), .ZN(new_n4447_));
  XOR2_X1    g01998(.A1(new_n4447_), .A2(new_n3604_), .Z(new_n4448_));
  OAI21_X1   g01999(.A1(new_n4448_), .A2(new_n4414_), .B(new_n3219_), .ZN(new_n4449_));
  NOR2_X1    g02000(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4450_));
  NAND2_X1   g02001(.A1(new_n4449_), .A2(new_n4450_), .ZN(new_n4451_));
  AOI21_X1   g02002(.A1(new_n4446_), .A2(new_n4416_), .B(new_n4451_), .ZN(new_n4452_));
  NAND2_X1   g02003(.A1(new_n4411_), .A2(pi0056), .ZN(new_n4453_));
  XOR2_X1    g02004(.A1(new_n4453_), .A2(new_n3599_), .Z(new_n4454_));
  OAI21_X1   g02005(.A1(new_n4454_), .A2(new_n4414_), .B(new_n3201_), .ZN(new_n4455_));
  AOI21_X1   g02006(.A1(new_n4444_), .A2(new_n4452_), .B(new_n4455_), .ZN(new_n4456_));
  NAND2_X1   g02007(.A1(new_n4411_), .A2(pi0062), .ZN(new_n4457_));
  XOR2_X1    g02008(.A1(new_n4457_), .A2(new_n3972_), .Z(new_n4458_));
  INV_X1     g02009(.I(pi0247), .ZN(new_n4459_));
  NOR2_X1    g02010(.A1(new_n3426_), .A2(new_n4459_), .ZN(new_n4460_));
  OAI21_X1   g02011(.A1(new_n4458_), .A2(new_n4414_), .B(new_n4460_), .ZN(new_n4461_));
  OAI22_X1   g02012(.A1(new_n4400_), .A2(new_n4405_), .B1(new_n4456_), .B2(new_n4461_), .ZN(po0160));
  NAND2_X1   g02013(.A1(new_n2820_), .A2(pi0877), .ZN(new_n4463_));
  AOI21_X1   g02014(.A1(pi0224), .A2(pi0269), .B(pi0222), .ZN(new_n4464_));
  INV_X1     g02015(.I(pi1138), .ZN(new_n4465_));
  NAND3_X1   g02016(.A1(new_n3103_), .A2(pi0222), .A3(pi0940), .ZN(new_n4466_));
  INV_X1     g02017(.I(pi0940), .ZN(new_n4467_));
  NAND3_X1   g02018(.A1(new_n3344_), .A2(pi0222), .A3(new_n4467_), .ZN(new_n4468_));
  AOI21_X1   g02019(.A1(new_n4468_), .A2(new_n4466_), .B(new_n4465_), .ZN(new_n4469_));
  AOI21_X1   g02020(.A1(new_n4469_), .A2(new_n4464_), .B(pi0224), .ZN(new_n4470_));
  OAI21_X1   g02021(.A1(new_n4470_), .A2(new_n4463_), .B(pi0223), .ZN(new_n4471_));
  XOR2_X1    g02022(.A1(new_n4471_), .A2(new_n3565_), .Z(new_n4472_));
  NAND2_X1   g02023(.A1(new_n4472_), .A2(pi1138), .ZN(new_n4473_));
  INV_X1     g02024(.I(pi0169), .ZN(new_n4474_));
  NAND3_X1   g02025(.A1(new_n3160_), .A2(pi0228), .A3(pi0877), .ZN(new_n4475_));
  INV_X1     g02026(.I(pi0877), .ZN(new_n4476_));
  NAND3_X1   g02027(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n4476_), .ZN(new_n4477_));
  AOI21_X1   g02028(.A1(new_n4475_), .A2(new_n4477_), .B(new_n4474_), .ZN(new_n4478_));
  NAND4_X1   g02029(.A1(new_n2820_), .A2(pi0105), .A3(pi0228), .A4(pi0877), .ZN(new_n4479_));
  NAND3_X1   g02030(.A1(new_n4463_), .A2(new_n3004_), .A3(pi0228), .ZN(new_n4480_));
  AOI21_X1   g02031(.A1(new_n4480_), .A2(new_n4479_), .B(new_n4474_), .ZN(new_n4481_));
  NOR2_X1    g02032(.A1(new_n4481_), .A2(pi0216), .ZN(new_n4482_));
  INV_X1     g02033(.I(new_n4482_), .ZN(new_n4483_));
  NOR2_X1    g02034(.A1(new_n3121_), .A2(pi0940), .ZN(new_n4484_));
  XOR2_X1    g02035(.A1(new_n3356_), .A2(new_n4484_), .Z(new_n4485_));
  AOI21_X1   g02036(.A1(pi0216), .A2(pi0269), .B(pi0221), .ZN(new_n4486_));
  NAND3_X1   g02037(.A1(new_n4485_), .A2(pi1138), .A3(new_n4486_), .ZN(new_n4487_));
  NAND2_X1   g02038(.A1(new_n4483_), .A2(new_n4487_), .ZN(new_n4488_));
  NAND3_X1   g02039(.A1(new_n4488_), .A2(new_n4478_), .A3(new_n3111_), .ZN(new_n4489_));
  OAI21_X1   g02040(.A1(new_n3111_), .A2(pi1138), .B(new_n4489_), .ZN(new_n4490_));
  OAI21_X1   g02041(.A1(new_n4490_), .A2(new_n3098_), .B(new_n4473_), .ZN(new_n4491_));
  INV_X1     g02042(.I(new_n4473_), .ZN(new_n4492_));
  NAND2_X1   g02043(.A1(new_n4485_), .A2(pi1138), .ZN(new_n4493_));
  NAND2_X1   g02044(.A1(new_n4493_), .A2(pi0215), .ZN(new_n4494_));
  NAND2_X1   g02045(.A1(new_n4482_), .A2(new_n4486_), .ZN(new_n4495_));
  NAND2_X1   g02046(.A1(new_n4495_), .A2(new_n3005_), .ZN(new_n4496_));
  NAND4_X1   g02047(.A1(new_n4496_), .A2(pi0169), .A3(pi0215), .A4(pi1138), .ZN(new_n4497_));
  XNOR2_X1   g02048(.A1(new_n4497_), .A2(new_n4494_), .ZN(new_n4498_));
  AOI21_X1   g02049(.A1(new_n4498_), .A2(pi0299), .B(new_n4492_), .ZN(new_n4499_));
  NOR2_X1    g02050(.A1(new_n4499_), .A2(new_n3134_), .ZN(new_n4500_));
  AOI21_X1   g02051(.A1(new_n3134_), .A2(new_n4491_), .B(new_n4500_), .ZN(new_n4501_));
  NAND2_X1   g02052(.A1(new_n3307_), .A2(pi0877), .ZN(new_n4502_));
  AOI21_X1   g02053(.A1(new_n3459_), .A2(new_n4474_), .B(new_n4502_), .ZN(new_n4503_));
  NAND3_X1   g02054(.A1(new_n3330_), .A2(pi0169), .A3(pi0877), .ZN(new_n4504_));
  NAND3_X1   g02055(.A1(new_n3862_), .A2(new_n4474_), .A3(pi0877), .ZN(new_n4505_));
  AOI21_X1   g02056(.A1(new_n4505_), .A2(new_n4504_), .B(new_n3308_), .ZN(new_n4506_));
  NAND2_X1   g02057(.A1(new_n3931_), .A2(new_n4481_), .ZN(new_n4507_));
  NAND2_X1   g02058(.A1(new_n4507_), .A2(new_n3011_), .ZN(new_n4508_));
  AOI21_X1   g02059(.A1(new_n4508_), .A2(new_n4487_), .B(pi0228), .ZN(new_n4509_));
  OAI21_X1   g02060(.A1(new_n4506_), .A2(new_n4503_), .B(new_n4509_), .ZN(new_n4510_));
  OR3_X2     g02061(.A1(new_n4510_), .A2(new_n3111_), .A3(new_n3098_), .Z(new_n4511_));
  NAND3_X1   g02062(.A1(new_n4510_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n4512_));
  AOI21_X1   g02063(.A1(new_n4511_), .A2(new_n4512_), .B(new_n4465_), .ZN(new_n4513_));
  AOI21_X1   g02064(.A1(pi0223), .A2(pi1138), .B(pi0299), .ZN(new_n4514_));
  AOI21_X1   g02065(.A1(new_n4464_), .A2(pi0224), .B(pi0877), .ZN(new_n4515_));
  NOR2_X1    g02066(.A1(new_n3702_), .A2(new_n4515_), .ZN(new_n4516_));
  NOR3_X1    g02067(.A1(new_n4516_), .A2(new_n3090_), .A3(new_n4469_), .ZN(new_n4517_));
  OAI21_X1   g02068(.A1(new_n4517_), .A2(new_n4464_), .B(new_n3306_), .ZN(new_n4518_));
  AOI21_X1   g02069(.A1(new_n4518_), .A2(new_n4514_), .B(pi0039), .ZN(new_n4519_));
  INV_X1     g02070(.I(new_n4514_), .ZN(new_n4520_));
  NOR3_X1    g02071(.A1(new_n4516_), .A2(new_n4469_), .A3(new_n4520_), .ZN(new_n4521_));
  OAI21_X1   g02072(.A1(new_n4513_), .A2(new_n4519_), .B(new_n4521_), .ZN(new_n4522_));
  OR2_X2     g02073(.A1(new_n4491_), .A2(new_n3183_), .Z(new_n4523_));
  AOI21_X1   g02074(.A1(new_n4522_), .A2(new_n3259_), .B(new_n4523_), .ZN(new_n4524_));
  INV_X1     g02075(.I(new_n4499_), .ZN(new_n4525_));
  NOR2_X1    g02076(.A1(new_n4525_), .A2(new_n3259_), .ZN(new_n4526_));
  OAI21_X1   g02077(.A1(new_n4524_), .A2(pi0100), .B(new_n4526_), .ZN(new_n4527_));
  NAND3_X1   g02078(.A1(new_n3400_), .A2(pi0228), .A3(pi0877), .ZN(new_n4528_));
  NAND3_X1   g02079(.A1(new_n3400_), .A2(new_n3005_), .A3(new_n4476_), .ZN(new_n4529_));
  AOI21_X1   g02080(.A1(new_n4528_), .A2(new_n4529_), .B(new_n4474_), .ZN(new_n4530_));
  AOI21_X1   g02081(.A1(new_n4530_), .A2(new_n4488_), .B(new_n3098_), .ZN(new_n4531_));
  XOR2_X1    g02082(.A1(new_n4531_), .A2(new_n3855_), .Z(new_n4532_));
  NOR2_X1    g02083(.A1(new_n4532_), .A2(new_n4465_), .ZN(new_n4533_));
  NAND2_X1   g02084(.A1(new_n4473_), .A2(new_n3211_), .ZN(new_n4534_));
  AOI21_X1   g02085(.A1(new_n4499_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4535_));
  OAI21_X1   g02086(.A1(new_n4533_), .A2(new_n4534_), .B(new_n4535_), .ZN(new_n4536_));
  NAND4_X1   g02087(.A1(new_n4527_), .A2(pi0075), .A3(pi0087), .A4(new_n4536_), .ZN(new_n4537_));
  NAND2_X1   g02088(.A1(new_n4527_), .A2(new_n4536_), .ZN(new_n4538_));
  NAND3_X1   g02089(.A1(new_n4538_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4539_));
  AOI21_X1   g02090(.A1(new_n4539_), .A2(new_n4537_), .B(new_n4501_), .ZN(new_n4540_));
  NOR2_X1    g02091(.A1(new_n4525_), .A2(new_n3235_), .ZN(new_n4541_));
  OAI21_X1   g02092(.A1(new_n4540_), .A2(pi0092), .B(new_n4541_), .ZN(new_n4542_));
  NAND2_X1   g02093(.A1(new_n4501_), .A2(pi0092), .ZN(new_n4543_));
  XNOR2_X1   g02094(.A1(new_n4543_), .A2(new_n3172_), .ZN(new_n4544_));
  NOR2_X1    g02095(.A1(new_n4544_), .A2(new_n4525_), .ZN(new_n4545_));
  INV_X1     g02096(.I(new_n4498_), .ZN(new_n4546_));
  NOR2_X1    g02097(.A1(new_n4490_), .A2(new_n3201_), .ZN(new_n4547_));
  XOR2_X1    g02098(.A1(new_n4547_), .A2(new_n3972_), .Z(new_n4548_));
  INV_X1     g02099(.I(pi0246), .ZN(new_n4549_));
  NAND2_X1   g02100(.A1(new_n3230_), .A2(new_n4549_), .ZN(new_n4550_));
  AOI21_X1   g02101(.A1(new_n4548_), .A2(new_n4546_), .B(new_n4550_), .ZN(new_n4551_));
  NOR2_X1    g02102(.A1(new_n4490_), .A2(new_n3219_), .ZN(new_n4552_));
  XOR2_X1    g02103(.A1(new_n4552_), .A2(new_n3797_), .Z(new_n4553_));
  OAI21_X1   g02104(.A1(new_n4553_), .A2(new_n4498_), .B(new_n3201_), .ZN(new_n4554_));
  NOR2_X1    g02105(.A1(new_n4551_), .A2(new_n4554_), .ZN(new_n4555_));
  NOR2_X1    g02106(.A1(new_n4490_), .A2(new_n3258_), .ZN(new_n4556_));
  XOR2_X1    g02107(.A1(new_n4556_), .A2(new_n3604_), .Z(new_n4557_));
  AOI21_X1   g02108(.A1(new_n4557_), .A2(new_n4546_), .B(pi0056), .ZN(new_n4558_));
  NAND2_X1   g02109(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n4559_));
  NOR4_X1    g02110(.A1(new_n4545_), .A2(new_n4555_), .A3(new_n4558_), .A4(new_n4559_), .ZN(new_n4560_));
  NOR2_X1    g02111(.A1(new_n4546_), .A2(new_n3230_), .ZN(new_n4561_));
  AOI21_X1   g02112(.A1(pi0216), .A2(pi0269), .B(new_n3612_), .ZN(new_n4562_));
  NAND2_X1   g02113(.A1(new_n4562_), .A2(pi0246), .ZN(new_n4563_));
  NOR2_X1    g02114(.A1(new_n4492_), .A2(new_n3385_), .ZN(new_n4564_));
  NOR2_X1    g02115(.A1(new_n4482_), .A2(new_n4486_), .ZN(new_n4565_));
  INV_X1     g02116(.I(new_n4565_), .ZN(new_n4566_));
  NOR3_X1    g02117(.A1(new_n3370_), .A2(new_n3111_), .A3(new_n4465_), .ZN(new_n4567_));
  OAI21_X1   g02118(.A1(new_n4566_), .A2(new_n4478_), .B(new_n4567_), .ZN(new_n4568_));
  XNOR2_X1   g02119(.A1(new_n4568_), .A2(new_n4494_), .ZN(new_n4569_));
  NAND2_X1   g02120(.A1(new_n4569_), .A2(pi0299), .ZN(new_n4570_));
  NAND2_X1   g02121(.A1(new_n4570_), .A2(new_n4564_), .ZN(new_n4571_));
  NOR2_X1    g02122(.A1(new_n4498_), .A2(new_n4562_), .ZN(new_n4572_));
  OAI21_X1   g02123(.A1(new_n4572_), .A2(new_n3098_), .B(new_n4564_), .ZN(new_n4573_));
  INV_X1     g02124(.I(new_n4573_), .ZN(new_n4574_));
  NOR2_X1    g02125(.A1(new_n4574_), .A2(new_n3134_), .ZN(new_n4575_));
  AOI21_X1   g02126(.A1(new_n4571_), .A2(new_n3134_), .B(new_n4575_), .ZN(new_n4576_));
  INV_X1     g02127(.I(new_n4576_), .ZN(new_n4577_));
  NAND3_X1   g02128(.A1(new_n3696_), .A2(pi0169), .A3(pi0877), .ZN(new_n4578_));
  NAND3_X1   g02129(.A1(new_n3459_), .A2(pi0169), .A3(new_n4476_), .ZN(new_n4579_));
  NAND2_X1   g02130(.A1(new_n3307_), .A2(pi0169), .ZN(new_n4580_));
  AOI21_X1   g02131(.A1(new_n4578_), .A2(new_n4579_), .B(new_n4580_), .ZN(new_n4581_));
  NAND2_X1   g02132(.A1(pi0228), .A2(pi0877), .ZN(new_n4582_));
  AOI21_X1   g02133(.A1(new_n3703_), .A2(new_n4483_), .B(new_n4582_), .ZN(new_n4583_));
  OAI21_X1   g02134(.A1(new_n4581_), .A2(new_n3330_), .B(new_n4583_), .ZN(new_n4584_));
  NAND2_X1   g02135(.A1(new_n4584_), .A2(new_n4486_), .ZN(new_n4585_));
  AOI21_X1   g02136(.A1(new_n4585_), .A2(new_n4493_), .B(new_n3098_), .ZN(new_n4586_));
  XOR2_X1    g02137(.A1(new_n4586_), .A2(new_n3855_), .Z(new_n4587_));
  NOR2_X1    g02138(.A1(pi0038), .A2(pi0100), .ZN(new_n4588_));
  INV_X1     g02139(.I(new_n4588_), .ZN(new_n4589_));
  AOI21_X1   g02140(.A1(new_n4571_), .A2(pi0039), .B(new_n4589_), .ZN(new_n4590_));
  OAI21_X1   g02141(.A1(new_n4519_), .A2(new_n4590_), .B(pi1138), .ZN(new_n4591_));
  NOR2_X1    g02142(.A1(new_n4587_), .A2(new_n4591_), .ZN(new_n4592_));
  OAI21_X1   g02143(.A1(new_n4530_), .A2(new_n4566_), .B(new_n4567_), .ZN(new_n4593_));
  XOR2_X1    g02144(.A1(new_n4593_), .A2(new_n4494_), .Z(new_n4594_));
  NOR2_X1    g02145(.A1(new_n4564_), .A2(new_n3211_), .ZN(new_n4595_));
  NOR2_X1    g02146(.A1(new_n4595_), .A2(new_n3098_), .ZN(new_n4596_));
  OAI21_X1   g02147(.A1(new_n4573_), .A2(new_n3211_), .B(pi0100), .ZN(new_n4597_));
  AOI21_X1   g02148(.A1(new_n4594_), .A2(new_n4596_), .B(new_n4597_), .ZN(new_n4598_));
  NOR4_X1    g02149(.A1(new_n4592_), .A2(new_n3235_), .A3(new_n3455_), .A4(new_n4598_), .ZN(new_n4599_));
  OAI21_X1   g02150(.A1(new_n4592_), .A2(new_n4598_), .B(pi0087), .ZN(new_n4600_));
  NOR2_X1    g02151(.A1(new_n4600_), .A2(new_n3694_), .ZN(new_n4601_));
  OAI21_X1   g02152(.A1(new_n4601_), .A2(new_n4599_), .B(new_n4577_), .ZN(new_n4602_));
  NAND2_X1   g02153(.A1(new_n4574_), .A2(pi0075), .ZN(new_n4603_));
  AOI21_X1   g02154(.A1(new_n4602_), .A2(new_n3303_), .B(new_n4603_), .ZN(new_n4604_));
  NAND2_X1   g02155(.A1(new_n4576_), .A2(pi0092), .ZN(new_n4605_));
  XOR2_X1    g02156(.A1(new_n4605_), .A2(new_n3172_), .Z(new_n4606_));
  NAND2_X1   g02157(.A1(new_n4606_), .A2(new_n4574_), .ZN(new_n4607_));
  NAND2_X1   g02158(.A1(new_n4569_), .A2(pi0062), .ZN(new_n4608_));
  XOR2_X1    g02159(.A1(new_n4608_), .A2(new_n3594_), .Z(new_n4609_));
  NAND2_X1   g02160(.A1(new_n4609_), .A2(new_n4572_), .ZN(new_n4610_));
  NAND3_X1   g02161(.A1(new_n4610_), .A2(pi0246), .A3(new_n3230_), .ZN(new_n4611_));
  NAND2_X1   g02162(.A1(new_n4569_), .A2(pi0056), .ZN(new_n4612_));
  XOR2_X1    g02163(.A1(new_n4612_), .A2(new_n3797_), .Z(new_n4613_));
  AOI21_X1   g02164(.A1(new_n4613_), .A2(new_n4572_), .B(pi0062), .ZN(new_n4614_));
  NAND2_X1   g02165(.A1(new_n4611_), .A2(new_n4614_), .ZN(new_n4615_));
  NAND2_X1   g02166(.A1(new_n4569_), .A2(pi0055), .ZN(new_n4616_));
  XOR2_X1    g02167(.A1(new_n4616_), .A2(new_n3605_), .Z(new_n4617_));
  NAND2_X1   g02168(.A1(new_n4617_), .A2(new_n4572_), .ZN(new_n4618_));
  NAND2_X1   g02169(.A1(new_n4618_), .A2(new_n3219_), .ZN(new_n4619_));
  NOR2_X1    g02170(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4620_));
  NAND4_X1   g02171(.A1(new_n4607_), .A2(new_n4615_), .A3(new_n4619_), .A4(new_n4620_), .ZN(new_n4621_));
  OAI22_X1   g02172(.A1(new_n4604_), .A2(new_n4621_), .B1(new_n4561_), .B2(new_n4563_), .ZN(new_n4622_));
  AOI21_X1   g02173(.A1(new_n4542_), .A2(new_n4560_), .B(new_n4622_), .ZN(po0161));
  NAND2_X1   g02174(.A1(new_n2820_), .A2(pi0878), .ZN(new_n4624_));
  AOI21_X1   g02175(.A1(pi0224), .A2(pi0280), .B(pi0222), .ZN(new_n4625_));
  INV_X1     g02176(.I(pi1137), .ZN(new_n4626_));
  NAND3_X1   g02177(.A1(new_n3103_), .A2(pi0222), .A3(pi0933), .ZN(new_n4627_));
  INV_X1     g02178(.I(pi0933), .ZN(new_n4628_));
  NAND3_X1   g02179(.A1(new_n3344_), .A2(pi0222), .A3(new_n4628_), .ZN(new_n4629_));
  AOI21_X1   g02180(.A1(new_n4629_), .A2(new_n4627_), .B(new_n4626_), .ZN(new_n4630_));
  AOI21_X1   g02181(.A1(new_n4630_), .A2(new_n4625_), .B(pi0224), .ZN(new_n4631_));
  OAI21_X1   g02182(.A1(new_n4631_), .A2(new_n4624_), .B(pi0223), .ZN(new_n4632_));
  XOR2_X1    g02183(.A1(new_n4632_), .A2(new_n3565_), .Z(new_n4633_));
  NAND2_X1   g02184(.A1(new_n4633_), .A2(pi1137), .ZN(new_n4634_));
  INV_X1     g02185(.I(pi0168), .ZN(new_n4635_));
  NAND3_X1   g02186(.A1(new_n3160_), .A2(pi0228), .A3(pi0878), .ZN(new_n4636_));
  INV_X1     g02187(.I(pi0878), .ZN(new_n4637_));
  NAND3_X1   g02188(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n4637_), .ZN(new_n4638_));
  AOI21_X1   g02189(.A1(new_n4636_), .A2(new_n4638_), .B(new_n4635_), .ZN(new_n4639_));
  NAND4_X1   g02190(.A1(new_n2820_), .A2(pi0105), .A3(pi0228), .A4(pi0878), .ZN(new_n4640_));
  NAND3_X1   g02191(.A1(new_n4624_), .A2(new_n3004_), .A3(pi0228), .ZN(new_n4641_));
  AOI21_X1   g02192(.A1(new_n4641_), .A2(new_n4640_), .B(new_n4635_), .ZN(new_n4642_));
  NOR2_X1    g02193(.A1(new_n4642_), .A2(pi0216), .ZN(new_n4643_));
  INV_X1     g02194(.I(new_n4643_), .ZN(new_n4644_));
  NOR2_X1    g02195(.A1(new_n3121_), .A2(pi0933), .ZN(new_n4645_));
  XOR2_X1    g02196(.A1(new_n3356_), .A2(new_n4645_), .Z(new_n4646_));
  AOI21_X1   g02197(.A1(pi0216), .A2(pi0280), .B(pi0221), .ZN(new_n4647_));
  NAND3_X1   g02198(.A1(new_n4646_), .A2(pi1137), .A3(new_n4647_), .ZN(new_n4648_));
  NAND2_X1   g02199(.A1(new_n4644_), .A2(new_n4648_), .ZN(new_n4649_));
  NAND3_X1   g02200(.A1(new_n4649_), .A2(new_n4639_), .A3(new_n3111_), .ZN(new_n4650_));
  OAI21_X1   g02201(.A1(new_n3111_), .A2(pi1137), .B(new_n4650_), .ZN(new_n4651_));
  OAI21_X1   g02202(.A1(new_n4651_), .A2(new_n3098_), .B(new_n4634_), .ZN(new_n4652_));
  INV_X1     g02203(.I(new_n4634_), .ZN(new_n4653_));
  NAND2_X1   g02204(.A1(new_n4646_), .A2(pi1137), .ZN(new_n4654_));
  NAND2_X1   g02205(.A1(new_n4654_), .A2(pi0215), .ZN(new_n4655_));
  NAND2_X1   g02206(.A1(new_n4643_), .A2(new_n4647_), .ZN(new_n4656_));
  NAND2_X1   g02207(.A1(new_n4656_), .A2(new_n3005_), .ZN(new_n4657_));
  NAND4_X1   g02208(.A1(new_n4657_), .A2(pi0168), .A3(pi0215), .A4(pi1137), .ZN(new_n4658_));
  XNOR2_X1   g02209(.A1(new_n4658_), .A2(new_n4655_), .ZN(new_n4659_));
  AOI21_X1   g02210(.A1(new_n4659_), .A2(pi0299), .B(new_n4653_), .ZN(new_n4660_));
  NOR2_X1    g02211(.A1(new_n4660_), .A2(new_n3134_), .ZN(new_n4661_));
  AOI21_X1   g02212(.A1(new_n3134_), .A2(new_n4652_), .B(new_n4661_), .ZN(new_n4662_));
  NAND2_X1   g02213(.A1(new_n3307_), .A2(pi0878), .ZN(new_n4663_));
  AOI21_X1   g02214(.A1(new_n3459_), .A2(new_n4635_), .B(new_n4663_), .ZN(new_n4664_));
  NAND3_X1   g02215(.A1(new_n3330_), .A2(pi0168), .A3(pi0878), .ZN(new_n4665_));
  NAND3_X1   g02216(.A1(new_n3862_), .A2(new_n4635_), .A3(pi0878), .ZN(new_n4666_));
  AOI21_X1   g02217(.A1(new_n4666_), .A2(new_n4665_), .B(new_n3308_), .ZN(new_n4667_));
  NAND2_X1   g02218(.A1(new_n3931_), .A2(new_n4642_), .ZN(new_n4668_));
  NAND2_X1   g02219(.A1(new_n4668_), .A2(new_n3011_), .ZN(new_n4669_));
  AOI21_X1   g02220(.A1(new_n4669_), .A2(new_n4648_), .B(pi0228), .ZN(new_n4670_));
  OAI21_X1   g02221(.A1(new_n4667_), .A2(new_n4664_), .B(new_n4670_), .ZN(new_n4671_));
  OR3_X2     g02222(.A1(new_n4671_), .A2(new_n3111_), .A3(new_n3098_), .Z(new_n4672_));
  NAND3_X1   g02223(.A1(new_n4671_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n4673_));
  AOI21_X1   g02224(.A1(new_n4672_), .A2(new_n4673_), .B(new_n4626_), .ZN(new_n4674_));
  AOI21_X1   g02225(.A1(pi0223), .A2(pi1137), .B(pi0299), .ZN(new_n4675_));
  AOI21_X1   g02226(.A1(new_n4625_), .A2(pi0224), .B(pi0878), .ZN(new_n4676_));
  NOR2_X1    g02227(.A1(new_n3702_), .A2(new_n4676_), .ZN(new_n4677_));
  NOR3_X1    g02228(.A1(new_n4677_), .A2(new_n3090_), .A3(new_n4630_), .ZN(new_n4678_));
  OAI21_X1   g02229(.A1(new_n4678_), .A2(new_n4625_), .B(new_n3306_), .ZN(new_n4679_));
  AOI21_X1   g02230(.A1(new_n4679_), .A2(new_n4675_), .B(pi0039), .ZN(new_n4680_));
  INV_X1     g02231(.I(new_n4675_), .ZN(new_n4681_));
  NOR3_X1    g02232(.A1(new_n4677_), .A2(new_n4630_), .A3(new_n4681_), .ZN(new_n4682_));
  OAI21_X1   g02233(.A1(new_n4674_), .A2(new_n4680_), .B(new_n4682_), .ZN(new_n4683_));
  OR2_X2     g02234(.A1(new_n4652_), .A2(new_n3183_), .Z(new_n4684_));
  AOI21_X1   g02235(.A1(new_n4683_), .A2(new_n3259_), .B(new_n4684_), .ZN(new_n4685_));
  INV_X1     g02236(.I(new_n4660_), .ZN(new_n4686_));
  NOR2_X1    g02237(.A1(new_n4686_), .A2(new_n3259_), .ZN(new_n4687_));
  OAI21_X1   g02238(.A1(new_n4685_), .A2(pi0100), .B(new_n4687_), .ZN(new_n4688_));
  NAND3_X1   g02239(.A1(new_n3400_), .A2(pi0228), .A3(pi0878), .ZN(new_n4689_));
  NAND3_X1   g02240(.A1(new_n3400_), .A2(new_n3005_), .A3(new_n4637_), .ZN(new_n4690_));
  AOI21_X1   g02241(.A1(new_n4689_), .A2(new_n4690_), .B(new_n4635_), .ZN(new_n4691_));
  AOI21_X1   g02242(.A1(new_n4691_), .A2(new_n4649_), .B(new_n3098_), .ZN(new_n4692_));
  XOR2_X1    g02243(.A1(new_n4692_), .A2(new_n3855_), .Z(new_n4693_));
  NOR2_X1    g02244(.A1(new_n4693_), .A2(new_n4626_), .ZN(new_n4694_));
  NAND2_X1   g02245(.A1(new_n4634_), .A2(new_n3211_), .ZN(new_n4695_));
  AOI21_X1   g02246(.A1(new_n4660_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4696_));
  OAI21_X1   g02247(.A1(new_n4694_), .A2(new_n4695_), .B(new_n4696_), .ZN(new_n4697_));
  NAND4_X1   g02248(.A1(new_n4688_), .A2(pi0075), .A3(pi0087), .A4(new_n4697_), .ZN(new_n4698_));
  NAND2_X1   g02249(.A1(new_n4688_), .A2(new_n4697_), .ZN(new_n4699_));
  NAND3_X1   g02250(.A1(new_n4699_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4700_));
  AOI21_X1   g02251(.A1(new_n4700_), .A2(new_n4698_), .B(new_n4662_), .ZN(new_n4701_));
  NOR2_X1    g02252(.A1(new_n4686_), .A2(new_n3235_), .ZN(new_n4702_));
  OAI21_X1   g02253(.A1(new_n4701_), .A2(pi0092), .B(new_n4702_), .ZN(new_n4703_));
  NAND2_X1   g02254(.A1(new_n4662_), .A2(pi0092), .ZN(new_n4704_));
  XNOR2_X1   g02255(.A1(new_n4704_), .A2(new_n3172_), .ZN(new_n4705_));
  NOR2_X1    g02256(.A1(new_n4705_), .A2(new_n4686_), .ZN(new_n4706_));
  INV_X1     g02257(.I(new_n4659_), .ZN(new_n4707_));
  NOR2_X1    g02258(.A1(new_n4651_), .A2(new_n3201_), .ZN(new_n4708_));
  XOR2_X1    g02259(.A1(new_n4708_), .A2(new_n3972_), .Z(new_n4709_));
  INV_X1     g02260(.I(pi0240), .ZN(new_n4710_));
  NAND2_X1   g02261(.A1(new_n3230_), .A2(new_n4710_), .ZN(new_n4711_));
  AOI21_X1   g02262(.A1(new_n4709_), .A2(new_n4707_), .B(new_n4711_), .ZN(new_n4712_));
  NOR2_X1    g02263(.A1(new_n4651_), .A2(new_n3219_), .ZN(new_n4713_));
  XOR2_X1    g02264(.A1(new_n4713_), .A2(new_n3797_), .Z(new_n4714_));
  OAI21_X1   g02265(.A1(new_n4714_), .A2(new_n4659_), .B(new_n3201_), .ZN(new_n4715_));
  NOR2_X1    g02266(.A1(new_n4712_), .A2(new_n4715_), .ZN(new_n4716_));
  NOR2_X1    g02267(.A1(new_n4651_), .A2(new_n3258_), .ZN(new_n4717_));
  XOR2_X1    g02268(.A1(new_n4717_), .A2(new_n3604_), .Z(new_n4718_));
  AOI21_X1   g02269(.A1(new_n4718_), .A2(new_n4707_), .B(pi0056), .ZN(new_n4719_));
  NAND2_X1   g02270(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n4720_));
  NOR4_X1    g02271(.A1(new_n4706_), .A2(new_n4716_), .A3(new_n4719_), .A4(new_n4720_), .ZN(new_n4721_));
  NOR2_X1    g02272(.A1(new_n4707_), .A2(new_n3230_), .ZN(new_n4722_));
  AOI21_X1   g02273(.A1(pi0216), .A2(pi0280), .B(new_n3612_), .ZN(new_n4723_));
  NAND2_X1   g02274(.A1(new_n4723_), .A2(pi0240), .ZN(new_n4724_));
  NOR2_X1    g02275(.A1(new_n4653_), .A2(new_n3385_), .ZN(new_n4725_));
  NOR2_X1    g02276(.A1(new_n4643_), .A2(new_n4647_), .ZN(new_n4726_));
  INV_X1     g02277(.I(new_n4726_), .ZN(new_n4727_));
  NOR3_X1    g02278(.A1(new_n3370_), .A2(new_n3111_), .A3(new_n4626_), .ZN(new_n4728_));
  OAI21_X1   g02279(.A1(new_n4727_), .A2(new_n4639_), .B(new_n4728_), .ZN(new_n4729_));
  XNOR2_X1   g02280(.A1(new_n4729_), .A2(new_n4655_), .ZN(new_n4730_));
  NAND2_X1   g02281(.A1(new_n4730_), .A2(pi0299), .ZN(new_n4731_));
  NAND2_X1   g02282(.A1(new_n4731_), .A2(new_n4725_), .ZN(new_n4732_));
  NOR2_X1    g02283(.A1(new_n4659_), .A2(new_n4723_), .ZN(new_n4733_));
  OAI21_X1   g02284(.A1(new_n4733_), .A2(new_n3098_), .B(new_n4725_), .ZN(new_n4734_));
  INV_X1     g02285(.I(new_n4734_), .ZN(new_n4735_));
  NOR2_X1    g02286(.A1(new_n4735_), .A2(new_n3134_), .ZN(new_n4736_));
  AOI21_X1   g02287(.A1(new_n4732_), .A2(new_n3134_), .B(new_n4736_), .ZN(new_n4737_));
  INV_X1     g02288(.I(new_n4737_), .ZN(new_n4738_));
  NAND3_X1   g02289(.A1(new_n3696_), .A2(pi0168), .A3(pi0878), .ZN(new_n4739_));
  NAND3_X1   g02290(.A1(new_n3459_), .A2(pi0168), .A3(new_n4637_), .ZN(new_n4740_));
  NAND2_X1   g02291(.A1(new_n3307_), .A2(pi0168), .ZN(new_n4741_));
  AOI21_X1   g02292(.A1(new_n4739_), .A2(new_n4740_), .B(new_n4741_), .ZN(new_n4742_));
  NAND2_X1   g02293(.A1(pi0228), .A2(pi0878), .ZN(new_n4743_));
  AOI21_X1   g02294(.A1(new_n3703_), .A2(new_n4644_), .B(new_n4743_), .ZN(new_n4744_));
  OAI21_X1   g02295(.A1(new_n4742_), .A2(new_n3330_), .B(new_n4744_), .ZN(new_n4745_));
  NAND2_X1   g02296(.A1(new_n4745_), .A2(new_n4647_), .ZN(new_n4746_));
  AOI21_X1   g02297(.A1(new_n4746_), .A2(new_n4654_), .B(new_n3098_), .ZN(new_n4747_));
  XOR2_X1    g02298(.A1(new_n4747_), .A2(new_n3855_), .Z(new_n4748_));
  NOR2_X1    g02299(.A1(pi0038), .A2(pi0100), .ZN(new_n4749_));
  INV_X1     g02300(.I(new_n4749_), .ZN(new_n4750_));
  AOI21_X1   g02301(.A1(new_n4732_), .A2(pi0039), .B(new_n4750_), .ZN(new_n4751_));
  OAI21_X1   g02302(.A1(new_n4680_), .A2(new_n4751_), .B(pi1137), .ZN(new_n4752_));
  NOR2_X1    g02303(.A1(new_n4748_), .A2(new_n4752_), .ZN(new_n4753_));
  OAI21_X1   g02304(.A1(new_n4691_), .A2(new_n4727_), .B(new_n4728_), .ZN(new_n4754_));
  XOR2_X1    g02305(.A1(new_n4754_), .A2(new_n4655_), .Z(new_n4755_));
  NOR2_X1    g02306(.A1(new_n4725_), .A2(new_n3211_), .ZN(new_n4756_));
  NOR2_X1    g02307(.A1(new_n4756_), .A2(new_n3098_), .ZN(new_n4757_));
  OAI21_X1   g02308(.A1(new_n4734_), .A2(new_n3211_), .B(pi0100), .ZN(new_n4758_));
  AOI21_X1   g02309(.A1(new_n4755_), .A2(new_n4757_), .B(new_n4758_), .ZN(new_n4759_));
  NOR4_X1    g02310(.A1(new_n4753_), .A2(new_n3235_), .A3(new_n3455_), .A4(new_n4759_), .ZN(new_n4760_));
  OAI21_X1   g02311(.A1(new_n4753_), .A2(new_n4759_), .B(pi0087), .ZN(new_n4761_));
  NOR2_X1    g02312(.A1(new_n4761_), .A2(new_n3694_), .ZN(new_n4762_));
  OAI21_X1   g02313(.A1(new_n4762_), .A2(new_n4760_), .B(new_n4738_), .ZN(new_n4763_));
  NAND2_X1   g02314(.A1(new_n4735_), .A2(pi0075), .ZN(new_n4764_));
  AOI21_X1   g02315(.A1(new_n4763_), .A2(new_n3303_), .B(new_n4764_), .ZN(new_n4765_));
  NAND2_X1   g02316(.A1(new_n4737_), .A2(pi0092), .ZN(new_n4766_));
  XOR2_X1    g02317(.A1(new_n4766_), .A2(new_n3172_), .Z(new_n4767_));
  NAND2_X1   g02318(.A1(new_n4767_), .A2(new_n4735_), .ZN(new_n4768_));
  NAND2_X1   g02319(.A1(new_n4730_), .A2(pi0062), .ZN(new_n4769_));
  XOR2_X1    g02320(.A1(new_n4769_), .A2(new_n3594_), .Z(new_n4770_));
  NAND2_X1   g02321(.A1(new_n4770_), .A2(new_n4733_), .ZN(new_n4771_));
  NAND3_X1   g02322(.A1(new_n4771_), .A2(pi0240), .A3(new_n3230_), .ZN(new_n4772_));
  NAND2_X1   g02323(.A1(new_n4730_), .A2(pi0056), .ZN(new_n4773_));
  XOR2_X1    g02324(.A1(new_n4773_), .A2(new_n3797_), .Z(new_n4774_));
  AOI21_X1   g02325(.A1(new_n4774_), .A2(new_n4733_), .B(pi0062), .ZN(new_n4775_));
  NAND2_X1   g02326(.A1(new_n4772_), .A2(new_n4775_), .ZN(new_n4776_));
  NAND2_X1   g02327(.A1(new_n4730_), .A2(pi0055), .ZN(new_n4777_));
  XOR2_X1    g02328(.A1(new_n4777_), .A2(new_n3605_), .Z(new_n4778_));
  NAND2_X1   g02329(.A1(new_n4778_), .A2(new_n4733_), .ZN(new_n4779_));
  NAND2_X1   g02330(.A1(new_n4779_), .A2(new_n3219_), .ZN(new_n4780_));
  NOR2_X1    g02331(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4781_));
  NAND4_X1   g02332(.A1(new_n4768_), .A2(new_n4776_), .A3(new_n4780_), .A4(new_n4781_), .ZN(new_n4782_));
  OAI22_X1   g02333(.A1(new_n4765_), .A2(new_n4782_), .B1(new_n4722_), .B2(new_n4724_), .ZN(new_n4783_));
  AOI21_X1   g02334(.A1(new_n4703_), .A2(new_n4721_), .B(new_n4783_), .ZN(po0162));
  INV_X1     g02335(.I(pi1136), .ZN(new_n4785_));
  INV_X1     g02336(.I(pi0266), .ZN(new_n4786_));
  AOI21_X1   g02337(.A1(new_n4786_), .A2(pi0224), .B(pi0222), .ZN(new_n4787_));
  INV_X1     g02338(.I(new_n4787_), .ZN(new_n4788_));
  NOR2_X1    g02339(.A1(pi0224), .A2(pi0875), .ZN(new_n4789_));
  AOI21_X1   g02340(.A1(new_n4788_), .A2(new_n4789_), .B(new_n2820_), .ZN(new_n4790_));
  NAND3_X1   g02341(.A1(new_n3103_), .A2(pi0222), .A3(pi0928), .ZN(new_n4791_));
  INV_X1     g02342(.I(pi0928), .ZN(new_n4792_));
  NAND3_X1   g02343(.A1(new_n3344_), .A2(pi0222), .A3(new_n4792_), .ZN(new_n4793_));
  AOI21_X1   g02344(.A1(new_n4793_), .A2(new_n4791_), .B(new_n4785_), .ZN(new_n4794_));
  NOR2_X1    g02345(.A1(new_n4794_), .A2(new_n4790_), .ZN(new_n4795_));
  NOR2_X1    g02346(.A1(new_n4795_), .A2(new_n3090_), .ZN(new_n4796_));
  XOR2_X1    g02347(.A1(new_n4796_), .A2(new_n3565_), .Z(new_n4797_));
  NOR2_X1    g02348(.A1(new_n4797_), .A2(new_n4785_), .ZN(new_n4798_));
  NOR2_X1    g02349(.A1(new_n3121_), .A2(pi0928), .ZN(new_n4799_));
  XOR2_X1    g02350(.A1(new_n3356_), .A2(new_n4799_), .Z(new_n4800_));
  NAND2_X1   g02351(.A1(new_n4800_), .A2(pi1136), .ZN(new_n4801_));
  NAND2_X1   g02352(.A1(new_n4801_), .A2(pi0215), .ZN(new_n4802_));
  NOR3_X1    g02353(.A1(new_n3111_), .A2(new_n4786_), .A3(new_n4785_), .ZN(new_n4803_));
  NOR2_X1    g02354(.A1(new_n3145_), .A2(new_n3005_), .ZN(new_n4804_));
  NOR2_X1    g02355(.A1(new_n3145_), .A2(pi0875), .ZN(new_n4805_));
  XOR2_X1    g02356(.A1(new_n4804_), .A2(new_n4805_), .Z(new_n4806_));
  NAND2_X1   g02357(.A1(new_n4806_), .A2(pi0166), .ZN(new_n4807_));
  INV_X1     g02358(.I(pi0166), .ZN(new_n4808_));
  INV_X1     g02359(.I(pi0875), .ZN(new_n4809_));
  NOR4_X1    g02360(.A1(new_n2820_), .A2(new_n3004_), .A3(new_n4808_), .A4(new_n4809_), .ZN(new_n4810_));
  NOR2_X1    g02361(.A1(new_n4808_), .A2(new_n4809_), .ZN(new_n4811_));
  NOR3_X1    g02362(.A1(new_n4811_), .A2(new_n2753_), .A3(new_n3004_), .ZN(new_n4812_));
  NOR2_X1    g02363(.A1(new_n4810_), .A2(new_n4812_), .ZN(new_n4813_));
  INV_X1     g02364(.I(new_n4813_), .ZN(new_n4814_));
  AOI21_X1   g02365(.A1(new_n4814_), .A2(pi0228), .B(new_n3369_), .ZN(new_n4815_));
  AOI21_X1   g02366(.A1(new_n4807_), .A2(new_n4815_), .B(new_n3011_), .ZN(new_n4816_));
  XOR2_X1    g02367(.A1(new_n4816_), .A2(new_n3373_), .Z(new_n4817_));
  NAND2_X1   g02368(.A1(new_n4817_), .A2(new_n4803_), .ZN(new_n4818_));
  XNOR2_X1   g02369(.A1(new_n4818_), .A2(new_n4802_), .ZN(new_n4819_));
  AOI21_X1   g02370(.A1(new_n4819_), .A2(pi0299), .B(new_n4798_), .ZN(new_n4820_));
  NOR2_X1    g02371(.A1(new_n4820_), .A2(new_n3474_), .ZN(new_n4821_));
  INV_X1     g02372(.I(new_n3373_), .ZN(new_n4822_));
  AOI21_X1   g02373(.A1(new_n4808_), .A2(new_n3005_), .B(new_n3011_), .ZN(new_n4823_));
  OAI21_X1   g02374(.A1(new_n4814_), .A2(new_n3005_), .B(new_n4823_), .ZN(new_n4824_));
  XOR2_X1    g02375(.A1(new_n4824_), .A2(new_n4822_), .Z(new_n4825_));
  NAND2_X1   g02376(.A1(new_n4825_), .A2(new_n4803_), .ZN(new_n4826_));
  XNOR2_X1   g02377(.A1(new_n4826_), .A2(new_n4802_), .ZN(new_n4827_));
  NOR2_X1    g02378(.A1(new_n4827_), .A2(new_n3913_), .ZN(new_n4828_));
  INV_X1     g02379(.I(new_n4828_), .ZN(new_n4829_));
  AOI21_X1   g02380(.A1(new_n4829_), .A2(pi0299), .B(new_n4798_), .ZN(new_n4830_));
  INV_X1     g02381(.I(new_n4830_), .ZN(new_n4831_));
  AOI21_X1   g02382(.A1(new_n3474_), .A2(new_n4831_), .B(new_n4821_), .ZN(new_n4832_));
  INV_X1     g02383(.I(new_n4801_), .ZN(new_n4833_));
  NOR2_X1    g02384(.A1(new_n3330_), .A2(new_n4808_), .ZN(new_n4834_));
  XOR2_X1    g02385(.A1(new_n4834_), .A2(new_n4811_), .Z(new_n4835_));
  NOR2_X1    g02386(.A1(new_n3005_), .A2(new_n4809_), .ZN(new_n4836_));
  OAI21_X1   g02387(.A1(new_n3696_), .A2(new_n4836_), .B(pi0166), .ZN(new_n4837_));
  NOR3_X1    g02388(.A1(new_n3309_), .A2(pi0216), .A3(pi0228), .ZN(new_n4838_));
  NOR2_X1    g02389(.A1(new_n4838_), .A2(new_n4813_), .ZN(new_n4839_));
  NOR2_X1    g02390(.A1(new_n3011_), .A2(new_n4786_), .ZN(new_n4840_));
  NAND2_X1   g02391(.A1(new_n4839_), .A2(new_n4840_), .ZN(new_n4841_));
  AOI21_X1   g02392(.A1(new_n4837_), .A2(new_n4841_), .B(new_n3308_), .ZN(new_n4842_));
  AOI21_X1   g02393(.A1(new_n4835_), .A2(new_n4842_), .B(pi0221), .ZN(new_n4843_));
  OAI21_X1   g02394(.A1(new_n4843_), .A2(new_n4833_), .B(pi0299), .ZN(new_n4844_));
  XOR2_X1    g02395(.A1(new_n4844_), .A2(new_n3855_), .Z(new_n4845_));
  NOR2_X1    g02396(.A1(new_n3306_), .A2(new_n3092_), .ZN(new_n4846_));
  INV_X1     g02397(.I(new_n4846_), .ZN(new_n4847_));
  OAI21_X1   g02398(.A1(new_n3183_), .A2(pi0299), .B(new_n3090_), .ZN(new_n4848_));
  NAND3_X1   g02399(.A1(new_n4847_), .A2(new_n4795_), .A3(new_n4848_), .ZN(new_n4849_));
  NOR2_X1    g02400(.A1(pi0038), .A2(pi0100), .ZN(new_n4850_));
  OAI21_X1   g02401(.A1(new_n4820_), .A2(new_n3183_), .B(new_n4850_), .ZN(new_n4851_));
  AOI21_X1   g02402(.A1(new_n4851_), .A2(new_n4849_), .B(new_n4785_), .ZN(new_n4852_));
  NAND2_X1   g02403(.A1(new_n4845_), .A2(new_n4852_), .ZN(new_n4853_));
  NOR3_X1    g02404(.A1(new_n3396_), .A2(new_n4809_), .A3(new_n2786_), .ZN(new_n4854_));
  NOR3_X1    g02405(.A1(new_n3393_), .A2(new_n4809_), .A3(new_n2785_), .ZN(new_n4855_));
  NOR2_X1    g02406(.A1(new_n3392_), .A2(new_n3005_), .ZN(new_n4856_));
  OAI21_X1   g02407(.A1(new_n4854_), .A2(new_n4855_), .B(new_n4856_), .ZN(new_n4857_));
  NAND2_X1   g02408(.A1(new_n4857_), .A2(new_n4808_), .ZN(new_n4858_));
  NAND3_X1   g02409(.A1(new_n4858_), .A2(new_n4809_), .A3(new_n3391_), .ZN(new_n4859_));
  AOI21_X1   g02410(.A1(new_n4859_), .A2(new_n4815_), .B(new_n3011_), .ZN(new_n4860_));
  XOR2_X1    g02411(.A1(new_n4860_), .A2(new_n3373_), .Z(new_n4861_));
  NAND2_X1   g02412(.A1(new_n4861_), .A2(new_n4803_), .ZN(new_n4862_));
  XNOR2_X1   g02413(.A1(new_n4862_), .A2(new_n4802_), .ZN(new_n4863_));
  OAI21_X1   g02414(.A1(new_n4798_), .A2(new_n3211_), .B(pi0299), .ZN(new_n4864_));
  AOI21_X1   g02415(.A1(new_n4830_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4865_));
  OAI21_X1   g02416(.A1(new_n4863_), .A2(new_n4864_), .B(new_n4865_), .ZN(new_n4866_));
  NAND4_X1   g02417(.A1(new_n4853_), .A2(pi0075), .A3(pi0087), .A4(new_n4866_), .ZN(new_n4867_));
  NAND2_X1   g02418(.A1(new_n4853_), .A2(new_n4866_), .ZN(new_n4868_));
  NAND3_X1   g02419(.A1(new_n4868_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4869_));
  AOI21_X1   g02420(.A1(new_n4869_), .A2(new_n4867_), .B(new_n4832_), .ZN(new_n4870_));
  NOR2_X1    g02421(.A1(new_n4831_), .A2(new_n3235_), .ZN(new_n4871_));
  OAI21_X1   g02422(.A1(new_n4870_), .A2(pi0092), .B(new_n4871_), .ZN(new_n4872_));
  NAND2_X1   g02423(.A1(new_n4832_), .A2(pi0092), .ZN(new_n4873_));
  XOR2_X1    g02424(.A1(new_n4873_), .A2(new_n3172_), .Z(new_n4874_));
  NAND2_X1   g02425(.A1(new_n4819_), .A2(pi0055), .ZN(new_n4875_));
  XOR2_X1    g02426(.A1(new_n4875_), .A2(new_n3604_), .Z(new_n4876_));
  OAI21_X1   g02427(.A1(new_n4876_), .A2(new_n4829_), .B(new_n3219_), .ZN(new_n4877_));
  NOR2_X1    g02428(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4878_));
  NAND2_X1   g02429(.A1(new_n4877_), .A2(new_n4878_), .ZN(new_n4879_));
  AOI21_X1   g02430(.A1(new_n4874_), .A2(new_n4830_), .B(new_n4879_), .ZN(new_n4880_));
  NAND2_X1   g02431(.A1(new_n4819_), .A2(pi0056), .ZN(new_n4881_));
  XOR2_X1    g02432(.A1(new_n4881_), .A2(new_n3599_), .Z(new_n4882_));
  OAI21_X1   g02433(.A1(new_n4882_), .A2(new_n4829_), .B(new_n3201_), .ZN(new_n4883_));
  AOI21_X1   g02434(.A1(new_n4872_), .A2(new_n4880_), .B(new_n4883_), .ZN(new_n4884_));
  NAND2_X1   g02435(.A1(new_n4819_), .A2(pi0062), .ZN(new_n4885_));
  XOR2_X1    g02436(.A1(new_n4885_), .A2(new_n3972_), .Z(new_n4886_));
  NOR2_X1    g02437(.A1(new_n3426_), .A2(pi0245), .ZN(new_n4887_));
  OAI21_X1   g02438(.A1(new_n4886_), .A2(new_n4829_), .B(new_n4887_), .ZN(new_n4888_));
  NAND2_X1   g02439(.A1(new_n4798_), .A2(new_n3128_), .ZN(new_n4889_));
  AOI21_X1   g02440(.A1(new_n4889_), .A2(new_n4809_), .B(new_n2820_), .ZN(new_n4890_));
  OAI21_X1   g02441(.A1(new_n4813_), .A2(new_n3005_), .B(pi0216), .ZN(new_n4891_));
  INV_X1     g02442(.I(new_n4840_), .ZN(new_n4892_));
  NOR2_X1    g02443(.A1(new_n4807_), .A2(new_n4892_), .ZN(new_n4893_));
  NOR2_X1    g02444(.A1(new_n4893_), .A2(new_n4891_), .ZN(new_n4894_));
  NAND2_X1   g02445(.A1(new_n4893_), .A2(new_n4891_), .ZN(new_n4895_));
  NAND2_X1   g02446(.A1(new_n4895_), .A2(new_n3121_), .ZN(new_n4896_));
  NOR2_X1    g02447(.A1(new_n4896_), .A2(new_n4894_), .ZN(new_n4897_));
  NAND2_X1   g02448(.A1(new_n4801_), .A2(new_n3111_), .ZN(new_n4898_));
  OAI22_X1   g02449(.A1(new_n4897_), .A2(new_n4898_), .B1(new_n3111_), .B2(pi1136), .ZN(new_n4899_));
  NOR2_X1    g02450(.A1(new_n4899_), .A2(new_n3098_), .ZN(new_n4900_));
  NOR2_X1    g02451(.A1(new_n4900_), .A2(new_n4890_), .ZN(new_n4901_));
  INV_X1     g02452(.I(new_n4901_), .ZN(new_n4902_));
  AOI21_X1   g02453(.A1(new_n4827_), .A2(pi0299), .B(new_n4890_), .ZN(new_n4903_));
  NOR2_X1    g02454(.A1(new_n4903_), .A2(new_n3134_), .ZN(new_n4904_));
  AOI21_X1   g02455(.A1(new_n4902_), .A2(new_n3134_), .B(new_n4904_), .ZN(new_n4905_));
  NOR2_X1    g02456(.A1(pi0166), .A2(pi0875), .ZN(new_n4906_));
  OAI21_X1   g02457(.A1(new_n3459_), .A2(new_n4906_), .B(new_n4839_), .ZN(new_n4907_));
  NAND2_X1   g02458(.A1(new_n4839_), .A2(pi0228), .ZN(new_n4908_));
  XNOR2_X1   g02459(.A1(new_n4907_), .A2(new_n4908_), .ZN(new_n4909_));
  OAI22_X1   g02460(.A1(new_n4909_), .A2(new_n3931_), .B1(new_n3121_), .B2(new_n4801_), .ZN(new_n4910_));
  NAND4_X1   g02461(.A1(new_n4910_), .A2(pi0215), .A3(pi0299), .A4(new_n4840_), .ZN(new_n4911_));
  NAND2_X1   g02462(.A1(new_n4910_), .A2(new_n4840_), .ZN(new_n4912_));
  NAND3_X1   g02463(.A1(new_n4912_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n4913_));
  AOI21_X1   g02464(.A1(new_n4902_), .A2(pi0039), .B(pi0038), .ZN(new_n4914_));
  AOI21_X1   g02465(.A1(pi0223), .A2(pi1136), .B(pi0299), .ZN(new_n4915_));
  OR2_X2     g02466(.A1(new_n4794_), .A2(new_n4915_), .Z(new_n4916_));
  NAND3_X1   g02467(.A1(new_n4846_), .A2(new_n4790_), .A3(new_n4916_), .ZN(new_n4917_));
  NAND2_X1   g02468(.A1(new_n4849_), .A2(new_n4917_), .ZN(new_n4918_));
  OAI21_X1   g02469(.A1(new_n4914_), .A2(new_n4918_), .B(pi1136), .ZN(new_n4919_));
  AOI21_X1   g02470(.A1(new_n4913_), .A2(new_n4911_), .B(new_n4919_), .ZN(new_n4920_));
  INV_X1     g02471(.I(new_n4903_), .ZN(new_n4921_));
  NOR2_X1    g02472(.A1(new_n4921_), .A2(new_n3259_), .ZN(new_n4922_));
  OAI21_X1   g02473(.A1(new_n4920_), .A2(pi0100), .B(new_n4922_), .ZN(new_n4923_));
  NOR2_X1    g02474(.A1(new_n4859_), .A2(new_n4892_), .ZN(new_n4924_));
  NOR2_X1    g02475(.A1(new_n4924_), .A2(new_n4891_), .ZN(new_n4925_));
  NAND2_X1   g02476(.A1(new_n4924_), .A2(new_n4891_), .ZN(new_n4926_));
  NAND2_X1   g02477(.A1(new_n4926_), .A2(new_n3121_), .ZN(new_n4927_));
  OAI21_X1   g02478(.A1(new_n4927_), .A2(new_n4925_), .B(new_n4801_), .ZN(new_n4928_));
  NAND2_X1   g02479(.A1(new_n4928_), .A2(pi0299), .ZN(new_n4929_));
  XOR2_X1    g02480(.A1(new_n4929_), .A2(new_n3695_), .Z(new_n4930_));
  NOR2_X1    g02481(.A1(new_n4930_), .A2(new_n4785_), .ZN(new_n4931_));
  OR2_X2     g02482(.A1(new_n4890_), .A2(new_n3212_), .Z(new_n4932_));
  AOI21_X1   g02483(.A1(new_n4903_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n4933_));
  OAI21_X1   g02484(.A1(new_n4931_), .A2(new_n4932_), .B(new_n4933_), .ZN(new_n4934_));
  NAND4_X1   g02485(.A1(new_n4923_), .A2(pi0075), .A3(pi0087), .A4(new_n4934_), .ZN(new_n4935_));
  NAND2_X1   g02486(.A1(new_n4923_), .A2(new_n4934_), .ZN(new_n4936_));
  NAND3_X1   g02487(.A1(new_n4936_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n4937_));
  AOI21_X1   g02488(.A1(new_n4937_), .A2(new_n4935_), .B(new_n4905_), .ZN(new_n4938_));
  NOR2_X1    g02489(.A1(new_n4921_), .A2(new_n3235_), .ZN(new_n4939_));
  OAI21_X1   g02490(.A1(new_n4938_), .A2(pi0092), .B(new_n4939_), .ZN(new_n4940_));
  NAND2_X1   g02491(.A1(new_n4905_), .A2(pi0092), .ZN(new_n4941_));
  XOR2_X1    g02492(.A1(new_n4941_), .A2(new_n3172_), .Z(new_n4942_));
  NOR2_X1    g02493(.A1(new_n4899_), .A2(new_n3258_), .ZN(new_n4943_));
  XOR2_X1    g02494(.A1(new_n4943_), .A2(new_n3605_), .Z(new_n4944_));
  OAI21_X1   g02495(.A1(new_n4944_), .A2(new_n4827_), .B(new_n3219_), .ZN(new_n4945_));
  NOR2_X1    g02496(.A1(new_n3203_), .A2(pi0055), .ZN(new_n4946_));
  NAND2_X1   g02497(.A1(new_n4945_), .A2(new_n4946_), .ZN(new_n4947_));
  AOI21_X1   g02498(.A1(new_n4942_), .A2(new_n4903_), .B(new_n4947_), .ZN(new_n4948_));
  NOR2_X1    g02499(.A1(new_n4899_), .A2(new_n3219_), .ZN(new_n4949_));
  XOR2_X1    g02500(.A1(new_n4949_), .A2(new_n3797_), .Z(new_n4950_));
  OAI21_X1   g02501(.A1(new_n4950_), .A2(new_n4827_), .B(new_n3201_), .ZN(new_n4951_));
  AOI21_X1   g02502(.A1(new_n4940_), .A2(new_n4948_), .B(new_n4951_), .ZN(new_n4952_));
  NOR2_X1    g02503(.A1(new_n4899_), .A2(new_n3201_), .ZN(new_n4953_));
  XOR2_X1    g02504(.A1(new_n4953_), .A2(new_n3594_), .Z(new_n4954_));
  INV_X1     g02505(.I(pi0245), .ZN(new_n4955_));
  NOR2_X1    g02506(.A1(new_n3426_), .A2(new_n4955_), .ZN(new_n4956_));
  OAI21_X1   g02507(.A1(new_n4954_), .A2(new_n4827_), .B(new_n4956_), .ZN(new_n4957_));
  OAI22_X1   g02508(.A1(new_n4884_), .A2(new_n4888_), .B1(new_n4952_), .B2(new_n4957_), .ZN(po0163));
  INV_X1     g02509(.I(pi1135), .ZN(new_n4959_));
  NAND3_X1   g02510(.A1(new_n3103_), .A2(pi0222), .A3(pi0938), .ZN(new_n4960_));
  INV_X1     g02511(.I(pi0938), .ZN(new_n4961_));
  NAND3_X1   g02512(.A1(new_n3344_), .A2(pi0222), .A3(new_n4961_), .ZN(new_n4962_));
  AOI21_X1   g02513(.A1(new_n4962_), .A2(new_n4960_), .B(new_n4959_), .ZN(new_n4963_));
  INV_X1     g02514(.I(pi0279), .ZN(new_n4964_));
  AOI21_X1   g02515(.A1(new_n4964_), .A2(pi0224), .B(pi0222), .ZN(new_n4965_));
  INV_X1     g02516(.I(new_n4965_), .ZN(new_n4966_));
  NOR2_X1    g02517(.A1(pi0224), .A2(pi0879), .ZN(new_n4967_));
  AOI21_X1   g02518(.A1(new_n4966_), .A2(new_n4967_), .B(new_n2820_), .ZN(new_n4968_));
  NOR2_X1    g02519(.A1(new_n4963_), .A2(new_n4968_), .ZN(new_n4969_));
  NOR2_X1    g02520(.A1(new_n4969_), .A2(new_n3090_), .ZN(new_n4970_));
  XOR2_X1    g02521(.A1(new_n4970_), .A2(new_n3565_), .Z(new_n4971_));
  NOR2_X1    g02522(.A1(new_n4971_), .A2(new_n4959_), .ZN(new_n4972_));
  NOR2_X1    g02523(.A1(new_n3121_), .A2(pi0938), .ZN(new_n4973_));
  XOR2_X1    g02524(.A1(new_n3356_), .A2(new_n4973_), .Z(new_n4974_));
  NAND2_X1   g02525(.A1(new_n4974_), .A2(pi1135), .ZN(new_n4975_));
  NAND2_X1   g02526(.A1(new_n4975_), .A2(pi0215), .ZN(new_n4976_));
  NOR3_X1    g02527(.A1(new_n3111_), .A2(new_n4964_), .A3(new_n4959_), .ZN(new_n4977_));
  NOR2_X1    g02528(.A1(new_n3145_), .A2(pi0879), .ZN(new_n4978_));
  XOR2_X1    g02529(.A1(new_n4804_), .A2(new_n4978_), .Z(new_n4979_));
  NAND2_X1   g02530(.A1(new_n4979_), .A2(pi0161), .ZN(new_n4980_));
  INV_X1     g02531(.I(pi0161), .ZN(new_n4981_));
  INV_X1     g02532(.I(pi0879), .ZN(new_n4982_));
  NOR4_X1    g02533(.A1(new_n2820_), .A2(new_n3004_), .A3(new_n4981_), .A4(new_n4982_), .ZN(new_n4983_));
  NOR2_X1    g02534(.A1(new_n4981_), .A2(new_n4982_), .ZN(new_n4984_));
  NOR3_X1    g02535(.A1(new_n4984_), .A2(new_n2753_), .A3(new_n3004_), .ZN(new_n4985_));
  NOR2_X1    g02536(.A1(new_n4983_), .A2(new_n4985_), .ZN(new_n4986_));
  INV_X1     g02537(.I(new_n4986_), .ZN(new_n4987_));
  AOI21_X1   g02538(.A1(new_n4987_), .A2(pi0228), .B(new_n3369_), .ZN(new_n4988_));
  AOI21_X1   g02539(.A1(new_n4980_), .A2(new_n4988_), .B(new_n3011_), .ZN(new_n4989_));
  XOR2_X1    g02540(.A1(new_n4989_), .A2(new_n3373_), .Z(new_n4990_));
  NAND2_X1   g02541(.A1(new_n4990_), .A2(new_n4977_), .ZN(new_n4991_));
  XNOR2_X1   g02542(.A1(new_n4991_), .A2(new_n4976_), .ZN(new_n4992_));
  AOI21_X1   g02543(.A1(new_n4992_), .A2(pi0299), .B(new_n4972_), .ZN(new_n4993_));
  NOR2_X1    g02544(.A1(new_n4993_), .A2(new_n3474_), .ZN(new_n4994_));
  AOI21_X1   g02545(.A1(new_n4981_), .A2(new_n3005_), .B(new_n3011_), .ZN(new_n4995_));
  OAI21_X1   g02546(.A1(new_n4987_), .A2(new_n3005_), .B(new_n4995_), .ZN(new_n4996_));
  XOR2_X1    g02547(.A1(new_n4996_), .A2(new_n4822_), .Z(new_n4997_));
  NAND2_X1   g02548(.A1(new_n4997_), .A2(new_n4977_), .ZN(new_n4998_));
  XNOR2_X1   g02549(.A1(new_n4998_), .A2(new_n4976_), .ZN(new_n4999_));
  NOR2_X1    g02550(.A1(new_n4999_), .A2(new_n3913_), .ZN(new_n5000_));
  INV_X1     g02551(.I(new_n5000_), .ZN(new_n5001_));
  AOI21_X1   g02552(.A1(new_n5001_), .A2(pi0299), .B(new_n4972_), .ZN(new_n5002_));
  INV_X1     g02553(.I(new_n5002_), .ZN(new_n5003_));
  AOI21_X1   g02554(.A1(new_n3474_), .A2(new_n5003_), .B(new_n4994_), .ZN(new_n5004_));
  NAND3_X1   g02555(.A1(new_n3330_), .A2(pi0161), .A3(pi0879), .ZN(new_n5005_));
  NAND3_X1   g02556(.A1(new_n3862_), .A2(pi0161), .A3(new_n4982_), .ZN(new_n5006_));
  NAND2_X1   g02557(.A1(pi0228), .A2(pi0879), .ZN(new_n5007_));
  AOI21_X1   g02558(.A1(new_n3459_), .A2(new_n5007_), .B(new_n4981_), .ZN(new_n5008_));
  NOR2_X1    g02559(.A1(new_n3011_), .A2(new_n4964_), .ZN(new_n5009_));
  INV_X1     g02560(.I(new_n5009_), .ZN(new_n5010_));
  NOR3_X1    g02561(.A1(new_n4838_), .A2(new_n4986_), .A3(new_n5010_), .ZN(new_n5011_));
  OAI21_X1   g02562(.A1(new_n5008_), .A2(new_n5011_), .B(new_n3307_), .ZN(new_n5012_));
  AOI21_X1   g02563(.A1(new_n5006_), .A2(new_n5005_), .B(new_n5012_), .ZN(new_n5013_));
  OAI21_X1   g02564(.A1(new_n5013_), .A2(pi0221), .B(new_n4975_), .ZN(new_n5014_));
  OR3_X2     g02565(.A1(new_n5014_), .A2(new_n3111_), .A3(new_n3098_), .Z(new_n5015_));
  NAND3_X1   g02566(.A1(new_n5014_), .A2(new_n3111_), .A3(pi0299), .ZN(new_n5016_));
  AOI21_X1   g02567(.A1(new_n5015_), .A2(new_n5016_), .B(new_n4959_), .ZN(new_n5017_));
  NAND2_X1   g02568(.A1(new_n3090_), .A2(new_n3098_), .ZN(new_n5018_));
  AOI21_X1   g02569(.A1(new_n4847_), .A2(new_n4969_), .B(new_n5018_), .ZN(new_n5019_));
  OAI21_X1   g02570(.A1(new_n5017_), .A2(pi0039), .B(new_n5019_), .ZN(new_n5020_));
  NAND2_X1   g02571(.A1(new_n4993_), .A2(pi0039), .ZN(new_n5021_));
  AOI21_X1   g02572(.A1(new_n5020_), .A2(new_n3259_), .B(new_n5021_), .ZN(new_n5022_));
  NOR2_X1    g02573(.A1(new_n5003_), .A2(new_n3259_), .ZN(new_n5023_));
  OAI21_X1   g02574(.A1(new_n5022_), .A2(pi0100), .B(new_n5023_), .ZN(new_n5024_));
  NOR4_X1    g02575(.A1(new_n3396_), .A2(pi0152), .A3(pi0166), .A4(new_n4982_), .ZN(new_n5025_));
  NOR2_X1    g02576(.A1(pi0152), .A2(pi0166), .ZN(new_n5026_));
  NOR3_X1    g02577(.A1(new_n3393_), .A2(new_n4982_), .A3(new_n5026_), .ZN(new_n5027_));
  OAI21_X1   g02578(.A1(new_n5027_), .A2(new_n5025_), .B(new_n4856_), .ZN(new_n5028_));
  NAND2_X1   g02579(.A1(new_n5028_), .A2(new_n4981_), .ZN(new_n5029_));
  NAND3_X1   g02580(.A1(new_n5029_), .A2(new_n4982_), .A3(new_n3391_), .ZN(new_n5030_));
  AOI21_X1   g02581(.A1(new_n5030_), .A2(new_n4988_), .B(new_n3011_), .ZN(new_n5031_));
  XOR2_X1    g02582(.A1(new_n5031_), .A2(new_n3373_), .Z(new_n5032_));
  NAND2_X1   g02583(.A1(new_n5032_), .A2(new_n4977_), .ZN(new_n5033_));
  XNOR2_X1   g02584(.A1(new_n5033_), .A2(new_n4976_), .ZN(new_n5034_));
  OAI21_X1   g02585(.A1(new_n4972_), .A2(new_n3211_), .B(pi0299), .ZN(new_n5035_));
  AOI21_X1   g02586(.A1(new_n5002_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n5036_));
  OAI21_X1   g02587(.A1(new_n5034_), .A2(new_n5035_), .B(new_n5036_), .ZN(new_n5037_));
  NAND4_X1   g02588(.A1(new_n5024_), .A2(pi0075), .A3(pi0087), .A4(new_n5037_), .ZN(new_n5038_));
  NAND2_X1   g02589(.A1(new_n5024_), .A2(new_n5037_), .ZN(new_n5039_));
  NAND3_X1   g02590(.A1(new_n5039_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n5040_));
  AOI21_X1   g02591(.A1(new_n5040_), .A2(new_n5038_), .B(new_n5004_), .ZN(new_n5041_));
  NOR2_X1    g02592(.A1(new_n5003_), .A2(new_n3235_), .ZN(new_n5042_));
  OAI21_X1   g02593(.A1(new_n5041_), .A2(pi0092), .B(new_n5042_), .ZN(new_n5043_));
  NAND2_X1   g02594(.A1(new_n5004_), .A2(pi0092), .ZN(new_n5044_));
  XOR2_X1    g02595(.A1(new_n5044_), .A2(new_n3172_), .Z(new_n5045_));
  NAND2_X1   g02596(.A1(new_n4992_), .A2(pi0055), .ZN(new_n5046_));
  XOR2_X1    g02597(.A1(new_n5046_), .A2(new_n3604_), .Z(new_n5047_));
  OAI21_X1   g02598(.A1(new_n5047_), .A2(new_n5001_), .B(new_n3219_), .ZN(new_n5048_));
  NOR2_X1    g02599(.A1(new_n3203_), .A2(pi0055), .ZN(new_n5049_));
  NAND2_X1   g02600(.A1(new_n5048_), .A2(new_n5049_), .ZN(new_n5050_));
  AOI21_X1   g02601(.A1(new_n5045_), .A2(new_n5002_), .B(new_n5050_), .ZN(new_n5051_));
  NAND2_X1   g02602(.A1(new_n4992_), .A2(pi0056), .ZN(new_n5052_));
  XOR2_X1    g02603(.A1(new_n5052_), .A2(new_n3599_), .Z(new_n5053_));
  OAI21_X1   g02604(.A1(new_n5053_), .A2(new_n5001_), .B(new_n3201_), .ZN(new_n5054_));
  AOI21_X1   g02605(.A1(new_n5043_), .A2(new_n5051_), .B(new_n5054_), .ZN(new_n5055_));
  NAND2_X1   g02606(.A1(new_n4992_), .A2(pi0062), .ZN(new_n5056_));
  XOR2_X1    g02607(.A1(new_n5056_), .A2(new_n3972_), .Z(new_n5057_));
  NOR2_X1    g02608(.A1(new_n3426_), .A2(pi0244), .ZN(new_n5058_));
  OAI21_X1   g02609(.A1(new_n5057_), .A2(new_n5001_), .B(new_n5058_), .ZN(new_n5059_));
  NAND2_X1   g02610(.A1(new_n4972_), .A2(new_n3128_), .ZN(new_n5060_));
  AOI21_X1   g02611(.A1(new_n5060_), .A2(new_n4982_), .B(new_n2820_), .ZN(new_n5061_));
  AOI21_X1   g02612(.A1(new_n4999_), .A2(pi0299), .B(new_n5061_), .ZN(new_n5062_));
  INV_X1     g02613(.I(new_n5062_), .ZN(new_n5063_));
  INV_X1     g02614(.I(new_n5061_), .ZN(new_n5064_));
  OAI21_X1   g02615(.A1(new_n4986_), .A2(new_n3005_), .B(pi0216), .ZN(new_n5065_));
  NOR2_X1    g02616(.A1(new_n4980_), .A2(new_n5010_), .ZN(new_n5066_));
  NOR2_X1    g02617(.A1(new_n5066_), .A2(new_n5065_), .ZN(new_n5067_));
  NAND2_X1   g02618(.A1(new_n5066_), .A2(new_n5065_), .ZN(new_n5068_));
  NAND2_X1   g02619(.A1(new_n5068_), .A2(new_n3121_), .ZN(new_n5069_));
  NOR2_X1    g02620(.A1(new_n5069_), .A2(new_n5067_), .ZN(new_n5070_));
  NAND2_X1   g02621(.A1(new_n4975_), .A2(new_n3111_), .ZN(new_n5071_));
  OAI22_X1   g02622(.A1(new_n5070_), .A2(new_n5071_), .B1(new_n3111_), .B2(pi1135), .ZN(new_n5072_));
  OAI21_X1   g02623(.A1(new_n5072_), .A2(new_n3098_), .B(new_n5064_), .ZN(new_n5073_));
  NOR2_X1    g02624(.A1(new_n5062_), .A2(new_n3134_), .ZN(new_n5074_));
  AOI21_X1   g02625(.A1(new_n5073_), .A2(new_n3134_), .B(new_n5074_), .ZN(new_n5075_));
  NOR2_X1    g02626(.A1(new_n4838_), .A2(new_n4986_), .ZN(new_n5076_));
  NAND2_X1   g02627(.A1(new_n4981_), .A2(new_n4982_), .ZN(new_n5077_));
  NAND4_X1   g02628(.A1(new_n3696_), .A2(pi0228), .A3(new_n5076_), .A4(new_n5077_), .ZN(new_n5078_));
  NAND2_X1   g02629(.A1(new_n3696_), .A2(new_n5077_), .ZN(new_n5079_));
  NAND3_X1   g02630(.A1(new_n5079_), .A2(new_n3005_), .A3(new_n5076_), .ZN(new_n5080_));
  AOI21_X1   g02631(.A1(new_n5080_), .A2(new_n5078_), .B(new_n3931_), .ZN(new_n5081_));
  NOR2_X1    g02632(.A1(new_n4975_), .A2(new_n3121_), .ZN(new_n5082_));
  OAI21_X1   g02633(.A1(new_n5081_), .A2(new_n5082_), .B(new_n5009_), .ZN(new_n5083_));
  OR3_X2     g02634(.A1(new_n5083_), .A2(new_n3111_), .A3(new_n3098_), .Z(new_n5084_));
  NAND3_X1   g02635(.A1(new_n5083_), .A2(pi0299), .A3(new_n3855_), .ZN(new_n5085_));
  AOI21_X1   g02636(.A1(new_n5084_), .A2(new_n5085_), .B(new_n4959_), .ZN(new_n5086_));
  NOR2_X1    g02637(.A1(new_n3090_), .A2(new_n4959_), .ZN(new_n5087_));
  AOI21_X1   g02638(.A1(new_n4963_), .A2(pi0223), .B(new_n4968_), .ZN(new_n5088_));
  NOR4_X1    g02639(.A1(new_n4847_), .A2(pi0299), .A3(new_n5087_), .A4(new_n5088_), .ZN(new_n5089_));
  OAI21_X1   g02640(.A1(new_n5086_), .A2(pi0039), .B(new_n5089_), .ZN(new_n5090_));
  OR2_X2     g02641(.A1(new_n5073_), .A2(new_n3183_), .Z(new_n5091_));
  AOI21_X1   g02642(.A1(new_n5090_), .A2(new_n3259_), .B(new_n5091_), .ZN(new_n5092_));
  NOR2_X1    g02643(.A1(new_n5063_), .A2(new_n3259_), .ZN(new_n5093_));
  OAI21_X1   g02644(.A1(new_n5092_), .A2(pi0100), .B(new_n5093_), .ZN(new_n5094_));
  NOR2_X1    g02645(.A1(new_n5030_), .A2(new_n5010_), .ZN(new_n5095_));
  NOR2_X1    g02646(.A1(new_n5095_), .A2(new_n5065_), .ZN(new_n5096_));
  NAND2_X1   g02647(.A1(new_n5095_), .A2(new_n5065_), .ZN(new_n5097_));
  NAND2_X1   g02648(.A1(new_n5097_), .A2(new_n3121_), .ZN(new_n5098_));
  OAI21_X1   g02649(.A1(new_n5098_), .A2(new_n5096_), .B(new_n4975_), .ZN(new_n5099_));
  NAND2_X1   g02650(.A1(new_n5099_), .A2(pi0299), .ZN(new_n5100_));
  XOR2_X1    g02651(.A1(new_n5100_), .A2(new_n3695_), .Z(new_n5101_));
  NOR2_X1    g02652(.A1(new_n5101_), .A2(new_n4959_), .ZN(new_n5102_));
  NAND2_X1   g02653(.A1(new_n5064_), .A2(new_n3211_), .ZN(new_n5103_));
  AOI21_X1   g02654(.A1(new_n5062_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n5104_));
  OAI21_X1   g02655(.A1(new_n5102_), .A2(new_n5103_), .B(new_n5104_), .ZN(new_n5105_));
  NAND4_X1   g02656(.A1(new_n5094_), .A2(pi0075), .A3(pi0087), .A4(new_n5105_), .ZN(new_n5106_));
  NAND2_X1   g02657(.A1(new_n5094_), .A2(new_n5105_), .ZN(new_n5107_));
  NAND3_X1   g02658(.A1(new_n5107_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n5108_));
  AOI21_X1   g02659(.A1(new_n5108_), .A2(new_n5106_), .B(new_n5075_), .ZN(new_n5109_));
  NOR2_X1    g02660(.A1(new_n5109_), .A2(pi0092), .ZN(new_n5110_));
  NOR3_X1    g02661(.A1(new_n5110_), .A2(new_n3235_), .A3(new_n5063_), .ZN(new_n5111_));
  NAND2_X1   g02662(.A1(new_n5075_), .A2(pi0092), .ZN(new_n5112_));
  XNOR2_X1   g02663(.A1(new_n5112_), .A2(new_n3172_), .ZN(new_n5113_));
  INV_X1     g02664(.I(new_n4999_), .ZN(new_n5114_));
  NOR2_X1    g02665(.A1(new_n5072_), .A2(new_n3201_), .ZN(new_n5115_));
  XOR2_X1    g02666(.A1(new_n5115_), .A2(new_n3972_), .Z(new_n5116_));
  AOI21_X1   g02667(.A1(new_n5116_), .A2(new_n5114_), .B(new_n3426_), .ZN(new_n5117_));
  NOR2_X1    g02668(.A1(new_n5072_), .A2(new_n3219_), .ZN(new_n5118_));
  XOR2_X1    g02669(.A1(new_n5118_), .A2(new_n3797_), .Z(new_n5119_));
  OAI21_X1   g02670(.A1(new_n5119_), .A2(new_n4999_), .B(new_n3201_), .ZN(new_n5120_));
  NOR2_X1    g02671(.A1(new_n5117_), .A2(new_n5120_), .ZN(new_n5121_));
  NOR2_X1    g02672(.A1(new_n5072_), .A2(new_n3258_), .ZN(new_n5122_));
  XOR2_X1    g02673(.A1(new_n5122_), .A2(new_n3605_), .Z(new_n5123_));
  OAI21_X1   g02674(.A1(new_n5123_), .A2(new_n4999_), .B(new_n3219_), .ZN(new_n5124_));
  NAND2_X1   g02675(.A1(new_n5000_), .A2(new_n3426_), .ZN(new_n5125_));
  NAND4_X1   g02676(.A1(new_n5125_), .A2(new_n3258_), .A3(pi0244), .A4(new_n3202_), .ZN(new_n5126_));
  AOI21_X1   g02677(.A1(new_n3203_), .A2(new_n5062_), .B(new_n5126_), .ZN(new_n5127_));
  NAND2_X1   g02678(.A1(new_n5124_), .A2(new_n5127_), .ZN(new_n5128_));
  NOR2_X1    g02679(.A1(new_n5121_), .A2(new_n5128_), .ZN(new_n5129_));
  OAI21_X1   g02680(.A1(new_n5063_), .A2(new_n5113_), .B(new_n5129_), .ZN(new_n5130_));
  OAI22_X1   g02681(.A1(new_n5055_), .A2(new_n5059_), .B1(new_n5111_), .B2(new_n5130_), .ZN(po0164));
  INV_X1     g02682(.I(pi1134), .ZN(new_n5132_));
  AOI21_X1   g02683(.A1(pi0224), .A2(pi0278), .B(pi0222), .ZN(new_n5133_));
  INV_X1     g02684(.I(new_n5133_), .ZN(new_n5134_));
  INV_X1     g02685(.I(pi0846), .ZN(new_n5135_));
  NOR2_X1    g02686(.A1(new_n2753_), .A2(new_n5135_), .ZN(new_n5136_));
  AOI21_X1   g02687(.A1(new_n5136_), .A2(new_n3100_), .B(new_n5134_), .ZN(new_n5137_));
  NOR2_X1    g02688(.A1(new_n3099_), .A2(pi0224), .ZN(new_n5138_));
  INV_X1     g02689(.I(new_n5138_), .ZN(new_n5139_));
  NOR3_X1    g02690(.A1(new_n5139_), .A2(new_n3058_), .A3(pi0930), .ZN(new_n5140_));
  INV_X1     g02691(.I(new_n5137_), .ZN(new_n5141_));
  NOR2_X1    g02692(.A1(new_n3109_), .A2(pi0299), .ZN(new_n5142_));
  NAND2_X1   g02693(.A1(new_n5142_), .A2(new_n5141_), .ZN(new_n5143_));
  AND2_X2    g02694(.A1(new_n5143_), .A2(new_n5140_), .Z(new_n5144_));
  INV_X1     g02695(.I(new_n5144_), .ZN(new_n5145_));
  NOR2_X1    g02696(.A1(new_n5145_), .A2(new_n3660_), .ZN(new_n5146_));
  AOI21_X1   g02697(.A1(new_n5146_), .A2(new_n3109_), .B(pi0299), .ZN(new_n5147_));
  INV_X1     g02698(.I(new_n5147_), .ZN(new_n5148_));
  AOI21_X1   g02699(.A1(new_n3090_), .A2(new_n5137_), .B(new_n5148_), .ZN(new_n5149_));
  INV_X1     g02700(.I(pi0930), .ZN(new_n5150_));
  NOR4_X1    g02701(.A1(new_n3011_), .A2(new_n3121_), .A3(new_n3058_), .A4(new_n5150_), .ZN(new_n5151_));
  INV_X1     g02702(.I(new_n5151_), .ZN(new_n5152_));
  INV_X1     g02703(.I(new_n5136_), .ZN(new_n5153_));
  AOI21_X1   g02704(.A1(new_n5153_), .A2(pi0228), .B(new_n3009_), .ZN(new_n5154_));
  NOR3_X1    g02705(.A1(new_n5136_), .A2(pi0105), .A3(new_n3005_), .ZN(new_n5155_));
  OAI21_X1   g02706(.A1(new_n5154_), .A2(new_n5155_), .B(pi0152), .ZN(new_n5156_));
  INV_X1     g02707(.I(new_n5156_), .ZN(new_n5157_));
  INV_X1     g02708(.I(pi0152), .ZN(new_n5158_));
  NAND3_X1   g02709(.A1(new_n3160_), .A2(pi0228), .A3(pi0846), .ZN(new_n5159_));
  NAND3_X1   g02710(.A1(new_n3160_), .A2(new_n3005_), .A3(new_n5135_), .ZN(new_n5160_));
  AOI21_X1   g02711(.A1(new_n5159_), .A2(new_n5160_), .B(new_n5158_), .ZN(new_n5161_));
  AOI21_X1   g02712(.A1(pi0216), .A2(pi0278), .B(pi0221), .ZN(new_n5162_));
  INV_X1     g02713(.I(new_n5162_), .ZN(new_n5163_));
  NOR2_X1    g02714(.A1(new_n5163_), .A2(new_n3011_), .ZN(new_n5164_));
  OAI21_X1   g02715(.A1(new_n5161_), .A2(new_n5164_), .B(new_n5157_), .ZN(new_n5165_));
  AOI21_X1   g02716(.A1(new_n5165_), .A2(new_n5152_), .B(pi0215), .ZN(new_n5166_));
  NOR2_X1    g02717(.A1(new_n5166_), .A2(new_n3098_), .ZN(new_n5167_));
  NOR2_X1    g02718(.A1(new_n5149_), .A2(new_n5167_), .ZN(new_n5168_));
  INV_X1     g02719(.I(new_n5168_), .ZN(new_n5169_));
  NOR2_X1    g02720(.A1(new_n5158_), .A2(pi0228), .ZN(new_n5170_));
  OAI21_X1   g02721(.A1(new_n5157_), .A2(new_n5170_), .B(new_n3011_), .ZN(new_n5171_));
  NAND2_X1   g02722(.A1(new_n5171_), .A2(new_n5162_), .ZN(new_n5172_));
  AOI21_X1   g02723(.A1(new_n5172_), .A2(new_n5152_), .B(pi0215), .ZN(new_n5173_));
  INV_X1     g02724(.I(new_n5173_), .ZN(new_n5174_));
  AOI21_X1   g02725(.A1(pi0299), .A2(new_n5174_), .B(new_n5149_), .ZN(new_n5175_));
  NOR2_X1    g02726(.A1(new_n5175_), .A2(new_n3134_), .ZN(new_n5176_));
  AOI21_X1   g02727(.A1(new_n5169_), .A2(new_n3134_), .B(new_n5176_), .ZN(new_n5177_));
  NAND3_X1   g02728(.A1(new_n3330_), .A2(pi0152), .A3(pi0846), .ZN(new_n5178_));
  NAND3_X1   g02729(.A1(new_n3862_), .A2(new_n5158_), .A3(pi0846), .ZN(new_n5179_));
  NOR2_X1    g02730(.A1(new_n3004_), .A2(new_n5158_), .ZN(new_n5180_));
  OAI21_X1   g02731(.A1(new_n3306_), .A2(pi0228), .B(new_n5180_), .ZN(new_n5181_));
  AOI21_X1   g02732(.A1(new_n3306_), .A2(new_n5135_), .B(new_n3005_), .ZN(new_n5182_));
  XOR2_X1    g02733(.A1(new_n5182_), .A2(new_n3009_), .Z(new_n5183_));
  OAI21_X1   g02734(.A1(new_n5183_), .A2(new_n5158_), .B(new_n3011_), .ZN(new_n5184_));
  NAND2_X1   g02735(.A1(new_n5184_), .A2(new_n5181_), .ZN(new_n5185_));
  NAND3_X1   g02736(.A1(new_n5158_), .A2(new_n3005_), .A3(new_n5135_), .ZN(new_n5186_));
  NAND4_X1   g02737(.A1(new_n3696_), .A2(new_n3307_), .A3(new_n5185_), .A4(new_n5186_), .ZN(new_n5187_));
  AOI21_X1   g02738(.A1(new_n5179_), .A2(new_n5178_), .B(new_n5187_), .ZN(new_n5188_));
  OAI21_X1   g02739(.A1(new_n5188_), .A2(new_n5163_), .B(new_n5152_), .ZN(new_n5189_));
  NOR2_X1    g02740(.A1(new_n3098_), .A2(pi0215), .ZN(new_n5190_));
  NAND2_X1   g02741(.A1(new_n5169_), .A2(pi0039), .ZN(new_n5191_));
  AOI21_X1   g02742(.A1(new_n5140_), .A2(new_n5133_), .B(pi0224), .ZN(new_n5192_));
  NOR3_X1    g02743(.A1(new_n3702_), .A2(pi0846), .A3(new_n5192_), .ZN(new_n5193_));
  NOR2_X1    g02744(.A1(new_n5193_), .A2(new_n3382_), .ZN(new_n5194_));
  NAND3_X1   g02745(.A1(new_n5153_), .A2(new_n3100_), .A3(new_n5134_), .ZN(new_n5195_));
  NAND2_X1   g02746(.A1(new_n3305_), .A2(new_n5195_), .ZN(new_n5196_));
  NOR2_X1    g02747(.A1(new_n5196_), .A2(new_n3382_), .ZN(new_n5197_));
  NOR4_X1    g02748(.A1(new_n5194_), .A2(pi0038), .A3(pi0039), .A4(new_n5197_), .ZN(new_n5198_));
  AOI21_X1   g02749(.A1(new_n5198_), .A2(new_n5191_), .B(new_n5190_), .ZN(new_n5199_));
  OAI21_X1   g02750(.A1(new_n5189_), .A2(new_n5199_), .B(new_n3462_), .ZN(new_n5200_));
  NAND3_X1   g02751(.A1(new_n5200_), .A2(pi0038), .A3(new_n5175_), .ZN(new_n5201_));
  AOI21_X1   g02752(.A1(new_n3391_), .A2(pi0846), .B(pi0228), .ZN(new_n5202_));
  INV_X1     g02753(.I(new_n5202_), .ZN(new_n5203_));
  AOI21_X1   g02754(.A1(new_n3399_), .A2(pi0152), .B(new_n5203_), .ZN(new_n5204_));
  OAI21_X1   g02755(.A1(new_n5204_), .A2(new_n5164_), .B(new_n5157_), .ZN(new_n5205_));
  AOI21_X1   g02756(.A1(new_n5205_), .A2(new_n3855_), .B(new_n5152_), .ZN(new_n5206_));
  OR2_X2     g02757(.A1(new_n5149_), .A2(new_n3212_), .Z(new_n5207_));
  AOI21_X1   g02758(.A1(new_n5175_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n5208_));
  OAI21_X1   g02759(.A1(new_n5206_), .A2(new_n5207_), .B(new_n5208_), .ZN(new_n5209_));
  NAND4_X1   g02760(.A1(new_n5201_), .A2(pi0075), .A3(pi0087), .A4(new_n5209_), .ZN(new_n5210_));
  NAND2_X1   g02761(.A1(new_n5201_), .A2(new_n5209_), .ZN(new_n5211_));
  NAND3_X1   g02762(.A1(new_n5211_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n5212_));
  AOI21_X1   g02763(.A1(new_n5212_), .A2(new_n5210_), .B(new_n5177_), .ZN(new_n5213_));
  AND2_X2    g02764(.A1(new_n5175_), .A2(pi0075), .Z(new_n5214_));
  OAI21_X1   g02765(.A1(new_n5213_), .A2(pi0092), .B(new_n5214_), .ZN(new_n5215_));
  NAND2_X1   g02766(.A1(new_n5177_), .A2(pi0092), .ZN(new_n5216_));
  XOR2_X1    g02767(.A1(new_n5216_), .A2(new_n3172_), .Z(new_n5217_));
  NOR2_X1    g02768(.A1(new_n5166_), .A2(new_n3258_), .ZN(new_n5218_));
  XOR2_X1    g02769(.A1(new_n5218_), .A2(new_n3605_), .Z(new_n5219_));
  OAI21_X1   g02770(.A1(new_n5219_), .A2(new_n5174_), .B(new_n3219_), .ZN(new_n5220_));
  NOR2_X1    g02771(.A1(new_n3203_), .A2(pi0055), .ZN(new_n5221_));
  NAND2_X1   g02772(.A1(new_n5220_), .A2(new_n5221_), .ZN(new_n5222_));
  AOI21_X1   g02773(.A1(new_n5217_), .A2(new_n5175_), .B(new_n5222_), .ZN(new_n5223_));
  NOR2_X1    g02774(.A1(new_n5166_), .A2(new_n3219_), .ZN(new_n5224_));
  XOR2_X1    g02775(.A1(new_n5224_), .A2(new_n3797_), .Z(new_n5225_));
  OAI21_X1   g02776(.A1(new_n5225_), .A2(new_n5174_), .B(new_n3201_), .ZN(new_n5226_));
  AOI21_X1   g02777(.A1(new_n5215_), .A2(new_n5223_), .B(new_n5226_), .ZN(new_n5227_));
  OAI21_X1   g02778(.A1(new_n5173_), .A2(pi0242), .B(new_n3426_), .ZN(new_n5228_));
  NOR2_X1    g02779(.A1(new_n5166_), .A2(new_n3201_), .ZN(new_n5229_));
  XOR2_X1    g02780(.A1(new_n5229_), .A2(new_n3594_), .Z(new_n5230_));
  NOR2_X1    g02781(.A1(new_n5230_), .A2(new_n5174_), .ZN(new_n5231_));
  OAI21_X1   g02782(.A1(new_n5227_), .A2(new_n5228_), .B(new_n5231_), .ZN(new_n5232_));
  NOR2_X1    g02783(.A1(new_n5174_), .A2(new_n3913_), .ZN(new_n5233_));
  OAI21_X1   g02784(.A1(new_n5233_), .A2(new_n3098_), .B(new_n5148_), .ZN(new_n5234_));
  AOI21_X1   g02785(.A1(new_n5156_), .A2(new_n3370_), .B(new_n5164_), .ZN(new_n5235_));
  INV_X1     g02786(.I(new_n5235_), .ZN(new_n5236_));
  NAND2_X1   g02787(.A1(new_n5161_), .A2(new_n5236_), .ZN(new_n5237_));
  NAND2_X1   g02788(.A1(new_n5237_), .A2(new_n5152_), .ZN(new_n5238_));
  NAND2_X1   g02789(.A1(new_n5238_), .A2(new_n3111_), .ZN(new_n5239_));
  AOI21_X1   g02790(.A1(new_n5239_), .A2(pi0299), .B(new_n5147_), .ZN(new_n5240_));
  NAND2_X1   g02791(.A1(new_n5234_), .A2(new_n3474_), .ZN(new_n5241_));
  OAI21_X1   g02792(.A1(new_n5240_), .A2(new_n3474_), .B(new_n5241_), .ZN(new_n5242_));
  INV_X1     g02793(.I(new_n5234_), .ZN(new_n5243_));
  NAND2_X1   g02794(.A1(new_n5158_), .A2(new_n5135_), .ZN(new_n5244_));
  OAI21_X1   g02795(.A1(new_n5184_), .A2(new_n5163_), .B(new_n3005_), .ZN(new_n5245_));
  NAND3_X1   g02796(.A1(new_n3696_), .A2(new_n5244_), .A3(new_n5245_), .ZN(new_n5246_));
  NAND2_X1   g02797(.A1(new_n5246_), .A2(new_n5152_), .ZN(new_n5247_));
  NOR3_X1    g02798(.A1(new_n5194_), .A2(pi0038), .A3(pi0039), .ZN(new_n5248_));
  NOR2_X1    g02799(.A1(new_n5248_), .A2(new_n5190_), .ZN(new_n5249_));
  OAI21_X1   g02800(.A1(new_n5247_), .A2(new_n5249_), .B(new_n3462_), .ZN(new_n5250_));
  AND3_X2    g02801(.A1(new_n5250_), .A2(pi0038), .A3(new_n5243_), .Z(new_n5251_));
  NAND2_X1   g02802(.A1(new_n5204_), .A2(new_n5236_), .ZN(new_n5252_));
  NAND2_X1   g02803(.A1(new_n5252_), .A2(new_n3855_), .ZN(new_n5253_));
  NAND2_X1   g02804(.A1(new_n5253_), .A2(new_n5151_), .ZN(new_n5254_));
  NOR2_X1    g02805(.A1(new_n5147_), .A2(new_n3212_), .ZN(new_n5255_));
  OAI21_X1   g02806(.A1(new_n5234_), .A2(new_n3211_), .B(pi0100), .ZN(new_n5256_));
  AOI21_X1   g02807(.A1(new_n5254_), .A2(new_n5255_), .B(new_n5256_), .ZN(new_n5257_));
  OAI21_X1   g02808(.A1(new_n5251_), .A2(new_n5257_), .B(pi0087), .ZN(new_n5258_));
  XOR2_X1    g02809(.A1(new_n5258_), .A2(new_n3953_), .Z(new_n5259_));
  AOI21_X1   g02810(.A1(new_n5259_), .A2(new_n5242_), .B(pi0092), .ZN(new_n5260_));
  NOR3_X1    g02811(.A1(new_n5260_), .A2(new_n3235_), .A3(new_n5234_), .ZN(new_n5261_));
  NOR2_X1    g02812(.A1(new_n5242_), .A2(new_n3303_), .ZN(new_n5262_));
  XOR2_X1    g02813(.A1(new_n5262_), .A2(new_n3172_), .Z(new_n5263_));
  NAND2_X1   g02814(.A1(new_n5239_), .A2(pi0055), .ZN(new_n5264_));
  XOR2_X1    g02815(.A1(new_n5264_), .A2(new_n3605_), .Z(new_n5265_));
  NAND2_X1   g02816(.A1(new_n5265_), .A2(new_n5233_), .ZN(new_n5266_));
  NAND2_X1   g02817(.A1(new_n3202_), .A2(new_n3258_), .ZN(new_n5267_));
  AOI21_X1   g02818(.A1(new_n5266_), .A2(new_n3219_), .B(new_n5267_), .ZN(new_n5268_));
  OAI21_X1   g02819(.A1(new_n5263_), .A2(new_n5234_), .B(new_n5268_), .ZN(new_n5269_));
  NAND2_X1   g02820(.A1(new_n5239_), .A2(pi0056), .ZN(new_n5270_));
  XOR2_X1    g02821(.A1(new_n5270_), .A2(new_n3797_), .Z(new_n5271_));
  AOI21_X1   g02822(.A1(new_n5271_), .A2(new_n5233_), .B(pi0062), .ZN(new_n5272_));
  OAI21_X1   g02823(.A1(new_n5261_), .A2(new_n5269_), .B(new_n5272_), .ZN(new_n5273_));
  NAND2_X1   g02824(.A1(new_n5239_), .A2(pi0062), .ZN(new_n5274_));
  XOR2_X1    g02825(.A1(new_n5274_), .A2(new_n3594_), .Z(new_n5275_));
  NAND2_X1   g02826(.A1(new_n3230_), .A2(pi0242), .ZN(new_n5276_));
  AOI21_X1   g02827(.A1(new_n5275_), .A2(new_n5233_), .B(new_n5276_), .ZN(new_n5277_));
  NAND2_X1   g02828(.A1(new_n5273_), .A2(new_n5277_), .ZN(new_n5278_));
  AOI21_X1   g02829(.A1(new_n5232_), .A2(new_n5132_), .B(new_n5278_), .ZN(new_n5279_));
  AOI21_X1   g02830(.A1(new_n3355_), .A2(pi0221), .B(pi0215), .ZN(new_n5280_));
  INV_X1     g02831(.I(new_n5280_), .ZN(new_n5281_));
  NOR2_X1    g02832(.A1(new_n5281_), .A2(new_n5151_), .ZN(new_n5282_));
  NAND2_X1   g02833(.A1(new_n5172_), .A2(new_n5282_), .ZN(new_n5283_));
  INV_X1     g02834(.I(new_n5283_), .ZN(new_n5284_));
  NOR2_X1    g02835(.A1(new_n5284_), .A2(new_n3913_), .ZN(new_n5285_));
  AOI21_X1   g02836(.A1(new_n5285_), .A2(pi0299), .B(new_n5146_), .ZN(new_n5286_));
  INV_X1     g02837(.I(new_n5146_), .ZN(new_n5287_));
  NAND2_X1   g02838(.A1(new_n5237_), .A2(new_n5282_), .ZN(new_n5288_));
  NAND2_X1   g02839(.A1(new_n5288_), .A2(pi0299), .ZN(new_n5289_));
  NAND2_X1   g02840(.A1(new_n5289_), .A2(new_n5287_), .ZN(new_n5290_));
  NOR2_X1    g02841(.A1(new_n5286_), .A2(new_n3134_), .ZN(new_n5291_));
  AOI21_X1   g02842(.A1(new_n5290_), .A2(new_n3134_), .B(new_n5291_), .ZN(new_n5292_));
  INV_X1     g02843(.I(new_n5190_), .ZN(new_n5293_));
  AOI21_X1   g02844(.A1(pi0221), .A2(new_n3355_), .B(new_n5293_), .ZN(new_n5294_));
  NAND2_X1   g02845(.A1(new_n5290_), .A2(pi0039), .ZN(new_n5295_));
  NOR2_X1    g02846(.A1(new_n3108_), .A2(new_n3382_), .ZN(new_n5296_));
  AOI21_X1   g02847(.A1(new_n5193_), .A2(new_n5296_), .B(new_n3212_), .ZN(new_n5297_));
  AOI21_X1   g02848(.A1(new_n5297_), .A2(new_n5295_), .B(new_n5294_), .ZN(new_n5298_));
  OAI21_X1   g02849(.A1(new_n5247_), .A2(new_n5298_), .B(new_n3462_), .ZN(new_n5299_));
  NAND3_X1   g02850(.A1(new_n5299_), .A2(pi0038), .A3(new_n5286_), .ZN(new_n5300_));
  AOI21_X1   g02851(.A1(new_n5252_), .A2(new_n5282_), .B(new_n3098_), .ZN(new_n5301_));
  NAND2_X1   g02852(.A1(new_n5287_), .A2(new_n3211_), .ZN(new_n5302_));
  AOI21_X1   g02853(.A1(new_n5286_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n5303_));
  OAI21_X1   g02854(.A1(new_n5301_), .A2(new_n5302_), .B(new_n5303_), .ZN(new_n5304_));
  AOI21_X1   g02855(.A1(new_n5300_), .A2(new_n5304_), .B(new_n3455_), .ZN(new_n5305_));
  XOR2_X1    g02856(.A1(new_n5305_), .A2(new_n3953_), .Z(new_n5306_));
  OAI21_X1   g02857(.A1(new_n5306_), .A2(new_n5292_), .B(new_n3303_), .ZN(new_n5307_));
  NAND3_X1   g02858(.A1(new_n5307_), .A2(pi0075), .A3(new_n5286_), .ZN(new_n5308_));
  INV_X1     g02859(.I(new_n5286_), .ZN(new_n5309_));
  AOI21_X1   g02860(.A1(new_n5309_), .A2(new_n3258_), .B(new_n3202_), .ZN(new_n5310_));
  NAND2_X1   g02861(.A1(new_n5308_), .A2(new_n5310_), .ZN(new_n5311_));
  NAND2_X1   g02862(.A1(new_n5292_), .A2(pi0092), .ZN(new_n5312_));
  XNOR2_X1   g02863(.A1(new_n5312_), .A2(new_n3172_), .ZN(new_n5313_));
  INV_X1     g02864(.I(new_n5285_), .ZN(new_n5314_));
  NAND2_X1   g02865(.A1(new_n5288_), .A2(pi0056), .ZN(new_n5315_));
  XOR2_X1    g02866(.A1(new_n5315_), .A2(new_n3599_), .Z(new_n5316_));
  OAI21_X1   g02867(.A1(new_n5316_), .A2(new_n5314_), .B(new_n3201_), .ZN(new_n5317_));
  NAND2_X1   g02868(.A1(new_n5288_), .A2(pi0055), .ZN(new_n5318_));
  XOR2_X1    g02869(.A1(new_n5318_), .A2(new_n3605_), .Z(new_n5319_));
  NAND2_X1   g02870(.A1(new_n5319_), .A2(new_n5285_), .ZN(new_n5320_));
  NAND4_X1   g02871(.A1(new_n5317_), .A2(new_n5320_), .A3(new_n3219_), .A4(new_n5286_), .ZN(new_n5321_));
  NOR2_X1    g02872(.A1(new_n5313_), .A2(new_n5321_), .ZN(new_n5322_));
  NAND2_X1   g02873(.A1(new_n5288_), .A2(pi0062), .ZN(new_n5323_));
  XNOR2_X1   g02874(.A1(new_n5323_), .A2(new_n3594_), .ZN(new_n5324_));
  NOR2_X1    g02875(.A1(new_n3426_), .A2(pi0242), .ZN(new_n5325_));
  OAI21_X1   g02876(.A1(new_n5324_), .A2(new_n5314_), .B(new_n5325_), .ZN(new_n5326_));
  AOI21_X1   g02877(.A1(new_n5311_), .A2(new_n5322_), .B(new_n5326_), .ZN(new_n5327_));
  NAND2_X1   g02878(.A1(new_n5165_), .A2(new_n5282_), .ZN(new_n5328_));
  AOI21_X1   g02879(.A1(new_n5328_), .A2(pi0299), .B(new_n5144_), .ZN(new_n5329_));
  INV_X1     g02880(.I(new_n5329_), .ZN(new_n5330_));
  AOI21_X1   g02881(.A1(new_n5283_), .A2(pi0299), .B(new_n5144_), .ZN(new_n5331_));
  NOR2_X1    g02882(.A1(new_n5331_), .A2(new_n3134_), .ZN(new_n5332_));
  AOI21_X1   g02883(.A1(new_n5330_), .A2(new_n3134_), .B(new_n5332_), .ZN(new_n5333_));
  NAND2_X1   g02884(.A1(new_n5330_), .A2(pi0039), .ZN(new_n5334_));
  NOR2_X1    g02885(.A1(new_n5296_), .A2(pi0039), .ZN(new_n5335_));
  NAND2_X1   g02886(.A1(new_n5140_), .A2(new_n3259_), .ZN(new_n5336_));
  AOI21_X1   g02887(.A1(new_n5196_), .A2(new_n5335_), .B(new_n5336_), .ZN(new_n5337_));
  AOI21_X1   g02888(.A1(new_n5337_), .A2(new_n5334_), .B(new_n5294_), .ZN(new_n5338_));
  OAI21_X1   g02889(.A1(new_n5189_), .A2(new_n5338_), .B(new_n3462_), .ZN(new_n5339_));
  NAND3_X1   g02890(.A1(new_n5339_), .A2(pi0038), .A3(new_n5331_), .ZN(new_n5340_));
  AOI21_X1   g02891(.A1(new_n5205_), .A2(new_n5282_), .B(new_n3098_), .ZN(new_n5341_));
  NAND2_X1   g02892(.A1(new_n5145_), .A2(new_n3211_), .ZN(new_n5342_));
  AOI21_X1   g02893(.A1(new_n5331_), .A2(new_n3212_), .B(new_n3462_), .ZN(new_n5343_));
  OAI21_X1   g02894(.A1(new_n5341_), .A2(new_n5342_), .B(new_n5343_), .ZN(new_n5344_));
  NAND4_X1   g02895(.A1(new_n5340_), .A2(pi0075), .A3(pi0087), .A4(new_n5344_), .ZN(new_n5345_));
  NAND2_X1   g02896(.A1(new_n5340_), .A2(new_n5344_), .ZN(new_n5346_));
  NAND3_X1   g02897(.A1(new_n5346_), .A2(pi0087), .A3(new_n3953_), .ZN(new_n5347_));
  AOI21_X1   g02898(.A1(new_n5347_), .A2(new_n5345_), .B(new_n5333_), .ZN(new_n5348_));
  AND2_X2    g02899(.A1(new_n5331_), .A2(pi0075), .Z(new_n5349_));
  OAI21_X1   g02900(.A1(new_n5348_), .A2(pi0092), .B(new_n5349_), .ZN(new_n5350_));
  NAND2_X1   g02901(.A1(new_n5333_), .A2(pi0092), .ZN(new_n5351_));
  XOR2_X1    g02902(.A1(new_n5351_), .A2(new_n3172_), .Z(new_n5352_));
  NAND2_X1   g02903(.A1(new_n5352_), .A2(new_n5331_), .ZN(new_n5353_));
  NAND2_X1   g02904(.A1(new_n5328_), .A2(pi0055), .ZN(new_n5354_));
  XOR2_X1    g02905(.A1(new_n5354_), .A2(new_n3604_), .Z(new_n5355_));
  OAI21_X1   g02906(.A1(new_n5355_), .A2(new_n5283_), .B(new_n3219_), .ZN(new_n5356_));
  NOR2_X1    g02907(.A1(new_n3203_), .A2(pi0055), .ZN(new_n5357_));
  NAND4_X1   g02908(.A1(new_n5350_), .A2(new_n5353_), .A3(new_n5356_), .A4(new_n5357_), .ZN(new_n5358_));
  NAND2_X1   g02909(.A1(new_n5328_), .A2(pi0056), .ZN(new_n5359_));
  XOR2_X1    g02910(.A1(new_n5359_), .A2(new_n3797_), .Z(new_n5360_));
  AOI21_X1   g02911(.A1(new_n5360_), .A2(new_n5284_), .B(pi0062), .ZN(new_n5361_));
  NAND2_X1   g02912(.A1(new_n5328_), .A2(pi0062), .ZN(new_n5362_));
  XNOR2_X1   g02913(.A1(new_n5362_), .A2(new_n3594_), .ZN(new_n5363_));
  INV_X1     g02914(.I(pi0242), .ZN(new_n5364_));
  NOR2_X1    g02915(.A1(new_n3426_), .A2(new_n5364_), .ZN(new_n5365_));
  OAI21_X1   g02916(.A1(new_n5363_), .A2(new_n5283_), .B(new_n5365_), .ZN(new_n5366_));
  AOI21_X1   g02917(.A1(new_n5358_), .A2(new_n5361_), .B(new_n5366_), .ZN(new_n5367_));
  NOR3_X1    g02918(.A1(new_n5367_), .A2(pi1134), .A3(new_n5327_), .ZN(new_n5368_));
  NOR2_X1    g02919(.A1(new_n5368_), .A2(new_n5279_), .ZN(po0165));
  INV_X1     g02920(.I(pi0057), .ZN(new_n5371_));
  NAND2_X1   g02921(.A1(new_n3145_), .A2(new_n3565_), .ZN(new_n5372_));
  NOR2_X1    g02922(.A1(pi0332), .A2(pi0468), .ZN(new_n5373_));
  INV_X1     g02923(.I(pi0661), .ZN(new_n5374_));
  INV_X1     g02924(.I(pi0680), .ZN(new_n5375_));
  NOR2_X1    g02925(.A1(new_n5375_), .A2(pi0662), .ZN(new_n5376_));
  NAND2_X1   g02926(.A1(new_n5376_), .A2(new_n5374_), .ZN(new_n5377_));
  NOR2_X1    g02927(.A1(new_n5377_), .A2(pi0681), .ZN(new_n5378_));
  INV_X1     g02928(.I(pi0642), .ZN(new_n5379_));
  NAND2_X1   g02929(.A1(new_n5379_), .A2(pi0603), .ZN(new_n5380_));
  NOR2_X1    g02930(.A1(pi0614), .A2(pi0616), .ZN(new_n5381_));
  INV_X1     g02931(.I(new_n5381_), .ZN(new_n5382_));
  NOR2_X1    g02932(.A1(new_n5382_), .A2(new_n5380_), .ZN(new_n5383_));
  NOR2_X1    g02933(.A1(new_n5378_), .A2(new_n5383_), .ZN(new_n5384_));
  NOR2_X1    g02934(.A1(new_n5384_), .A2(new_n5373_), .ZN(new_n5385_));
  INV_X1     g02935(.I(new_n5373_), .ZN(new_n5386_));
  INV_X1     g02936(.I(pi0969), .ZN(new_n5387_));
  INV_X1     g02937(.I(pi0971), .ZN(new_n5388_));
  INV_X1     g02938(.I(pi0974), .ZN(new_n5389_));
  INV_X1     g02939(.I(pi0977), .ZN(new_n5390_));
  NOR4_X1    g02940(.A1(new_n5387_), .A2(new_n5388_), .A3(new_n5389_), .A4(new_n5390_), .ZN(new_n5391_));
  INV_X1     g02941(.I(pi0587), .ZN(new_n5392_));
  INV_X1     g02942(.I(pi0602), .ZN(new_n5393_));
  INV_X1     g02943(.I(pi0961), .ZN(new_n5394_));
  INV_X1     g02944(.I(pi0967), .ZN(new_n5395_));
  NOR4_X1    g02945(.A1(new_n5392_), .A2(new_n5393_), .A3(new_n5394_), .A4(new_n5395_), .ZN(new_n5396_));
  NAND2_X1   g02946(.A1(new_n5391_), .A2(new_n5396_), .ZN(new_n5397_));
  INV_X1     g02947(.I(new_n5397_), .ZN(new_n5398_));
  NOR2_X1    g02948(.A1(new_n5398_), .A2(new_n5386_), .ZN(new_n5399_));
  NOR2_X1    g02949(.A1(new_n5385_), .A2(new_n5399_), .ZN(new_n5400_));
  INV_X1     g02950(.I(pi0287), .ZN(new_n5401_));
  INV_X1     g02951(.I(pi0835), .ZN(new_n5402_));
  INV_X1     g02952(.I(pi0984), .ZN(new_n5403_));
  NOR2_X1    g02953(.A1(new_n5402_), .A2(new_n5403_), .ZN(new_n5404_));
  INV_X1     g02954(.I(pi0979), .ZN(new_n5405_));
  OAI21_X1   g02955(.A1(pi0252), .A2(pi1001), .B(new_n5405_), .ZN(new_n5406_));
  NOR2_X1    g02956(.A1(new_n5406_), .A2(new_n5404_), .ZN(new_n5407_));
  INV_X1     g02957(.I(new_n5407_), .ZN(new_n5408_));
  NOR4_X1    g02958(.A1(new_n5408_), .A2(new_n5401_), .A3(new_n5402_), .A4(new_n2722_), .ZN(new_n5409_));
  INV_X1     g02959(.I(new_n5409_), .ZN(new_n5410_));
  NOR2_X1    g02960(.A1(new_n5410_), .A2(new_n2745_), .ZN(new_n5411_));
  NAND4_X1   g02961(.A1(new_n5411_), .A2(new_n5372_), .A3(new_n3101_), .A4(new_n5400_), .ZN(new_n5412_));
  INV_X1     g02962(.I(new_n2666_), .ZN(new_n5413_));
  INV_X1     g02963(.I(new_n2877_), .ZN(new_n5414_));
  NOR2_X1    g02964(.A1(new_n2520_), .A2(new_n2897_), .ZN(new_n5415_));
  INV_X1     g02965(.I(new_n2876_), .ZN(new_n5416_));
  AOI21_X1   g02966(.A1(pi0108), .A2(new_n2524_), .B(new_n2550_), .ZN(new_n5417_));
  AOI21_X1   g02967(.A1(new_n2665_), .A2(new_n5416_), .B(new_n5417_), .ZN(new_n5418_));
  NAND4_X1   g02968(.A1(new_n2656_), .A2(new_n2526_), .A3(new_n5415_), .A4(new_n5418_), .ZN(new_n5419_));
  INV_X1     g02969(.I(new_n2468_), .ZN(new_n5420_));
  NOR2_X1    g02970(.A1(new_n5420_), .A2(new_n2673_), .ZN(new_n5421_));
  OAI21_X1   g02971(.A1(new_n2458_), .A2(new_n5421_), .B(new_n2672_), .ZN(new_n5422_));
  NOR2_X1    g02972(.A1(new_n2869_), .A2(pi0090), .ZN(new_n5423_));
  INV_X1     g02973(.I(new_n5423_), .ZN(new_n5424_));
  OAI21_X1   g02974(.A1(new_n5424_), .A2(new_n5422_), .B(new_n2673_), .ZN(new_n5425_));
  NAND4_X1   g02975(.A1(new_n5419_), .A2(new_n5413_), .A3(new_n5414_), .A4(new_n5425_), .ZN(new_n5426_));
  AOI21_X1   g02976(.A1(new_n2508_), .A2(new_n2732_), .B(new_n2509_), .ZN(new_n5427_));
  INV_X1     g02977(.I(new_n5427_), .ZN(new_n5428_));
  OAI21_X1   g02978(.A1(new_n2509_), .A2(new_n5428_), .B(new_n5426_), .ZN(new_n5429_));
  AOI21_X1   g02979(.A1(new_n5429_), .A2(new_n2680_), .B(new_n2692_), .ZN(new_n5430_));
  NAND2_X1   g02980(.A1(pi0035), .A2(pi0070), .ZN(new_n5431_));
  XOR2_X1    g02981(.A1(new_n5430_), .A2(new_n5431_), .Z(new_n5432_));
  INV_X1     g02982(.I(new_n5384_), .ZN(po1101));
  NOR2_X1    g02983(.A1(po1101), .A2(new_n5373_), .ZN(new_n5434_));
  AOI21_X1   g02984(.A1(new_n2726_), .A2(new_n2984_), .B(new_n2721_), .ZN(new_n5435_));
  AOI21_X1   g02985(.A1(pi0824), .A2(pi1091), .B(new_n5435_), .ZN(new_n5436_));
  INV_X1     g02986(.I(new_n5436_), .ZN(new_n5437_));
  NAND3_X1   g02987(.A1(new_n5409_), .A2(new_n5437_), .A3(pi1092), .ZN(new_n5438_));
  OAI21_X1   g02988(.A1(new_n5438_), .A2(new_n5434_), .B(new_n3160_), .ZN(new_n5439_));
  NOR2_X1    g02989(.A1(new_n3140_), .A2(new_n5386_), .ZN(new_n5440_));
  INV_X1     g02990(.I(new_n5440_), .ZN(new_n5441_));
  NAND2_X1   g02991(.A1(new_n5438_), .A2(new_n5386_), .ZN(new_n5442_));
  NAND4_X1   g02992(.A1(new_n5441_), .A2(new_n3145_), .A3(po1101), .A4(new_n5442_), .ZN(new_n5443_));
  NAND2_X1   g02993(.A1(new_n5443_), .A2(pi0215), .ZN(new_n5444_));
  NOR2_X1    g02994(.A1(pi0960), .A2(pi0963), .ZN(new_n5445_));
  INV_X1     g02995(.I(pi0970), .ZN(new_n5446_));
  INV_X1     g02996(.I(pi0972), .ZN(new_n5447_));
  INV_X1     g02997(.I(pi0975), .ZN(new_n5448_));
  INV_X1     g02998(.I(pi0978), .ZN(new_n5449_));
  NOR4_X1    g02999(.A1(new_n5446_), .A2(new_n5447_), .A3(new_n5448_), .A4(new_n5449_), .ZN(new_n5450_));
  NAND2_X1   g03000(.A1(new_n5450_), .A2(new_n5445_), .ZN(new_n5451_));
  NOR2_X1    g03001(.A1(pi0907), .A2(pi0947), .ZN(new_n5452_));
  INV_X1     g03002(.I(new_n5452_), .ZN(new_n5453_));
  NOR2_X1    g03003(.A1(new_n5451_), .A2(new_n5453_), .ZN(new_n5454_));
  INV_X1     g03004(.I(new_n5454_), .ZN(new_n5455_));
  NOR2_X1    g03005(.A1(new_n5455_), .A2(new_n3111_), .ZN(new_n5456_));
  XOR2_X1    g03006(.A1(new_n5444_), .A2(new_n5456_), .Z(new_n5457_));
  NOR2_X1    g03007(.A1(new_n5457_), .A2(new_n5439_), .ZN(new_n5458_));
  NAND2_X1   g03008(.A1(new_n3145_), .A2(new_n3855_), .ZN(new_n5459_));
  AOI21_X1   g03009(.A1(new_n5373_), .A2(new_n5454_), .B(new_n5434_), .ZN(new_n5460_));
  INV_X1     g03010(.I(new_n5460_), .ZN(new_n5461_));
  NAND4_X1   g03011(.A1(new_n5461_), .A2(new_n3373_), .A3(new_n5411_), .A4(new_n5459_), .ZN(new_n5462_));
  NOR2_X1    g03012(.A1(new_n2499_), .A2(pi0035), .ZN(new_n5463_));
  INV_X1     g03013(.I(new_n5463_), .ZN(new_n5464_));
  NOR3_X1    g03014(.A1(new_n2916_), .A2(pi0040), .A3(new_n5464_), .ZN(new_n5465_));
  INV_X1     g03015(.I(new_n5465_), .ZN(new_n5466_));
  NOR2_X1    g03016(.A1(new_n3072_), .A2(pi0299), .ZN(new_n5467_));
  AOI21_X1   g03017(.A1(pi0210), .A2(pi0299), .B(new_n5467_), .ZN(new_n5468_));
  INV_X1     g03018(.I(new_n5468_), .ZN(new_n5469_));
  NAND2_X1   g03019(.A1(new_n5469_), .A2(pi0032), .ZN(new_n5470_));
  XOR2_X1    g03020(.A1(new_n3325_), .A2(new_n5470_), .Z(new_n5471_));
  NOR2_X1    g03021(.A1(new_n5471_), .A2(new_n5466_), .ZN(new_n5472_));
  NAND2_X1   g03022(.A1(new_n5472_), .A2(new_n2503_), .ZN(new_n5473_));
  OAI21_X1   g03023(.A1(new_n2793_), .A2(new_n3183_), .B(new_n2436_), .ZN(new_n5474_));
  OAI21_X1   g03024(.A1(pi0072), .A2(pi0096), .B(new_n2702_), .ZN(new_n5475_));
  NAND4_X1   g03025(.A1(new_n5474_), .A2(pi0039), .A3(new_n5475_), .A4(new_n2696_), .ZN(new_n5476_));
  AOI21_X1   g03026(.A1(new_n5473_), .A2(new_n2485_), .B(new_n5476_), .ZN(new_n5477_));
  OAI21_X1   g03027(.A1(new_n5458_), .A2(new_n5462_), .B(new_n5477_), .ZN(new_n5478_));
  OAI21_X1   g03028(.A1(new_n5432_), .A2(new_n5478_), .B(new_n5412_), .ZN(new_n5479_));
  NAND2_X1   g03029(.A1(new_n5443_), .A2(pi0223), .ZN(new_n5480_));
  NOR2_X1    g03030(.A1(new_n5397_), .A2(new_n3090_), .ZN(new_n5481_));
  XOR2_X1    g03031(.A1(new_n5480_), .A2(new_n5481_), .Z(new_n5482_));
  NOR2_X1    g03032(.A1(new_n5482_), .A2(new_n5439_), .ZN(new_n5483_));
  AOI21_X1   g03033(.A1(new_n5479_), .A2(new_n5483_), .B(new_n3259_), .ZN(new_n5484_));
  NOR2_X1    g03034(.A1(new_n3259_), .A2(new_n3462_), .ZN(new_n5485_));
  INV_X1     g03035(.I(new_n5485_), .ZN(new_n5486_));
  XOR2_X1    g03036(.A1(new_n5484_), .A2(new_n5486_), .Z(new_n5487_));
  NOR2_X1    g03037(.A1(new_n3140_), .A2(new_n3474_), .ZN(new_n5488_));
  NAND2_X1   g03038(.A1(new_n3206_), .A2(new_n3175_), .ZN(new_n5489_));
  OAI21_X1   g03039(.A1(new_n5488_), .A2(new_n5489_), .B(pi0054), .ZN(new_n5490_));
  NAND2_X1   g03040(.A1(new_n5490_), .A2(new_n3258_), .ZN(new_n5491_));
  NOR2_X1    g03041(.A1(new_n3140_), .A2(pi0039), .ZN(new_n5492_));
  NAND3_X1   g03042(.A1(new_n5491_), .A2(pi0074), .A3(new_n5492_), .ZN(new_n5493_));
  INV_X1     g03043(.I(new_n5488_), .ZN(new_n5494_));
  NOR2_X1    g03044(.A1(new_n5494_), .A2(new_n3210_), .ZN(new_n5495_));
  OAI21_X1   g03045(.A1(new_n5495_), .A2(new_n3221_), .B(new_n3219_), .ZN(new_n5496_));
  INV_X1     g03046(.I(new_n5496_), .ZN(new_n5497_));
  AOI21_X1   g03047(.A1(new_n5494_), .A2(pi0087), .B(pi0075), .ZN(new_n5498_));
  NOR2_X1    g03048(.A1(pi0054), .A2(pi0092), .ZN(new_n5499_));
  NOR2_X1    g03049(.A1(new_n3079_), .A2(pi0142), .ZN(new_n5500_));
  NOR2_X1    g03050(.A1(new_n5500_), .A2(pi0299), .ZN(new_n5501_));
  AOI21_X1   g03051(.A1(new_n3044_), .A2(pi0299), .B(new_n5501_), .ZN(new_n5502_));
  NOR2_X1    g03052(.A1(new_n3145_), .A2(pi0039), .ZN(new_n5503_));
  INV_X1     g03053(.I(new_n5503_), .ZN(new_n5504_));
  NOR2_X1    g03054(.A1(new_n3462_), .A2(pi0038), .ZN(new_n5505_));
  INV_X1     g03055(.I(new_n5505_), .ZN(new_n5506_));
  NOR2_X1    g03056(.A1(new_n5504_), .A2(new_n5506_), .ZN(new_n5507_));
  INV_X1     g03057(.I(new_n5502_), .ZN(new_n5508_));
  INV_X1     g03058(.I(pi0042), .ZN(new_n5509_));
  INV_X1     g03059(.I(pi0043), .ZN(new_n5510_));
  INV_X1     g03060(.I(pi0052), .ZN(new_n5511_));
  INV_X1     g03061(.I(pi0113), .ZN(new_n5512_));
  INV_X1     g03062(.I(pi0114), .ZN(new_n5513_));
  INV_X1     g03063(.I(pi0115), .ZN(new_n5514_));
  INV_X1     g03064(.I(pi0116), .ZN(new_n5515_));
  NOR4_X1    g03065(.A1(new_n5512_), .A2(new_n5513_), .A3(new_n5514_), .A4(new_n5515_), .ZN(new_n5516_));
  INV_X1     g03066(.I(new_n5516_), .ZN(new_n5517_));
  NOR4_X1    g03067(.A1(new_n5517_), .A2(new_n5509_), .A3(new_n5510_), .A4(new_n5511_), .ZN(new_n5518_));
  INV_X1     g03068(.I(new_n5518_), .ZN(new_n5519_));
  NOR2_X1    g03069(.A1(pi0041), .A2(pi0099), .ZN(new_n5520_));
  INV_X1     g03070(.I(new_n5520_), .ZN(new_n5521_));
  NOR2_X1    g03071(.A1(new_n5521_), .A2(pi0101), .ZN(new_n5522_));
  INV_X1     g03072(.I(new_n5522_), .ZN(new_n5523_));
  NOR2_X1    g03073(.A1(new_n5519_), .A2(new_n5523_), .ZN(new_n5524_));
  INV_X1     g03074(.I(new_n5524_), .ZN(new_n5525_));
  NOR2_X1    g03075(.A1(new_n5525_), .A2(pi0044), .ZN(new_n5526_));
  NOR2_X1    g03076(.A1(new_n5526_), .A2(new_n5508_), .ZN(new_n5527_));
  INV_X1     g03077(.I(pi0683), .ZN(new_n5528_));
  INV_X1     g03078(.I(new_n5526_), .ZN(po1057));
  INV_X1     g03079(.I(pi0250), .ZN(new_n5530_));
  NOR2_X1    g03080(.A1(pi0824), .A2(pi0829), .ZN(new_n5531_));
  NOR2_X1    g03081(.A1(new_n2981_), .A2(new_n5531_), .ZN(new_n5532_));
  INV_X1     g03082(.I(new_n5532_), .ZN(new_n5533_));
  NOR2_X1    g03083(.A1(new_n5533_), .A2(pi1093), .ZN(po0740));
  NOR2_X1    g03084(.A1(new_n5530_), .A2(pi0129), .ZN(new_n5535_));
  AOI21_X1   g03085(.A1(po0740), .A2(new_n5530_), .B(new_n5535_), .ZN(new_n5536_));
  INV_X1     g03086(.I(new_n5536_), .ZN(new_n5537_));
  AOI21_X1   g03087(.A1(po1057), .A2(new_n5528_), .B(new_n5537_), .ZN(new_n5538_));
  NAND2_X1   g03088(.A1(new_n5538_), .A2(new_n5527_), .ZN(new_n5539_));
  NAND3_X1   g03089(.A1(new_n5539_), .A2(pi0087), .A3(new_n5507_), .ZN(new_n5540_));
  AOI21_X1   g03090(.A1(new_n5540_), .A2(new_n5502_), .B(new_n3396_), .ZN(new_n5541_));
  OAI21_X1   g03091(.A1(new_n5498_), .A2(new_n5499_), .B(new_n5541_), .ZN(new_n5542_));
  NOR4_X1    g03092(.A1(new_n5487_), .A2(new_n5493_), .A3(new_n5497_), .A4(new_n5542_), .ZN(new_n5543_));
  OAI21_X1   g03093(.A1(new_n5494_), .A2(new_n3431_), .B(pi0062), .ZN(new_n5544_));
  NAND2_X1   g03094(.A1(new_n5544_), .A2(new_n3230_), .ZN(new_n5545_));
  NOR2_X1    g03095(.A1(new_n5371_), .A2(new_n3229_), .ZN(new_n5546_));
  NOR3_X1    g03096(.A1(new_n3224_), .A2(new_n3226_), .A3(new_n5546_), .ZN(new_n5547_));
  AOI21_X1   g03097(.A1(new_n5547_), .A2(new_n3160_), .B(new_n3230_), .ZN(new_n5548_));
  OAI22_X1   g03098(.A1(new_n5543_), .A2(new_n5545_), .B1(new_n5371_), .B2(new_n5548_), .ZN(po0167));
  INV_X1     g03099(.I(pi1090), .ZN(po0170));
  INV_X1     g03100(.I(pi0232), .ZN(new_n5551_));
  INV_X1     g03101(.I(pi0030), .ZN(new_n5552_));
  NAND2_X1   g03102(.A1(new_n5373_), .A2(pi0602), .ZN(new_n5553_));
  NAND2_X1   g03103(.A1(new_n5378_), .A2(new_n5386_), .ZN(new_n5554_));
  NAND2_X1   g03104(.A1(new_n5554_), .A2(new_n5553_), .ZN(new_n5555_));
  NAND4_X1   g03105(.A1(new_n2495_), .A2(pi0093), .A3(pi0841), .A4(new_n2487_), .ZN(new_n5556_));
  NOR3_X1    g03106(.A1(new_n5556_), .A2(new_n2796_), .A3(new_n2989_), .ZN(new_n5557_));
  INV_X1     g03107(.I(new_n5557_), .ZN(new_n5558_));
  NOR4_X1    g03108(.A1(new_n5558_), .A2(new_n2794_), .A3(new_n2436_), .A4(new_n3072_), .ZN(new_n5559_));
  INV_X1     g03109(.I(new_n5559_), .ZN(new_n5560_));
  NOR2_X1    g03110(.A1(new_n2483_), .A2(new_n3138_), .ZN(new_n5561_));
  NOR2_X1    g03111(.A1(new_n2512_), .A2(pi0109), .ZN(new_n5562_));
  INV_X1     g03112(.I(new_n2861_), .ZN(new_n5563_));
  NOR2_X1    g03113(.A1(new_n2587_), .A2(new_n2575_), .ZN(new_n5564_));
  NAND2_X1   g03114(.A1(new_n5564_), .A2(pi0066), .ZN(new_n5565_));
  XOR2_X1    g03115(.A1(new_n5564_), .A2(new_n2591_), .Z(new_n5566_));
  NAND2_X1   g03116(.A1(new_n5566_), .A2(new_n2589_), .ZN(new_n5567_));
  XOR2_X1    g03117(.A1(new_n5567_), .A2(new_n5565_), .Z(new_n5568_));
  NAND2_X1   g03118(.A1(new_n5568_), .A2(pi0068), .ZN(new_n5569_));
  NOR2_X1    g03119(.A1(new_n2611_), .A2(new_n2598_), .ZN(new_n5570_));
  XOR2_X1    g03120(.A1(new_n5568_), .A2(new_n5570_), .Z(new_n5571_));
  NAND2_X1   g03121(.A1(new_n5571_), .A2(new_n2609_), .ZN(new_n5572_));
  XOR2_X1    g03122(.A1(new_n5572_), .A2(new_n5569_), .Z(new_n5573_));
  NAND2_X1   g03123(.A1(new_n2629_), .A2(pi0067), .ZN(new_n5574_));
  AOI21_X1   g03124(.A1(new_n2623_), .A2(new_n2630_), .B(new_n2633_), .ZN(new_n5575_));
  NAND2_X1   g03125(.A1(new_n5574_), .A2(new_n5575_), .ZN(new_n5576_));
  OAI21_X1   g03126(.A1(new_n2604_), .A2(new_n2607_), .B(new_n2610_), .ZN(new_n5577_));
  NAND3_X1   g03127(.A1(new_n2570_), .A2(new_n2644_), .A3(new_n2539_), .ZN(new_n5578_));
  NOR2_X1    g03128(.A1(new_n5578_), .A2(new_n2492_), .ZN(new_n5579_));
  NOR2_X1    g03129(.A1(new_n5579_), .A2(pi0071), .ZN(new_n5580_));
  INV_X1     g03130(.I(new_n5580_), .ZN(new_n5581_));
  NAND4_X1   g03131(.A1(new_n5573_), .A2(new_n5576_), .A3(new_n5577_), .A4(new_n5581_), .ZN(new_n5582_));
  INV_X1     g03132(.I(new_n2514_), .ZN(new_n5583_));
  AOI21_X1   g03133(.A1(new_n2454_), .A2(new_n2455_), .B(new_n5583_), .ZN(new_n5584_));
  INV_X1     g03134(.I(new_n5584_), .ZN(new_n5585_));
  OAI21_X1   g03135(.A1(new_n5582_), .A2(new_n5585_), .B(new_n2636_), .ZN(new_n5586_));
  AOI21_X1   g03136(.A1(new_n2552_), .A2(new_n2859_), .B(new_n2555_), .ZN(new_n5587_));
  NOR2_X1    g03137(.A1(new_n5587_), .A2(new_n5578_), .ZN(new_n5588_));
  INV_X1     g03138(.I(new_n2658_), .ZN(new_n5589_));
  NOR3_X1    g03139(.A1(new_n5589_), .A2(pi0046), .A3(new_n2873_), .ZN(new_n5590_));
  AOI22_X1   g03140(.A1(new_n5586_), .A2(new_n5588_), .B1(pi0086), .B2(new_n5590_), .ZN(new_n5591_));
  NOR2_X1    g03141(.A1(new_n5591_), .A2(new_n5563_), .ZN(new_n5592_));
  OAI21_X1   g03142(.A1(new_n5592_), .A2(new_n2875_), .B(new_n5562_), .ZN(new_n5593_));
  NOR2_X1    g03143(.A1(pi0091), .A2(pi0314), .ZN(new_n5594_));
  AOI21_X1   g03144(.A1(new_n2684_), .A2(pi0091), .B(pi0058), .ZN(new_n5595_));
  INV_X1     g03145(.I(new_n5595_), .ZN(new_n5596_));
  NAND2_X1   g03146(.A1(new_n5596_), .A2(new_n2679_), .ZN(new_n5597_));
  AOI21_X1   g03147(.A1(new_n5593_), .A2(new_n5594_), .B(new_n5597_), .ZN(new_n5598_));
  INV_X1     g03148(.I(new_n5590_), .ZN(new_n5599_));
  AOI21_X1   g03149(.A1(new_n2555_), .A2(new_n2552_), .B(new_n5584_), .ZN(new_n5600_));
  OAI21_X1   g03150(.A1(new_n5582_), .A2(new_n5600_), .B(new_n2859_), .ZN(new_n5601_));
  AOI21_X1   g03151(.A1(new_n5601_), .A2(new_n5563_), .B(pi0086), .ZN(new_n5602_));
  NOR2_X1    g03152(.A1(new_n5602_), .A2(new_n5599_), .ZN(new_n5603_));
  OAI21_X1   g03153(.A1(new_n5603_), .A2(new_n2875_), .B(new_n5562_), .ZN(new_n5604_));
  NAND3_X1   g03154(.A1(new_n5604_), .A2(new_n2674_), .A3(pi0314), .ZN(new_n5605_));
  INV_X1     g03155(.I(new_n2693_), .ZN(new_n5606_));
  AOI21_X1   g03156(.A1(new_n2732_), .A2(new_n5606_), .B(new_n2507_), .ZN(new_n5607_));
  INV_X1     g03157(.I(new_n5607_), .ZN(new_n5608_));
  OAI22_X1   g03158(.A1(new_n5598_), .A2(new_n5605_), .B1(new_n2509_), .B2(new_n5608_), .ZN(new_n5609_));
  OAI21_X1   g03159(.A1(new_n2758_), .A2(new_n2437_), .B(new_n2707_), .ZN(new_n5610_));
  NAND3_X1   g03160(.A1(new_n5609_), .A2(new_n2680_), .A3(new_n5610_), .ZN(new_n5611_));
  AOI21_X1   g03161(.A1(new_n5611_), .A2(new_n5561_), .B(new_n2827_), .ZN(new_n5612_));
  NAND2_X1   g03162(.A1(new_n5612_), .A2(new_n5560_), .ZN(new_n5613_));
  NAND2_X1   g03163(.A1(new_n5613_), .A2(new_n5373_), .ZN(new_n5614_));
  INV_X1     g03164(.I(new_n5594_), .ZN(new_n5615_));
  OAI21_X1   g03165(.A1(new_n5602_), .A2(new_n5599_), .B(new_n2876_), .ZN(new_n5616_));
  NOR2_X1    g03166(.A1(new_n2877_), .A2(new_n2512_), .ZN(new_n5617_));
  INV_X1     g03167(.I(new_n5617_), .ZN(new_n5618_));
  AOI21_X1   g03168(.A1(new_n5594_), .A2(new_n5596_), .B(new_n5618_), .ZN(new_n5619_));
  AOI21_X1   g03169(.A1(new_n5616_), .A2(new_n5619_), .B(new_n5615_), .ZN(new_n5620_));
  OAI21_X1   g03170(.A1(new_n5592_), .A2(new_n5416_), .B(new_n5617_), .ZN(new_n5621_));
  OAI21_X1   g03171(.A1(new_n5621_), .A2(new_n5620_), .B(pi0090), .ZN(new_n5622_));
  NAND2_X1   g03172(.A1(pi0090), .A2(pi0093), .ZN(new_n5623_));
  XOR2_X1    g03173(.A1(new_n5622_), .A2(new_n5623_), .Z(new_n5624_));
  INV_X1     g03174(.I(new_n5561_), .ZN(new_n5625_));
  OAI21_X1   g03175(.A1(new_n5625_), .A2(new_n2822_), .B(new_n2437_), .ZN(new_n5626_));
  OAI21_X1   g03176(.A1(new_n2758_), .A2(new_n2707_), .B(new_n5608_), .ZN(new_n5627_));
  NAND4_X1   g03177(.A1(new_n5624_), .A2(new_n2470_), .A3(new_n5626_), .A4(new_n5627_), .ZN(new_n5628_));
  NOR2_X1    g03178(.A1(new_n5628_), .A2(new_n5559_), .ZN(new_n5629_));
  OAI21_X1   g03179(.A1(new_n5373_), .A2(new_n5629_), .B(new_n5614_), .ZN(new_n5630_));
  NAND2_X1   g03180(.A1(new_n5630_), .A2(new_n5555_), .ZN(new_n5631_));
  INV_X1     g03181(.I(pi0681), .ZN(new_n5632_));
  INV_X1     g03182(.I(pi0662), .ZN(new_n5633_));
  NAND2_X1   g03183(.A1(new_n5633_), .A2(pi0680), .ZN(new_n5634_));
  NOR2_X1    g03184(.A1(new_n5634_), .A2(pi0661), .ZN(new_n5635_));
  NAND2_X1   g03185(.A1(new_n5635_), .A2(new_n5632_), .ZN(new_n5636_));
  NOR2_X1    g03186(.A1(new_n5636_), .A2(new_n5373_), .ZN(new_n5637_));
  AOI21_X1   g03187(.A1(pi0602), .A2(new_n5373_), .B(new_n5637_), .ZN(new_n5638_));
  NOR2_X1    g03188(.A1(new_n5638_), .A2(new_n3005_), .ZN(new_n5639_));
  XOR2_X1    g03189(.A1(new_n5631_), .A2(new_n5639_), .Z(new_n5640_));
  INV_X1     g03190(.I(pi0145), .ZN(new_n5641_));
  INV_X1     g03191(.I(pi0180), .ZN(new_n5642_));
  INV_X1     g03192(.I(pi0181), .ZN(new_n5643_));
  INV_X1     g03193(.I(pi0182), .ZN(new_n5644_));
  NOR4_X1    g03194(.A1(new_n5641_), .A2(new_n5642_), .A3(new_n5643_), .A4(new_n5644_), .ZN(new_n5645_));
  INV_X1     g03195(.I(new_n5645_), .ZN(new_n5646_));
  NOR3_X1    g03196(.A1(new_n5640_), .A2(new_n5552_), .A3(new_n5646_), .ZN(new_n5647_));
  NOR2_X1    g03197(.A1(new_n3005_), .A2(pi0030), .ZN(new_n5648_));
  AOI21_X1   g03198(.A1(new_n5629_), .A2(new_n3005_), .B(new_n5648_), .ZN(new_n5649_));
  NAND4_X1   g03199(.A1(new_n5649_), .A2(new_n3098_), .A3(new_n5555_), .A4(new_n5645_), .ZN(new_n5650_));
  OAI21_X1   g03200(.A1(new_n5647_), .A2(new_n5650_), .B(new_n5551_), .ZN(new_n5651_));
  AOI21_X1   g03201(.A1(pi0907), .A2(new_n5373_), .B(new_n5637_), .ZN(new_n5652_));
  NOR4_X1    g03202(.A1(new_n5558_), .A2(new_n2794_), .A3(new_n2436_), .A4(new_n2777_), .ZN(new_n5653_));
  NOR2_X1    g03203(.A1(new_n5628_), .A2(new_n5653_), .ZN(new_n5654_));
  NAND2_X1   g03204(.A1(new_n5373_), .A2(pi0907), .ZN(new_n5655_));
  NAND2_X1   g03205(.A1(new_n5554_), .A2(new_n5655_), .ZN(new_n5656_));
  INV_X1     g03206(.I(new_n5653_), .ZN(new_n5657_));
  NAND2_X1   g03207(.A1(new_n5612_), .A2(new_n5657_), .ZN(new_n5658_));
  NAND2_X1   g03208(.A1(new_n5658_), .A2(new_n5373_), .ZN(new_n5659_));
  OAI21_X1   g03209(.A1(new_n5373_), .A2(new_n5654_), .B(new_n5659_), .ZN(new_n5660_));
  INV_X1     g03210(.I(pi0158), .ZN(new_n5661_));
  INV_X1     g03211(.I(pi0159), .ZN(new_n5662_));
  NOR2_X1    g03212(.A1(new_n5661_), .A2(new_n5662_), .ZN(new_n5663_));
  INV_X1     g03213(.I(pi0160), .ZN(new_n5664_));
  INV_X1     g03214(.I(pi0197), .ZN(new_n5665_));
  NOR2_X1    g03215(.A1(new_n5664_), .A2(new_n5665_), .ZN(new_n5666_));
  NAND2_X1   g03216(.A1(new_n5663_), .A2(new_n5666_), .ZN(new_n5667_));
  AOI21_X1   g03217(.A1(new_n5660_), .A2(new_n5656_), .B(new_n5667_), .ZN(new_n5668_));
  NOR2_X1    g03218(.A1(new_n5667_), .A2(new_n3005_), .ZN(new_n5669_));
  XNOR2_X1   g03219(.A1(new_n5668_), .A2(new_n5669_), .ZN(new_n5670_));
  NOR2_X1    g03220(.A1(new_n5552_), .A2(new_n3005_), .ZN(new_n5671_));
  AOI21_X1   g03221(.A1(new_n5656_), .A2(new_n5671_), .B(new_n3098_), .ZN(new_n5672_));
  INV_X1     g03222(.I(new_n5672_), .ZN(new_n5673_));
  NOR4_X1    g03223(.A1(new_n5670_), .A2(new_n5652_), .A3(new_n5654_), .A4(new_n5673_), .ZN(new_n5674_));
  AOI21_X1   g03224(.A1(new_n5649_), .A2(new_n5555_), .B(pi0299), .ZN(new_n5675_));
  OAI22_X1   g03225(.A1(new_n5654_), .A2(new_n5652_), .B1(new_n5551_), .B2(new_n5673_), .ZN(new_n5676_));
  NAND2_X1   g03226(.A1(new_n5676_), .A2(pi0228), .ZN(new_n5677_));
  INV_X1     g03227(.I(new_n5671_), .ZN(new_n5678_));
  NOR2_X1    g03228(.A1(new_n3145_), .A2(pi0287), .ZN(new_n5679_));
  NOR2_X1    g03229(.A1(new_n5408_), .A2(new_n5402_), .ZN(new_n5680_));
  NAND2_X1   g03230(.A1(new_n5679_), .A2(new_n5680_), .ZN(new_n5681_));
  INV_X1     g03231(.I(new_n5681_), .ZN(new_n5682_));
  INV_X1     g03232(.I(pi0824), .ZN(new_n5683_));
  NOR2_X1    g03233(.A1(new_n5683_), .A2(new_n2984_), .ZN(new_n5684_));
  NAND2_X1   g03234(.A1(new_n2980_), .A2(new_n5684_), .ZN(new_n5685_));
  NOR2_X1    g03235(.A1(new_n2728_), .A2(pi0829), .ZN(new_n5686_));
  NOR2_X1    g03236(.A1(new_n5686_), .A2(new_n2726_), .ZN(new_n5687_));
  NOR2_X1    g03237(.A1(new_n5687_), .A2(new_n5685_), .ZN(new_n5688_));
  NAND2_X1   g03238(.A1(new_n5682_), .A2(new_n5688_), .ZN(new_n5689_));
  INV_X1     g03239(.I(new_n5685_), .ZN(new_n5690_));
  NOR2_X1    g03240(.A1(new_n2983_), .A2(new_n2726_), .ZN(new_n5691_));
  INV_X1     g03241(.I(new_n5691_), .ZN(new_n5692_));
  NAND2_X1   g03242(.A1(new_n5692_), .A2(new_n5690_), .ZN(new_n5693_));
  NAND2_X1   g03243(.A1(new_n2745_), .A2(new_n5693_), .ZN(new_n5694_));
  NAND2_X1   g03244(.A1(new_n5682_), .A2(new_n5694_), .ZN(new_n5695_));
  NOR2_X1    g03245(.A1(new_n5681_), .A2(new_n2726_), .ZN(new_n5696_));
  XNOR2_X1   g03246(.A1(new_n5695_), .A2(new_n5696_), .ZN(new_n5697_));
  NAND2_X1   g03247(.A1(new_n5697_), .A2(new_n5690_), .ZN(new_n5698_));
  INV_X1     g03248(.I(new_n5698_), .ZN(new_n5699_));
  NOR2_X1    g03249(.A1(new_n3099_), .A2(pi0223), .ZN(new_n5700_));
  NAND3_X1   g03250(.A1(new_n5699_), .A2(pi0224), .A3(new_n5700_), .ZN(new_n5701_));
  NAND3_X1   g03251(.A1(new_n5698_), .A2(new_n3100_), .A3(new_n5700_), .ZN(new_n5702_));
  AOI21_X1   g03252(.A1(new_n5701_), .A2(new_n5702_), .B(new_n5689_), .ZN(new_n5703_));
  INV_X1     g03253(.I(new_n5703_), .ZN(new_n5704_));
  AOI21_X1   g03254(.A1(new_n5704_), .A2(new_n3005_), .B(new_n5648_), .ZN(new_n5705_));
  OAI21_X1   g03255(.A1(new_n5555_), .A2(pi0039), .B(pi0299), .ZN(new_n5706_));
  OAI21_X1   g03256(.A1(new_n5705_), .A2(new_n5706_), .B(new_n5652_), .ZN(new_n5707_));
  AOI21_X1   g03257(.A1(new_n5689_), .A2(new_n3011_), .B(new_n3362_), .ZN(new_n5708_));
  OAI21_X1   g03258(.A1(new_n5698_), .A2(new_n3011_), .B(new_n5708_), .ZN(new_n5709_));
  NAND2_X1   g03259(.A1(new_n3361_), .A2(pi0228), .ZN(new_n5710_));
  XOR2_X1    g03260(.A1(new_n5709_), .A2(new_n5710_), .Z(new_n5711_));
  NAND2_X1   g03261(.A1(new_n5711_), .A2(pi0030), .ZN(new_n5712_));
  NAND3_X1   g03262(.A1(new_n5707_), .A2(new_n5678_), .A3(new_n5712_), .ZN(new_n5713_));
  AOI21_X1   g03263(.A1(new_n5713_), .A2(new_n3259_), .B(new_n3183_), .ZN(new_n5714_));
  OAI21_X1   g03264(.A1(new_n5675_), .A2(new_n5677_), .B(new_n5714_), .ZN(new_n5715_));
  AOI21_X1   g03265(.A1(new_n5651_), .A2(new_n5674_), .B(new_n5715_), .ZN(new_n5716_));
  NAND2_X1   g03266(.A1(new_n5671_), .A2(pi0299), .ZN(new_n5717_));
  AOI21_X1   g03267(.A1(new_n5652_), .A2(new_n5671_), .B(new_n5717_), .ZN(new_n5718_));
  NOR3_X1    g03268(.A1(new_n5656_), .A2(pi0299), .A3(new_n5678_), .ZN(new_n5719_));
  OAI21_X1   g03269(.A1(new_n5718_), .A2(new_n5719_), .B(new_n5555_), .ZN(new_n5720_));
  INV_X1     g03270(.I(new_n5720_), .ZN(new_n5721_));
  NOR3_X1    g03271(.A1(new_n5716_), .A2(pi0038), .A3(new_n5721_), .ZN(new_n5722_));
  INV_X1     g03272(.I(new_n5500_), .ZN(new_n5723_));
  NOR3_X1    g03273(.A1(new_n5441_), .A2(new_n3721_), .A3(new_n5636_), .ZN(new_n5724_));
  NOR3_X1    g03274(.A1(new_n5440_), .A2(new_n3721_), .A3(new_n5378_), .ZN(new_n5725_));
  OAI21_X1   g03275(.A1(new_n5724_), .A2(new_n5725_), .B(new_n3160_), .ZN(new_n5726_));
  INV_X1     g03276(.I(new_n5726_), .ZN(new_n5727_));
  NOR2_X1    g03277(.A1(new_n5727_), .A2(new_n5723_), .ZN(new_n5728_));
  NOR3_X1    g03278(.A1(new_n5526_), .A2(new_n5528_), .A3(new_n5536_), .ZN(new_n5729_));
  NAND2_X1   g03279(.A1(new_n5729_), .A2(new_n3160_), .ZN(new_n5730_));
  AOI21_X1   g03280(.A1(new_n5386_), .A2(new_n5636_), .B(new_n5730_), .ZN(new_n5731_));
  INV_X1     g03281(.I(new_n5731_), .ZN(new_n5732_));
  NOR3_X1    g03282(.A1(new_n5732_), .A2(new_n3721_), .A3(new_n5723_), .ZN(new_n5733_));
  INV_X1     g03283(.I(new_n5733_), .ZN(new_n5734_));
  NAND2_X1   g03284(.A1(new_n5728_), .A2(new_n5734_), .ZN(new_n5735_));
  NOR2_X1    g03285(.A1(new_n5728_), .A2(new_n5734_), .ZN(new_n5736_));
  NOR2_X1    g03286(.A1(new_n5736_), .A2(pi0228), .ZN(new_n5737_));
  AOI21_X1   g03287(.A1(new_n5737_), .A2(new_n5735_), .B(new_n5553_), .ZN(new_n5738_));
  NOR2_X1    g03288(.A1(new_n5638_), .A2(new_n5678_), .ZN(new_n5739_));
  OAI21_X1   g03289(.A1(new_n5738_), .A2(pi0299), .B(new_n5739_), .ZN(new_n5740_));
  INV_X1     g03290(.I(pi0907), .ZN(new_n5741_));
  AOI21_X1   g03291(.A1(new_n5373_), .A2(new_n5741_), .B(pi0228), .ZN(new_n5742_));
  NAND3_X1   g03292(.A1(new_n5731_), .A2(new_n3030_), .A3(new_n5742_), .ZN(new_n5743_));
  NAND3_X1   g03293(.A1(new_n5732_), .A2(new_n3044_), .A3(new_n5742_), .ZN(new_n5744_));
  NAND2_X1   g03294(.A1(new_n5744_), .A2(new_n5743_), .ZN(new_n5745_));
  NAND3_X1   g03295(.A1(new_n5745_), .A2(new_n5672_), .A3(new_n5727_), .ZN(new_n5746_));
  AOI21_X1   g03296(.A1(new_n5740_), .A2(new_n3212_), .B(new_n5746_), .ZN(new_n5747_));
  NOR2_X1    g03297(.A1(new_n5720_), .A2(new_n3212_), .ZN(new_n5748_));
  OAI21_X1   g03298(.A1(new_n5747_), .A2(pi0100), .B(new_n5748_), .ZN(new_n5749_));
  NAND2_X1   g03299(.A1(new_n5749_), .A2(new_n3455_), .ZN(new_n5750_));
  AOI21_X1   g03300(.A1(new_n3412_), .A2(new_n5678_), .B(pi0039), .ZN(new_n5751_));
  NAND3_X1   g03301(.A1(new_n5751_), .A2(pi0299), .A3(new_n5656_), .ZN(new_n5752_));
  NAND3_X1   g03302(.A1(new_n5751_), .A2(new_n3098_), .A3(new_n5652_), .ZN(new_n5753_));
  NAND2_X1   g03303(.A1(new_n5752_), .A2(new_n5753_), .ZN(new_n5754_));
  NAND4_X1   g03304(.A1(new_n5750_), .A2(pi0100), .A3(new_n5555_), .A4(new_n5754_), .ZN(new_n5755_));
  OAI21_X1   g03305(.A1(new_n5722_), .A2(new_n5755_), .B(new_n3235_), .ZN(new_n5756_));
  NOR2_X1    g03306(.A1(new_n5720_), .A2(new_n3455_), .ZN(new_n5757_));
  AOI21_X1   g03307(.A1(new_n5756_), .A2(new_n5757_), .B(pi0092), .ZN(new_n5758_));
  NAND2_X1   g03308(.A1(new_n5754_), .A2(new_n5555_), .ZN(new_n5759_));
  OAI22_X1   g03309(.A1(new_n5759_), .A2(new_n5720_), .B1(new_n3187_), .B2(new_n3194_), .ZN(new_n5760_));
  NAND2_X1   g03310(.A1(new_n5760_), .A2(pi0075), .ZN(new_n5761_));
  NOR2_X1    g03311(.A1(new_n5760_), .A2(new_n3115_), .ZN(new_n5762_));
  NAND2_X1   g03312(.A1(new_n3188_), .A2(pi0054), .ZN(new_n5763_));
  XNOR2_X1   g03313(.A1(new_n5762_), .A2(new_n5763_), .ZN(new_n5764_));
  NOR2_X1    g03314(.A1(new_n3189_), .A2(pi0054), .ZN(new_n5765_));
  NOR2_X1    g03315(.A1(pi0055), .A2(pi0074), .ZN(new_n5766_));
  INV_X1     g03316(.I(new_n5766_), .ZN(new_n5767_));
  AOI21_X1   g03317(.A1(new_n5760_), .A2(new_n5765_), .B(new_n5767_), .ZN(new_n5768_));
  INV_X1     g03318(.I(new_n5765_), .ZN(new_n5769_));
  NAND2_X1   g03319(.A1(new_n5720_), .A2(new_n5769_), .ZN(new_n5770_));
  OAI21_X1   g03320(.A1(new_n5768_), .A2(new_n5770_), .B(new_n3175_), .ZN(new_n5771_));
  AOI21_X1   g03321(.A1(new_n5764_), .A2(new_n5721_), .B(new_n5771_), .ZN(new_n5772_));
  NOR2_X1    g03322(.A1(new_n5760_), .A2(new_n3303_), .ZN(new_n5773_));
  XOR2_X1    g03323(.A1(new_n5773_), .A2(new_n3483_), .Z(new_n5774_));
  OAI21_X1   g03324(.A1(new_n5774_), .A2(new_n5720_), .B(new_n3115_), .ZN(new_n5775_));
  NOR2_X1    g03325(.A1(new_n5772_), .A2(new_n5775_), .ZN(new_n5776_));
  OAI21_X1   g03326(.A1(new_n5758_), .A2(new_n5761_), .B(new_n5776_), .ZN(new_n5777_));
  NOR2_X1    g03327(.A1(new_n3291_), .A2(new_n3005_), .ZN(new_n5778_));
  NAND2_X1   g03328(.A1(new_n3160_), .A2(new_n5671_), .ZN(new_n5779_));
  XOR2_X1    g03329(.A1(new_n5778_), .A2(new_n5779_), .Z(new_n5780_));
  NOR2_X1    g03330(.A1(new_n5780_), .A2(new_n5652_), .ZN(new_n5781_));
  NAND2_X1   g03331(.A1(new_n5678_), .A2(new_n3229_), .ZN(new_n5782_));
  NOR2_X1    g03332(.A1(new_n5656_), .A2(new_n5782_), .ZN(new_n5783_));
  NOR2_X1    g03333(.A1(new_n5781_), .A2(pi0057), .ZN(new_n5784_));
  NAND2_X1   g03334(.A1(new_n3225_), .A2(new_n3258_), .ZN(new_n5785_));
  NAND2_X1   g03335(.A1(new_n5785_), .A2(new_n3005_), .ZN(new_n5786_));
  NOR2_X1    g03336(.A1(new_n5785_), .A2(pi0059), .ZN(new_n5787_));
  INV_X1     g03337(.I(new_n5787_), .ZN(new_n5788_));
  NOR3_X1    g03338(.A1(new_n5788_), .A2(new_n3005_), .A3(new_n5786_), .ZN(new_n5789_));
  OAI21_X1   g03339(.A1(new_n5781_), .A2(new_n5546_), .B(new_n5789_), .ZN(new_n5790_));
  OAI22_X1   g03340(.A1(new_n5790_), .A2(new_n5784_), .B1(new_n3226_), .B2(new_n5783_), .ZN(new_n5791_));
  NAND3_X1   g03341(.A1(new_n5791_), .A2(pi0055), .A3(new_n5781_), .ZN(new_n5792_));
  AOI21_X1   g03342(.A1(new_n5777_), .A2(new_n3226_), .B(new_n5792_), .ZN(po0171));
  INV_X1     g03343(.I(pi0603), .ZN(new_n5794_));
  NOR2_X1    g03344(.A1(new_n5794_), .A2(pi0642), .ZN(new_n5795_));
  NAND2_X1   g03345(.A1(new_n5795_), .A2(new_n5381_), .ZN(new_n5796_));
  NOR2_X1    g03346(.A1(new_n5796_), .A2(new_n5373_), .ZN(new_n5797_));
  AOI21_X1   g03347(.A1(pi0947), .A2(new_n5373_), .B(new_n5797_), .ZN(new_n5798_));
  NOR2_X1    g03348(.A1(new_n5654_), .A2(new_n5798_), .ZN(new_n5799_));
  INV_X1     g03349(.I(pi0947), .ZN(new_n5800_));
  NAND2_X1   g03350(.A1(new_n5383_), .A2(new_n5386_), .ZN(new_n5801_));
  OAI21_X1   g03351(.A1(new_n5800_), .A2(new_n5386_), .B(new_n5801_), .ZN(new_n5802_));
  AOI21_X1   g03352(.A1(new_n5802_), .A2(new_n5671_), .B(new_n3098_), .ZN(new_n5803_));
  AOI21_X1   g03353(.A1(pi0232), .A2(new_n5803_), .B(new_n5799_), .ZN(new_n5804_));
  NOR2_X1    g03354(.A1(new_n5804_), .A2(new_n3005_), .ZN(new_n5805_));
  INV_X1     g03355(.I(new_n5649_), .ZN(new_n5806_));
  AOI21_X1   g03356(.A1(pi0587), .A2(new_n5373_), .B(new_n5797_), .ZN(new_n5807_));
  NOR2_X1    g03357(.A1(new_n5806_), .A2(new_n5807_), .ZN(new_n5808_));
  OAI21_X1   g03358(.A1(new_n5392_), .A2(new_n5386_), .B(new_n5801_), .ZN(new_n5809_));
  NAND2_X1   g03359(.A1(new_n5630_), .A2(new_n5809_), .ZN(new_n5810_));
  NOR2_X1    g03360(.A1(new_n5807_), .A2(new_n3005_), .ZN(new_n5811_));
  XOR2_X1    g03361(.A1(new_n5810_), .A2(new_n5811_), .Z(new_n5812_));
  OAI21_X1   g03362(.A1(new_n5812_), .A2(new_n5552_), .B(new_n5645_), .ZN(new_n5813_));
  NAND2_X1   g03363(.A1(new_n5645_), .A2(pi0299), .ZN(new_n5814_));
  XOR2_X1    g03364(.A1(new_n5813_), .A2(new_n5814_), .Z(new_n5815_));
  NAND2_X1   g03365(.A1(new_n5815_), .A2(new_n5808_), .ZN(new_n5816_));
  AOI21_X1   g03366(.A1(new_n5660_), .A2(new_n5802_), .B(new_n5667_), .ZN(new_n5817_));
  XOR2_X1    g03367(.A1(new_n5817_), .A2(new_n5669_), .Z(new_n5818_));
  NAND4_X1   g03368(.A1(new_n5818_), .A2(pi0039), .A3(new_n5799_), .A4(new_n5803_), .ZN(new_n5819_));
  AOI21_X1   g03369(.A1(new_n5816_), .A2(new_n5551_), .B(new_n5819_), .ZN(new_n5820_));
  NOR2_X1    g03370(.A1(new_n5808_), .A2(pi0299), .ZN(new_n5821_));
  OAI21_X1   g03371(.A1(new_n5820_), .A2(new_n5805_), .B(new_n5821_), .ZN(new_n5822_));
  NAND2_X1   g03372(.A1(new_n5822_), .A2(new_n3259_), .ZN(new_n5823_));
  INV_X1     g03373(.I(new_n5712_), .ZN(new_n5824_));
  NOR2_X1    g03374(.A1(new_n3362_), .A2(new_n3098_), .ZN(new_n5825_));
  AOI22_X1   g03375(.A1(new_n5824_), .A2(new_n5825_), .B1(new_n5802_), .B2(new_n5803_), .ZN(new_n5826_));
  NOR2_X1    g03376(.A1(new_n3183_), .A2(new_n3098_), .ZN(new_n5827_));
  NOR2_X1    g03377(.A1(new_n5809_), .A2(new_n5827_), .ZN(new_n5828_));
  NOR3_X1    g03378(.A1(new_n5826_), .A2(new_n5705_), .A3(new_n5828_), .ZN(new_n5829_));
  NAND3_X1   g03379(.A1(new_n5802_), .A2(pi0299), .A3(new_n5671_), .ZN(new_n5830_));
  NAND3_X1   g03380(.A1(new_n5798_), .A2(new_n5671_), .A3(new_n5717_), .ZN(new_n5831_));
  AOI21_X1   g03381(.A1(new_n5830_), .A2(new_n5831_), .B(new_n5807_), .ZN(new_n5832_));
  INV_X1     g03382(.I(new_n5832_), .ZN(new_n5833_));
  NAND2_X1   g03383(.A1(new_n5833_), .A2(new_n3259_), .ZN(new_n5834_));
  AOI21_X1   g03384(.A1(new_n5823_), .A2(new_n5829_), .B(new_n5834_), .ZN(new_n5835_));
  INV_X1     g03385(.I(new_n5730_), .ZN(new_n5836_));
  OAI21_X1   g03386(.A1(new_n5373_), .A2(new_n5383_), .B(new_n5836_), .ZN(new_n5837_));
  NOR3_X1    g03387(.A1(new_n5441_), .A2(new_n3721_), .A3(new_n5796_), .ZN(new_n5838_));
  NOR3_X1    g03388(.A1(new_n5440_), .A2(new_n3721_), .A3(new_n5383_), .ZN(new_n5839_));
  OAI21_X1   g03389(.A1(new_n5838_), .A2(new_n5839_), .B(new_n3160_), .ZN(new_n5840_));
  NOR2_X1    g03390(.A1(new_n3005_), .A2(new_n5392_), .ZN(new_n5841_));
  OAI21_X1   g03391(.A1(new_n5383_), .A2(new_n5841_), .B(new_n5373_), .ZN(new_n5842_));
  INV_X1     g03392(.I(new_n5842_), .ZN(new_n5843_));
  NAND2_X1   g03393(.A1(new_n5840_), .A2(new_n5843_), .ZN(new_n5844_));
  NOR2_X1    g03394(.A1(new_n5842_), .A2(new_n3089_), .ZN(new_n5845_));
  XOR2_X1    g03395(.A1(new_n5844_), .A2(new_n5845_), .Z(new_n5846_));
  OAI22_X1   g03396(.A1(new_n5846_), .A2(new_n5837_), .B1(new_n5678_), .B2(new_n5807_), .ZN(new_n5847_));
  NOR2_X1    g03397(.A1(new_n5386_), .A2(pi0587), .ZN(new_n5848_));
  NOR2_X1    g03398(.A1(new_n3080_), .A2(pi0228), .ZN(new_n5849_));
  OAI21_X1   g03399(.A1(new_n5840_), .A2(new_n5848_), .B(new_n5849_), .ZN(new_n5850_));
  NAND3_X1   g03400(.A1(new_n3030_), .A2(pi0947), .A3(new_n5373_), .ZN(new_n5851_));
  OAI21_X1   g03401(.A1(new_n5840_), .A2(new_n5837_), .B(new_n5851_), .ZN(new_n5852_));
  NAND2_X1   g03402(.A1(new_n5803_), .A2(new_n3211_), .ZN(new_n5853_));
  AOI21_X1   g03403(.A1(new_n5853_), .A2(new_n3005_), .B(new_n3098_), .ZN(new_n5854_));
  NAND2_X1   g03404(.A1(new_n5852_), .A2(new_n5854_), .ZN(new_n5855_));
  NAND2_X1   g03405(.A1(new_n3079_), .A2(pi0228), .ZN(new_n5856_));
  AOI21_X1   g03406(.A1(new_n5855_), .A2(new_n5850_), .B(new_n5856_), .ZN(new_n5857_));
  AOI21_X1   g03407(.A1(new_n5847_), .A2(new_n5857_), .B(pi0100), .ZN(new_n5858_));
  NAND2_X1   g03408(.A1(new_n5832_), .A2(new_n3211_), .ZN(new_n5859_));
  OAI21_X1   g03409(.A1(new_n5858_), .A2(new_n5859_), .B(new_n3455_), .ZN(new_n5860_));
  NAND3_X1   g03410(.A1(new_n5751_), .A2(pi0299), .A3(new_n5802_), .ZN(new_n5861_));
  NAND3_X1   g03411(.A1(new_n5751_), .A2(new_n3098_), .A3(new_n5798_), .ZN(new_n5862_));
  AOI21_X1   g03412(.A1(new_n5861_), .A2(new_n5862_), .B(new_n5807_), .ZN(new_n5863_));
  NAND3_X1   g03413(.A1(new_n5860_), .A2(pi0100), .A3(new_n5863_), .ZN(new_n5864_));
  OAI21_X1   g03414(.A1(new_n5835_), .A2(new_n5864_), .B(new_n3235_), .ZN(new_n5865_));
  NOR2_X1    g03415(.A1(new_n5833_), .A2(new_n3455_), .ZN(new_n5866_));
  AOI21_X1   g03416(.A1(new_n5865_), .A2(new_n5866_), .B(pi0092), .ZN(new_n5867_));
  NOR2_X1    g03417(.A1(new_n3194_), .A2(new_n3187_), .ZN(new_n5868_));
  AOI21_X1   g03418(.A1(new_n5863_), .A2(new_n5832_), .B(new_n5868_), .ZN(new_n5869_));
  OR2_X2     g03419(.A1(new_n5869_), .A2(new_n3235_), .Z(new_n5870_));
  NAND2_X1   g03420(.A1(new_n5869_), .A2(pi0054), .ZN(new_n5871_));
  XOR2_X1    g03421(.A1(new_n5871_), .A2(new_n5763_), .Z(new_n5872_));
  NAND3_X1   g03422(.A1(new_n5833_), .A2(new_n5769_), .A3(new_n5767_), .ZN(new_n5873_));
  NAND2_X1   g03423(.A1(new_n5873_), .A2(new_n3175_), .ZN(new_n5874_));
  AOI21_X1   g03424(.A1(new_n5872_), .A2(new_n5832_), .B(new_n5874_), .ZN(new_n5875_));
  NAND2_X1   g03425(.A1(new_n5869_), .A2(pi0092), .ZN(new_n5876_));
  XNOR2_X1   g03426(.A1(new_n5876_), .A2(new_n3483_), .ZN(new_n5877_));
  OAI21_X1   g03427(.A1(new_n5877_), .A2(new_n5833_), .B(new_n3115_), .ZN(new_n5878_));
  NOR2_X1    g03428(.A1(new_n5878_), .A2(new_n5875_), .ZN(new_n5879_));
  OAI21_X1   g03429(.A1(new_n5867_), .A2(new_n5870_), .B(new_n5879_), .ZN(new_n5880_));
  NOR2_X1    g03430(.A1(new_n5780_), .A2(new_n5798_), .ZN(new_n5881_));
  NOR2_X1    g03431(.A1(new_n5802_), .A2(new_n5782_), .ZN(new_n5882_));
  NOR2_X1    g03432(.A1(new_n5881_), .A2(pi0057), .ZN(new_n5883_));
  OAI21_X1   g03433(.A1(new_n5881_), .A2(new_n5546_), .B(new_n5789_), .ZN(new_n5884_));
  OAI22_X1   g03434(.A1(new_n5884_), .A2(new_n5883_), .B1(new_n3226_), .B2(new_n5882_), .ZN(new_n5885_));
  NAND3_X1   g03435(.A1(new_n5885_), .A2(pi0055), .A3(new_n5881_), .ZN(new_n5886_));
  AOI21_X1   g03436(.A1(new_n5880_), .A2(new_n3226_), .B(new_n5886_), .ZN(po0172));
  NOR2_X1    g03437(.A1(new_n5678_), .A2(new_n5386_), .ZN(new_n5888_));
  INV_X1     g03438(.I(new_n5888_), .ZN(new_n5889_));
  NOR2_X1    g03439(.A1(new_n5889_), .A2(new_n5446_), .ZN(new_n5890_));
  NAND2_X1   g03440(.A1(new_n5659_), .A2(new_n5666_), .ZN(new_n5891_));
  NAND2_X1   g03441(.A1(new_n5654_), .A2(new_n5666_), .ZN(new_n5892_));
  XOR2_X1    g03442(.A1(new_n5891_), .A2(new_n5892_), .Z(new_n5893_));
  NAND2_X1   g03443(.A1(new_n5893_), .A2(new_n5373_), .ZN(new_n5894_));
  INV_X1     g03444(.I(new_n5894_), .ZN(new_n5895_));
  INV_X1     g03445(.I(new_n5663_), .ZN(new_n5896_));
  NOR2_X1    g03446(.A1(new_n5896_), .A2(new_n3005_), .ZN(new_n5897_));
  OAI21_X1   g03447(.A1(new_n5895_), .A2(new_n5890_), .B(new_n5897_), .ZN(new_n5898_));
  INV_X1     g03448(.I(new_n5654_), .ZN(new_n5899_));
  NAND2_X1   g03449(.A1(new_n5899_), .A2(new_n5373_), .ZN(new_n5900_));
  NOR2_X1    g03450(.A1(pi0299), .A2(pi0970), .ZN(new_n5901_));
  NAND2_X1   g03451(.A1(new_n5900_), .A2(new_n5901_), .ZN(new_n5902_));
  NAND2_X1   g03452(.A1(new_n5902_), .A2(pi0228), .ZN(new_n5903_));
  NOR2_X1    g03453(.A1(new_n5614_), .A2(pi0228), .ZN(new_n5904_));
  INV_X1     g03454(.I(new_n5904_), .ZN(new_n5905_));
  INV_X1     g03455(.I(new_n5629_), .ZN(new_n5906_));
  AOI21_X1   g03456(.A1(new_n5906_), .A2(new_n5646_), .B(new_n5888_), .ZN(new_n5907_));
  NOR2_X1    g03457(.A1(new_n5806_), .A2(new_n5386_), .ZN(new_n5908_));
  INV_X1     g03458(.I(new_n5908_), .ZN(new_n5909_));
  AOI22_X1   g03459(.A1(new_n5909_), .A2(new_n5646_), .B1(new_n5907_), .B2(new_n5905_), .ZN(new_n5910_));
  INV_X1     g03460(.I(new_n5910_), .ZN(new_n5911_));
  NOR2_X1    g03461(.A1(new_n5551_), .A2(new_n3098_), .ZN(new_n5912_));
  NOR2_X1    g03462(.A1(new_n5912_), .A2(pi0967), .ZN(new_n5913_));
  AOI21_X1   g03463(.A1(new_n5908_), .A2(pi0967), .B(pi0299), .ZN(new_n5914_));
  NOR2_X1    g03464(.A1(new_n3183_), .A2(pi0232), .ZN(new_n5915_));
  NAND2_X1   g03465(.A1(new_n5903_), .A2(new_n5915_), .ZN(new_n5916_));
  OAI22_X1   g03466(.A1(new_n5911_), .A2(new_n5913_), .B1(new_n5914_), .B2(new_n5916_), .ZN(new_n5917_));
  NOR2_X1    g03467(.A1(new_n5896_), .A2(pi0299), .ZN(new_n5918_));
  NAND4_X1   g03468(.A1(new_n5917_), .A2(new_n5898_), .A3(new_n5903_), .A4(new_n5918_), .ZN(new_n5919_));
  OAI21_X1   g03469(.A1(new_n5709_), .A2(new_n5386_), .B(new_n3005_), .ZN(new_n5920_));
  NAND2_X1   g03470(.A1(new_n5920_), .A2(pi0299), .ZN(new_n5921_));
  INV_X1     g03471(.I(new_n5921_), .ZN(new_n5922_));
  AOI21_X1   g03472(.A1(pi0039), .A2(pi0228), .B(new_n5373_), .ZN(new_n5923_));
  NOR3_X1    g03473(.A1(new_n5923_), .A2(new_n5552_), .A3(new_n3259_), .ZN(new_n5924_));
  AOI21_X1   g03474(.A1(new_n5922_), .A2(pi0970), .B(new_n5924_), .ZN(new_n5925_));
  OAI21_X1   g03475(.A1(new_n5704_), .A2(new_n5386_), .B(new_n3005_), .ZN(new_n5926_));
  NAND2_X1   g03476(.A1(new_n5926_), .A2(new_n3098_), .ZN(new_n5927_));
  NOR3_X1    g03477(.A1(new_n5927_), .A2(new_n5395_), .A3(new_n5925_), .ZN(new_n5928_));
  NOR2_X1    g03478(.A1(new_n5441_), .A2(new_n3721_), .ZN(new_n5929_));
  INV_X1     g03479(.I(new_n5929_), .ZN(new_n5930_));
  NOR2_X1    g03480(.A1(new_n5730_), .A2(new_n5386_), .ZN(new_n5931_));
  INV_X1     g03481(.I(new_n5931_), .ZN(new_n5932_));
  NOR4_X1    g03482(.A1(new_n5930_), .A2(new_n5932_), .A3(new_n3005_), .A4(new_n5723_), .ZN(new_n5933_));
  OAI21_X1   g03483(.A1(new_n5933_), .A2(pi0030), .B(new_n5373_), .ZN(new_n5934_));
  INV_X1     g03484(.I(new_n5934_), .ZN(new_n5935_));
  NOR3_X1    g03485(.A1(new_n5930_), .A2(new_n3005_), .A3(new_n3044_), .ZN(new_n5936_));
  NOR3_X1    g03486(.A1(new_n5929_), .A2(pi0228), .A3(new_n3044_), .ZN(new_n5937_));
  OAI21_X1   g03487(.A1(new_n5936_), .A2(new_n5937_), .B(new_n5931_), .ZN(new_n5938_));
  OAI21_X1   g03488(.A1(new_n3211_), .A2(pi0970), .B(pi0299), .ZN(new_n5939_));
  OAI21_X1   g03489(.A1(new_n5938_), .A2(new_n5939_), .B(new_n5395_), .ZN(new_n5940_));
  AOI21_X1   g03490(.A1(new_n5940_), .A2(new_n5935_), .B(pi0100), .ZN(new_n5941_));
  NAND2_X1   g03491(.A1(new_n5888_), .A2(new_n5446_), .ZN(new_n5942_));
  NAND2_X1   g03492(.A1(new_n5888_), .A2(pi0299), .ZN(new_n5943_));
  XOR2_X1    g03493(.A1(new_n5942_), .A2(new_n5943_), .Z(new_n5944_));
  NAND2_X1   g03494(.A1(new_n5944_), .A2(pi0967), .ZN(new_n5945_));
  INV_X1     g03495(.I(new_n5945_), .ZN(new_n5946_));
  NAND2_X1   g03496(.A1(new_n5946_), .A2(new_n3211_), .ZN(new_n5947_));
  OAI21_X1   g03497(.A1(new_n5941_), .A2(new_n5947_), .B(new_n3455_), .ZN(new_n5948_));
  NOR2_X1    g03498(.A1(new_n3139_), .A2(new_n5386_), .ZN(new_n5949_));
  NOR2_X1    g03499(.A1(new_n5386_), .A2(new_n3005_), .ZN(new_n5950_));
  XOR2_X1    g03500(.A1(new_n5949_), .A2(new_n5950_), .Z(new_n5951_));
  NAND2_X1   g03501(.A1(new_n5951_), .A2(pi0030), .ZN(new_n5952_));
  OAI21_X1   g03502(.A1(new_n5952_), .A2(new_n5395_), .B(new_n3098_), .ZN(new_n5953_));
  NOR2_X1    g03503(.A1(new_n5890_), .A2(new_n3098_), .ZN(new_n5954_));
  NOR2_X1    g03504(.A1(new_n5441_), .A2(pi0228), .ZN(new_n5955_));
  INV_X1     g03505(.I(new_n5955_), .ZN(new_n5956_));
  NOR2_X1    g03506(.A1(new_n5956_), .A2(new_n5446_), .ZN(new_n5957_));
  NAND2_X1   g03507(.A1(new_n5957_), .A2(new_n5954_), .ZN(new_n5958_));
  AOI21_X1   g03508(.A1(new_n5953_), .A2(new_n3183_), .B(new_n5958_), .ZN(new_n5959_));
  NOR2_X1    g03509(.A1(new_n5945_), .A2(new_n3183_), .ZN(new_n5960_));
  OAI21_X1   g03510(.A1(new_n5959_), .A2(pi0038), .B(new_n5960_), .ZN(new_n5961_));
  NAND3_X1   g03511(.A1(new_n5948_), .A2(pi0100), .A3(new_n5961_), .ZN(new_n5962_));
  AOI21_X1   g03512(.A1(new_n5919_), .A2(new_n5928_), .B(new_n5962_), .ZN(new_n5963_));
  NOR2_X1    g03513(.A1(new_n5945_), .A2(new_n3455_), .ZN(new_n5964_));
  OAI21_X1   g03514(.A1(new_n5963_), .A2(pi0075), .B(new_n5964_), .ZN(new_n5965_));
  AOI21_X1   g03515(.A1(new_n5959_), .A2(new_n5946_), .B(new_n5868_), .ZN(new_n5966_));
  NAND2_X1   g03516(.A1(new_n5966_), .A2(pi0092), .ZN(new_n5967_));
  XNOR2_X1   g03517(.A1(new_n5967_), .A2(new_n3483_), .ZN(new_n5968_));
  NOR2_X1    g03518(.A1(new_n5968_), .A2(new_n5945_), .ZN(new_n5969_));
  NAND2_X1   g03519(.A1(new_n3115_), .A2(pi0074), .ZN(new_n5970_));
  NOR2_X1    g03520(.A1(new_n5966_), .A2(new_n3235_), .ZN(new_n5971_));
  OAI21_X1   g03521(.A1(new_n5969_), .A2(new_n5970_), .B(new_n5971_), .ZN(new_n5972_));
  AOI21_X1   g03522(.A1(new_n5965_), .A2(new_n3303_), .B(new_n5972_), .ZN(new_n5973_));
  INV_X1     g03523(.I(new_n5890_), .ZN(new_n5974_));
  NOR2_X1    g03524(.A1(new_n3225_), .A2(pi0055), .ZN(new_n5975_));
  INV_X1     g03525(.I(new_n5975_), .ZN(new_n5976_));
  AOI21_X1   g03526(.A1(new_n5957_), .A2(new_n3291_), .B(new_n5976_), .ZN(new_n5977_));
  OAI21_X1   g03527(.A1(new_n5977_), .A2(new_n5974_), .B(new_n3258_), .ZN(new_n5978_));
  NAND2_X1   g03528(.A1(new_n5945_), .A2(new_n5769_), .ZN(new_n5979_));
  AOI21_X1   g03529(.A1(new_n5979_), .A2(pi0074), .B(new_n3188_), .ZN(new_n5980_));
  AOI21_X1   g03530(.A1(new_n5966_), .A2(new_n5980_), .B(new_n3115_), .ZN(new_n5981_));
  OAI21_X1   g03531(.A1(new_n5973_), .A2(new_n5978_), .B(new_n5981_), .ZN(new_n5982_));
  NAND2_X1   g03532(.A1(new_n5982_), .A2(new_n3229_), .ZN(new_n5983_));
  NOR2_X1    g03533(.A1(new_n5974_), .A2(new_n3226_), .ZN(new_n5984_));
  AOI21_X1   g03534(.A1(new_n5983_), .A2(new_n5984_), .B(new_n5371_), .ZN(new_n5985_));
  NAND2_X1   g03535(.A1(new_n5957_), .A2(new_n3291_), .ZN(new_n5986_));
  NOR2_X1    g03536(.A1(new_n5785_), .A2(new_n5371_), .ZN(new_n5987_));
  NAND3_X1   g03537(.A1(new_n5974_), .A2(pi0059), .A3(new_n5987_), .ZN(new_n5988_));
  NOR3_X1    g03538(.A1(new_n5986_), .A2(new_n5787_), .A3(new_n5988_), .ZN(new_n5989_));
  XOR2_X1    g03539(.A1(new_n5985_), .A2(new_n5989_), .Z(po0173));
  NOR2_X1    g03540(.A1(new_n5889_), .A2(new_n5447_), .ZN(new_n5991_));
  OAI21_X1   g03541(.A1(new_n5895_), .A2(new_n5991_), .B(new_n5897_), .ZN(new_n5992_));
  NOR2_X1    g03542(.A1(pi0299), .A2(pi0972), .ZN(new_n5993_));
  NAND2_X1   g03543(.A1(new_n5900_), .A2(new_n5993_), .ZN(new_n5994_));
  NAND2_X1   g03544(.A1(new_n5994_), .A2(pi0228), .ZN(new_n5995_));
  NOR2_X1    g03545(.A1(new_n5912_), .A2(pi0961), .ZN(new_n5996_));
  AOI21_X1   g03546(.A1(new_n5908_), .A2(pi0961), .B(pi0299), .ZN(new_n5997_));
  NAND2_X1   g03547(.A1(new_n5995_), .A2(new_n5915_), .ZN(new_n5998_));
  OAI22_X1   g03548(.A1(new_n5911_), .A2(new_n5996_), .B1(new_n5997_), .B2(new_n5998_), .ZN(new_n5999_));
  NAND4_X1   g03549(.A1(new_n5999_), .A2(new_n5992_), .A3(new_n5918_), .A4(new_n5995_), .ZN(new_n6000_));
  AOI21_X1   g03550(.A1(new_n5922_), .A2(pi0972), .B(new_n5924_), .ZN(new_n6001_));
  NOR3_X1    g03551(.A1(new_n5927_), .A2(new_n5394_), .A3(new_n6001_), .ZN(new_n6002_));
  OAI21_X1   g03552(.A1(new_n3211_), .A2(pi0972), .B(pi0299), .ZN(new_n6003_));
  OAI21_X1   g03553(.A1(new_n5938_), .A2(new_n6003_), .B(new_n5394_), .ZN(new_n6004_));
  AOI21_X1   g03554(.A1(new_n6004_), .A2(new_n5935_), .B(pi0100), .ZN(new_n6005_));
  NAND2_X1   g03555(.A1(new_n5888_), .A2(new_n5447_), .ZN(new_n6006_));
  XOR2_X1    g03556(.A1(new_n5943_), .A2(new_n6006_), .Z(new_n6007_));
  NAND2_X1   g03557(.A1(new_n6007_), .A2(pi0961), .ZN(new_n6008_));
  INV_X1     g03558(.I(new_n6008_), .ZN(new_n6009_));
  NAND2_X1   g03559(.A1(new_n6009_), .A2(new_n3211_), .ZN(new_n6010_));
  OAI21_X1   g03560(.A1(new_n6005_), .A2(new_n6010_), .B(new_n3455_), .ZN(new_n6011_));
  OAI21_X1   g03561(.A1(new_n5952_), .A2(new_n5394_), .B(new_n3098_), .ZN(new_n6012_));
  NOR2_X1    g03562(.A1(new_n5991_), .A2(new_n3098_), .ZN(new_n6013_));
  NOR2_X1    g03563(.A1(new_n5956_), .A2(new_n5447_), .ZN(new_n6014_));
  NAND2_X1   g03564(.A1(new_n6014_), .A2(new_n6013_), .ZN(new_n6015_));
  AOI21_X1   g03565(.A1(new_n6012_), .A2(new_n3183_), .B(new_n6015_), .ZN(new_n6016_));
  NOR2_X1    g03566(.A1(new_n6008_), .A2(new_n3183_), .ZN(new_n6017_));
  OAI21_X1   g03567(.A1(new_n6016_), .A2(pi0038), .B(new_n6017_), .ZN(new_n6018_));
  NAND3_X1   g03568(.A1(new_n6011_), .A2(pi0100), .A3(new_n6018_), .ZN(new_n6019_));
  AOI21_X1   g03569(.A1(new_n6000_), .A2(new_n6002_), .B(new_n6019_), .ZN(new_n6020_));
  NOR2_X1    g03570(.A1(new_n6008_), .A2(new_n3455_), .ZN(new_n6021_));
  OAI21_X1   g03571(.A1(new_n6020_), .A2(pi0075), .B(new_n6021_), .ZN(new_n6022_));
  AOI21_X1   g03572(.A1(new_n6016_), .A2(new_n6009_), .B(new_n5868_), .ZN(new_n6023_));
  NAND2_X1   g03573(.A1(new_n6023_), .A2(pi0092), .ZN(new_n6024_));
  XNOR2_X1   g03574(.A1(new_n6024_), .A2(new_n3483_), .ZN(new_n6025_));
  NOR2_X1    g03575(.A1(new_n6025_), .A2(new_n6008_), .ZN(new_n6026_));
  NAND2_X1   g03576(.A1(new_n3115_), .A2(pi0074), .ZN(new_n6027_));
  NOR2_X1    g03577(.A1(new_n6023_), .A2(new_n3235_), .ZN(new_n6028_));
  OAI21_X1   g03578(.A1(new_n6026_), .A2(new_n6027_), .B(new_n6028_), .ZN(new_n6029_));
  AOI21_X1   g03579(.A1(new_n6022_), .A2(new_n3303_), .B(new_n6029_), .ZN(new_n6030_));
  INV_X1     g03580(.I(new_n5991_), .ZN(new_n6031_));
  AOI21_X1   g03581(.A1(new_n6014_), .A2(new_n3291_), .B(new_n5976_), .ZN(new_n6032_));
  OAI21_X1   g03582(.A1(new_n6032_), .A2(new_n6031_), .B(new_n3258_), .ZN(new_n6033_));
  NAND2_X1   g03583(.A1(new_n6008_), .A2(new_n5769_), .ZN(new_n6034_));
  AOI21_X1   g03584(.A1(new_n6034_), .A2(pi0074), .B(new_n3188_), .ZN(new_n6035_));
  AOI21_X1   g03585(.A1(new_n6023_), .A2(new_n6035_), .B(new_n3115_), .ZN(new_n6036_));
  OAI21_X1   g03586(.A1(new_n6030_), .A2(new_n6033_), .B(new_n6036_), .ZN(new_n6037_));
  NAND2_X1   g03587(.A1(new_n6037_), .A2(new_n3229_), .ZN(new_n6038_));
  NOR2_X1    g03588(.A1(new_n6031_), .A2(new_n3226_), .ZN(new_n6039_));
  AOI21_X1   g03589(.A1(new_n6038_), .A2(new_n6039_), .B(new_n5371_), .ZN(new_n6040_));
  NAND2_X1   g03590(.A1(new_n6014_), .A2(new_n3291_), .ZN(new_n6041_));
  NAND3_X1   g03591(.A1(new_n6031_), .A2(pi0059), .A3(new_n5987_), .ZN(new_n6042_));
  NOR3_X1    g03592(.A1(new_n6041_), .A2(new_n5787_), .A3(new_n6042_), .ZN(new_n6043_));
  XOR2_X1    g03593(.A1(new_n6040_), .A2(new_n6043_), .Z(po0174));
  INV_X1     g03594(.I(pi0960), .ZN(new_n6045_));
  NOR2_X1    g03595(.A1(new_n5889_), .A2(new_n6045_), .ZN(new_n6046_));
  OAI21_X1   g03596(.A1(new_n5895_), .A2(new_n6046_), .B(new_n5897_), .ZN(new_n6047_));
  NOR2_X1    g03597(.A1(pi0299), .A2(pi0960), .ZN(new_n6048_));
  NAND2_X1   g03598(.A1(new_n5900_), .A2(new_n6048_), .ZN(new_n6049_));
  NAND2_X1   g03599(.A1(new_n6049_), .A2(pi0228), .ZN(new_n6050_));
  NOR2_X1    g03600(.A1(new_n5912_), .A2(pi0977), .ZN(new_n6051_));
  AOI21_X1   g03601(.A1(new_n5908_), .A2(pi0977), .B(pi0299), .ZN(new_n6052_));
  NAND2_X1   g03602(.A1(new_n6050_), .A2(new_n5915_), .ZN(new_n6053_));
  OAI22_X1   g03603(.A1(new_n5911_), .A2(new_n6051_), .B1(new_n6052_), .B2(new_n6053_), .ZN(new_n6054_));
  NAND4_X1   g03604(.A1(new_n6054_), .A2(new_n6047_), .A3(new_n5918_), .A4(new_n6050_), .ZN(new_n6055_));
  AOI21_X1   g03605(.A1(new_n5922_), .A2(pi0960), .B(new_n5924_), .ZN(new_n6056_));
  NOR3_X1    g03606(.A1(new_n5927_), .A2(new_n5390_), .A3(new_n6056_), .ZN(new_n6057_));
  OAI21_X1   g03607(.A1(new_n3211_), .A2(pi0960), .B(pi0299), .ZN(new_n6058_));
  OAI21_X1   g03608(.A1(new_n5938_), .A2(new_n6058_), .B(new_n5390_), .ZN(new_n6059_));
  AOI21_X1   g03609(.A1(new_n6059_), .A2(new_n5935_), .B(pi0100), .ZN(new_n6060_));
  NAND2_X1   g03610(.A1(new_n5888_), .A2(new_n6045_), .ZN(new_n6061_));
  XOR2_X1    g03611(.A1(new_n5943_), .A2(new_n6061_), .Z(new_n6062_));
  NAND2_X1   g03612(.A1(new_n6062_), .A2(pi0977), .ZN(new_n6063_));
  INV_X1     g03613(.I(new_n6063_), .ZN(new_n6064_));
  NAND2_X1   g03614(.A1(new_n6064_), .A2(new_n3211_), .ZN(new_n6065_));
  OAI21_X1   g03615(.A1(new_n6060_), .A2(new_n6065_), .B(new_n3455_), .ZN(new_n6066_));
  OAI21_X1   g03616(.A1(new_n5952_), .A2(new_n5390_), .B(new_n3098_), .ZN(new_n6067_));
  NOR2_X1    g03617(.A1(new_n6046_), .A2(new_n3098_), .ZN(new_n6068_));
  NOR2_X1    g03618(.A1(new_n5956_), .A2(new_n6045_), .ZN(new_n6069_));
  NAND2_X1   g03619(.A1(new_n6069_), .A2(new_n6068_), .ZN(new_n6070_));
  AOI21_X1   g03620(.A1(new_n6067_), .A2(new_n3183_), .B(new_n6070_), .ZN(new_n6071_));
  NOR2_X1    g03621(.A1(new_n6063_), .A2(new_n3183_), .ZN(new_n6072_));
  OAI21_X1   g03622(.A1(new_n6071_), .A2(pi0038), .B(new_n6072_), .ZN(new_n6073_));
  NAND3_X1   g03623(.A1(new_n6066_), .A2(pi0100), .A3(new_n6073_), .ZN(new_n6074_));
  AOI21_X1   g03624(.A1(new_n6055_), .A2(new_n6057_), .B(new_n6074_), .ZN(new_n6075_));
  NOR2_X1    g03625(.A1(new_n6063_), .A2(new_n3455_), .ZN(new_n6076_));
  OAI21_X1   g03626(.A1(new_n6075_), .A2(pi0075), .B(new_n6076_), .ZN(new_n6077_));
  AOI21_X1   g03627(.A1(new_n6071_), .A2(new_n6064_), .B(new_n5868_), .ZN(new_n6078_));
  NAND2_X1   g03628(.A1(new_n6078_), .A2(pi0092), .ZN(new_n6079_));
  XNOR2_X1   g03629(.A1(new_n6079_), .A2(new_n3483_), .ZN(new_n6080_));
  NOR2_X1    g03630(.A1(new_n6080_), .A2(new_n6063_), .ZN(new_n6081_));
  NAND2_X1   g03631(.A1(new_n3115_), .A2(pi0074), .ZN(new_n6082_));
  NOR2_X1    g03632(.A1(new_n6078_), .A2(new_n3235_), .ZN(new_n6083_));
  OAI21_X1   g03633(.A1(new_n6081_), .A2(new_n6082_), .B(new_n6083_), .ZN(new_n6084_));
  AOI21_X1   g03634(.A1(new_n6077_), .A2(new_n3303_), .B(new_n6084_), .ZN(new_n6085_));
  INV_X1     g03635(.I(new_n6046_), .ZN(new_n6086_));
  AOI21_X1   g03636(.A1(new_n6069_), .A2(new_n3291_), .B(new_n5976_), .ZN(new_n6087_));
  OAI21_X1   g03637(.A1(new_n6087_), .A2(new_n6086_), .B(new_n3258_), .ZN(new_n6088_));
  NAND2_X1   g03638(.A1(new_n6063_), .A2(new_n5769_), .ZN(new_n6089_));
  AOI21_X1   g03639(.A1(new_n6089_), .A2(pi0074), .B(new_n3188_), .ZN(new_n6090_));
  AOI21_X1   g03640(.A1(new_n6078_), .A2(new_n6090_), .B(new_n3115_), .ZN(new_n6091_));
  OAI21_X1   g03641(.A1(new_n6085_), .A2(new_n6088_), .B(new_n6091_), .ZN(new_n6092_));
  NAND2_X1   g03642(.A1(new_n6092_), .A2(new_n3229_), .ZN(new_n6093_));
  NOR2_X1    g03643(.A1(new_n6086_), .A2(new_n3226_), .ZN(new_n6094_));
  AOI21_X1   g03644(.A1(new_n6093_), .A2(new_n6094_), .B(new_n5371_), .ZN(new_n6095_));
  NAND2_X1   g03645(.A1(new_n6069_), .A2(new_n3291_), .ZN(new_n6096_));
  NAND3_X1   g03646(.A1(new_n6086_), .A2(pi0059), .A3(new_n5987_), .ZN(new_n6097_));
  NOR3_X1    g03647(.A1(new_n6096_), .A2(new_n5787_), .A3(new_n6097_), .ZN(new_n6098_));
  XOR2_X1    g03648(.A1(new_n6095_), .A2(new_n6098_), .Z(po0175));
  INV_X1     g03649(.I(pi0963), .ZN(new_n6100_));
  NOR2_X1    g03650(.A1(new_n5889_), .A2(new_n6100_), .ZN(new_n6101_));
  OAI21_X1   g03651(.A1(new_n5895_), .A2(new_n6101_), .B(new_n5897_), .ZN(new_n6102_));
  NOR2_X1    g03652(.A1(pi0299), .A2(pi0963), .ZN(new_n6103_));
  NAND2_X1   g03653(.A1(new_n5900_), .A2(new_n6103_), .ZN(new_n6104_));
  NAND2_X1   g03654(.A1(new_n6104_), .A2(pi0228), .ZN(new_n6105_));
  NOR2_X1    g03655(.A1(new_n5912_), .A2(pi0969), .ZN(new_n6106_));
  AOI21_X1   g03656(.A1(new_n5908_), .A2(pi0969), .B(pi0299), .ZN(new_n6107_));
  NAND2_X1   g03657(.A1(new_n6105_), .A2(new_n5915_), .ZN(new_n6108_));
  OAI22_X1   g03658(.A1(new_n5911_), .A2(new_n6106_), .B1(new_n6107_), .B2(new_n6108_), .ZN(new_n6109_));
  NAND4_X1   g03659(.A1(new_n6109_), .A2(new_n6102_), .A3(new_n5918_), .A4(new_n6105_), .ZN(new_n6110_));
  AOI21_X1   g03660(.A1(new_n5922_), .A2(pi0963), .B(new_n5924_), .ZN(new_n6111_));
  NOR3_X1    g03661(.A1(new_n5927_), .A2(new_n5387_), .A3(new_n6111_), .ZN(new_n6112_));
  OAI21_X1   g03662(.A1(new_n3211_), .A2(pi0963), .B(pi0299), .ZN(new_n6113_));
  OAI21_X1   g03663(.A1(new_n5938_), .A2(new_n6113_), .B(new_n5387_), .ZN(new_n6114_));
  AOI21_X1   g03664(.A1(new_n6114_), .A2(new_n5935_), .B(pi0100), .ZN(new_n6115_));
  NAND2_X1   g03665(.A1(new_n5888_), .A2(new_n6100_), .ZN(new_n6116_));
  XOR2_X1    g03666(.A1(new_n5943_), .A2(new_n6116_), .Z(new_n6117_));
  NAND2_X1   g03667(.A1(new_n6117_), .A2(pi0969), .ZN(new_n6118_));
  INV_X1     g03668(.I(new_n6118_), .ZN(new_n6119_));
  NAND2_X1   g03669(.A1(new_n6119_), .A2(new_n3211_), .ZN(new_n6120_));
  OAI21_X1   g03670(.A1(new_n6115_), .A2(new_n6120_), .B(new_n3455_), .ZN(new_n6121_));
  OAI21_X1   g03671(.A1(new_n5952_), .A2(new_n5387_), .B(new_n3098_), .ZN(new_n6122_));
  NOR2_X1    g03672(.A1(new_n6101_), .A2(new_n3098_), .ZN(new_n6123_));
  NOR2_X1    g03673(.A1(new_n5956_), .A2(new_n6100_), .ZN(new_n6124_));
  NAND2_X1   g03674(.A1(new_n6124_), .A2(new_n6123_), .ZN(new_n6125_));
  AOI21_X1   g03675(.A1(new_n6122_), .A2(new_n3183_), .B(new_n6125_), .ZN(new_n6126_));
  NOR2_X1    g03676(.A1(new_n6118_), .A2(new_n3183_), .ZN(new_n6127_));
  OAI21_X1   g03677(.A1(new_n6126_), .A2(pi0038), .B(new_n6127_), .ZN(new_n6128_));
  NAND3_X1   g03678(.A1(new_n6121_), .A2(pi0100), .A3(new_n6128_), .ZN(new_n6129_));
  AOI21_X1   g03679(.A1(new_n6110_), .A2(new_n6112_), .B(new_n6129_), .ZN(new_n6130_));
  NOR2_X1    g03680(.A1(new_n6118_), .A2(new_n3455_), .ZN(new_n6131_));
  OAI21_X1   g03681(.A1(new_n6130_), .A2(pi0075), .B(new_n6131_), .ZN(new_n6132_));
  AOI21_X1   g03682(.A1(new_n6126_), .A2(new_n6119_), .B(new_n5868_), .ZN(new_n6133_));
  NAND2_X1   g03683(.A1(new_n6133_), .A2(pi0092), .ZN(new_n6134_));
  XNOR2_X1   g03684(.A1(new_n6134_), .A2(new_n3483_), .ZN(new_n6135_));
  NOR2_X1    g03685(.A1(new_n6135_), .A2(new_n6118_), .ZN(new_n6136_));
  NAND2_X1   g03686(.A1(new_n3115_), .A2(pi0074), .ZN(new_n6137_));
  NOR2_X1    g03687(.A1(new_n6133_), .A2(new_n3235_), .ZN(new_n6138_));
  OAI21_X1   g03688(.A1(new_n6136_), .A2(new_n6137_), .B(new_n6138_), .ZN(new_n6139_));
  AOI21_X1   g03689(.A1(new_n6132_), .A2(new_n3303_), .B(new_n6139_), .ZN(new_n6140_));
  INV_X1     g03690(.I(new_n6101_), .ZN(new_n6141_));
  AOI21_X1   g03691(.A1(new_n6124_), .A2(new_n3291_), .B(new_n5976_), .ZN(new_n6142_));
  OAI21_X1   g03692(.A1(new_n6142_), .A2(new_n6141_), .B(new_n3258_), .ZN(new_n6143_));
  NAND2_X1   g03693(.A1(new_n6118_), .A2(new_n5769_), .ZN(new_n6144_));
  AOI21_X1   g03694(.A1(new_n6144_), .A2(pi0074), .B(new_n3188_), .ZN(new_n6145_));
  AOI21_X1   g03695(.A1(new_n6133_), .A2(new_n6145_), .B(new_n3115_), .ZN(new_n6146_));
  OAI21_X1   g03696(.A1(new_n6140_), .A2(new_n6143_), .B(new_n6146_), .ZN(new_n6147_));
  NAND2_X1   g03697(.A1(new_n6147_), .A2(new_n3229_), .ZN(new_n6148_));
  NOR2_X1    g03698(.A1(new_n6141_), .A2(new_n3226_), .ZN(new_n6149_));
  AOI21_X1   g03699(.A1(new_n6148_), .A2(new_n6149_), .B(new_n5371_), .ZN(new_n6150_));
  NAND2_X1   g03700(.A1(new_n6124_), .A2(new_n3291_), .ZN(new_n6151_));
  NAND3_X1   g03701(.A1(new_n6141_), .A2(pi0059), .A3(new_n5987_), .ZN(new_n6152_));
  NOR3_X1    g03702(.A1(new_n6151_), .A2(new_n5787_), .A3(new_n6152_), .ZN(new_n6153_));
  XOR2_X1    g03703(.A1(new_n6150_), .A2(new_n6153_), .Z(po0176));
  NOR2_X1    g03704(.A1(new_n5889_), .A2(new_n5448_), .ZN(new_n6155_));
  OAI21_X1   g03705(.A1(new_n5895_), .A2(new_n6155_), .B(new_n5897_), .ZN(new_n6156_));
  NOR2_X1    g03706(.A1(pi0299), .A2(pi0975), .ZN(new_n6157_));
  NAND2_X1   g03707(.A1(new_n5900_), .A2(new_n6157_), .ZN(new_n6158_));
  NAND2_X1   g03708(.A1(new_n6158_), .A2(pi0228), .ZN(new_n6159_));
  NOR2_X1    g03709(.A1(new_n5912_), .A2(pi0971), .ZN(new_n6160_));
  AOI21_X1   g03710(.A1(new_n5908_), .A2(pi0971), .B(pi0299), .ZN(new_n6161_));
  NAND2_X1   g03711(.A1(new_n6159_), .A2(new_n5915_), .ZN(new_n6162_));
  OAI22_X1   g03712(.A1(new_n5911_), .A2(new_n6160_), .B1(new_n6161_), .B2(new_n6162_), .ZN(new_n6163_));
  NAND4_X1   g03713(.A1(new_n6163_), .A2(new_n6156_), .A3(new_n5918_), .A4(new_n6159_), .ZN(new_n6164_));
  AOI21_X1   g03714(.A1(new_n5922_), .A2(pi0975), .B(new_n5924_), .ZN(new_n6165_));
  NOR3_X1    g03715(.A1(new_n5927_), .A2(new_n5388_), .A3(new_n6165_), .ZN(new_n6166_));
  OAI21_X1   g03716(.A1(new_n3211_), .A2(pi0975), .B(pi0299), .ZN(new_n6167_));
  OAI21_X1   g03717(.A1(new_n5938_), .A2(new_n6167_), .B(new_n5388_), .ZN(new_n6168_));
  AOI21_X1   g03718(.A1(new_n6168_), .A2(new_n5935_), .B(pi0100), .ZN(new_n6169_));
  NAND2_X1   g03719(.A1(new_n5888_), .A2(new_n5448_), .ZN(new_n6170_));
  XOR2_X1    g03720(.A1(new_n5943_), .A2(new_n6170_), .Z(new_n6171_));
  NAND2_X1   g03721(.A1(new_n6171_), .A2(pi0971), .ZN(new_n6172_));
  INV_X1     g03722(.I(new_n6172_), .ZN(new_n6173_));
  NAND2_X1   g03723(.A1(new_n6173_), .A2(new_n3211_), .ZN(new_n6174_));
  OAI21_X1   g03724(.A1(new_n6169_), .A2(new_n6174_), .B(new_n3455_), .ZN(new_n6175_));
  OAI21_X1   g03725(.A1(new_n5952_), .A2(new_n5388_), .B(new_n3098_), .ZN(new_n6176_));
  NOR2_X1    g03726(.A1(new_n6155_), .A2(new_n3098_), .ZN(new_n6177_));
  NOR2_X1    g03727(.A1(new_n5956_), .A2(new_n5448_), .ZN(new_n6178_));
  NAND2_X1   g03728(.A1(new_n6178_), .A2(new_n6177_), .ZN(new_n6179_));
  AOI21_X1   g03729(.A1(new_n6176_), .A2(new_n3183_), .B(new_n6179_), .ZN(new_n6180_));
  NOR2_X1    g03730(.A1(new_n6172_), .A2(new_n3183_), .ZN(new_n6181_));
  OAI21_X1   g03731(.A1(new_n6180_), .A2(pi0038), .B(new_n6181_), .ZN(new_n6182_));
  NAND3_X1   g03732(.A1(new_n6175_), .A2(pi0100), .A3(new_n6182_), .ZN(new_n6183_));
  AOI21_X1   g03733(.A1(new_n6164_), .A2(new_n6166_), .B(new_n6183_), .ZN(new_n6184_));
  NOR2_X1    g03734(.A1(new_n6172_), .A2(new_n3455_), .ZN(new_n6185_));
  OAI21_X1   g03735(.A1(new_n6184_), .A2(pi0075), .B(new_n6185_), .ZN(new_n6186_));
  AOI21_X1   g03736(.A1(new_n6180_), .A2(new_n6173_), .B(new_n5868_), .ZN(new_n6187_));
  NAND2_X1   g03737(.A1(new_n6187_), .A2(pi0092), .ZN(new_n6188_));
  XNOR2_X1   g03738(.A1(new_n6188_), .A2(new_n3483_), .ZN(new_n6189_));
  NOR2_X1    g03739(.A1(new_n6189_), .A2(new_n6172_), .ZN(new_n6190_));
  NAND2_X1   g03740(.A1(new_n3115_), .A2(pi0074), .ZN(new_n6191_));
  NOR2_X1    g03741(.A1(new_n6187_), .A2(new_n3235_), .ZN(new_n6192_));
  OAI21_X1   g03742(.A1(new_n6190_), .A2(new_n6191_), .B(new_n6192_), .ZN(new_n6193_));
  AOI21_X1   g03743(.A1(new_n6186_), .A2(new_n3303_), .B(new_n6193_), .ZN(new_n6194_));
  INV_X1     g03744(.I(new_n6155_), .ZN(new_n6195_));
  AOI21_X1   g03745(.A1(new_n6178_), .A2(new_n3291_), .B(new_n5976_), .ZN(new_n6196_));
  OAI21_X1   g03746(.A1(new_n6196_), .A2(new_n6195_), .B(new_n3258_), .ZN(new_n6197_));
  NAND2_X1   g03747(.A1(new_n6172_), .A2(new_n5769_), .ZN(new_n6198_));
  AOI21_X1   g03748(.A1(new_n6198_), .A2(pi0074), .B(new_n3188_), .ZN(new_n6199_));
  AOI21_X1   g03749(.A1(new_n6187_), .A2(new_n6199_), .B(new_n3115_), .ZN(new_n6200_));
  OAI21_X1   g03750(.A1(new_n6194_), .A2(new_n6197_), .B(new_n6200_), .ZN(new_n6201_));
  NAND2_X1   g03751(.A1(new_n6201_), .A2(new_n3229_), .ZN(new_n6202_));
  NOR2_X1    g03752(.A1(new_n6195_), .A2(new_n3226_), .ZN(new_n6203_));
  AOI21_X1   g03753(.A1(new_n6202_), .A2(new_n6203_), .B(new_n5371_), .ZN(new_n6204_));
  NAND2_X1   g03754(.A1(new_n6178_), .A2(new_n3291_), .ZN(new_n6205_));
  NAND3_X1   g03755(.A1(new_n6195_), .A2(pi0059), .A3(new_n5987_), .ZN(new_n6206_));
  NOR3_X1    g03756(.A1(new_n6205_), .A2(new_n5787_), .A3(new_n6206_), .ZN(new_n6207_));
  XOR2_X1    g03757(.A1(new_n6204_), .A2(new_n6207_), .Z(po0177));
  INV_X1     g03758(.I(new_n5918_), .ZN(new_n6209_));
  INV_X1     g03759(.I(new_n5897_), .ZN(new_n6210_));
  NOR2_X1    g03760(.A1(new_n5889_), .A2(new_n5449_), .ZN(new_n6211_));
  INV_X1     g03761(.I(new_n6211_), .ZN(new_n6212_));
  AOI21_X1   g03762(.A1(new_n5894_), .A2(new_n6212_), .B(new_n6210_), .ZN(new_n6213_));
  NOR2_X1    g03763(.A1(pi0299), .A2(pi0978), .ZN(new_n6214_));
  AOI21_X1   g03764(.A1(new_n5900_), .A2(new_n6214_), .B(new_n3005_), .ZN(new_n6215_));
  INV_X1     g03765(.I(new_n5912_), .ZN(new_n6216_));
  NAND2_X1   g03766(.A1(new_n6216_), .A2(new_n5389_), .ZN(new_n6217_));
  OAI21_X1   g03767(.A1(new_n5909_), .A2(new_n5389_), .B(new_n3098_), .ZN(new_n6218_));
  NOR3_X1    g03768(.A1(new_n6215_), .A2(new_n3183_), .A3(pi0232), .ZN(new_n6219_));
  AOI22_X1   g03769(.A1(new_n5910_), .A2(new_n6217_), .B1(new_n6218_), .B2(new_n6219_), .ZN(new_n6220_));
  NOR4_X1    g03770(.A1(new_n6220_), .A2(new_n6209_), .A3(new_n6213_), .A4(new_n6215_), .ZN(new_n6221_));
  AOI21_X1   g03771(.A1(new_n5922_), .A2(pi0978), .B(new_n5924_), .ZN(new_n6222_));
  OR3_X2     g03772(.A1(new_n5927_), .A2(new_n5389_), .A3(new_n6222_), .Z(new_n6223_));
  NAND3_X1   g03773(.A1(new_n5888_), .A2(pi0299), .A3(pi0978), .ZN(new_n6224_));
  NAND3_X1   g03774(.A1(new_n5888_), .A2(new_n3098_), .A3(new_n5449_), .ZN(new_n6225_));
  AOI21_X1   g03775(.A1(new_n6224_), .A2(new_n6225_), .B(new_n5389_), .ZN(new_n6226_));
  INV_X1     g03776(.I(new_n6226_), .ZN(new_n6227_));
  NOR3_X1    g03777(.A1(new_n5952_), .A2(new_n3098_), .A3(new_n5449_), .ZN(new_n6228_));
  NOR3_X1    g03778(.A1(new_n5952_), .A2(pi0299), .A3(pi0978), .ZN(new_n6229_));
  OAI21_X1   g03779(.A1(new_n6228_), .A2(new_n6229_), .B(pi0974), .ZN(new_n6230_));
  NAND2_X1   g03780(.A1(new_n6230_), .A2(pi0038), .ZN(new_n6231_));
  XOR2_X1    g03781(.A1(new_n6231_), .A2(new_n3262_), .Z(new_n6232_));
  NOR2_X1    g03782(.A1(new_n6232_), .A2(new_n6227_), .ZN(new_n6233_));
  INV_X1     g03783(.I(new_n5938_), .ZN(new_n6234_));
  AOI21_X1   g03784(.A1(new_n3212_), .A2(new_n5449_), .B(new_n3098_), .ZN(new_n6235_));
  AOI21_X1   g03785(.A1(new_n6234_), .A2(new_n6235_), .B(pi0974), .ZN(new_n6236_));
  OAI21_X1   g03786(.A1(new_n6236_), .A2(new_n5934_), .B(new_n3462_), .ZN(new_n6237_));
  NOR2_X1    g03787(.A1(new_n6227_), .A2(new_n3212_), .ZN(new_n6238_));
  AOI21_X1   g03788(.A1(new_n6237_), .A2(new_n6238_), .B(pi0087), .ZN(new_n6239_));
  NOR3_X1    g03789(.A1(new_n6233_), .A2(new_n3462_), .A3(new_n6239_), .ZN(new_n6240_));
  OAI21_X1   g03790(.A1(new_n6221_), .A2(new_n6223_), .B(new_n6240_), .ZN(new_n6241_));
  NAND2_X1   g03791(.A1(new_n6226_), .A2(pi0087), .ZN(new_n6242_));
  AOI21_X1   g03792(.A1(new_n6241_), .A2(new_n3235_), .B(new_n6242_), .ZN(new_n6243_));
  AOI21_X1   g03793(.A1(new_n3005_), .A2(new_n3194_), .B(new_n6230_), .ZN(new_n6244_));
  NOR2_X1    g03794(.A1(new_n6244_), .A2(new_n3303_), .ZN(new_n6245_));
  XNOR2_X1   g03795(.A1(new_n6245_), .A2(new_n3483_), .ZN(new_n6246_));
  NAND2_X1   g03796(.A1(new_n6246_), .A2(new_n6226_), .ZN(new_n6247_));
  NOR2_X1    g03797(.A1(new_n3175_), .A2(pi0054), .ZN(new_n6248_));
  NAND2_X1   g03798(.A1(new_n6244_), .A2(pi0075), .ZN(new_n6249_));
  AOI21_X1   g03799(.A1(new_n6247_), .A2(new_n6248_), .B(new_n6249_), .ZN(new_n6250_));
  OAI21_X1   g03800(.A1(new_n6243_), .A2(pi0092), .B(new_n6250_), .ZN(new_n6251_));
  NAND4_X1   g03801(.A1(new_n5440_), .A2(pi0228), .A3(pi0978), .A4(new_n3291_), .ZN(new_n6252_));
  NAND2_X1   g03802(.A1(new_n6252_), .A2(new_n5975_), .ZN(new_n6253_));
  AOI21_X1   g03803(.A1(new_n6253_), .A2(new_n6211_), .B(pi0055), .ZN(new_n6254_));
  OAI21_X1   g03804(.A1(new_n6226_), .A2(new_n5765_), .B(pi0074), .ZN(new_n6255_));
  NAND3_X1   g03805(.A1(new_n6255_), .A2(new_n3115_), .A3(new_n3189_), .ZN(new_n6256_));
  NAND2_X1   g03806(.A1(new_n6244_), .A2(new_n6256_), .ZN(new_n6257_));
  AOI21_X1   g03807(.A1(new_n6251_), .A2(new_n6254_), .B(new_n6257_), .ZN(new_n6258_));
  NOR2_X1    g03808(.A1(new_n6212_), .A2(new_n3226_), .ZN(new_n6259_));
  OAI21_X1   g03809(.A1(new_n6258_), .A2(pi0059), .B(new_n6259_), .ZN(new_n6260_));
  NAND2_X1   g03810(.A1(new_n6260_), .A2(pi0057), .ZN(new_n6261_));
  NAND3_X1   g03811(.A1(new_n6212_), .A2(pi0059), .A3(new_n5987_), .ZN(new_n6262_));
  NOR3_X1    g03812(.A1(new_n6252_), .A2(new_n5787_), .A3(new_n6262_), .ZN(new_n6263_));
  XNOR2_X1   g03813(.A1(new_n6261_), .A2(new_n6263_), .ZN(po0178));
  INV_X1     g03814(.I(pi0954), .ZN(po1110));
  NAND2_X1   g03815(.A1(new_n5896_), .A2(pi0299), .ZN(new_n6266_));
  OAI21_X1   g03816(.A1(new_n5899_), .A2(new_n6266_), .B(new_n5551_), .ZN(new_n6267_));
  OAI21_X1   g03817(.A1(new_n5906_), .A2(new_n3098_), .B(new_n5646_), .ZN(new_n6268_));
  NOR4_X1    g03818(.A1(new_n5386_), .A2(new_n5661_), .A3(new_n5662_), .A4(new_n3098_), .ZN(new_n6269_));
  NAND4_X1   g03819(.A1(new_n5893_), .A2(new_n6267_), .A3(new_n6268_), .A4(new_n6269_), .ZN(new_n6270_));
  AOI21_X1   g03820(.A1(new_n6270_), .A2(new_n5646_), .B(new_n5614_), .ZN(new_n6271_));
  INV_X1     g03821(.I(new_n5400_), .ZN(new_n6272_));
  AOI21_X1   g03822(.A1(new_n5704_), .A2(new_n3097_), .B(new_n6272_), .ZN(new_n6273_));
  NAND2_X1   g03823(.A1(new_n5709_), .A2(new_n3098_), .ZN(new_n6274_));
  OAI21_X1   g03824(.A1(new_n6273_), .A2(new_n6274_), .B(new_n5461_), .ZN(new_n6275_));
  NAND2_X1   g03825(.A1(new_n6275_), .A2(new_n3183_), .ZN(new_n6276_));
  NOR2_X1    g03826(.A1(new_n5654_), .A2(new_n3098_), .ZN(new_n6277_));
  XOR2_X1    g03827(.A1(new_n6277_), .A2(new_n6216_), .Z(new_n6278_));
  NOR3_X1    g03828(.A1(new_n6278_), .A2(pi0038), .A3(new_n5906_), .ZN(new_n6279_));
  OAI21_X1   g03829(.A1(new_n6271_), .A2(new_n6276_), .B(new_n6279_), .ZN(new_n6280_));
  NAND2_X1   g03830(.A1(new_n5492_), .A2(pi0038), .ZN(new_n6281_));
  NAND3_X1   g03831(.A1(new_n6280_), .A2(new_n5541_), .A3(new_n6281_), .ZN(new_n6282_));
  NAND2_X1   g03832(.A1(new_n5541_), .A2(pi0100), .ZN(new_n6283_));
  XNOR2_X1   g03833(.A1(new_n6282_), .A2(new_n6283_), .ZN(new_n6284_));
  NOR2_X1    g03834(.A1(new_n5504_), .A2(pi0038), .ZN(new_n6285_));
  NOR2_X1    g03835(.A1(new_n5504_), .A2(new_n3187_), .ZN(new_n6286_));
  NOR2_X1    g03836(.A1(new_n6286_), .A2(new_n3235_), .ZN(new_n6287_));
  NOR3_X1    g03837(.A1(new_n5504_), .A2(new_n3133_), .A3(new_n3204_), .ZN(new_n6288_));
  NOR2_X1    g03838(.A1(new_n6288_), .A2(new_n3303_), .ZN(new_n6289_));
  NOR2_X1    g03839(.A1(new_n6289_), .A2(new_n6287_), .ZN(new_n6290_));
  INV_X1     g03840(.I(new_n6290_), .ZN(new_n6291_));
  OAI21_X1   g03841(.A1(new_n6291_), .A2(new_n3115_), .B(new_n3189_), .ZN(new_n6292_));
  NAND2_X1   g03842(.A1(new_n6292_), .A2(new_n6285_), .ZN(new_n6293_));
  OAI22_X1   g03843(.A1(new_n6284_), .A2(new_n6293_), .B1(new_n3175_), .B2(new_n5490_), .ZN(new_n6294_));
  NOR2_X1    g03844(.A1(new_n5488_), .A2(new_n3294_), .ZN(new_n6295_));
  OAI21_X1   g03845(.A1(new_n6295_), .A2(new_n3208_), .B(new_n3201_), .ZN(new_n6296_));
  AOI21_X1   g03846(.A1(new_n6288_), .A2(new_n3303_), .B(new_n3115_), .ZN(new_n6297_));
  NAND3_X1   g03847(.A1(new_n6296_), .A2(pi0055), .A3(new_n6297_), .ZN(new_n6298_));
  INV_X1     g03848(.I(new_n6298_), .ZN(new_n6299_));
  AOI21_X1   g03849(.A1(new_n6294_), .A2(new_n6299_), .B(new_n3426_), .ZN(new_n6300_));
  NOR2_X1    g03850(.A1(new_n6300_), .A2(new_n5548_), .ZN(po0195));
  NAND2_X1   g03851(.A1(po0195), .A2(po1110), .ZN(new_n6302_));
  OAI21_X1   g03852(.A1(pi0024), .A2(po1110), .B(new_n6302_), .ZN(po0182));
  AOI21_X1   g03853(.A1(new_n5723_), .A2(pi0252), .B(pi0299), .ZN(new_n6304_));
  AOI22_X1   g03854(.A1(new_n3400_), .A2(pi0299), .B1(new_n3160_), .B2(new_n6304_), .ZN(new_n6305_));
  INV_X1     g03855(.I(new_n6305_), .ZN(new_n6306_));
  NAND2_X1   g03856(.A1(new_n3183_), .A2(new_n3462_), .ZN(new_n6307_));
  OAI21_X1   g03857(.A1(new_n6306_), .A2(new_n6307_), .B(new_n3411_), .ZN(new_n6308_));
  NOR2_X1    g03858(.A1(new_n3412_), .A2(new_n3214_), .ZN(new_n6309_));
  INV_X1     g03859(.I(new_n6309_), .ZN(new_n6310_));
  AOI21_X1   g03860(.A1(new_n6310_), .A2(new_n3953_), .B(new_n3009_), .ZN(new_n6311_));
  NOR2_X1    g03861(.A1(new_n3412_), .A2(new_n3495_), .ZN(new_n6312_));
  NOR2_X1    g03862(.A1(new_n3203_), .A2(new_n3303_), .ZN(new_n6313_));
  NOR2_X1    g03863(.A1(new_n6312_), .A2(new_n6313_), .ZN(new_n6314_));
  NOR2_X1    g03864(.A1(new_n3006_), .A2(new_n3235_), .ZN(new_n6315_));
  NOR4_X1    g03865(.A1(new_n6314_), .A2(pi0092), .A3(new_n3009_), .A4(new_n6315_), .ZN(new_n6316_));
  NOR2_X1    g03866(.A1(new_n3411_), .A2(new_n3262_), .ZN(new_n6317_));
  NAND2_X1   g03867(.A1(new_n3006_), .A2(pi0087), .ZN(new_n6318_));
  AOI21_X1   g03868(.A1(new_n6317_), .A2(new_n6318_), .B(new_n3462_), .ZN(new_n6319_));
  OAI21_X1   g03869(.A1(new_n6316_), .A2(new_n6311_), .B(new_n6319_), .ZN(new_n6320_));
  AOI21_X1   g03870(.A1(new_n4359_), .A2(new_n6308_), .B(new_n6320_), .ZN(new_n6321_));
  NOR2_X1    g03871(.A1(new_n6321_), .A2(pi0055), .ZN(new_n6322_));
  NAND2_X1   g03872(.A1(new_n3006_), .A2(new_n3202_), .ZN(new_n6323_));
  OAI21_X1   g03873(.A1(new_n6322_), .A2(new_n6323_), .B(new_n3219_), .ZN(new_n6324_));
  NOR3_X1    g03874(.A1(new_n3206_), .A2(new_n3214_), .A3(pi0054), .ZN(new_n6325_));
  NOR2_X1    g03875(.A1(new_n6325_), .A2(new_n3006_), .ZN(new_n6326_));
  NOR2_X1    g03876(.A1(new_n3258_), .A2(new_n3175_), .ZN(new_n6327_));
  INV_X1     g03877(.I(new_n6327_), .ZN(new_n6328_));
  AOI21_X1   g03878(.A1(new_n3412_), .A2(new_n6326_), .B(new_n6328_), .ZN(new_n6329_));
  AOI21_X1   g03879(.A1(new_n6324_), .A2(new_n6329_), .B(new_n3201_), .ZN(new_n6330_));
  NOR2_X1    g03880(.A1(new_n6310_), .A2(new_n3431_), .ZN(new_n6331_));
  INV_X1     g03881(.I(new_n6331_), .ZN(new_n6332_));
  NOR2_X1    g03882(.A1(new_n3224_), .A2(new_n3412_), .ZN(new_n6333_));
  NOR3_X1    g03883(.A1(new_n3006_), .A2(new_n3219_), .A3(new_n3201_), .ZN(new_n6334_));
  NAND3_X1   g03884(.A1(new_n6332_), .A2(new_n6333_), .A3(new_n6334_), .ZN(new_n6335_));
  AND2_X2    g03885(.A1(new_n6330_), .A2(new_n6335_), .Z(new_n6336_));
  OAI21_X1   g03886(.A1(new_n6330_), .A2(new_n6335_), .B(new_n3230_), .ZN(new_n6337_));
  OAI22_X1   g03887(.A1(new_n6336_), .A2(new_n6337_), .B1(new_n3009_), .B2(new_n3230_), .ZN(po0183));
  NAND2_X1   g03888(.A1(pi0119), .A2(pi0468), .ZN(new_n6339_));
  AOI21_X1   g03889(.A1(new_n6339_), .A2(new_n3721_), .B(new_n3005_), .ZN(new_n6340_));
  NAND2_X1   g03890(.A1(pi0119), .A2(pi1056), .ZN(new_n6341_));
  NAND2_X1   g03891(.A1(new_n6340_), .A2(new_n6341_), .ZN(po0184));
  NAND2_X1   g03892(.A1(pi0119), .A2(pi1077), .ZN(new_n6343_));
  NAND2_X1   g03893(.A1(new_n6340_), .A2(new_n6343_), .ZN(po0185));
  NAND2_X1   g03894(.A1(pi0119), .A2(pi1073), .ZN(new_n6345_));
  NAND2_X1   g03895(.A1(new_n6340_), .A2(new_n6345_), .ZN(po0186));
  NAND2_X1   g03896(.A1(pi0119), .A2(pi1041), .ZN(new_n6347_));
  NAND2_X1   g03897(.A1(new_n6340_), .A2(new_n6347_), .ZN(po0187));
  INV_X1     g03898(.I(pi0031), .ZN(new_n6349_));
  INV_X1     g03899(.I(pi0591), .ZN(new_n6350_));
  INV_X1     g03900(.I(pi0461), .ZN(new_n6351_));
  NOR2_X1    g03901(.A1(new_n6351_), .A2(pi0357), .ZN(new_n6352_));
  NAND2_X1   g03902(.A1(new_n6351_), .A2(pi0357), .ZN(new_n6353_));
  INV_X1     g03903(.I(new_n6353_), .ZN(new_n6354_));
  INV_X1     g03904(.I(pi1199), .ZN(new_n6356_));
  INV_X1     g03905(.I(pi0592), .ZN(new_n6358_));
  NOR2_X1    g03906(.A1(new_n2721_), .A2(pi0122), .ZN(new_n6359_));
  INV_X1     g03907(.I(pi0088), .ZN(new_n6360_));
  NOR2_X1    g03908(.A1(pi0050), .A2(pi0077), .ZN(new_n6361_));
  NAND3_X1   g03909(.A1(new_n2557_), .A2(new_n2530_), .A3(new_n6361_), .ZN(new_n6362_));
  NOR4_X1    g03910(.A1(new_n6362_), .A2(new_n6360_), .A3(new_n2558_), .A4(new_n2460_), .ZN(new_n6363_));
  NOR2_X1    g03911(.A1(new_n6363_), .A2(pi0097), .ZN(new_n6364_));
  NOR2_X1    g03912(.A1(new_n6364_), .A2(new_n2903_), .ZN(new_n6365_));
  INV_X1     g03913(.I(new_n6365_), .ZN(new_n6366_));
  NOR2_X1    g03914(.A1(new_n2479_), .A2(pi0035), .ZN(new_n6367_));
  INV_X1     g03915(.I(new_n6367_), .ZN(new_n6368_));
  NOR2_X1    g03916(.A1(new_n6368_), .A2(pi0070), .ZN(new_n6369_));
  AOI21_X1   g03917(.A1(new_n2471_), .A2(new_n2478_), .B(new_n2732_), .ZN(new_n6370_));
  INV_X1     g03918(.I(new_n6370_), .ZN(new_n6371_));
  NAND2_X1   g03919(.A1(new_n5428_), .A2(new_n2698_), .ZN(new_n6372_));
  INV_X1     g03920(.I(new_n6372_), .ZN(new_n6373_));
  AOI21_X1   g03921(.A1(new_n6371_), .A2(new_n6373_), .B(pi0051), .ZN(new_n6374_));
  AOI21_X1   g03922(.A1(new_n6374_), .A2(new_n2712_), .B(new_n6369_), .ZN(new_n6375_));
  NOR2_X1    g03923(.A1(new_n6375_), .A2(new_n6366_), .ZN(new_n6376_));
  NOR2_X1    g03924(.A1(new_n6376_), .A2(pi0096), .ZN(new_n6377_));
  INV_X1     g03925(.I(new_n6359_), .ZN(new_n6378_));
  NOR2_X1    g03926(.A1(new_n2981_), .A2(new_n6378_), .ZN(new_n6379_));
  INV_X1     g03927(.I(new_n6379_), .ZN(new_n6380_));
  NOR4_X1    g03928(.A1(new_n2706_), .A2(new_n2509_), .A3(new_n2732_), .A4(new_n2678_), .ZN(new_n6381_));
  AOI21_X1   g03929(.A1(new_n6381_), .A2(new_n2795_), .B(new_n2755_), .ZN(new_n6382_));
  NOR2_X1    g03930(.A1(new_n6382_), .A2(new_n3304_), .ZN(new_n6383_));
  INV_X1     g03931(.I(new_n6383_), .ZN(new_n6384_));
  NOR3_X1    g03932(.A1(new_n6377_), .A2(new_n6380_), .A3(new_n6384_), .ZN(new_n6385_));
  NOR2_X1    g03933(.A1(new_n3304_), .A2(pi0096), .ZN(new_n6386_));
  NAND2_X1   g03934(.A1(new_n6376_), .A2(new_n6386_), .ZN(new_n6387_));
  INV_X1     g03935(.I(new_n6387_), .ZN(new_n6388_));
  OR3_X2     g03936(.A1(new_n6385_), .A2(new_n5532_), .A3(new_n6388_), .Z(new_n6389_));
  NAND2_X1   g03937(.A1(new_n6389_), .A2(new_n6359_), .ZN(new_n6390_));
  INV_X1     g03938(.I(new_n6390_), .ZN(new_n6391_));
  NOR2_X1    g03939(.A1(new_n6391_), .A2(pi1093), .ZN(new_n6392_));
  INV_X1     g03940(.I(new_n6392_), .ZN(new_n6393_));
  NAND2_X1   g03941(.A1(new_n3213_), .A2(new_n3235_), .ZN(new_n6394_));
  OAI21_X1   g03942(.A1(new_n3455_), .A2(new_n6394_), .B(new_n3145_), .ZN(new_n6395_));
  NAND3_X1   g03943(.A1(new_n6395_), .A2(pi0567), .A3(po0740), .ZN(new_n6396_));
  AOI21_X1   g03944(.A1(new_n3455_), .A2(new_n6396_), .B(new_n6393_), .ZN(new_n6397_));
  INV_X1     g03945(.I(new_n5499_), .ZN(new_n6398_));
  NOR2_X1    g03946(.A1(new_n6398_), .A2(pi0074), .ZN(new_n6399_));
  INV_X1     g03947(.I(new_n6399_), .ZN(new_n6400_));
  NOR2_X1    g03948(.A1(new_n6397_), .A2(new_n6400_), .ZN(new_n6401_));
  NOR2_X1    g03949(.A1(new_n2981_), .A2(new_n5683_), .ZN(new_n6402_));
  INV_X1     g03950(.I(new_n6402_), .ZN(new_n6403_));
  NOR2_X1    g03951(.A1(new_n2984_), .A2(pi0122), .ZN(new_n6404_));
  INV_X1     g03952(.I(new_n6404_), .ZN(new_n6405_));
  NOR2_X1    g03953(.A1(new_n6403_), .A2(new_n6405_), .ZN(new_n6406_));
  NAND2_X1   g03954(.A1(new_n6406_), .A2(new_n2726_), .ZN(new_n6407_));
  NOR2_X1    g03955(.A1(new_n6407_), .A2(pi0098), .ZN(new_n6408_));
  INV_X1     g03956(.I(new_n6408_), .ZN(new_n6409_));
  INV_X1     g03957(.I(pi0122), .ZN(new_n6410_));
  NOR2_X1    g03958(.A1(new_n2714_), .A2(new_n3304_), .ZN(new_n6411_));
  INV_X1     g03959(.I(new_n6411_), .ZN(new_n6412_));
  NOR2_X1    g03960(.A1(new_n6374_), .A2(new_n6412_), .ZN(new_n6413_));
  INV_X1     g03961(.I(new_n6413_), .ZN(new_n6414_));
  NOR2_X1    g03962(.A1(new_n6414_), .A2(new_n6403_), .ZN(new_n6415_));
  NOR2_X1    g03963(.A1(new_n6415_), .A2(new_n6410_), .ZN(new_n6416_));
  NOR2_X1    g03964(.A1(new_n6403_), .A2(pi0098), .ZN(new_n6417_));
  NOR2_X1    g03965(.A1(new_n6417_), .A2(pi0122), .ZN(new_n6418_));
  NOR2_X1    g03966(.A1(new_n6413_), .A2(new_n6410_), .ZN(new_n6419_));
  INV_X1     g03967(.I(new_n6419_), .ZN(new_n6420_));
  AOI21_X1   g03968(.A1(pi0096), .A2(new_n2712_), .B(new_n6374_), .ZN(new_n6421_));
  NOR2_X1    g03969(.A1(new_n2868_), .A2(pi0024), .ZN(new_n6422_));
  NAND4_X1   g03970(.A1(new_n5562_), .A2(pi0046), .A3(pi0097), .A4(pi0108), .ZN(new_n6423_));
  NOR2_X1    g03971(.A1(new_n2874_), .A2(new_n6423_), .ZN(new_n6424_));
  AOI21_X1   g03972(.A1(new_n2674_), .A2(new_n6424_), .B(new_n6422_), .ZN(new_n6425_));
  NOR4_X1    g03973(.A1(new_n6421_), .A2(new_n2678_), .A3(new_n6372_), .A4(new_n6425_), .ZN(new_n6426_));
  INV_X1     g03974(.I(new_n2982_), .ZN(new_n6427_));
  NOR2_X1    g03975(.A1(new_n6384_), .A2(new_n6427_), .ZN(new_n6428_));
  AOI22_X1   g03976(.A1(new_n6426_), .A2(new_n6415_), .B1(pi0829), .B2(new_n6428_), .ZN(new_n6429_));
  NOR3_X1    g03977(.A1(new_n6429_), .A2(new_n6410_), .A3(new_n5533_), .ZN(new_n6430_));
  NOR2_X1    g03978(.A1(new_n2728_), .A2(new_n2984_), .ZN(new_n6431_));
  INV_X1     g03979(.I(new_n6431_), .ZN(new_n6432_));
  AOI21_X1   g03980(.A1(new_n6430_), .A2(new_n6420_), .B(new_n6432_), .ZN(new_n6433_));
  OAI21_X1   g03981(.A1(new_n6420_), .A2(new_n6430_), .B(new_n6433_), .ZN(new_n6434_));
  NAND2_X1   g03982(.A1(new_n6434_), .A2(pi1091), .ZN(new_n6435_));
  NOR2_X1    g03983(.A1(new_n6435_), .A2(new_n6392_), .ZN(new_n6436_));
  NOR4_X1    g03984(.A1(new_n6436_), .A2(pi0039), .A3(pi1091), .A4(new_n6392_), .ZN(new_n6437_));
  OAI22_X1   g03985(.A1(new_n6437_), .A2(pi1093), .B1(new_n6416_), .B2(new_n6418_), .ZN(new_n6438_));
  NOR4_X1    g03986(.A1(new_n5681_), .A2(new_n2721_), .A3(new_n2722_), .A4(new_n2983_), .ZN(new_n6439_));
  OR2_X2     g03987(.A1(new_n6439_), .A2(new_n2726_), .Z(new_n6440_));
  INV_X1     g03988(.I(new_n6417_), .ZN(new_n6441_));
  NOR2_X1    g03989(.A1(new_n6441_), .A2(new_n6405_), .ZN(new_n6442_));
  NOR2_X1    g03990(.A1(new_n2723_), .A2(new_n2726_), .ZN(new_n6443_));
  NAND2_X1   g03991(.A1(new_n6442_), .A2(new_n6443_), .ZN(new_n6444_));
  XOR2_X1    g03992(.A1(new_n6440_), .A2(new_n6444_), .Z(new_n6445_));
  NOR2_X1    g03993(.A1(new_n6445_), .A2(new_n5434_), .ZN(new_n6446_));
  AOI21_X1   g03994(.A1(new_n5434_), .A2(new_n6409_), .B(new_n6446_), .ZN(new_n6447_));
  INV_X1     g03995(.I(new_n5385_), .ZN(new_n6448_));
  NOR2_X1    g03996(.A1(new_n6445_), .A2(new_n6448_), .ZN(new_n6449_));
  AOI21_X1   g03997(.A1(new_n6448_), .A2(new_n6409_), .B(new_n6449_), .ZN(new_n6450_));
  NOR2_X1    g03998(.A1(new_n3362_), .A2(pi0216), .ZN(new_n6451_));
  NAND2_X1   g03999(.A1(new_n6450_), .A2(new_n6451_), .ZN(new_n6452_));
  INV_X1     g04000(.I(new_n6451_), .ZN(new_n6453_));
  NOR2_X1    g04001(.A1(new_n5455_), .A2(new_n6453_), .ZN(new_n6454_));
  XOR2_X1    g04002(.A1(new_n6452_), .A2(new_n6454_), .Z(new_n6455_));
  OAI21_X1   g04003(.A1(new_n6455_), .A2(new_n6447_), .B(new_n3098_), .ZN(new_n6456_));
  NOR2_X1    g04004(.A1(new_n6409_), .A2(new_n6453_), .ZN(new_n6457_));
  AOI21_X1   g04005(.A1(new_n6456_), .A2(new_n6457_), .B(pi0039), .ZN(new_n6458_));
  NOR2_X1    g04006(.A1(new_n5139_), .A2(pi0223), .ZN(new_n6459_));
  NAND2_X1   g04007(.A1(new_n6450_), .A2(new_n6459_), .ZN(new_n6460_));
  INV_X1     g04008(.I(new_n6459_), .ZN(new_n6461_));
  NOR2_X1    g04009(.A1(new_n6461_), .A2(new_n5397_), .ZN(new_n6462_));
  XOR2_X1    g04010(.A1(new_n6460_), .A2(new_n6462_), .Z(new_n6463_));
  OAI21_X1   g04011(.A1(new_n6463_), .A2(new_n6447_), .B(new_n3098_), .ZN(new_n6464_));
  NAND3_X1   g04012(.A1(new_n6464_), .A2(new_n6408_), .A3(new_n6459_), .ZN(new_n6465_));
  AOI21_X1   g04013(.A1(new_n6438_), .A2(new_n6458_), .B(new_n6465_), .ZN(new_n6466_));
  NOR2_X1    g04014(.A1(new_n6466_), .A2(new_n3259_), .ZN(new_n6467_));
  XOR2_X1    g04015(.A1(new_n6467_), .A2(new_n5486_), .Z(new_n6468_));
  OAI21_X1   g04016(.A1(new_n6468_), .A2(new_n6409_), .B(new_n3455_), .ZN(new_n6469_));
  NOR2_X1    g04017(.A1(new_n3145_), .A2(new_n6403_), .ZN(new_n6470_));
  NOR2_X1    g04018(.A1(new_n6470_), .A2(new_n2984_), .ZN(new_n6471_));
  NOR2_X1    g04019(.A1(new_n6410_), .A2(new_n2984_), .ZN(new_n6472_));
  XNOR2_X1   g04020(.A1(new_n6471_), .A2(new_n6472_), .ZN(new_n6473_));
  NOR2_X1    g04021(.A1(new_n2983_), .A2(new_n2984_), .ZN(new_n6474_));
  INV_X1     g04022(.I(new_n6474_), .ZN(new_n6475_));
  NOR2_X1    g04023(.A1(new_n3160_), .A2(new_n5532_), .ZN(new_n6476_));
  AOI21_X1   g04024(.A1(new_n6476_), .A2(new_n2726_), .B(new_n6475_), .ZN(new_n6477_));
  NOR2_X1    g04025(.A1(new_n6477_), .A2(new_n3134_), .ZN(new_n6478_));
  AOI21_X1   g04026(.A1(new_n3160_), .A2(po0740), .B(pi1091), .ZN(new_n6479_));
  INV_X1     g04027(.I(new_n6479_), .ZN(new_n6480_));
  NOR4_X1    g04028(.A1(new_n6473_), .A2(new_n6441_), .A3(new_n6478_), .A4(new_n6480_), .ZN(new_n6481_));
  OAI21_X1   g04029(.A1(new_n6481_), .A2(new_n3694_), .B(new_n6408_), .ZN(new_n6482_));
  NOR2_X1    g04030(.A1(new_n5526_), .A2(new_n2728_), .ZN(new_n6483_));
  INV_X1     g04031(.I(new_n6483_), .ZN(new_n6484_));
  NOR3_X1    g04032(.A1(new_n3145_), .A2(pi0024), .A3(new_n3721_), .ZN(new_n6485_));
  NOR2_X1    g04033(.A1(new_n6380_), .A2(new_n2984_), .ZN(new_n6486_));
  NOR3_X1    g04034(.A1(new_n6485_), .A2(pi1091), .A3(new_n6486_), .ZN(new_n6487_));
  NOR2_X1    g04035(.A1(new_n6484_), .A2(new_n6487_), .ZN(new_n6488_));
  NOR2_X1    g04036(.A1(new_n2787_), .A2(new_n3098_), .ZN(new_n6489_));
  NOR2_X1    g04037(.A1(new_n3079_), .A2(pi0299), .ZN(new_n6490_));
  NOR2_X1    g04038(.A1(new_n6489_), .A2(new_n6490_), .ZN(new_n6491_));
  INV_X1     g04039(.I(new_n6491_), .ZN(new_n6492_));
  NOR2_X1    g04040(.A1(new_n5386_), .A2(new_n5551_), .ZN(new_n6493_));
  INV_X1     g04041(.I(new_n6493_), .ZN(new_n6494_));
  NOR2_X1    g04042(.A1(new_n6492_), .A2(new_n6494_), .ZN(new_n6495_));
  NOR2_X1    g04043(.A1(new_n6495_), .A2(new_n3194_), .ZN(new_n6496_));
  INV_X1     g04044(.I(new_n6496_), .ZN(new_n6497_));
  NOR2_X1    g04045(.A1(new_n6488_), .A2(new_n6497_), .ZN(new_n6498_));
  INV_X1     g04046(.I(new_n6498_), .ZN(new_n6499_));
  OAI21_X1   g04047(.A1(new_n6409_), .A2(new_n6496_), .B(pi0075), .ZN(new_n6500_));
  OAI21_X1   g04048(.A1(new_n6499_), .A2(new_n6500_), .B(new_n2726_), .ZN(new_n6501_));
  NAND3_X1   g04049(.A1(new_n6501_), .A2(pi0567), .A3(new_n6442_), .ZN(new_n6502_));
  NAND2_X1   g04050(.A1(new_n6502_), .A2(new_n6482_), .ZN(new_n6503_));
  INV_X1     g04051(.I(new_n6486_), .ZN(new_n6504_));
  NOR2_X1    g04052(.A1(new_n6484_), .A2(new_n6504_), .ZN(new_n6505_));
  NAND2_X1   g04053(.A1(new_n6505_), .A2(new_n3160_), .ZN(new_n6506_));
  NOR2_X1    g04054(.A1(new_n6506_), .A2(new_n2726_), .ZN(new_n6507_));
  INV_X1     g04055(.I(new_n6442_), .ZN(new_n6508_));
  NOR2_X1    g04056(.A1(new_n6508_), .A2(pi1091), .ZN(new_n6509_));
  NOR3_X1    g04057(.A1(new_n6507_), .A2(new_n3212_), .A3(new_n6509_), .ZN(new_n6510_));
  NOR2_X1    g04058(.A1(new_n6495_), .A2(new_n3005_), .ZN(new_n6511_));
  NAND2_X1   g04059(.A1(new_n6511_), .A2(new_n3211_), .ZN(new_n6512_));
  XNOR2_X1   g04060(.A1(new_n6510_), .A2(new_n6512_), .ZN(new_n6513_));
  INV_X1     g04061(.I(pi0567), .ZN(new_n6514_));
  NAND2_X1   g04062(.A1(new_n6399_), .A2(pi0100), .ZN(new_n6515_));
  NOR4_X1    g04063(.A1(new_n6409_), .A2(new_n6514_), .A3(new_n3212_), .A4(new_n6515_), .ZN(new_n6516_));
  NAND4_X1   g04064(.A1(new_n6469_), .A2(new_n6503_), .A3(new_n6513_), .A4(new_n6516_), .ZN(new_n6517_));
  OR2_X2     g04065(.A1(new_n6517_), .A2(new_n6401_), .Z(new_n6518_));
  NAND2_X1   g04066(.A1(new_n6517_), .A2(new_n6401_), .ZN(new_n6519_));
  NAND2_X1   g04067(.A1(new_n6518_), .A2(new_n6519_), .ZN(new_n6520_));
  INV_X1     g04068(.I(new_n6520_), .ZN(new_n6521_));
  NOR2_X1    g04069(.A1(new_n6521_), .A2(new_n6358_), .ZN(new_n6522_));
  INV_X1     g04070(.I(new_n6485_), .ZN(new_n6523_));
  NOR3_X1    g04071(.A1(new_n6484_), .A2(new_n2726_), .A3(new_n6380_), .ZN(new_n6524_));
  INV_X1     g04072(.I(new_n6524_), .ZN(new_n6525_));
  NOR2_X1    g04073(.A1(new_n6525_), .A2(new_n6523_), .ZN(new_n6526_));
  INV_X1     g04074(.I(new_n6526_), .ZN(new_n6527_));
  NOR2_X1    g04075(.A1(new_n6527_), .A2(new_n2984_), .ZN(new_n6528_));
  AOI21_X1   g04076(.A1(new_n6528_), .A2(new_n6496_), .B(new_n3235_), .ZN(new_n6529_));
  INV_X1     g04077(.I(new_n6401_), .ZN(new_n6530_));
  INV_X1     g04078(.I(new_n6495_), .ZN(new_n6531_));
  INV_X1     g04079(.I(new_n6507_), .ZN(new_n6532_));
  NAND3_X1   g04080(.A1(new_n6532_), .A2(new_n3462_), .A3(new_n3005_), .ZN(new_n6533_));
  NAND3_X1   g04081(.A1(new_n6533_), .A2(new_n3211_), .A3(new_n6531_), .ZN(new_n6534_));
  NAND2_X1   g04082(.A1(new_n6534_), .A2(new_n3455_), .ZN(new_n6535_));
  NOR2_X1    g04083(.A1(new_n6392_), .A2(pi1091), .ZN(new_n6536_));
  NAND2_X1   g04084(.A1(new_n6439_), .A2(new_n6443_), .ZN(new_n6537_));
  NOR2_X1    g04085(.A1(new_n6537_), .A2(new_n5461_), .ZN(new_n6538_));
  INV_X1     g04086(.I(new_n6538_), .ZN(new_n6539_));
  INV_X1     g04087(.I(new_n5825_), .ZN(new_n6540_));
  NOR2_X1    g04088(.A1(new_n6540_), .A2(pi0216), .ZN(new_n6541_));
  NOR2_X1    g04089(.A1(new_n6537_), .A2(new_n5400_), .ZN(new_n6542_));
  INV_X1     g04090(.I(new_n6542_), .ZN(new_n6543_));
  INV_X1     g04091(.I(new_n5700_), .ZN(new_n6544_));
  NOR2_X1    g04092(.A1(new_n6544_), .A2(pi0299), .ZN(new_n6545_));
  NOR2_X1    g04093(.A1(new_n6545_), .A2(pi0039), .ZN(new_n6546_));
  NAND2_X1   g04094(.A1(new_n6543_), .A2(new_n6546_), .ZN(new_n6547_));
  NOR2_X1    g04095(.A1(new_n3259_), .A2(new_n3100_), .ZN(new_n6548_));
  AOI21_X1   g04096(.A1(new_n6547_), .A2(new_n6548_), .B(new_n6541_), .ZN(new_n6549_));
  NOR2_X1    g04097(.A1(new_n6549_), .A2(new_n6539_), .ZN(new_n6550_));
  INV_X1     g04098(.I(new_n6550_), .ZN(new_n6551_));
  OAI22_X1   g04099(.A1(new_n6435_), .A2(new_n6392_), .B1(new_n3183_), .B2(new_n6551_), .ZN(new_n6552_));
  AOI21_X1   g04100(.A1(new_n6552_), .A2(new_n6536_), .B(pi0100), .ZN(new_n6553_));
  NOR3_X1    g04101(.A1(new_n3212_), .A2(new_n3455_), .A3(pi0100), .ZN(new_n6554_));
  NOR3_X1    g04102(.A1(new_n6477_), .A2(pi0075), .A3(new_n6554_), .ZN(new_n6555_));
  NOR2_X1    g04103(.A1(new_n6555_), .A2(new_n6480_), .ZN(new_n6556_));
  OAI21_X1   g04104(.A1(new_n6553_), .A2(new_n6535_), .B(new_n6556_), .ZN(new_n6557_));
  OAI21_X1   g04105(.A1(new_n6530_), .A2(new_n6514_), .B(new_n6557_), .ZN(new_n6558_));
  NAND2_X1   g04106(.A1(new_n6558_), .A2(new_n6529_), .ZN(new_n6559_));
  INV_X1     g04107(.I(new_n6559_), .ZN(new_n6560_));
  NOR2_X1    g04108(.A1(new_n6560_), .A2(pi0592), .ZN(new_n6561_));
  NOR2_X1    g04109(.A1(new_n6522_), .A2(new_n6561_), .ZN(new_n6562_));
  INV_X1     g04110(.I(pi1198), .ZN(new_n6577_));
  INV_X1     g04111(.I(pi0342), .ZN(new_n6581_));
  INV_X1     g04112(.I(pi0320), .ZN(new_n6584_));
  INV_X1     g04113(.I(pi1196), .ZN(new_n6595_));
  INV_X1     g04114(.I(pi0452), .ZN(new_n6596_));
  INV_X1     g04115(.I(pi0348), .ZN(new_n6604_));
  INV_X1     g04116(.I(pi0322), .ZN(new_n6606_));
  NOR2_X1    g04117(.A1(new_n6521_), .A2(pi1196), .ZN(new_n6643_));
  NOR2_X1    g04118(.A1(new_n6354_), .A2(new_n6352_), .ZN(new_n6648_));
  NOR2_X1    g04119(.A1(new_n6648_), .A2(pi0356), .ZN(new_n6649_));
  INV_X1     g04120(.I(pi0356), .ZN(new_n6650_));
  NOR2_X1    g04121(.A1(new_n6648_), .A2(new_n6650_), .ZN(new_n6651_));
  NOR2_X1    g04122(.A1(new_n6649_), .A2(new_n6651_), .ZN(new_n6652_));
  INV_X1     g04123(.I(pi0354), .ZN(new_n6653_));
  INV_X1     g04124(.I(pi0353), .ZN(new_n6654_));
  XOR2_X1    g04125(.A1(pi0352), .A2(pi0360), .Z(new_n6655_));
  XOR2_X1    g04126(.A1(new_n6655_), .A2(new_n6654_), .Z(new_n6656_));
  XOR2_X1    g04127(.A1(new_n6656_), .A2(pi0462), .Z(new_n6657_));
  XOR2_X1    g04128(.A1(new_n6657_), .A2(new_n6653_), .Z(new_n6658_));
  NOR3_X1    g04129(.A1(new_n6658_), .A2(new_n6350_), .A3(new_n6652_), .ZN(new_n6659_));
  NOR2_X1    g04130(.A1(new_n6659_), .A2(pi0590), .ZN(new_n6660_));
  NAND2_X1   g04131(.A1(new_n6520_), .A2(pi0591), .ZN(new_n6661_));
  INV_X1     g04132(.I(pi0285), .ZN(new_n6662_));
  INV_X1     g04133(.I(pi0286), .ZN(new_n6663_));
  INV_X1     g04134(.I(pi0288), .ZN(new_n6664_));
  INV_X1     g04135(.I(pi0289), .ZN(new_n6665_));
  NOR2_X1    g04136(.A1(new_n6664_), .A2(new_n6665_), .ZN(new_n6666_));
  INV_X1     g04137(.I(new_n6666_), .ZN(new_n6667_));
  NOR3_X1    g04138(.A1(new_n6667_), .A2(new_n6662_), .A3(new_n6663_), .ZN(new_n6668_));
  NOR2_X1    g04139(.A1(new_n6668_), .A2(pi0588), .ZN(new_n6669_));
  OAI21_X1   g04140(.A1(new_n6661_), .A2(new_n6660_), .B(new_n6669_), .ZN(new_n6670_));
  INV_X1     g04141(.I(pi0371), .ZN(new_n6671_));
  NAND2_X1   g04142(.A1(pi0374), .A2(pi1198), .ZN(new_n6675_));
  INV_X1     g04143(.I(pi0377), .ZN(new_n6677_));
  INV_X1     g04144(.I(pi0381), .ZN(new_n6678_));
  INV_X1     g04145(.I(pi0317), .ZN(new_n6679_));
  NOR2_X1    g04146(.A1(pi0378), .A2(pi0385), .ZN(new_n6680_));
  INV_X1     g04147(.I(pi0378), .ZN(new_n6681_));
  INV_X1     g04148(.I(pi0385), .ZN(new_n6682_));
  NOR2_X1    g04149(.A1(new_n6681_), .A2(new_n6682_), .ZN(new_n6683_));
  OAI21_X1   g04150(.A1(new_n6683_), .A2(new_n6680_), .B(new_n6679_), .ZN(new_n6684_));
  NOR2_X1    g04151(.A1(new_n6681_), .A2(pi0385), .ZN(new_n6685_));
  NOR2_X1    g04152(.A1(new_n6682_), .A2(pi0378), .ZN(new_n6686_));
  OAI21_X1   g04153(.A1(new_n6685_), .A2(new_n6686_), .B(pi0317), .ZN(new_n6687_));
  NAND2_X1   g04154(.A1(new_n6684_), .A2(new_n6687_), .ZN(new_n6688_));
  XOR2_X1    g04155(.A1(new_n6688_), .A2(new_n6678_), .Z(new_n6689_));
  XOR2_X1    g04156(.A1(new_n6689_), .A2(pi0376), .Z(new_n6690_));
  XOR2_X1    g04157(.A1(new_n6690_), .A2(pi0439), .Z(new_n6691_));
  XNOR2_X1   g04158(.A1(pi0379), .A2(pi0382), .ZN(new_n6692_));
  NAND2_X1   g04159(.A1(new_n6691_), .A2(new_n6692_), .ZN(new_n6693_));
  XNOR2_X1   g04160(.A1(pi0379), .A2(pi0382), .ZN(new_n6694_));
  OAI21_X1   g04161(.A1(new_n6691_), .A2(new_n6694_), .B(new_n6693_), .ZN(new_n6695_));
  INV_X1     g04162(.I(pi0388), .ZN(new_n6699_));
  INV_X1     g04163(.I(pi0387), .ZN(new_n6700_));
  INV_X1     g04164(.I(pi0339), .ZN(new_n6701_));
  XOR2_X1    g04165(.A1(pi0337), .A2(pi0380), .Z(new_n6702_));
  XOR2_X1    g04166(.A1(new_n6702_), .A2(new_n6701_), .Z(new_n6703_));
  XOR2_X1    g04167(.A1(new_n6703_), .A2(new_n6700_), .Z(new_n6704_));
  INV_X1     g04168(.I(pi0363), .ZN(new_n6705_));
  NOR2_X1    g04169(.A1(pi0372), .A2(pi0386), .ZN(new_n6706_));
  INV_X1     g04170(.I(pi0372), .ZN(new_n6707_));
  INV_X1     g04171(.I(pi0386), .ZN(new_n6708_));
  NOR2_X1    g04172(.A1(new_n6707_), .A2(new_n6708_), .ZN(new_n6709_));
  OAI21_X1   g04173(.A1(new_n6709_), .A2(new_n6706_), .B(new_n6705_), .ZN(new_n6710_));
  NOR2_X1    g04174(.A1(new_n6707_), .A2(pi0386), .ZN(new_n6711_));
  NOR2_X1    g04175(.A1(new_n6708_), .A2(pi0372), .ZN(new_n6712_));
  OAI21_X1   g04176(.A1(new_n6711_), .A2(new_n6712_), .B(pi0363), .ZN(new_n6713_));
  NAND2_X1   g04177(.A1(new_n6710_), .A2(new_n6713_), .ZN(new_n6714_));
  XOR2_X1    g04178(.A1(new_n6714_), .A2(pi0338), .Z(new_n6715_));
  XOR2_X1    g04179(.A1(new_n6704_), .A2(new_n6715_), .Z(new_n6716_));
  XOR2_X1    g04180(.A1(new_n6716_), .A2(new_n6699_), .Z(new_n6717_));
  NAND2_X1   g04181(.A1(new_n6717_), .A2(pi1196), .ZN(new_n6718_));
  INV_X1     g04182(.I(new_n6718_), .ZN(new_n6719_));
  XOR2_X1    g04183(.A1(pi0365), .A2(pi0447), .Z(new_n6720_));
  INV_X1     g04184(.I(new_n6720_), .ZN(new_n6721_));
  INV_X1     g04185(.I(pi0364), .ZN(new_n6722_));
  XOR2_X1    g04186(.A1(pi0336), .A2(pi0366), .Z(new_n6723_));
  XOR2_X1    g04187(.A1(new_n6723_), .A2(new_n6722_), .Z(new_n6724_));
  XOR2_X1    g04188(.A1(new_n6724_), .A2(pi0383), .Z(new_n6725_));
  XOR2_X1    g04189(.A1(new_n6725_), .A2(new_n6721_), .Z(new_n6726_));
  INV_X1     g04190(.I(new_n6726_), .ZN(new_n6727_));
  INV_X1     g04191(.I(pi1197), .ZN(new_n6728_));
  INV_X1     g04192(.I(pi0367), .ZN(new_n6729_));
  XOR2_X1    g04193(.A1(pi0368), .A2(pi0389), .Z(new_n6730_));
  XOR2_X1    g04194(.A1(new_n6730_), .A2(new_n6729_), .Z(new_n6731_));
  XOR2_X1    g04195(.A1(new_n6731_), .A2(new_n6728_), .Z(new_n6732_));
  NAND2_X1   g04196(.A1(new_n6727_), .A2(new_n6732_), .ZN(new_n6733_));
  INV_X1     g04197(.I(new_n6733_), .ZN(new_n6734_));
  NOR2_X1    g04198(.A1(new_n6719_), .A2(new_n6734_), .ZN(new_n6735_));
  INV_X1     g04199(.I(new_n6735_), .ZN(new_n6736_));
  XNOR2_X1   g04200(.A1(pi0369), .A2(pi0370), .ZN(new_n6742_));
  INV_X1     g04201(.I(pi0384), .ZN(new_n6743_));
  INV_X1     g04202(.I(pi0440), .ZN(new_n6744_));
  NOR2_X1    g04203(.A1(new_n6744_), .A2(pi0442), .ZN(new_n6745_));
  INV_X1     g04204(.I(pi0442), .ZN(new_n6746_));
  NOR2_X1    g04205(.A1(new_n6746_), .A2(pi0440), .ZN(new_n6747_));
  OAI21_X1   g04206(.A1(new_n6745_), .A2(new_n6747_), .B(new_n6743_), .ZN(new_n6748_));
  NOR2_X1    g04207(.A1(pi0440), .A2(pi0442), .ZN(new_n6749_));
  NOR2_X1    g04208(.A1(new_n6744_), .A2(new_n6746_), .ZN(new_n6750_));
  OAI21_X1   g04209(.A1(new_n6750_), .A2(new_n6749_), .B(pi0384), .ZN(new_n6751_));
  NAND2_X1   g04210(.A1(new_n6751_), .A2(new_n6748_), .ZN(new_n6752_));
  XOR2_X1    g04211(.A1(pi0373), .A2(pi0375), .Z(new_n6753_));
  NOR2_X1    g04212(.A1(new_n6752_), .A2(new_n6753_), .ZN(new_n6754_));
  XOR2_X1    g04213(.A1(pi0373), .A2(pi0375), .Z(new_n6755_));
  AOI21_X1   g04214(.A1(new_n6752_), .A2(new_n6755_), .B(new_n6754_), .ZN(new_n6756_));
  INV_X1     g04215(.I(pi0333), .ZN(new_n6757_));
  XNOR2_X1   g04216(.A1(pi0328), .A2(pi0396), .ZN(new_n6759_));
  XOR2_X1    g04217(.A1(new_n6759_), .A2(pi0394), .Z(new_n6760_));
  XOR2_X1    g04218(.A1(new_n6760_), .A2(pi0408), .Z(new_n6761_));
  INV_X1     g04219(.I(pi0400), .ZN(new_n6762_));
  XNOR2_X1   g04220(.A1(pi0329), .A2(pi0398), .ZN(new_n6763_));
  XOR2_X1    g04221(.A1(new_n6763_), .A2(pi0395), .Z(new_n6764_));
  XOR2_X1    g04222(.A1(new_n6764_), .A2(pi0399), .Z(new_n6765_));
  XOR2_X1    g04223(.A1(new_n6765_), .A2(new_n6762_), .Z(new_n6766_));
  XOR2_X1    g04224(.A1(new_n6765_), .A2(pi0400), .Z(new_n6767_));
  MUX2_X1    g04225(.I0(new_n6767_), .I1(new_n6766_), .S(new_n6761_), .Z(new_n6768_));
  INV_X1     g04226(.I(new_n6768_), .ZN(new_n6769_));
  NOR2_X1    g04227(.A1(new_n6769_), .A2(new_n6577_), .ZN(new_n6770_));
  INV_X1     g04228(.I(pi0404), .ZN(new_n6773_));
  INV_X1     g04229(.I(pi0319), .ZN(new_n6774_));
  INV_X1     g04230(.I(pi0324), .ZN(new_n6775_));
  NOR2_X1    g04231(.A1(new_n6775_), .A2(pi0456), .ZN(new_n6776_));
  INV_X1     g04232(.I(pi0456), .ZN(new_n6777_));
  NOR2_X1    g04233(.A1(new_n6777_), .A2(pi0324), .ZN(new_n6778_));
  OAI21_X1   g04234(.A1(new_n6776_), .A2(new_n6778_), .B(new_n6774_), .ZN(new_n6779_));
  NOR2_X1    g04235(.A1(pi0324), .A2(pi0456), .ZN(new_n6780_));
  NOR2_X1    g04236(.A1(new_n6775_), .A2(new_n6777_), .ZN(new_n6781_));
  OAI21_X1   g04237(.A1(new_n6781_), .A2(new_n6780_), .B(pi0319), .ZN(new_n6782_));
  NAND2_X1   g04238(.A1(new_n6782_), .A2(new_n6779_), .ZN(new_n6783_));
  XOR2_X1    g04239(.A1(new_n6783_), .A2(new_n6773_), .Z(new_n6784_));
  XOR2_X1    g04240(.A1(new_n6784_), .A2(pi0397), .Z(new_n6785_));
  XOR2_X1    g04241(.A1(new_n6785_), .A2(pi0412), .Z(new_n6786_));
  XOR2_X1    g04242(.A1(pi0390), .A2(pi0410), .Z(new_n6787_));
  INV_X1     g04243(.I(new_n6787_), .ZN(new_n6788_));
  XNOR2_X1   g04244(.A1(pi0390), .A2(pi0410), .ZN(new_n6789_));
  NOR2_X1    g04245(.A1(new_n6786_), .A2(new_n6789_), .ZN(new_n6790_));
  AOI21_X1   g04246(.A1(new_n6786_), .A2(new_n6788_), .B(new_n6790_), .ZN(new_n6791_));
  XOR2_X1    g04247(.A1(new_n6791_), .A2(pi0411), .Z(new_n6792_));
  NOR2_X1    g04248(.A1(new_n6537_), .A2(new_n6448_), .ZN(new_n6796_));
  NOR2_X1    g04249(.A1(new_n6537_), .A2(new_n5434_), .ZN(new_n6797_));
  INV_X1     g04250(.I(new_n6796_), .ZN(new_n6803_));
  NOR2_X1    g04251(.A1(new_n6595_), .A2(pi0592), .ZN(new_n6815_));
  INV_X1     g04252(.I(new_n6815_), .ZN(new_n6816_));
  INV_X1     g04253(.I(pi0326), .ZN(new_n6820_));
  XOR2_X1    g04254(.A1(pi0325), .A2(pi0403), .Z(new_n6821_));
  XOR2_X1    g04255(.A1(new_n6821_), .A2(new_n6820_), .Z(new_n6822_));
  XOR2_X1    g04256(.A1(new_n6822_), .A2(pi0405), .Z(new_n6823_));
  XOR2_X1    g04257(.A1(new_n6823_), .A2(pi0402), .Z(new_n6824_));
  XOR2_X1    g04258(.A1(new_n6824_), .A2(pi0401), .Z(new_n6825_));
  XOR2_X1    g04259(.A1(new_n6825_), .A2(pi0406), .Z(new_n6826_));
  INV_X1     g04260(.I(new_n6826_), .ZN(new_n6827_));
  XOR2_X1    g04261(.A1(pi0318), .A2(pi0409), .Z(new_n6828_));
  NOR2_X1    g04262(.A1(new_n6827_), .A2(new_n6828_), .ZN(new_n6829_));
  XNOR2_X1   g04263(.A1(pi0318), .A2(pi0409), .ZN(new_n6830_));
  NOR2_X1    g04264(.A1(new_n6826_), .A2(new_n6830_), .ZN(new_n6831_));
  NOR2_X1    g04265(.A1(new_n6829_), .A2(new_n6831_), .ZN(new_n6832_));
  INV_X1     g04266(.I(new_n6832_), .ZN(new_n6833_));
  INV_X1     g04267(.I(new_n6792_), .ZN(new_n6845_));
  INV_X1     g04268(.I(new_n6490_), .ZN(new_n6878_));
  INV_X1     g04269(.I(new_n6488_), .ZN(new_n6894_));
  INV_X1     g04270(.I(pi0334), .ZN(new_n6925_));
  XNOR2_X1   g04271(.A1(pi0335), .A2(pi0413), .ZN(new_n6926_));
  XOR2_X1    g04272(.A1(new_n6926_), .A2(pi0407), .Z(new_n6927_));
  XOR2_X1    g04273(.A1(new_n6927_), .A2(pi0463), .Z(new_n6928_));
  NOR2_X1    g04274(.A1(new_n6928_), .A2(new_n6925_), .ZN(new_n6929_));
  AND2_X2    g04275(.A1(new_n6928_), .A2(new_n6925_), .Z(new_n6930_));
  NOR2_X1    g04276(.A1(new_n6930_), .A2(new_n6929_), .ZN(new_n6931_));
  XOR2_X1    g04277(.A1(new_n6931_), .A2(pi0393), .Z(new_n6932_));
  INV_X1     g04278(.I(pi0590), .ZN(new_n6933_));
  NOR2_X1    g04279(.A1(new_n6933_), .A2(new_n6350_), .ZN(new_n6934_));
  INV_X1     g04280(.I(new_n6934_), .ZN(new_n6935_));
  NOR3_X1    g04281(.A1(new_n6756_), .A2(new_n6671_), .A3(new_n6742_), .ZN(new_n6938_));
  INV_X1     g04282(.I(new_n6668_), .ZN(new_n6939_));
  NOR2_X1    g04283(.A1(new_n2984_), .A2(pi1091), .ZN(new_n6940_));
  INV_X1     g04284(.I(new_n6940_), .ZN(new_n6941_));
  AOI21_X1   g04285(.A1(new_n6476_), .A2(new_n6941_), .B(new_n6475_), .ZN(new_n6942_));
  INV_X1     g04286(.I(new_n6942_), .ZN(new_n6943_));
  NOR2_X1    g04287(.A1(new_n6470_), .A2(new_n6941_), .ZN(new_n6944_));
  NOR3_X1    g04288(.A1(new_n6944_), .A2(pi0087), .A3(new_n3134_), .ZN(new_n6945_));
  NOR2_X1    g04289(.A1(new_n6945_), .A2(new_n6943_), .ZN(new_n6946_));
  INV_X1     g04290(.I(new_n6946_), .ZN(new_n6947_));
  NOR4_X1    g04291(.A1(new_n6435_), .A2(new_n5685_), .A3(new_n6414_), .A4(new_n6551_), .ZN(new_n6948_));
  NOR2_X1    g04292(.A1(new_n6534_), .A2(new_n3455_), .ZN(new_n6949_));
  OAI21_X1   g04293(.A1(new_n6553_), .A2(new_n6949_), .B(new_n6948_), .ZN(new_n6950_));
  AOI21_X1   g04294(.A1(new_n6950_), .A2(new_n6947_), .B(pi0075), .ZN(new_n6951_));
  NOR2_X1    g04295(.A1(new_n6951_), .A2(new_n6529_), .ZN(new_n6952_));
  OAI21_X1   g04296(.A1(new_n6952_), .A2(new_n6514_), .B(new_n6401_), .ZN(new_n6953_));
  XOR2_X1    g04297(.A1(pi0370), .A2(pi0371), .Z(new_n6976_));
  NOR2_X1    g04298(.A1(pi0590), .A2(pi0591), .ZN(new_n6977_));
  INV_X1     g04299(.I(new_n6770_), .ZN(new_n6983_));
  INV_X1     g04300(.I(new_n6554_), .ZN(new_n6989_));
  NOR2_X1    g04301(.A1(pi0075), .A2(pi0592), .ZN(new_n6991_));
  NAND3_X1   g04302(.A1(new_n6752_), .A2(pi0375), .A3(new_n6976_), .ZN(new_n7013_));
  NAND2_X1   g04303(.A1(new_n7013_), .A2(new_n6939_), .ZN(new_n7014_));
  AOI21_X1   g04304(.A1(new_n6670_), .A2(new_n6938_), .B(new_n7014_), .ZN(new_n7015_));
  NOR2_X1    g04305(.A1(new_n6354_), .A2(new_n6352_), .ZN(new_n7039_));
  NOR2_X1    g04306(.A1(new_n7039_), .A2(pi0356), .ZN(new_n7040_));
  NOR2_X1    g04307(.A1(new_n7039_), .A2(new_n6650_), .ZN(new_n7041_));
  NOR2_X1    g04308(.A1(new_n7040_), .A2(new_n7041_), .ZN(new_n7042_));
  NOR3_X1    g04309(.A1(new_n6658_), .A2(new_n6350_), .A3(new_n7042_), .ZN(new_n7043_));
  NOR2_X1    g04310(.A1(new_n7043_), .A2(pi0590), .ZN(new_n7044_));
  INV_X1     g04311(.I(pi0416), .ZN(new_n7046_));
  XOR2_X1    g04312(.A1(pi0415), .A2(pi0431), .Z(new_n7047_));
  XOR2_X1    g04313(.A1(new_n7047_), .A2(new_n7046_), .Z(new_n7048_));
  XOR2_X1    g04314(.A1(new_n7048_), .A2(pi0438), .Z(new_n7049_));
  INV_X1     g04315(.I(new_n7049_), .ZN(new_n7050_));
  XOR2_X1    g04316(.A1(pi0421), .A2(pi0454), .Z(new_n7051_));
  XOR2_X1    g04317(.A1(new_n7051_), .A2(pi0432), .Z(new_n7052_));
  XOR2_X1    g04318(.A1(new_n7052_), .A2(pi0459), .Z(new_n7053_));
  INV_X1     g04319(.I(pi0420), .ZN(new_n7054_));
  XOR2_X1    g04320(.A1(pi0419), .A2(pi0423), .Z(new_n7055_));
  XOR2_X1    g04321(.A1(new_n7055_), .A2(new_n7054_), .Z(new_n7056_));
  XOR2_X1    g04322(.A1(new_n7056_), .A2(pi0424), .Z(new_n7057_));
  XOR2_X1    g04323(.A1(new_n7057_), .A2(pi0425), .Z(new_n7058_));
  XOR2_X1    g04324(.A1(new_n7058_), .A2(new_n6577_), .Z(new_n7059_));
  NAND2_X1   g04325(.A1(new_n7059_), .A2(new_n7053_), .ZN(new_n7060_));
  NAND2_X1   g04326(.A1(new_n7060_), .A2(new_n7050_), .ZN(new_n7061_));
  NAND3_X1   g04327(.A1(new_n7059_), .A2(new_n7049_), .A3(new_n7053_), .ZN(new_n7062_));
  INV_X1     g04328(.I(pi0417), .ZN(new_n7063_));
  INV_X1     g04329(.I(pi0418), .ZN(new_n7064_));
  NOR2_X1    g04330(.A1(new_n7064_), .A2(pi0437), .ZN(new_n7065_));
  INV_X1     g04331(.I(pi0437), .ZN(new_n7066_));
  NOR2_X1    g04332(.A1(new_n7066_), .A2(pi0418), .ZN(new_n7067_));
  OAI21_X1   g04333(.A1(new_n7065_), .A2(new_n7067_), .B(new_n7063_), .ZN(new_n7068_));
  NOR2_X1    g04334(.A1(pi0418), .A2(pi0437), .ZN(new_n7069_));
  NOR2_X1    g04335(.A1(new_n7064_), .A2(new_n7066_), .ZN(new_n7070_));
  OAI21_X1   g04336(.A1(new_n7070_), .A2(new_n7069_), .B(pi0417), .ZN(new_n7071_));
  NAND2_X1   g04337(.A1(new_n7071_), .A2(new_n7068_), .ZN(new_n7072_));
  XOR2_X1    g04338(.A1(pi0453), .A2(pi0464), .Z(new_n7073_));
  NOR2_X1    g04339(.A1(new_n7072_), .A2(new_n7073_), .ZN(new_n7074_));
  XOR2_X1    g04340(.A1(pi0453), .A2(pi0464), .Z(new_n7075_));
  AOI21_X1   g04341(.A1(new_n7072_), .A2(new_n7075_), .B(new_n7074_), .ZN(new_n7076_));
  NAND3_X1   g04342(.A1(new_n7061_), .A2(new_n7062_), .A3(new_n7076_), .ZN(new_n7077_));
  NAND2_X1   g04343(.A1(new_n7077_), .A2(pi1197), .ZN(new_n7078_));
  NAND2_X1   g04344(.A1(new_n6358_), .A2(pi0443), .ZN(new_n7079_));
  INV_X1     g04345(.I(pi0444), .ZN(new_n7082_));
  NOR2_X1    g04346(.A1(pi0443), .A2(pi0592), .ZN(new_n7083_));
  INV_X1     g04347(.I(new_n7083_), .ZN(new_n7084_));
  XNOR2_X1   g04348(.A1(pi0414), .A2(pi0434), .ZN(new_n7089_));
  XOR2_X1    g04349(.A1(new_n7089_), .A2(pi0422), .Z(new_n7090_));
  XOR2_X1    g04350(.A1(new_n7090_), .A2(pi0446), .Z(new_n7091_));
  INV_X1     g04351(.I(new_n7091_), .ZN(new_n7092_));
  XNOR2_X1   g04352(.A1(pi0429), .A2(pi0435), .ZN(new_n7093_));
  NOR2_X1    g04353(.A1(new_n7092_), .A2(new_n7093_), .ZN(new_n7094_));
  XOR2_X1    g04354(.A1(pi0429), .A2(pi0435), .Z(new_n7095_));
  NOR2_X1    g04355(.A1(new_n7091_), .A2(new_n7095_), .ZN(new_n7096_));
  NOR2_X1    g04356(.A1(new_n7094_), .A2(new_n7096_), .ZN(new_n7097_));
  INV_X1     g04357(.I(new_n7078_), .ZN(new_n7110_));
  XOR2_X1    g04358(.A1(pi0426), .A2(pi0430), .Z(new_n7113_));
  INV_X1     g04359(.I(pi0448), .ZN(new_n7114_));
  INV_X1     g04360(.I(pi0433), .ZN(new_n7115_));
  NOR2_X1    g04361(.A1(pi0449), .A2(pi0451), .ZN(new_n7116_));
  INV_X1     g04362(.I(pi0449), .ZN(new_n7117_));
  INV_X1     g04363(.I(pi0451), .ZN(new_n7118_));
  NOR2_X1    g04364(.A1(new_n7117_), .A2(new_n7118_), .ZN(new_n7119_));
  OAI21_X1   g04365(.A1(new_n7119_), .A2(new_n7116_), .B(new_n7115_), .ZN(new_n7120_));
  NOR2_X1    g04366(.A1(new_n7117_), .A2(pi0451), .ZN(new_n7121_));
  NOR2_X1    g04367(.A1(new_n7118_), .A2(pi0449), .ZN(new_n7122_));
  OAI21_X1   g04368(.A1(new_n7121_), .A2(new_n7122_), .B(pi0433), .ZN(new_n7123_));
  NAND2_X1   g04369(.A1(new_n7120_), .A2(new_n7123_), .ZN(new_n7124_));
  XOR2_X1    g04370(.A1(new_n7124_), .A2(new_n7114_), .Z(new_n7125_));
  NAND3_X1   g04371(.A1(new_n7125_), .A2(pi0445), .A3(new_n7113_), .ZN(new_n7127_));
  NAND2_X1   g04372(.A1(new_n7127_), .A2(new_n6939_), .ZN(new_n7128_));
  INV_X1     g04373(.I(new_n6977_), .ZN(new_n7129_));
  NOR2_X1    g04374(.A1(new_n6953_), .A2(new_n7129_), .ZN(new_n7130_));
  NAND2_X1   g04375(.A1(new_n5787_), .A2(new_n5371_), .ZN(po1038));
  AOI22_X1   g04376(.A1(new_n7130_), .A2(new_n7128_), .B1(pi0588), .B2(po1038), .ZN(new_n7132_));
  NAND3_X1   g04377(.A1(new_n6559_), .A2(pi0443), .A3(new_n6358_), .ZN(new_n7134_));
  XOR2_X1    g04378(.A1(pi0436), .A2(pi0444), .Z(new_n7135_));
  XOR2_X1    g04379(.A1(new_n7097_), .A2(new_n7135_), .Z(new_n7136_));
  NAND3_X1   g04380(.A1(new_n7134_), .A2(pi1196), .A3(new_n7136_), .ZN(new_n7137_));
  NOR2_X1    g04381(.A1(new_n7136_), .A2(new_n7079_), .ZN(new_n7138_));
  OAI21_X1   g04382(.A1(new_n6560_), .A2(new_n7084_), .B(new_n7138_), .ZN(new_n7139_));
  OAI21_X1   g04383(.A1(new_n7137_), .A2(new_n7139_), .B(new_n6521_), .ZN(new_n7140_));
  AOI21_X1   g04384(.A1(new_n7140_), .A2(new_n7083_), .B(new_n7078_), .ZN(new_n7141_));
  NAND3_X1   g04385(.A1(new_n6562_), .A2(new_n6643_), .A3(new_n7110_), .ZN(new_n7142_));
  XOR2_X1    g04386(.A1(new_n7142_), .A2(new_n7141_), .Z(new_n7143_));
  XOR2_X1    g04387(.A1(new_n7124_), .A2(pi0448), .Z(new_n7147_));
  NOR2_X1    g04388(.A1(new_n6668_), .A2(new_n7129_), .ZN(new_n7148_));
  OAI21_X1   g04389(.A1(new_n6520_), .A2(new_n6977_), .B(new_n7148_), .ZN(new_n7149_));
  OAI21_X1   g04390(.A1(new_n7143_), .A2(new_n7149_), .B(new_n6356_), .ZN(new_n7150_));
  NOR2_X1    g04391(.A1(new_n6409_), .A2(new_n6514_), .ZN(new_n7152_));
  INV_X1     g04392(.I(new_n7152_), .ZN(new_n7153_));
  NOR2_X1    g04393(.A1(new_n7153_), .A2(new_n6358_), .ZN(new_n7154_));
  INV_X1     g04394(.I(new_n7154_), .ZN(new_n7164_));
  NAND2_X1   g04395(.A1(new_n6932_), .A2(pi0591), .ZN(new_n7175_));
  XOR2_X1    g04396(.A1(new_n7175_), .A2(new_n6935_), .Z(new_n7176_));
  INV_X1     g04397(.I(pi0375), .ZN(new_n7177_));
  INV_X1     g04398(.I(pi0374), .ZN(new_n7178_));
  INV_X1     g04399(.I(pi0370), .ZN(new_n7179_));
  XOR2_X1    g04400(.A1(pi0369), .A2(pi0371), .Z(new_n7180_));
  XOR2_X1    g04401(.A1(new_n7180_), .A2(new_n7179_), .Z(new_n7181_));
  XOR2_X1    g04402(.A1(new_n7181_), .A2(new_n7178_), .Z(new_n7182_));
  XOR2_X1    g04403(.A1(new_n6752_), .A2(pi0373), .Z(new_n7183_));
  XOR2_X1    g04404(.A1(new_n7182_), .A2(new_n7183_), .Z(new_n7184_));
  XOR2_X1    g04405(.A1(new_n7184_), .A2(new_n7177_), .Z(new_n7185_));
  XOR2_X1    g04406(.A1(new_n6695_), .A2(new_n6677_), .Z(new_n7186_));
  NAND2_X1   g04407(.A1(new_n7186_), .A2(new_n6735_), .ZN(new_n7187_));
  INV_X1     g04408(.I(new_n7187_), .ZN(new_n7188_));
  OAI21_X1   g04409(.A1(new_n7153_), .A2(new_n6356_), .B(new_n6358_), .ZN(new_n7189_));
  AOI22_X1   g04410(.A1(new_n7188_), .A2(new_n7189_), .B1(pi0592), .B2(new_n6736_), .ZN(new_n7190_));
  NOR2_X1    g04411(.A1(new_n7153_), .A2(pi0592), .ZN(new_n7191_));
  NAND3_X1   g04412(.A1(new_n7190_), .A2(new_n7154_), .A3(new_n7191_), .ZN(new_n7192_));
  AOI21_X1   g04413(.A1(new_n7192_), .A2(new_n6577_), .B(new_n7185_), .ZN(new_n7193_));
  NOR2_X1    g04414(.A1(new_n6354_), .A2(new_n6352_), .ZN(new_n7212_));
  XOR2_X1    g04415(.A1(new_n6658_), .A2(pi0356), .Z(new_n7213_));
  INV_X1     g04416(.I(new_n7213_), .ZN(new_n7214_));
  OAI21_X1   g04417(.A1(new_n7213_), .A2(new_n7212_), .B(pi0590), .ZN(new_n7215_));
  AOI21_X1   g04418(.A1(new_n7212_), .A2(new_n7214_), .B(new_n7215_), .ZN(new_n7216_));
  XOR2_X1    g04419(.A1(new_n7216_), .A2(new_n6934_), .Z(new_n7217_));
  INV_X1     g04420(.I(pi0436), .ZN(new_n7218_));
  INV_X1     g04421(.I(pi0443), .ZN(new_n7219_));
  NOR2_X1    g04422(.A1(new_n7219_), .A2(pi0444), .ZN(new_n7220_));
  NOR2_X1    g04423(.A1(new_n7082_), .A2(pi0443), .ZN(new_n7221_));
  OAI21_X1   g04424(.A1(new_n7220_), .A2(new_n7221_), .B(new_n7218_), .ZN(new_n7222_));
  XOR2_X1    g04425(.A1(pi0443), .A2(pi0444), .Z(new_n7223_));
  OAI21_X1   g04426(.A1(new_n7218_), .A2(new_n7223_), .B(new_n7222_), .ZN(new_n7224_));
  AND2_X2    g04427(.A1(new_n7078_), .A2(new_n7224_), .Z(new_n7225_));
  OAI21_X1   g04428(.A1(new_n7078_), .A2(new_n7224_), .B(new_n7097_), .ZN(new_n7226_));
  OAI21_X1   g04429(.A1(new_n7225_), .A2(new_n7226_), .B(new_n6815_), .ZN(new_n7227_));
  NOR3_X1    g04430(.A1(new_n7227_), .A2(pi0592), .A3(new_n7153_), .ZN(new_n7228_));
  NAND2_X1   g04431(.A1(new_n7164_), .A2(pi0448), .ZN(new_n7229_));
  NAND2_X1   g04432(.A1(new_n7154_), .A2(new_n7114_), .ZN(new_n7230_));
  INV_X1     g04433(.I(pi0427), .ZN(new_n7231_));
  XOR2_X1    g04434(.A1(pi0426), .A2(pi0428), .Z(new_n7232_));
  XOR2_X1    g04435(.A1(new_n7232_), .A2(new_n7231_), .Z(new_n7233_));
  XOR2_X1    g04436(.A1(new_n7233_), .A2(pi0430), .Z(new_n7234_));
  XOR2_X1    g04437(.A1(new_n7234_), .A2(pi0445), .Z(new_n7235_));
  NAND3_X1   g04438(.A1(new_n7229_), .A2(new_n7230_), .A3(new_n7235_), .ZN(new_n7236_));
  NAND4_X1   g04439(.A1(new_n7228_), .A2(pi1199), .A3(new_n7124_), .A4(new_n7236_), .ZN(new_n7237_));
  NOR3_X1    g04440(.A1(new_n7228_), .A2(pi1199), .A3(new_n7154_), .ZN(new_n7238_));
  NAND2_X1   g04441(.A1(new_n7152_), .A2(new_n7129_), .ZN(new_n7239_));
  INV_X1     g04442(.I(po1038), .ZN(new_n7240_));
  NAND2_X1   g04443(.A1(new_n7240_), .A2(new_n6939_), .ZN(new_n7241_));
  NAND4_X1   g04444(.A1(new_n7239_), .A2(pi0588), .A3(new_n6977_), .A4(new_n7241_), .ZN(new_n7242_));
  NOR2_X1    g04445(.A1(new_n7238_), .A2(new_n7242_), .ZN(new_n7243_));
  AOI22_X1   g04446(.A1(new_n7243_), .A2(new_n7237_), .B1(new_n7193_), .B2(new_n7217_), .ZN(new_n7244_));
  NOR2_X1    g04447(.A1(new_n7244_), .A2(new_n7153_), .ZN(new_n7245_));
  AOI21_X1   g04448(.A1(new_n7245_), .A2(new_n7176_), .B(pi0217), .ZN(new_n7246_));
  NOR3_X1    g04449(.A1(new_n6953_), .A2(new_n6350_), .A3(new_n7246_), .ZN(new_n7247_));
  NAND3_X1   g04450(.A1(new_n7150_), .A2(new_n7147_), .A3(new_n7247_), .ZN(new_n7248_));
  NOR4_X1    g04451(.A1(new_n7248_), .A2(new_n7015_), .A3(new_n7044_), .A4(new_n7132_), .ZN(new_n7249_));
  NOR3_X1    g04452(.A1(pi1161), .A2(pi1162), .A3(pi1163), .ZN(new_n7250_));
  NOR2_X1    g04453(.A1(new_n6520_), .A2(new_n6939_), .ZN(new_n7251_));
  NOR2_X1    g04454(.A1(new_n7240_), .A2(new_n6939_), .ZN(new_n7252_));
  INV_X1     g04455(.I(new_n7252_), .ZN(new_n7253_));
  XOR2_X1    g04456(.A1(new_n7251_), .A2(new_n7253_), .Z(new_n7254_));
  NOR3_X1    g04457(.A1(new_n7152_), .A2(pi0217), .A3(po1038), .ZN(new_n7255_));
  NOR4_X1    g04458(.A1(new_n7254_), .A2(new_n6939_), .A3(new_n6953_), .A4(new_n7255_), .ZN(new_n7256_));
  OAI21_X1   g04459(.A1(new_n7249_), .A2(new_n7250_), .B(new_n7256_), .ZN(new_n7257_));
  INV_X1     g04460(.I(pi1161), .ZN(new_n7258_));
  NOR3_X1    g04461(.A1(new_n2723_), .A2(new_n7258_), .A3(pi1163), .ZN(new_n7259_));
  NOR2_X1    g04462(.A1(new_n7259_), .A2(pi1162), .ZN(new_n7260_));
  AOI21_X1   g04463(.A1(new_n7257_), .A2(new_n7260_), .B(new_n6349_), .ZN(po0189));
  NAND2_X1   g04464(.A1(pi0024), .A2(pi0841), .ZN(new_n7262_));
  AOI21_X1   g04465(.A1(new_n2773_), .A2(new_n2794_), .B(new_n7262_), .ZN(new_n7263_));
  NOR2_X1    g04466(.A1(new_n2546_), .A2(new_n2517_), .ZN(new_n7264_));
  INV_X1     g04467(.I(new_n7264_), .ZN(new_n7265_));
  INV_X1     g04468(.I(new_n2900_), .ZN(new_n7266_));
  NOR2_X1    g04469(.A1(new_n2873_), .A2(pi0094), .ZN(new_n7267_));
  INV_X1     g04470(.I(new_n7267_), .ZN(new_n7268_));
  NOR4_X1    g04471(.A1(new_n7268_), .A2(pi0047), .A3(new_n5420_), .A4(new_n7266_), .ZN(new_n7269_));
  INV_X1     g04472(.I(new_n7269_), .ZN(new_n7270_));
  NOR4_X1    g04473(.A1(new_n7265_), .A2(new_n2509_), .A3(new_n2460_), .A4(new_n7270_), .ZN(new_n7271_));
  INV_X1     g04474(.I(pi0024), .ZN(new_n7272_));
  NOR4_X1    g04475(.A1(new_n5464_), .A2(new_n7272_), .A3(new_n2486_), .A4(new_n2679_), .ZN(new_n7273_));
  NAND2_X1   g04476(.A1(new_n7271_), .A2(new_n7273_), .ZN(new_n7274_));
  NOR2_X1    g04477(.A1(new_n2465_), .A2(new_n2469_), .ZN(new_n7275_));
  NAND3_X1   g04478(.A1(new_n2591_), .A2(pi0049), .A3(pi0064), .ZN(new_n7276_));
  INV_X1     g04479(.I(new_n6361_), .ZN(new_n7277_));
  NOR3_X1    g04480(.A1(new_n7277_), .A2(pi0089), .A3(pi0102), .ZN(new_n7278_));
  NAND4_X1   g04481(.A1(new_n7278_), .A2(pi0076), .A3(pi0081), .A4(new_n5570_), .ZN(new_n7279_));
  NOR4_X1    g04482(.A1(new_n7279_), .A2(new_n2610_), .A3(new_n2448_), .A4(new_n7276_), .ZN(new_n7280_));
  INV_X1     g04483(.I(new_n2513_), .ZN(new_n7281_));
  NOR2_X1    g04484(.A1(new_n7281_), .A2(new_n2607_), .ZN(new_n7282_));
  NAND4_X1   g04485(.A1(new_n7282_), .A2(new_n2575_), .A3(new_n2632_), .A4(new_n2576_), .ZN(new_n7283_));
  INV_X1     g04486(.I(new_n7283_), .ZN(new_n7284_));
  INV_X1     g04487(.I(pi0061), .ZN(new_n7285_));
  NOR2_X1    g04488(.A1(new_n2640_), .A2(new_n2631_), .ZN(new_n7286_));
  INV_X1     g04489(.I(new_n7286_), .ZN(new_n7287_));
  NOR2_X1    g04490(.A1(pi0045), .A2(pi0048), .ZN(new_n7288_));
  INV_X1     g04491(.I(new_n7288_), .ZN(new_n7289_));
  NOR4_X1    g04492(.A1(new_n7287_), .A2(new_n7285_), .A3(new_n2585_), .A4(new_n7289_), .ZN(new_n7290_));
  NAND3_X1   g04493(.A1(new_n7280_), .A2(new_n7284_), .A3(new_n7290_), .ZN(new_n7291_));
  NAND2_X1   g04494(.A1(new_n7265_), .A2(new_n7291_), .ZN(new_n7292_));
  NOR3_X1    g04495(.A1(new_n2981_), .A2(new_n2721_), .A3(pi1093), .ZN(new_n7293_));
  NOR2_X1    g04496(.A1(new_n2731_), .A2(new_n7293_), .ZN(new_n7294_));
  NAND2_X1   g04497(.A1(new_n2959_), .A2(new_n2498_), .ZN(new_n7295_));
  NOR3_X1    g04498(.A1(new_n7295_), .A2(new_n6368_), .A3(new_n2776_), .ZN(new_n7296_));
  NAND3_X1   g04499(.A1(new_n7294_), .A2(new_n6939_), .A3(new_n7296_), .ZN(new_n7297_));
  AOI21_X1   g04500(.A1(new_n7292_), .A2(new_n7275_), .B(new_n7297_), .ZN(new_n7298_));
  NOR2_X1    g04501(.A1(new_n7297_), .A2(new_n7272_), .ZN(new_n7299_));
  XOR2_X1    g04502(.A1(new_n7298_), .A2(new_n7299_), .Z(new_n7300_));
  NOR2_X1    g04503(.A1(new_n7291_), .A2(new_n2460_), .ZN(new_n7301_));
  INV_X1     g04504(.I(new_n7301_), .ZN(new_n7302_));
  NOR2_X1    g04505(.A1(new_n7302_), .A2(new_n7270_), .ZN(new_n7303_));
  NAND3_X1   g04506(.A1(new_n7300_), .A2(pi0032), .A3(new_n7303_), .ZN(new_n7304_));
  INV_X1     g04507(.I(new_n7294_), .ZN(po0840));
  OAI21_X1   g04508(.A1(po0840), .A2(new_n6668_), .B(new_n2776_), .ZN(new_n7306_));
  AOI21_X1   g04509(.A1(new_n7304_), .A2(new_n7274_), .B(new_n7306_), .ZN(new_n7307_));
  NAND2_X1   g04510(.A1(new_n7274_), .A2(new_n5469_), .ZN(new_n7308_));
  XNOR2_X1   g04511(.A1(new_n7308_), .A2(new_n5470_), .ZN(new_n7309_));
  NOR2_X1    g04512(.A1(new_n3213_), .A2(pi0095), .ZN(new_n7310_));
  NOR4_X1    g04513(.A1(new_n7309_), .A2(new_n5466_), .A3(new_n5469_), .A4(new_n7310_), .ZN(new_n7311_));
  OAI21_X1   g04514(.A1(new_n7263_), .A2(new_n7307_), .B(new_n7311_), .ZN(new_n7312_));
  NOR2_X1    g04515(.A1(new_n3211_), .A2(pi0100), .ZN(new_n7313_));
  NOR4_X1    g04516(.A1(new_n5526_), .A2(new_n3145_), .A3(new_n5502_), .A4(new_n5536_), .ZN(new_n7314_));
  NOR2_X1    g04517(.A1(new_n5526_), .A2(new_n6495_), .ZN(new_n7315_));
  NOR3_X1    g04518(.A1(new_n5502_), .A2(new_n2776_), .A3(new_n3721_), .ZN(new_n7316_));
  AND3_X2    g04519(.A1(new_n7314_), .A2(new_n7315_), .A3(new_n7316_), .Z(new_n7317_));
  INV_X1     g04520(.I(pi0129), .ZN(new_n7318_));
  NOR2_X1    g04521(.A1(new_n3145_), .A2(new_n7318_), .ZN(new_n7319_));
  INV_X1     g04522(.I(new_n7319_), .ZN(new_n7320_));
  NOR2_X1    g04523(.A1(new_n7320_), .A2(new_n2776_), .ZN(new_n7321_));
  NOR2_X1    g04524(.A1(new_n3304_), .A2(new_n2473_), .ZN(new_n7322_));
  INV_X1     g04525(.I(new_n7322_), .ZN(new_n7323_));
  NOR3_X1    g04526(.A1(new_n7323_), .A2(new_n7272_), .A3(new_n2702_), .ZN(new_n7324_));
  NAND2_X1   g04527(.A1(new_n2715_), .A2(new_n7324_), .ZN(new_n7325_));
  NOR2_X1    g04528(.A1(new_n7315_), .A2(new_n3721_), .ZN(new_n7326_));
  INV_X1     g04529(.I(new_n7326_), .ZN(new_n7327_));
  NOR2_X1    g04530(.A1(new_n3426_), .A2(new_n3226_), .ZN(new_n7328_));
  INV_X1     g04531(.I(new_n7328_), .ZN(new_n7329_));
  NOR2_X1    g04532(.A1(new_n7329_), .A2(new_n5767_), .ZN(new_n7330_));
  NAND2_X1   g04533(.A1(new_n7330_), .A2(new_n5499_), .ZN(new_n7331_));
  INV_X1     g04534(.I(new_n7331_), .ZN(new_n7332_));
  NOR2_X1    g04535(.A1(new_n3212_), .A2(pi0087), .ZN(new_n7333_));
  INV_X1     g04536(.I(new_n7333_), .ZN(new_n7334_));
  NOR2_X1    g04537(.A1(new_n3235_), .A2(pi0100), .ZN(new_n7335_));
  INV_X1     g04538(.I(new_n7335_), .ZN(new_n7336_));
  NOR2_X1    g04539(.A1(new_n7334_), .A2(new_n7336_), .ZN(new_n7337_));
  NAND4_X1   g04540(.A1(new_n7332_), .A2(new_n2776_), .A3(po0840), .A4(new_n7337_), .ZN(new_n7338_));
  NOR4_X1    g04541(.A1(new_n7327_), .A2(new_n5527_), .A3(new_n7325_), .A4(new_n7338_), .ZN(new_n7339_));
  OAI22_X1   g04542(.A1(new_n7339_), .A2(new_n3171_), .B1(new_n7317_), .B2(new_n7321_), .ZN(new_n7340_));
  AOI21_X1   g04543(.A1(new_n7312_), .A2(new_n7313_), .B(new_n7340_), .ZN(po0190));
  INV_X1     g04544(.I(pi0193), .ZN(new_n7342_));
  AOI21_X1   g04545(.A1(new_n7264_), .A2(new_n2519_), .B(new_n2896_), .ZN(new_n7343_));
  INV_X1     g04546(.I(new_n7343_), .ZN(new_n7344_));
  NOR4_X1    g04547(.A1(new_n2899_), .A2(new_n2679_), .A3(new_n2708_), .A4(new_n2903_), .ZN(new_n7345_));
  AOI21_X1   g04548(.A1(new_n7345_), .A2(new_n7344_), .B(pi0070), .ZN(new_n7346_));
  INV_X1     g04549(.I(new_n7346_), .ZN(new_n7347_));
  NOR2_X1    g04550(.A1(new_n2758_), .A2(new_n3304_), .ZN(new_n7348_));
  AOI21_X1   g04551(.A1(new_n7347_), .A2(new_n7348_), .B(new_n5559_), .ZN(new_n7349_));
  INV_X1     g04552(.I(new_n7348_), .ZN(new_n7350_));
  INV_X1     g04553(.I(new_n2456_), .ZN(new_n7351_));
  NOR3_X1    g04554(.A1(pi0064), .A2(pi0081), .A3(pi0102), .ZN(new_n7352_));
  INV_X1     g04555(.I(new_n7352_), .ZN(new_n7353_));
  NOR2_X1    g04556(.A1(new_n7353_), .A2(new_n2640_), .ZN(new_n7354_));
  INV_X1     g04557(.I(new_n7354_), .ZN(new_n7355_));
  NOR2_X1    g04558(.A1(new_n7355_), .A2(new_n7351_), .ZN(new_n7356_));
  INV_X1     g04559(.I(new_n7356_), .ZN(new_n7357_));
  NOR2_X1    g04560(.A1(new_n2569_), .A2(new_n7357_), .ZN(new_n7358_));
  NOR2_X1    g04561(.A1(new_n7344_), .A2(new_n2518_), .ZN(new_n7359_));
  OAI21_X1   g04562(.A1(new_n7359_), .A2(new_n7358_), .B(pi0060), .ZN(new_n7360_));
  INV_X1     g04563(.I(pi0082), .ZN(new_n7361_));
  INV_X1     g04564(.I(new_n2446_), .ZN(new_n7362_));
  NOR2_X1    g04565(.A1(new_n7362_), .A2(pi0111), .ZN(new_n7363_));
  NAND4_X1   g04566(.A1(new_n7363_), .A2(pi0036), .A3(pi0068), .A4(new_n2444_), .ZN(new_n7364_));
  NOR4_X1    g04567(.A1(new_n7364_), .A2(new_n7361_), .A3(new_n2598_), .A4(new_n2592_), .ZN(new_n7365_));
  NAND3_X1   g04568(.A1(new_n7365_), .A2(new_n2589_), .A3(new_n7356_), .ZN(new_n7366_));
  NAND3_X1   g04569(.A1(new_n7366_), .A2(new_n2519_), .A3(new_n2448_), .ZN(new_n7367_));
  NAND3_X1   g04570(.A1(new_n7360_), .A2(pi0053), .A3(new_n7367_), .ZN(new_n7368_));
  NAND2_X1   g04571(.A1(new_n7368_), .A2(new_n2516_), .ZN(new_n7369_));
  NAND3_X1   g04572(.A1(new_n7369_), .A2(new_n2707_), .A3(new_n2448_), .ZN(new_n7370_));
  NAND2_X1   g04573(.A1(new_n7370_), .A2(new_n7345_), .ZN(new_n7371_));
  INV_X1     g04574(.I(new_n7371_), .ZN(new_n7372_));
  NOR2_X1    g04575(.A1(new_n7372_), .A2(new_n7350_), .ZN(new_n7373_));
  NOR2_X1    g04576(.A1(new_n7373_), .A2(new_n5559_), .ZN(new_n7374_));
  INV_X1     g04577(.I(pi0183), .ZN(new_n7375_));
  NOR2_X1    g04578(.A1(new_n5386_), .A2(new_n7375_), .ZN(new_n7376_));
  NAND3_X1   g04579(.A1(new_n7374_), .A2(pi0174), .A3(new_n7376_), .ZN(new_n7377_));
  INV_X1     g04580(.I(pi0174), .ZN(new_n7378_));
  INV_X1     g04581(.I(new_n7374_), .ZN(new_n7379_));
  NAND3_X1   g04582(.A1(new_n7379_), .A2(new_n7378_), .A3(new_n7376_), .ZN(new_n7380_));
  NAND2_X1   g04583(.A1(new_n7380_), .A2(new_n7377_), .ZN(new_n7381_));
  AOI21_X1   g04584(.A1(new_n7381_), .A2(new_n7349_), .B(new_n7342_), .ZN(new_n7382_));
  NOR3_X1    g04585(.A1(new_n2471_), .A2(new_n2679_), .A3(pi0841), .ZN(new_n7383_));
  OAI21_X1   g04586(.A1(new_n2496_), .A2(new_n5423_), .B(new_n7383_), .ZN(new_n7384_));
  NAND2_X1   g04587(.A1(new_n7372_), .A2(new_n7384_), .ZN(new_n7385_));
  NAND2_X1   g04588(.A1(new_n7385_), .A2(new_n7348_), .ZN(new_n7386_));
  INV_X1     g04589(.I(new_n7386_), .ZN(new_n7387_));
  INV_X1     g04590(.I(new_n7373_), .ZN(new_n7388_));
  NAND3_X1   g04591(.A1(new_n7388_), .A2(new_n2794_), .A3(new_n5558_), .ZN(new_n7389_));
  NAND2_X1   g04592(.A1(new_n7389_), .A2(pi0095), .ZN(new_n7390_));
  INV_X1     g04593(.I(new_n7390_), .ZN(new_n7391_));
  NOR2_X1    g04594(.A1(new_n7391_), .A2(pi0198), .ZN(new_n7392_));
  NOR2_X1    g04595(.A1(new_n7392_), .A2(new_n7387_), .ZN(new_n7393_));
  NAND2_X1   g04596(.A1(new_n7346_), .A2(new_n7384_), .ZN(new_n7394_));
  NAND2_X1   g04597(.A1(new_n7394_), .A2(new_n7348_), .ZN(new_n7395_));
  INV_X1     g04598(.I(new_n7395_), .ZN(new_n7396_));
  OAI21_X1   g04599(.A1(new_n7396_), .A2(new_n5559_), .B(new_n5373_), .ZN(new_n7397_));
  NAND2_X1   g04600(.A1(new_n7397_), .A2(pi0174), .ZN(new_n7398_));
  NOR2_X1    g04601(.A1(new_n7378_), .A2(new_n7375_), .ZN(new_n7399_));
  XOR2_X1    g04602(.A1(new_n7398_), .A2(new_n7399_), .Z(new_n7400_));
  INV_X1     g04603(.I(new_n3142_), .ZN(new_n7401_));
  NOR2_X1    g04604(.A1(new_n7401_), .A2(new_n5386_), .ZN(new_n7402_));
  INV_X1     g04605(.I(new_n7402_), .ZN(new_n7403_));
  NOR2_X1    g04606(.A1(new_n7403_), .A2(pi0040), .ZN(new_n7404_));
  INV_X1     g04607(.I(new_n7404_), .ZN(new_n7405_));
  NOR2_X1    g04608(.A1(pi0072), .A2(pi0093), .ZN(new_n7406_));
  OAI21_X1   g04609(.A1(new_n2476_), .A2(new_n7406_), .B(new_n7383_), .ZN(new_n7407_));
  INV_X1     g04610(.I(new_n7275_), .ZN(new_n7408_));
  NOR2_X1    g04611(.A1(new_n7366_), .A2(new_n7408_), .ZN(new_n7409_));
  INV_X1     g04612(.I(new_n7409_), .ZN(new_n7410_));
  NOR2_X1    g04613(.A1(new_n7410_), .A2(new_n2448_), .ZN(new_n7411_));
  INV_X1     g04614(.I(new_n7411_), .ZN(new_n7412_));
  AOI21_X1   g04615(.A1(new_n5423_), .A2(new_n7412_), .B(new_n7407_), .ZN(new_n7413_));
  INV_X1     g04616(.I(new_n7413_), .ZN(new_n7414_));
  NOR3_X1    g04617(.A1(new_n7414_), .A2(pi0183), .A3(new_n7405_), .ZN(new_n7415_));
  NOR2_X1    g04618(.A1(new_n7407_), .A2(new_n5423_), .ZN(new_n7416_));
  INV_X1     g04619(.I(new_n7416_), .ZN(new_n7417_));
  NOR2_X1    g04620(.A1(new_n7417_), .A2(new_n7405_), .ZN(new_n7418_));
  INV_X1     g04621(.I(new_n7418_), .ZN(new_n7419_));
  NOR4_X1    g04622(.A1(new_n7400_), .A2(pi0174), .A3(new_n7415_), .A4(new_n7419_), .ZN(new_n7420_));
  OR2_X2     g04623(.A1(new_n7420_), .A2(new_n7376_), .Z(new_n7421_));
  NAND3_X1   g04624(.A1(new_n2476_), .A2(new_n2679_), .A3(new_n7406_), .ZN(new_n7422_));
  NOR2_X1    g04625(.A1(new_n7412_), .A2(new_n7422_), .ZN(new_n7423_));
  INV_X1     g04626(.I(new_n7423_), .ZN(new_n7424_));
  NOR2_X1    g04627(.A1(new_n7424_), .A2(new_n7401_), .ZN(new_n7425_));
  INV_X1     g04628(.I(new_n7425_), .ZN(new_n7426_));
  NOR2_X1    g04629(.A1(new_n5386_), .A2(pi0040), .ZN(new_n7427_));
  INV_X1     g04630(.I(new_n7427_), .ZN(new_n7428_));
  NOR2_X1    g04631(.A1(new_n7426_), .A2(new_n7428_), .ZN(new_n7429_));
  INV_X1     g04632(.I(new_n7429_), .ZN(new_n7430_));
  NOR4_X1    g04633(.A1(new_n7430_), .A2(pi0174), .A3(pi0183), .A4(new_n7342_), .ZN(new_n7431_));
  NAND3_X1   g04634(.A1(new_n7393_), .A2(new_n7421_), .A3(new_n7431_), .ZN(new_n7432_));
  AND2_X2    g04635(.A1(new_n7432_), .A2(new_n7382_), .Z(new_n7433_));
  OAI21_X1   g04636(.A1(new_n7432_), .A2(new_n7382_), .B(new_n3098_), .ZN(new_n7434_));
  NOR2_X1    g04637(.A1(new_n2822_), .A2(new_n5386_), .ZN(new_n7435_));
  INV_X1     g04638(.I(new_n7435_), .ZN(new_n7436_));
  NOR2_X1    g04639(.A1(new_n7436_), .A2(new_n5642_), .ZN(new_n7437_));
  OAI21_X1   g04640(.A1(new_n7433_), .A2(new_n7434_), .B(new_n7437_), .ZN(new_n7438_));
  NOR2_X1    g04641(.A1(new_n3362_), .A2(new_n3011_), .ZN(new_n7439_));
  INV_X1     g04642(.I(new_n7439_), .ZN(new_n7440_));
  INV_X1     g04643(.I(new_n6537_), .ZN(new_n7441_));
  NOR2_X1    g04644(.A1(new_n5454_), .A2(new_n5386_), .ZN(new_n7442_));
  NAND2_X1   g04645(.A1(new_n7441_), .A2(new_n7442_), .ZN(new_n7443_));
  INV_X1     g04646(.I(new_n7442_), .ZN(new_n7444_));
  NOR2_X1    g04647(.A1(new_n5689_), .A2(new_n7444_), .ZN(new_n7445_));
  NOR2_X1    g04648(.A1(new_n5699_), .A2(new_n7444_), .ZN(new_n7446_));
  AOI21_X1   g04649(.A1(new_n5158_), .A2(new_n3336_), .B(new_n7443_), .ZN(new_n7447_));
  OAI21_X1   g04650(.A1(new_n7447_), .A2(new_n7440_), .B(pi0299), .ZN(new_n7448_));
  INV_X1     g04651(.I(new_n5399_), .ZN(new_n7449_));
  NOR2_X1    g04652(.A1(new_n6544_), .A2(new_n3100_), .ZN(new_n7450_));
  INV_X1     g04653(.I(new_n7450_), .ZN(new_n7451_));
  NOR2_X1    g04654(.A1(new_n7449_), .A2(new_n7451_), .ZN(new_n7452_));
  NAND2_X1   g04655(.A1(new_n5698_), .A2(new_n7452_), .ZN(new_n7453_));
  NAND2_X1   g04656(.A1(new_n7441_), .A2(new_n7452_), .ZN(new_n7454_));
  NAND2_X1   g04657(.A1(new_n7454_), .A2(pi0174), .ZN(new_n7455_));
  NOR2_X1    g04658(.A1(new_n7378_), .A2(new_n3098_), .ZN(new_n7456_));
  XOR2_X1    g04659(.A1(new_n7455_), .A2(new_n7456_), .Z(new_n7457_));
  OAI21_X1   g04660(.A1(new_n7457_), .A2(new_n7453_), .B(pi0232), .ZN(new_n7458_));
  INV_X1     g04661(.I(pi0176), .ZN(new_n7459_));
  NOR2_X1    g04662(.A1(new_n7459_), .A2(new_n5551_), .ZN(new_n7460_));
  INV_X1     g04663(.I(new_n7460_), .ZN(new_n7461_));
  XOR2_X1    g04664(.A1(new_n7458_), .A2(new_n7461_), .Z(new_n7462_));
  NOR3_X1    g04665(.A1(new_n5689_), .A2(new_n7449_), .A3(new_n7451_), .ZN(new_n7463_));
  AOI21_X1   g04666(.A1(new_n7463_), .A2(new_n7378_), .B(pi0299), .ZN(new_n7464_));
  NAND2_X1   g04667(.A1(new_n7462_), .A2(new_n7464_), .ZN(new_n7465_));
  NAND3_X1   g04668(.A1(new_n7465_), .A2(pi0039), .A3(new_n7448_), .ZN(new_n7466_));
  NOR2_X1    g04669(.A1(new_n5551_), .A2(pi0039), .ZN(new_n7467_));
  INV_X1     g04670(.I(new_n7467_), .ZN(new_n7468_));
  NAND3_X1   g04671(.A1(new_n7438_), .A2(new_n7466_), .A3(new_n7468_), .ZN(new_n7469_));
  NAND2_X1   g04672(.A1(new_n7388_), .A2(new_n5657_), .ZN(new_n7470_));
  NAND2_X1   g04673(.A1(new_n7470_), .A2(new_n5158_), .ZN(new_n7471_));
  NAND2_X1   g04674(.A1(new_n7347_), .A2(new_n7348_), .ZN(new_n7472_));
  NAND2_X1   g04675(.A1(new_n7472_), .A2(new_n5657_), .ZN(new_n7473_));
  NAND2_X1   g04676(.A1(new_n7473_), .A2(new_n5158_), .ZN(new_n7474_));
  INV_X1     g04677(.I(pi0149), .ZN(new_n7475_));
  NOR4_X1    g04678(.A1(new_n7395_), .A2(new_n7475_), .A3(new_n3827_), .A4(new_n5386_), .ZN(new_n7476_));
  NAND4_X1   g04679(.A1(new_n7471_), .A2(new_n7387_), .A3(new_n7474_), .A4(new_n7476_), .ZN(new_n7477_));
  OAI21_X1   g04680(.A1(new_n7436_), .A2(new_n5661_), .B(pi0299), .ZN(new_n7478_));
  NAND2_X1   g04681(.A1(new_n5158_), .A2(pi0172), .ZN(new_n7479_));
  NOR2_X1    g04682(.A1(new_n7414_), .A2(new_n7405_), .ZN(new_n7480_));
  NAND2_X1   g04683(.A1(new_n7480_), .A2(new_n5158_), .ZN(new_n7481_));
  NAND4_X1   g04684(.A1(new_n7481_), .A2(pi0172), .A3(new_n7419_), .A4(new_n7429_), .ZN(new_n7482_));
  XOR2_X1    g04685(.A1(new_n7482_), .A2(new_n7479_), .Z(new_n7483_));
  NAND2_X1   g04686(.A1(new_n7483_), .A2(pi0149), .ZN(new_n7484_));
  AOI21_X1   g04687(.A1(new_n7477_), .A2(new_n7478_), .B(new_n7484_), .ZN(new_n7485_));
  AOI21_X1   g04688(.A1(new_n7469_), .A2(new_n7485_), .B(new_n3259_), .ZN(new_n7486_));
  NOR2_X1    g04689(.A1(new_n3259_), .A2(new_n3455_), .ZN(new_n7487_));
  XOR2_X1    g04690(.A1(new_n7486_), .A2(new_n7487_), .Z(new_n7488_));
  INV_X1     g04691(.I(pi0186), .ZN(new_n7489_));
  NOR2_X1    g04692(.A1(new_n5503_), .A2(new_n6494_), .ZN(new_n7490_));
  INV_X1     g04693(.I(pi0164), .ZN(new_n7491_));
  NOR2_X1    g04694(.A1(new_n6494_), .A2(new_n3098_), .ZN(new_n7492_));
  INV_X1     g04695(.I(new_n7492_), .ZN(new_n7493_));
  NOR2_X1    g04696(.A1(new_n5492_), .A2(new_n7493_), .ZN(new_n7494_));
  NOR2_X1    g04697(.A1(new_n7494_), .A2(new_n7491_), .ZN(new_n7495_));
  NOR2_X1    g04698(.A1(new_n7491_), .A2(new_n7489_), .ZN(new_n7496_));
  XOR2_X1    g04699(.A1(new_n7495_), .A2(new_n7496_), .Z(new_n7497_));
  NAND2_X1   g04700(.A1(new_n7497_), .A2(new_n7490_), .ZN(new_n7498_));
  INV_X1     g04701(.I(new_n5492_), .ZN(new_n7499_));
  NAND3_X1   g04702(.A1(new_n7499_), .A2(new_n3098_), .A3(new_n6493_), .ZN(new_n7500_));
  NAND3_X1   g04703(.A1(new_n7498_), .A2(new_n7489_), .A3(new_n7500_), .ZN(new_n7501_));
  NAND3_X1   g04704(.A1(new_n6493_), .A2(pi0164), .A3(pi0299), .ZN(new_n7502_));
  NAND3_X1   g04705(.A1(new_n6493_), .A2(new_n7491_), .A3(new_n3098_), .ZN(new_n7503_));
  AOI21_X1   g04706(.A1(new_n7503_), .A2(new_n7502_), .B(new_n7489_), .ZN(new_n7504_));
  NOR2_X1    g04707(.A1(new_n7504_), .A2(new_n3477_), .ZN(new_n7505_));
  XNOR2_X1   g04708(.A1(pi0149), .A2(pi0157), .ZN(new_n7506_));
  NOR2_X1    g04709(.A1(new_n7506_), .A2(new_n5386_), .ZN(new_n7507_));
  NOR2_X1    g04710(.A1(new_n7507_), .A2(new_n5551_), .ZN(new_n7508_));
  XOR2_X1    g04711(.A1(new_n7508_), .A2(new_n5912_), .Z(new_n7509_));
  INV_X1     g04712(.I(pi0178), .ZN(new_n7510_));
  NAND2_X1   g04713(.A1(new_n7510_), .A2(pi0183), .ZN(new_n7511_));
  NAND2_X1   g04714(.A1(new_n7375_), .A2(pi0178), .ZN(new_n7512_));
  AOI21_X1   g04715(.A1(new_n7511_), .A2(new_n7512_), .B(new_n5386_), .ZN(new_n7513_));
  NAND2_X1   g04716(.A1(new_n7509_), .A2(new_n7513_), .ZN(new_n7514_));
  NAND2_X1   g04717(.A1(new_n7514_), .A2(pi0100), .ZN(new_n7515_));
  OAI22_X1   g04718(.A1(new_n7515_), .A2(new_n3189_), .B1(new_n3259_), .B2(new_n7505_), .ZN(new_n7516_));
  AND4_X2    g04719(.A1(pi0164), .A2(new_n7488_), .A3(new_n7501_), .A4(new_n7516_), .Z(new_n7517_));
  NAND2_X1   g04720(.A1(new_n7514_), .A2(pi0075), .ZN(new_n7518_));
  NAND2_X1   g04721(.A1(new_n7518_), .A2(new_n3115_), .ZN(new_n7519_));
  AOI21_X1   g04722(.A1(new_n3336_), .A2(pi0299), .B(new_n5551_), .ZN(new_n7520_));
  NOR2_X1    g04723(.A1(new_n7520_), .A2(new_n5373_), .ZN(new_n7521_));
  NOR3_X1    g04724(.A1(new_n7521_), .A2(new_n7459_), .A3(new_n3098_), .ZN(new_n7522_));
  NOR2_X1    g04725(.A1(pi0038), .A2(pi0087), .ZN(new_n7523_));
  NAND3_X1   g04726(.A1(new_n7522_), .A2(new_n3462_), .A3(new_n7523_), .ZN(new_n7524_));
  NOR2_X1    g04727(.A1(new_n7504_), .A2(new_n3462_), .ZN(new_n7525_));
  NOR2_X1    g04728(.A1(new_n7514_), .A2(new_n5486_), .ZN(new_n7526_));
  XNOR2_X1   g04729(.A1(new_n7526_), .A2(new_n7525_), .ZN(new_n7527_));
  NOR2_X1    g04730(.A1(new_n3303_), .A2(pi0075), .ZN(new_n7528_));
  INV_X1     g04731(.I(new_n7528_), .ZN(new_n7529_));
  OR2_X2     g04732(.A1(new_n7527_), .A2(new_n7529_), .Z(new_n7530_));
  AOI21_X1   g04733(.A1(new_n7530_), .A2(new_n7524_), .B(new_n7499_), .ZN(new_n7531_));
  OAI21_X1   g04734(.A1(new_n7517_), .A2(new_n7519_), .B(new_n7531_), .ZN(new_n7532_));
  NAND2_X1   g04735(.A1(new_n7515_), .A2(new_n7518_), .ZN(new_n7533_));
  NAND2_X1   g04736(.A1(new_n7533_), .A2(new_n6328_), .ZN(new_n7534_));
  NOR2_X1    g04737(.A1(pi0191), .A2(pi0299), .ZN(new_n7535_));
  AOI21_X1   g04738(.A1(new_n4474_), .A2(pi0299), .B(new_n7535_), .ZN(new_n7536_));
  NOR2_X1    g04739(.A1(pi0075), .A2(pi0100), .ZN(new_n7537_));
  INV_X1     g04740(.I(new_n7537_), .ZN(new_n7538_));
  NOR2_X1    g04741(.A1(new_n6494_), .A2(new_n7538_), .ZN(new_n7539_));
  NAND4_X1   g04742(.A1(new_n7534_), .A2(pi0074), .A3(new_n7536_), .A4(new_n7539_), .ZN(new_n7540_));
  OAI21_X1   g04743(.A1(new_n7533_), .A2(new_n3115_), .B(new_n7538_), .ZN(new_n7541_));
  AND2_X2    g04744(.A1(new_n7541_), .A2(new_n7504_), .Z(new_n7542_));
  NAND2_X1   g04745(.A1(new_n7507_), .A2(pi0232), .ZN(new_n7543_));
  INV_X1     g04746(.I(new_n7543_), .ZN(new_n7544_));
  NOR2_X1    g04747(.A1(new_n7544_), .A2(new_n7537_), .ZN(new_n7545_));
  OAI21_X1   g04748(.A1(new_n7545_), .A2(new_n3175_), .B(new_n4474_), .ZN(new_n7546_));
  NAND2_X1   g04749(.A1(new_n7546_), .A2(new_n7539_), .ZN(new_n7547_));
  AOI21_X1   g04750(.A1(pi0164), .A2(new_n7539_), .B(new_n7545_), .ZN(new_n7548_));
  NOR2_X1    g04751(.A1(new_n7548_), .A2(new_n3115_), .ZN(new_n7549_));
  NOR2_X1    g04752(.A1(new_n6494_), .A2(new_n7491_), .ZN(new_n7550_));
  NOR2_X1    g04753(.A1(new_n7550_), .A2(new_n3259_), .ZN(new_n7551_));
  INV_X1     g04754(.I(new_n7550_), .ZN(new_n7552_));
  OAI21_X1   g04755(.A1(new_n7552_), .A2(new_n3259_), .B(pi0100), .ZN(new_n7553_));
  NOR2_X1    g04756(.A1(new_n7543_), .A2(new_n3455_), .ZN(new_n7554_));
  NOR4_X1    g04757(.A1(new_n7553_), .A2(pi0087), .A3(pi0100), .A4(new_n7551_), .ZN(new_n7555_));
  NOR2_X1    g04758(.A1(new_n6494_), .A2(new_n7475_), .ZN(new_n7556_));
  OAI21_X1   g04759(.A1(new_n7555_), .A2(pi0038), .B(new_n7556_), .ZN(new_n7557_));
  OAI21_X1   g04760(.A1(new_n7499_), .A2(new_n7557_), .B(pi0075), .ZN(new_n7558_));
  XOR2_X1    g04761(.A1(new_n7558_), .A2(new_n3483_), .Z(new_n7559_));
  AOI21_X1   g04762(.A1(new_n7559_), .A2(new_n7544_), .B(pi0054), .ZN(new_n7560_));
  NOR2_X1    g04763(.A1(new_n7552_), .A2(new_n3259_), .ZN(new_n7561_));
  AOI21_X1   g04764(.A1(new_n7537_), .A2(new_n7561_), .B(new_n7545_), .ZN(new_n7562_));
  INV_X1     g04765(.I(new_n7562_), .ZN(new_n7563_));
  NOR3_X1    g04766(.A1(new_n7560_), .A2(new_n3303_), .A3(new_n7563_), .ZN(new_n7564_));
  OAI21_X1   g04767(.A1(new_n7564_), .A2(new_n7549_), .B(new_n3175_), .ZN(new_n7565_));
  AOI21_X1   g04768(.A1(new_n7565_), .A2(new_n5975_), .B(new_n7547_), .ZN(new_n7566_));
  NOR2_X1    g04769(.A1(new_n7547_), .A2(new_n3175_), .ZN(new_n7567_));
  OAI21_X1   g04770(.A1(new_n7567_), .A2(new_n7562_), .B(new_n7549_), .ZN(new_n7568_));
  NAND2_X1   g04771(.A1(new_n7568_), .A2(new_n3226_), .ZN(new_n7569_));
  NAND2_X1   g04772(.A1(new_n7569_), .A2(new_n3230_), .ZN(new_n7570_));
  NAND2_X1   g04773(.A1(new_n7547_), .A2(new_n3426_), .ZN(new_n7571_));
  NAND3_X1   g04774(.A1(new_n7571_), .A2(pi0074), .A3(new_n7548_), .ZN(new_n7572_));
  NOR2_X1    g04775(.A1(new_n7570_), .A2(new_n7572_), .ZN(new_n7573_));
  OAI21_X1   g04776(.A1(new_n7566_), .A2(new_n7573_), .B(new_n7542_), .ZN(new_n7574_));
  AOI21_X1   g04777(.A1(new_n7532_), .A2(new_n7540_), .B(new_n7574_), .ZN(new_n7575_));
  NOR2_X1    g04778(.A1(new_n2448_), .A2(pi0040), .ZN(new_n7576_));
  INV_X1     g04779(.I(new_n7576_), .ZN(new_n7577_));
  INV_X1     g04780(.I(new_n7358_), .ZN(new_n7578_));
  NOR2_X1    g04781(.A1(new_n2901_), .A2(new_n2897_), .ZN(new_n7579_));
  INV_X1     g04782(.I(new_n7579_), .ZN(new_n7580_));
  NOR4_X1    g04783(.A1(new_n7578_), .A2(new_n2518_), .A3(new_n2519_), .A4(new_n7580_), .ZN(new_n7581_));
  INV_X1     g04784(.I(new_n7581_), .ZN(new_n7582_));
  NOR2_X1    g04785(.A1(new_n7582_), .A2(pi0058), .ZN(new_n7583_));
  INV_X1     g04786(.I(new_n7583_), .ZN(new_n7584_));
  NOR2_X1    g04787(.A1(new_n7584_), .A2(new_n6368_), .ZN(new_n7585_));
  NAND3_X1   g04788(.A1(new_n7585_), .A2(new_n2794_), .A3(new_n2500_), .ZN(new_n7586_));
  NOR2_X1    g04789(.A1(new_n7586_), .A2(pi0095), .ZN(new_n7587_));
  INV_X1     g04790(.I(new_n7587_), .ZN(new_n7588_));
  NAND4_X1   g04791(.A1(new_n5409_), .A2(pi1092), .A3(new_n5684_), .A4(new_n5687_), .ZN(new_n7589_));
  NOR2_X1    g04792(.A1(new_n7588_), .A2(new_n7589_), .ZN(new_n7590_));
  INV_X1     g04793(.I(new_n7590_), .ZN(new_n7591_));
  AOI21_X1   g04794(.A1(new_n5398_), .A2(new_n7576_), .B(new_n5373_), .ZN(new_n7592_));
  NOR2_X1    g04795(.A1(new_n7591_), .A2(new_n7592_), .ZN(new_n7593_));
  OAI21_X1   g04796(.A1(new_n7450_), .A2(new_n7577_), .B(new_n7593_), .ZN(new_n7594_));
  INV_X1     g04797(.I(new_n7594_), .ZN(new_n7595_));
  NOR2_X1    g04798(.A1(new_n7577_), .A2(new_n7450_), .ZN(new_n7596_));
  INV_X1     g04799(.I(new_n5411_), .ZN(new_n7597_));
  AOI21_X1   g04800(.A1(new_n7597_), .A2(new_n7589_), .B(new_n7588_), .ZN(new_n7598_));
  AOI21_X1   g04801(.A1(new_n7598_), .A2(new_n5385_), .B(new_n7577_), .ZN(new_n7599_));
  NOR2_X1    g04802(.A1(new_n7599_), .A2(new_n7596_), .ZN(new_n7600_));
  INV_X1     g04803(.I(new_n7600_), .ZN(new_n7601_));
  OAI21_X1   g04804(.A1(new_n7601_), .A2(new_n3098_), .B(new_n7378_), .ZN(new_n7602_));
  NAND2_X1   g04805(.A1(new_n7440_), .A2(new_n7576_), .ZN(new_n7603_));
  NAND2_X1   g04806(.A1(new_n7603_), .A2(pi0299), .ZN(new_n7604_));
  INV_X1     g04807(.I(new_n7604_), .ZN(new_n7605_));
  AOI21_X1   g04808(.A1(new_n5455_), .A2(new_n5386_), .B(new_n7577_), .ZN(new_n7606_));
  NAND2_X1   g04809(.A1(new_n7590_), .A2(new_n7606_), .ZN(new_n7607_));
  AOI21_X1   g04810(.A1(new_n7599_), .A2(pi0154), .B(pi0152), .ZN(new_n7608_));
  OAI21_X1   g04811(.A1(new_n7608_), .A2(new_n7607_), .B(new_n7440_), .ZN(new_n7609_));
  INV_X1     g04812(.I(new_n7599_), .ZN(new_n7610_));
  INV_X1     g04813(.I(new_n5434_), .ZN(new_n7611_));
  NOR2_X1    g04814(.A1(new_n7588_), .A2(new_n7597_), .ZN(new_n7612_));
  AOI21_X1   g04815(.A1(new_n7612_), .A2(new_n7611_), .B(new_n7577_), .ZN(new_n7613_));
  OR2_X2     g04816(.A1(new_n7613_), .A2(new_n5373_), .Z(new_n7614_));
  NOR2_X1    g04817(.A1(new_n7614_), .A2(pi0154), .ZN(new_n7615_));
  INV_X1     g04818(.I(new_n7598_), .ZN(new_n7616_));
  AOI21_X1   g04819(.A1(new_n5454_), .A2(new_n7576_), .B(new_n5373_), .ZN(new_n7617_));
  NOR2_X1    g04820(.A1(new_n7616_), .A2(new_n7617_), .ZN(new_n7618_));
  NOR4_X1    g04821(.A1(new_n7615_), .A2(new_n5158_), .A3(new_n7610_), .A4(new_n7618_), .ZN(new_n7619_));
  NAND2_X1   g04822(.A1(new_n7619_), .A2(new_n7609_), .ZN(new_n7620_));
  AOI22_X1   g04823(.A1(new_n7620_), .A2(new_n7605_), .B1(new_n7602_), .B2(new_n7595_), .ZN(new_n7621_));
  NOR2_X1    g04824(.A1(new_n7621_), .A2(new_n7461_), .ZN(new_n7622_));
  NOR2_X1    g04825(.A1(new_n7616_), .A2(new_n7592_), .ZN(new_n7623_));
  INV_X1     g04826(.I(new_n7623_), .ZN(new_n7624_));
  AOI21_X1   g04827(.A1(new_n7624_), .A2(new_n7599_), .B(new_n7596_), .ZN(new_n7625_));
  INV_X1     g04828(.I(new_n7625_), .ZN(new_n7626_));
  NOR2_X1    g04829(.A1(new_n7610_), .A2(new_n7618_), .ZN(new_n7627_));
  NOR3_X1    g04830(.A1(new_n7627_), .A2(new_n5551_), .A3(new_n7604_), .ZN(new_n7628_));
  OAI21_X1   g04831(.A1(new_n7628_), .A2(pi0299), .B(new_n7626_), .ZN(new_n7629_));
  NAND2_X1   g04832(.A1(new_n7629_), .A2(pi0039), .ZN(new_n7630_));
  NOR2_X1    g04833(.A1(pi0176), .A2(pi0232), .ZN(new_n7631_));
  OAI21_X1   g04834(.A1(new_n7622_), .A2(new_n7630_), .B(new_n7631_), .ZN(new_n7632_));
  INV_X1     g04835(.I(new_n7612_), .ZN(new_n7633_));
  NOR2_X1    g04836(.A1(new_n7633_), .A2(new_n7449_), .ZN(new_n7634_));
  AOI21_X1   g04837(.A1(new_n7634_), .A2(new_n7450_), .B(new_n7577_), .ZN(new_n7635_));
  OAI21_X1   g04838(.A1(pi0299), .A2(new_n7635_), .B(new_n7621_), .ZN(new_n7636_));
  INV_X1     g04839(.I(new_n7636_), .ZN(new_n7637_));
  AOI21_X1   g04840(.A1(new_n7637_), .A2(new_n7632_), .B(new_n3259_), .ZN(new_n7638_));
  OAI21_X1   g04841(.A1(new_n7585_), .A2(new_n2448_), .B(pi0070), .ZN(new_n7639_));
  INV_X1     g04842(.I(new_n7639_), .ZN(new_n7640_));
  AOI21_X1   g04843(.A1(new_n2708_), .A2(new_n2539_), .B(pi0070), .ZN(new_n7641_));
  AOI21_X1   g04844(.A1(new_n7582_), .A2(new_n2539_), .B(new_n2686_), .ZN(new_n7642_));
  NAND2_X1   g04845(.A1(new_n2539_), .A2(new_n2516_), .ZN(new_n7643_));
  AOI21_X1   g04846(.A1(new_n7369_), .A2(new_n2901_), .B(new_n7643_), .ZN(new_n7644_));
  NOR2_X1    g04847(.A1(new_n2901_), .A2(new_n2448_), .ZN(new_n7645_));
  OAI21_X1   g04848(.A1(new_n7644_), .A2(pi0058), .B(new_n7645_), .ZN(new_n7646_));
  NOR2_X1    g04849(.A1(new_n7584_), .A2(pi0841), .ZN(new_n7647_));
  AOI21_X1   g04850(.A1(new_n2708_), .A2(new_n2448_), .B(new_n2679_), .ZN(new_n7648_));
  NAND2_X1   g04851(.A1(new_n7647_), .A2(new_n7648_), .ZN(new_n7649_));
  NAND2_X1   g04852(.A1(new_n7646_), .A2(new_n7649_), .ZN(new_n7650_));
  NAND2_X1   g04853(.A1(new_n7650_), .A2(new_n7642_), .ZN(new_n7651_));
  AND2_X2    g04854(.A1(new_n7651_), .A2(new_n7641_), .Z(new_n7652_));
  NOR2_X1    g04855(.A1(new_n2958_), .A2(new_n2702_), .ZN(new_n7653_));
  OAI21_X1   g04856(.A1(new_n7652_), .A2(new_n7640_), .B(new_n7653_), .ZN(new_n7654_));
  INV_X1     g04857(.I(new_n7653_), .ZN(new_n7655_));
  NOR2_X1    g04858(.A1(new_n7655_), .A2(new_n2448_), .ZN(new_n7656_));
  AOI21_X1   g04859(.A1(new_n7654_), .A2(new_n7656_), .B(pi0040), .ZN(new_n7657_));
  OAI21_X1   g04860(.A1(new_n7654_), .A2(new_n7656_), .B(new_n7657_), .ZN(new_n7658_));
  NAND2_X1   g04861(.A1(new_n7658_), .A2(new_n2794_), .ZN(new_n7659_));
  OAI21_X1   g04862(.A1(new_n7659_), .A2(new_n2436_), .B(new_n2794_), .ZN(new_n7660_));
  NAND2_X1   g04863(.A1(new_n7660_), .A2(new_n7576_), .ZN(new_n7661_));
  NOR3_X1    g04864(.A1(new_n2436_), .A2(pi0040), .A3(pi0479), .ZN(new_n7662_));
  NOR2_X1    g04865(.A1(new_n7576_), .A2(new_n2436_), .ZN(new_n7663_));
  NAND2_X1   g04866(.A1(new_n7586_), .A2(new_n2539_), .ZN(new_n7664_));
  INV_X1     g04867(.I(new_n7664_), .ZN(new_n7665_));
  AOI21_X1   g04868(.A1(new_n7665_), .A2(new_n7663_), .B(new_n7662_), .ZN(new_n7666_));
  NAND2_X1   g04869(.A1(new_n7661_), .A2(new_n7666_), .ZN(new_n7667_));
  INV_X1     g04870(.I(new_n7422_), .ZN(new_n7668_));
  AOI21_X1   g04871(.A1(new_n7647_), .A2(new_n7668_), .B(new_n7577_), .ZN(new_n7669_));
  NOR2_X1    g04872(.A1(new_n7669_), .A2(new_n2794_), .ZN(new_n7670_));
  INV_X1     g04873(.I(new_n7670_), .ZN(new_n7671_));
  NAND2_X1   g04874(.A1(new_n7659_), .A2(new_n7671_), .ZN(new_n7672_));
  NAND2_X1   g04875(.A1(new_n7672_), .A2(new_n2436_), .ZN(new_n7673_));
  NOR2_X1    g04876(.A1(new_n7673_), .A2(pi0198), .ZN(new_n7674_));
  NOR2_X1    g04877(.A1(new_n7667_), .A2(new_n7674_), .ZN(new_n7675_));
  INV_X1     g04878(.I(new_n7675_), .ZN(new_n7676_));
  NOR2_X1    g04879(.A1(new_n7676_), .A2(new_n5373_), .ZN(new_n7677_));
  NAND2_X1   g04880(.A1(new_n5373_), .A2(pi0095), .ZN(new_n7678_));
  NOR3_X1    g04881(.A1(new_n7408_), .A2(new_n5464_), .A3(new_n2479_), .ZN(new_n7679_));
  INV_X1     g04882(.I(new_n7679_), .ZN(new_n7680_));
  NAND3_X1   g04883(.A1(new_n7680_), .A2(new_n7366_), .A3(new_n7577_), .ZN(new_n7681_));
  NAND2_X1   g04884(.A1(new_n7681_), .A2(pi0032), .ZN(new_n7682_));
  NAND2_X1   g04885(.A1(new_n7682_), .A2(new_n5373_), .ZN(new_n7683_));
  XNOR2_X1   g04886(.A1(new_n7683_), .A2(new_n7678_), .ZN(new_n7684_));
  NOR2_X1    g04887(.A1(new_n7684_), .A2(new_n7577_), .ZN(new_n7685_));
  NOR2_X1    g04888(.A1(new_n7677_), .A2(new_n7685_), .ZN(new_n7686_));
  NAND2_X1   g04889(.A1(new_n2487_), .A2(new_n2496_), .ZN(new_n7687_));
  NAND2_X1   g04890(.A1(new_n7687_), .A2(new_n2448_), .ZN(new_n7688_));
  OAI21_X1   g04891(.A1(new_n2707_), .A2(new_n7688_), .B(new_n7646_), .ZN(new_n7689_));
  NAND2_X1   g04892(.A1(new_n7689_), .A2(new_n6367_), .ZN(new_n7690_));
  NAND2_X1   g04893(.A1(new_n7690_), .A2(new_n7639_), .ZN(new_n7691_));
  NOR4_X1    g04894(.A1(new_n2486_), .A2(pi0051), .A3(pi0072), .A4(pi0096), .ZN(new_n7692_));
  NAND2_X1   g04895(.A1(new_n7691_), .A2(new_n7692_), .ZN(new_n7693_));
  NOR2_X1    g04896(.A1(new_n7693_), .A2(pi0032), .ZN(new_n7694_));
  NOR2_X1    g04897(.A1(new_n2539_), .A2(pi0040), .ZN(new_n7695_));
  AOI21_X1   g04898(.A1(pi0032), .A2(new_n7695_), .B(new_n7694_), .ZN(new_n7696_));
  OAI21_X1   g04899(.A1(new_n7696_), .A2(new_n2436_), .B(new_n7577_), .ZN(new_n7697_));
  NAND2_X1   g04900(.A1(new_n7697_), .A2(new_n2959_), .ZN(new_n7698_));
  INV_X1     g04901(.I(new_n7698_), .ZN(new_n7699_));
  NOR2_X1    g04902(.A1(new_n7699_), .A2(new_n7663_), .ZN(new_n7700_));
  INV_X1     g04903(.I(new_n7700_), .ZN(new_n7701_));
  OAI21_X1   g04904(.A1(new_n7669_), .A2(pi0040), .B(pi0032), .ZN(new_n7702_));
  NOR2_X1    g04905(.A1(new_n7702_), .A2(new_n2436_), .ZN(new_n7703_));
  NOR2_X1    g04906(.A1(new_n7703_), .A2(pi0032), .ZN(new_n7704_));
  NOR2_X1    g04907(.A1(new_n7693_), .A2(new_n7704_), .ZN(new_n7705_));
  NOR2_X1    g04908(.A1(new_n7695_), .A2(new_n2436_), .ZN(new_n7706_));
  NOR2_X1    g04909(.A1(new_n7705_), .A2(new_n7706_), .ZN(new_n7707_));
  NOR2_X1    g04910(.A1(new_n7701_), .A2(new_n7707_), .ZN(new_n7708_));
  NOR2_X1    g04911(.A1(new_n7708_), .A2(pi0198), .ZN(new_n7709_));
  NOR3_X1    g04912(.A1(new_n7709_), .A2(new_n5386_), .A3(new_n7701_), .ZN(new_n7710_));
  NOR2_X1    g04913(.A1(new_n7710_), .A2(new_n7677_), .ZN(new_n7711_));
  NOR2_X1    g04914(.A1(new_n7711_), .A2(new_n7378_), .ZN(new_n7712_));
  XNOR2_X1   g04915(.A1(new_n7712_), .A2(new_n7399_), .ZN(new_n7713_));
  INV_X1     g04916(.I(new_n7713_), .ZN(new_n7714_));
  NOR2_X1    g04917(.A1(pi0180), .A2(pi0193), .ZN(new_n7715_));
  INV_X1     g04918(.I(new_n7715_), .ZN(new_n7716_));
  AOI21_X1   g04919(.A1(new_n7714_), .A2(new_n7686_), .B(new_n7716_), .ZN(new_n7717_));
  NOR2_X1    g04920(.A1(new_n7577_), .A2(new_n5386_), .ZN(new_n7718_));
  NOR2_X1    g04921(.A1(new_n7677_), .A2(new_n7718_), .ZN(new_n7719_));
  INV_X1     g04922(.I(new_n7677_), .ZN(new_n7720_));
  INV_X1     g04923(.I(new_n7688_), .ZN(new_n7721_));
  NAND2_X1   g04924(.A1(new_n2539_), .A2(pi0058), .ZN(new_n7722_));
  AOI21_X1   g04925(.A1(new_n7360_), .A2(new_n7722_), .B(new_n7580_), .ZN(new_n7723_));
  INV_X1     g04926(.I(new_n7723_), .ZN(new_n7724_));
  OAI22_X1   g04927(.A1(new_n7639_), .A2(new_n2707_), .B1(new_n7724_), .B2(new_n6368_), .ZN(new_n7725_));
  AOI21_X1   g04928(.A1(new_n7725_), .A2(new_n7721_), .B(new_n7655_), .ZN(new_n7726_));
  XNOR2_X1   g04929(.A1(new_n7726_), .A2(new_n7656_), .ZN(new_n7727_));
  NOR2_X1    g04930(.A1(new_n7727_), .A2(pi0040), .ZN(new_n7728_));
  NOR2_X1    g04931(.A1(new_n7728_), .A2(pi0032), .ZN(new_n7729_));
  INV_X1     g04932(.I(new_n7729_), .ZN(new_n7730_));
  AOI21_X1   g04933(.A1(new_n7730_), .A2(new_n7702_), .B(pi0095), .ZN(new_n7731_));
  NOR2_X1    g04934(.A1(new_n7731_), .A2(new_n7706_), .ZN(new_n7732_));
  INV_X1     g04935(.I(new_n7732_), .ZN(new_n7733_));
  NOR2_X1    g04936(.A1(new_n7733_), .A2(pi0198), .ZN(new_n7734_));
  INV_X1     g04937(.I(new_n7706_), .ZN(new_n7735_));
  OAI21_X1   g04938(.A1(new_n7728_), .A2(new_n2436_), .B(new_n2794_), .ZN(new_n7736_));
  NAND2_X1   g04939(.A1(new_n7736_), .A2(new_n7695_), .ZN(new_n7737_));
  NAND2_X1   g04940(.A1(new_n7737_), .A2(new_n7735_), .ZN(new_n7738_));
  NOR2_X1    g04941(.A1(new_n7738_), .A2(new_n3072_), .ZN(new_n7739_));
  NOR2_X1    g04942(.A1(new_n7734_), .A2(new_n7739_), .ZN(new_n7740_));
  INV_X1     g04943(.I(new_n7740_), .ZN(new_n7741_));
  OAI21_X1   g04944(.A1(new_n7428_), .A2(new_n7741_), .B(new_n7720_), .ZN(new_n7742_));
  NAND2_X1   g04945(.A1(new_n7742_), .A2(pi0183), .ZN(new_n7743_));
  XOR2_X1    g04946(.A1(new_n7743_), .A2(new_n7399_), .Z(new_n7744_));
  NOR2_X1    g04947(.A1(new_n7744_), .A2(new_n7719_), .ZN(new_n7745_));
  INV_X1     g04948(.I(new_n7745_), .ZN(new_n7746_));
  INV_X1     g04949(.I(new_n7666_), .ZN(new_n7747_));
  AOI21_X1   g04950(.A1(new_n2436_), .A2(new_n7577_), .B(new_n7747_), .ZN(new_n7748_));
  NOR2_X1    g04951(.A1(new_n7748_), .A2(new_n5386_), .ZN(new_n7749_));
  NOR2_X1    g04952(.A1(new_n7675_), .A2(new_n5373_), .ZN(new_n7750_));
  NOR2_X1    g04953(.A1(new_n7750_), .A2(new_n7749_), .ZN(new_n7751_));
  INV_X1     g04954(.I(new_n7751_), .ZN(new_n7752_));
  AOI21_X1   g04955(.A1(new_n7727_), .A2(new_n2486_), .B(pi0032), .ZN(new_n7753_));
  NAND2_X1   g04956(.A1(new_n7753_), .A2(pi0095), .ZN(new_n7754_));
  NAND2_X1   g04957(.A1(new_n7754_), .A2(new_n2794_), .ZN(new_n7755_));
  NAND2_X1   g04958(.A1(new_n7755_), .A2(new_n7576_), .ZN(new_n7756_));
  NAND2_X1   g04959(.A1(new_n7756_), .A2(new_n7666_), .ZN(new_n7757_));
  NOR2_X1    g04960(.A1(new_n7753_), .A2(new_n7670_), .ZN(new_n7758_));
  NOR2_X1    g04961(.A1(new_n7758_), .A2(pi0095), .ZN(new_n7759_));
  AOI21_X1   g04962(.A1(new_n3072_), .A2(new_n7759_), .B(new_n7757_), .ZN(new_n7760_));
  AOI21_X1   g04963(.A1(new_n5373_), .A2(new_n7760_), .B(new_n7677_), .ZN(new_n7761_));
  NAND2_X1   g04964(.A1(new_n7761_), .A2(pi0183), .ZN(new_n7762_));
  XNOR2_X1   g04965(.A1(new_n7762_), .A2(new_n7399_), .ZN(new_n7763_));
  AOI21_X1   g04966(.A1(new_n7763_), .A2(new_n7752_), .B(pi0180), .ZN(new_n7764_));
  OAI21_X1   g04967(.A1(new_n7746_), .A2(new_n7717_), .B(new_n7764_), .ZN(new_n7765_));
  NOR2_X1    g04968(.A1(new_n7682_), .A2(new_n2436_), .ZN(new_n7766_));
  OAI21_X1   g04969(.A1(new_n7747_), .A2(new_n5373_), .B(new_n7766_), .ZN(new_n7767_));
  INV_X1     g04970(.I(new_n7767_), .ZN(new_n7768_));
  OAI21_X1   g04971(.A1(new_n5386_), .A2(new_n7577_), .B(new_n7720_), .ZN(new_n7770_));
  NAND2_X1   g04972(.A1(new_n7770_), .A2(pi0174), .ZN(new_n7771_));
  XOR2_X1    g04973(.A1(new_n7771_), .A2(new_n7399_), .Z(new_n7772_));
  NOR3_X1    g04974(.A1(new_n7772_), .A2(new_n7677_), .A3(new_n7768_), .ZN(new_n7773_));
  NOR2_X1    g04975(.A1(new_n7673_), .A2(pi0210), .ZN(new_n7774_));
  NOR2_X1    g04976(.A1(new_n7667_), .A2(new_n7774_), .ZN(new_n7775_));
  INV_X1     g04977(.I(new_n7775_), .ZN(new_n7776_));
  NOR2_X1    g04978(.A1(new_n7776_), .A2(new_n5373_), .ZN(new_n7777_));
  NOR2_X1    g04979(.A1(new_n7777_), .A2(new_n7718_), .ZN(new_n7778_));
  NOR2_X1    g04980(.A1(new_n5158_), .A2(new_n3827_), .ZN(new_n7779_));
  INV_X1     g04981(.I(new_n7777_), .ZN(new_n7780_));
  OAI21_X1   g04982(.A1(new_n7577_), .A2(new_n7684_), .B(new_n7780_), .ZN(new_n7781_));
  NAND2_X1   g04983(.A1(new_n7781_), .A2(pi0172), .ZN(new_n7782_));
  XOR2_X1    g04984(.A1(new_n7782_), .A2(new_n7779_), .Z(new_n7783_));
  NOR2_X1    g04985(.A1(new_n7783_), .A2(new_n7778_), .ZN(new_n7784_));
  NAND2_X1   g04986(.A1(new_n7776_), .A2(new_n5386_), .ZN(new_n7785_));
  OAI21_X1   g04987(.A1(new_n5386_), .A2(new_n7748_), .B(new_n7785_), .ZN(new_n7786_));
  INV_X1     g04988(.I(new_n7779_), .ZN(new_n7787_));
  NAND2_X1   g04989(.A1(new_n7780_), .A2(new_n7767_), .ZN(new_n7788_));
  NAND2_X1   g04990(.A1(new_n7788_), .A2(pi0172), .ZN(new_n7789_));
  XOR2_X1    g04991(.A1(new_n7789_), .A2(new_n7787_), .Z(new_n7790_));
  NAND2_X1   g04992(.A1(new_n7790_), .A2(new_n7786_), .ZN(new_n7791_));
  NOR2_X1    g04993(.A1(new_n3098_), .A2(pi0158), .ZN(new_n7792_));
  INV_X1     g04994(.I(new_n7792_), .ZN(new_n7793_));
  OAI21_X1   g04995(.A1(new_n7475_), .A2(new_n7793_), .B(new_n7791_), .ZN(new_n7794_));
  NOR2_X1    g04996(.A1(new_n7647_), .A2(new_n2448_), .ZN(new_n7795_));
  NOR2_X1    g04997(.A1(new_n2448_), .A2(new_n2679_), .ZN(new_n7796_));
  XOR2_X1    g04998(.A1(new_n7795_), .A2(new_n7796_), .Z(new_n7797_));
  NAND2_X1   g04999(.A1(new_n7797_), .A2(new_n7642_), .ZN(new_n7798_));
  AOI21_X1   g05000(.A1(pi0093), .A2(new_n2448_), .B(new_n5464_), .ZN(new_n7799_));
  AOI21_X1   g05001(.A1(new_n5464_), .A2(new_n2539_), .B(pi0032), .ZN(new_n7800_));
  AOI21_X1   g05002(.A1(new_n7799_), .A2(new_n7800_), .B(pi0093), .ZN(new_n7801_));
  AOI21_X1   g05003(.A1(new_n2448_), .A2(pi0032), .B(pi0040), .ZN(new_n7802_));
  OAI21_X1   g05004(.A1(new_n7798_), .A2(new_n7801_), .B(new_n7802_), .ZN(new_n7803_));
  AND2_X2    g05005(.A1(new_n7803_), .A2(new_n2436_), .Z(new_n7804_));
  INV_X1     g05006(.I(new_n7804_), .ZN(new_n7805_));
  AOI21_X1   g05007(.A1(new_n7805_), .A2(new_n7666_), .B(new_n5386_), .ZN(new_n7806_));
  INV_X1     g05008(.I(new_n7806_), .ZN(new_n7807_));
  NAND2_X1   g05009(.A1(new_n7785_), .A2(new_n7807_), .ZN(new_n7808_));
  NAND2_X1   g05010(.A1(new_n7808_), .A2(pi0152), .ZN(new_n7809_));
  XOR2_X1    g05011(.A1(new_n7809_), .A2(new_n7779_), .Z(new_n7810_));
  NOR2_X1    g05012(.A1(new_n5661_), .A2(new_n3098_), .ZN(new_n7811_));
  INV_X1     g05013(.I(new_n7811_), .ZN(new_n7812_));
  OAI21_X1   g05014(.A1(new_n7798_), .A2(new_n2509_), .B(new_n7410_), .ZN(new_n7813_));
  INV_X1     g05015(.I(new_n7799_), .ZN(new_n7814_));
  NAND2_X1   g05016(.A1(new_n7800_), .A2(new_n7802_), .ZN(new_n7815_));
  AOI21_X1   g05017(.A1(new_n7814_), .A2(new_n7815_), .B(new_n2679_), .ZN(new_n7816_));
  NAND2_X1   g05018(.A1(new_n7813_), .A2(new_n7816_), .ZN(new_n7817_));
  AOI21_X1   g05019(.A1(new_n7747_), .A2(new_n5373_), .B(pi0095), .ZN(new_n7818_));
  NOR2_X1    g05020(.A1(new_n7817_), .A2(new_n7818_), .ZN(new_n7819_));
  INV_X1     g05021(.I(new_n7819_), .ZN(new_n7820_));
  NAND2_X1   g05022(.A1(new_n7785_), .A2(new_n7820_), .ZN(new_n7821_));
  NOR3_X1    g05023(.A1(new_n7810_), .A2(new_n7812_), .A3(new_n7821_), .ZN(new_n7822_));
  AOI21_X1   g05024(.A1(new_n7794_), .A2(new_n7822_), .B(new_n7784_), .ZN(new_n7823_));
  NOR2_X1    g05025(.A1(new_n7663_), .A2(new_n5386_), .ZN(new_n7824_));
  NAND2_X1   g05026(.A1(new_n7805_), .A2(new_n7824_), .ZN(new_n7825_));
  INV_X1     g05027(.I(new_n7825_), .ZN(new_n7826_));
  NOR2_X1    g05028(.A1(new_n7777_), .A2(new_n7826_), .ZN(new_n7827_));
  NAND2_X1   g05029(.A1(new_n7817_), .A2(new_n5373_), .ZN(new_n7828_));
  XNOR2_X1   g05030(.A1(new_n7828_), .A2(new_n7678_), .ZN(new_n7829_));
  OAI21_X1   g05031(.A1(new_n7577_), .A2(new_n7829_), .B(new_n7780_), .ZN(new_n7830_));
  NAND2_X1   g05032(.A1(new_n7830_), .A2(pi0152), .ZN(new_n7831_));
  XOR2_X1    g05033(.A1(new_n7831_), .A2(new_n7787_), .Z(new_n7832_));
  NAND2_X1   g05034(.A1(new_n7832_), .A2(new_n7827_), .ZN(new_n7833_));
  NOR2_X1    g05035(.A1(new_n7708_), .A2(pi0210), .ZN(new_n7834_));
  NOR2_X1    g05036(.A1(new_n7577_), .A2(new_n5386_), .ZN(new_n7835_));
  NOR2_X1    g05037(.A1(new_n7835_), .A2(new_n3827_), .ZN(new_n7836_));
  XOR2_X1    g05038(.A1(new_n7836_), .A2(new_n7787_), .Z(new_n7837_));
  INV_X1     g05039(.I(new_n7837_), .ZN(new_n7838_));
  NOR2_X1    g05040(.A1(new_n7775_), .A2(new_n5158_), .ZN(new_n7839_));
  XOR2_X1    g05041(.A1(new_n7839_), .A2(new_n7787_), .Z(new_n7840_));
  NAND2_X1   g05042(.A1(new_n7649_), .A2(new_n7724_), .ZN(new_n7841_));
  NAND2_X1   g05043(.A1(new_n7841_), .A2(new_n7642_), .ZN(new_n7842_));
  NAND2_X1   g05044(.A1(new_n7842_), .A2(new_n7641_), .ZN(new_n7843_));
  AOI21_X1   g05045(.A1(new_n7843_), .A2(new_n7639_), .B(new_n7655_), .ZN(new_n7844_));
  XNOR2_X1   g05046(.A1(new_n7844_), .A2(new_n7656_), .ZN(new_n7845_));
  NAND2_X1   g05047(.A1(new_n7845_), .A2(new_n2486_), .ZN(new_n7846_));
  NAND2_X1   g05048(.A1(new_n7846_), .A2(new_n2794_), .ZN(new_n7847_));
  NAND2_X1   g05049(.A1(new_n7847_), .A2(new_n7671_), .ZN(new_n7848_));
  NAND2_X1   g05050(.A1(new_n7848_), .A2(new_n2436_), .ZN(new_n7849_));
  NOR2_X1    g05051(.A1(new_n7849_), .A2(pi0210), .ZN(new_n7850_));
  OAI21_X1   g05052(.A1(new_n7847_), .A2(new_n2436_), .B(new_n2794_), .ZN(new_n7851_));
  NAND2_X1   g05053(.A1(new_n7851_), .A2(new_n7576_), .ZN(new_n7852_));
  NAND2_X1   g05054(.A1(new_n7852_), .A2(new_n7666_), .ZN(new_n7853_));
  NOR2_X1    g05055(.A1(new_n7853_), .A2(new_n7850_), .ZN(new_n7854_));
  INV_X1     g05056(.I(new_n7854_), .ZN(new_n7855_));
  NOR2_X1    g05057(.A1(new_n7855_), .A2(new_n5386_), .ZN(new_n7856_));
  INV_X1     g05058(.I(new_n7856_), .ZN(new_n7857_));
  NOR2_X1    g05059(.A1(new_n5386_), .A2(new_n2777_), .ZN(new_n7858_));
  OAI21_X1   g05060(.A1(new_n7759_), .A2(new_n7858_), .B(new_n7663_), .ZN(new_n7859_));
  NOR2_X1    g05061(.A1(new_n7757_), .A2(new_n7859_), .ZN(new_n7860_));
  OAI21_X1   g05062(.A1(new_n7860_), .A2(new_n5373_), .B(new_n7576_), .ZN(new_n7861_));
  INV_X1     g05063(.I(new_n7861_), .ZN(new_n7862_));
  NAND2_X1   g05064(.A1(new_n7862_), .A2(new_n7792_), .ZN(new_n7863_));
  NOR4_X1    g05065(.A1(new_n7840_), .A2(new_n7780_), .A3(new_n7857_), .A4(new_n7863_), .ZN(new_n7864_));
  AOI21_X1   g05066(.A1(new_n7864_), .A2(new_n7838_), .B(pi0149), .ZN(new_n7865_));
  OAI21_X1   g05067(.A1(new_n7823_), .A2(new_n7833_), .B(new_n7865_), .ZN(new_n7866_));
  NAND2_X1   g05068(.A1(new_n7577_), .A2(pi0095), .ZN(new_n7867_));
  AOI21_X1   g05069(.A1(new_n7780_), .A2(new_n7867_), .B(new_n7756_), .ZN(new_n7868_));
  OR3_X2     g05070(.A1(new_n7834_), .A2(new_n5386_), .A3(new_n7701_), .Z(new_n7869_));
  NAND2_X1   g05071(.A1(new_n7869_), .A2(new_n7780_), .ZN(new_n7870_));
  NAND2_X1   g05072(.A1(new_n7870_), .A2(pi0172), .ZN(new_n7871_));
  XOR2_X1    g05073(.A1(new_n7871_), .A2(new_n7787_), .Z(new_n7872_));
  INV_X1     g05074(.I(new_n7663_), .ZN(new_n7873_));
  NAND2_X1   g05075(.A1(new_n7661_), .A2(new_n7873_), .ZN(new_n7874_));
  OR2_X2     g05076(.A1(new_n7874_), .A2(new_n7774_), .Z(new_n7875_));
  OAI21_X1   g05077(.A1(new_n5386_), .A2(new_n7875_), .B(new_n7780_), .ZN(new_n7876_));
  NAND2_X1   g05078(.A1(new_n7852_), .A2(new_n7824_), .ZN(new_n7877_));
  OAI21_X1   g05079(.A1(new_n7850_), .A2(new_n7877_), .B(new_n7780_), .ZN(new_n7878_));
  NAND2_X1   g05080(.A1(new_n7878_), .A2(pi0152), .ZN(new_n7879_));
  XOR2_X1    g05081(.A1(new_n7879_), .A2(new_n7787_), .Z(new_n7880_));
  AOI22_X1   g05082(.A1(new_n7880_), .A2(new_n7876_), .B1(new_n7872_), .B2(new_n7868_), .ZN(new_n7881_));
  NOR3_X1    g05083(.A1(new_n7881_), .A2(new_n3098_), .A3(new_n7812_), .ZN(new_n7882_));
  AOI22_X1   g05084(.A1(new_n7765_), .A2(new_n7773_), .B1(new_n7866_), .B2(new_n7882_), .ZN(new_n7883_));
  NOR2_X1    g05085(.A1(new_n7820_), .A2(new_n7375_), .ZN(new_n7884_));
  NOR2_X1    g05086(.A1(new_n7378_), .A2(new_n5642_), .ZN(new_n7885_));
  INV_X1     g05087(.I(new_n7885_), .ZN(new_n7886_));
  NOR2_X1    g05088(.A1(new_n7884_), .A2(new_n7886_), .ZN(new_n7887_));
  OAI21_X1   g05089(.A1(new_n7376_), .A2(new_n7887_), .B(new_n7675_), .ZN(new_n7888_));
  NOR2_X1    g05090(.A1(new_n7849_), .A2(pi0198), .ZN(new_n7889_));
  OAI21_X1   g05091(.A1(new_n7877_), .A2(new_n7889_), .B(new_n7720_), .ZN(new_n7890_));
  NOR2_X1    g05092(.A1(new_n7890_), .A2(pi0183), .ZN(new_n7891_));
  NOR2_X1    g05093(.A1(new_n7677_), .A2(new_n7826_), .ZN(new_n7892_));
  AOI21_X1   g05094(.A1(pi0183), .A2(new_n7892_), .B(new_n7891_), .ZN(new_n7893_));
  NAND2_X1   g05095(.A1(new_n7893_), .A2(pi0180), .ZN(new_n7894_));
  XOR2_X1    g05096(.A1(new_n7894_), .A2(new_n7885_), .Z(new_n7895_));
  NOR2_X1    g05097(.A1(new_n7874_), .A2(new_n7674_), .ZN(new_n7896_));
  AOI21_X1   g05098(.A1(new_n7427_), .A2(new_n7896_), .B(new_n7677_), .ZN(new_n7897_));
  AND2_X2    g05099(.A1(new_n7897_), .A2(new_n7375_), .Z(new_n7898_));
  NOR2_X1    g05100(.A1(new_n7829_), .A2(new_n7577_), .ZN(new_n7899_));
  NOR3_X1    g05101(.A1(new_n7677_), .A2(new_n7375_), .A3(new_n7899_), .ZN(new_n7900_));
  OAI21_X1   g05102(.A1(new_n7898_), .A2(new_n7900_), .B(pi0193), .ZN(new_n7901_));
  OAI21_X1   g05103(.A1(new_n7895_), .A2(new_n7901_), .B(new_n7888_), .ZN(new_n7902_));
  NAND2_X1   g05104(.A1(new_n7501_), .A2(pi0164), .ZN(new_n7903_));
  OAI21_X1   g05105(.A1(new_n7667_), .A2(new_n5551_), .B(new_n7673_), .ZN(new_n7904_));
  NAND2_X1   g05106(.A1(new_n7904_), .A2(new_n5469_), .ZN(new_n7905_));
  INV_X1     g05107(.I(new_n7905_), .ZN(new_n7906_));
  NOR2_X1    g05108(.A1(new_n7906_), .A2(pi0039), .ZN(new_n7907_));
  NAND2_X1   g05109(.A1(new_n7666_), .A2(new_n7378_), .ZN(new_n7908_));
  NAND4_X1   g05110(.A1(new_n7908_), .A2(pi0038), .A3(pi0095), .A4(pi0232), .ZN(new_n7909_));
  NOR4_X1    g05111(.A1(new_n7893_), .A2(new_n7903_), .A3(new_n7907_), .A4(new_n7909_), .ZN(new_n7910_));
  AND2_X2    g05112(.A1(new_n7902_), .A2(new_n7910_), .Z(new_n7911_));
  INV_X1     g05113(.I(new_n7911_), .ZN(new_n7912_));
  OAI21_X1   g05114(.A1(new_n7912_), .A2(new_n7883_), .B(new_n7638_), .ZN(new_n7913_));
  OR3_X2     g05115(.A1(new_n7912_), .A2(new_n7638_), .A3(new_n7883_), .Z(new_n7914_));
  NAND3_X1   g05116(.A1(new_n7914_), .A2(pi0100), .A3(new_n7913_), .ZN(new_n7915_));
  XOR2_X1    g05117(.A1(new_n7915_), .A2(new_n3477_), .Z(new_n7916_));
  NOR3_X1    g05118(.A1(new_n7552_), .A2(new_n3259_), .A3(new_n3185_), .ZN(new_n7917_));
  OAI21_X1   g05119(.A1(new_n7917_), .A2(new_n7576_), .B(new_n7556_), .ZN(new_n7918_));
  AOI21_X1   g05120(.A1(new_n7588_), .A2(new_n3183_), .B(new_n7918_), .ZN(new_n7919_));
  NAND3_X1   g05121(.A1(new_n7550_), .A2(pi0038), .A3(pi0100), .ZN(new_n7920_));
  NAND2_X1   g05122(.A1(new_n7551_), .A2(new_n5486_), .ZN(new_n7921_));
  AOI21_X1   g05123(.A1(new_n7921_), .A2(new_n7920_), .B(new_n7577_), .ZN(new_n7922_));
  AOI21_X1   g05124(.A1(new_n7922_), .A2(pi0100), .B(new_n7554_), .ZN(new_n7923_));
  OAI21_X1   g05125(.A1(new_n7919_), .A2(new_n7923_), .B(pi0075), .ZN(new_n7924_));
  XOR2_X1    g05126(.A1(new_n7924_), .A2(new_n3483_), .Z(new_n7925_));
  AOI21_X1   g05127(.A1(new_n7925_), .A2(new_n7544_), .B(new_n3115_), .ZN(new_n7926_));
  NAND2_X1   g05128(.A1(new_n7545_), .A2(new_n3303_), .ZN(new_n7927_));
  NOR2_X1    g05129(.A1(new_n3115_), .A2(new_n3235_), .ZN(new_n7928_));
  NAND4_X1   g05130(.A1(new_n7548_), .A2(new_n7922_), .A3(new_n7927_), .A4(new_n7928_), .ZN(new_n7929_));
  XNOR2_X1   g05131(.A1(new_n7926_), .A2(new_n7929_), .ZN(new_n7930_));
  AOI21_X1   g05132(.A1(new_n7547_), .A2(new_n3258_), .B(new_n3175_), .ZN(new_n7931_));
  AOI21_X1   g05133(.A1(new_n7930_), .A2(new_n7931_), .B(new_n3225_), .ZN(new_n7932_));
  NOR2_X1    g05134(.A1(new_n7588_), .A2(new_n3192_), .ZN(new_n7933_));
  OAI21_X1   g05135(.A1(new_n7518_), .A2(new_n7529_), .B(new_n7527_), .ZN(new_n7934_));
  NAND2_X1   g05136(.A1(new_n7577_), .A2(new_n3133_), .ZN(new_n7935_));
  NAND4_X1   g05137(.A1(new_n7933_), .A2(new_n7522_), .A3(new_n7934_), .A4(new_n7935_), .ZN(new_n7936_));
  NAND2_X1   g05138(.A1(new_n7527_), .A2(new_n3455_), .ZN(new_n7937_));
  NOR2_X1    g05139(.A1(new_n7577_), .A2(new_n3133_), .ZN(new_n7938_));
  AOI21_X1   g05140(.A1(new_n7937_), .A2(new_n7938_), .B(new_n3188_), .ZN(new_n7939_));
  NAND2_X1   g05141(.A1(new_n7936_), .A2(new_n7939_), .ZN(new_n7940_));
  NOR2_X1    g05142(.A1(new_n7577_), .A2(pi0038), .ZN(new_n7941_));
  INV_X1     g05143(.I(new_n7941_), .ZN(new_n7942_));
  NOR2_X1    g05144(.A1(new_n7942_), .A2(new_n7538_), .ZN(new_n7943_));
  NAND3_X1   g05145(.A1(new_n7943_), .A2(new_n3202_), .A3(new_n3226_), .ZN(new_n7944_));
  NAND3_X1   g05146(.A1(new_n7570_), .A2(new_n7572_), .A3(new_n7944_), .ZN(new_n7945_));
  NAND3_X1   g05147(.A1(new_n7534_), .A2(new_n7536_), .A3(new_n7539_), .ZN(new_n7946_));
  AOI21_X1   g05148(.A1(new_n7542_), .A2(pi0074), .B(pi0054), .ZN(new_n7947_));
  NOR3_X1    g05149(.A1(new_n7947_), .A2(new_n7946_), .A3(new_n7514_), .ZN(new_n7948_));
  NAND3_X1   g05150(.A1(new_n7940_), .A2(new_n7945_), .A3(new_n7948_), .ZN(new_n7949_));
  OR3_X2     g05151(.A1(new_n7916_), .A2(new_n7932_), .A3(new_n7949_), .Z(new_n7950_));
  INV_X1     g05152(.I(pi0034), .ZN(new_n7951_));
  INV_X1     g05153(.I(pi0079), .ZN(new_n7952_));
  INV_X1     g05154(.I(pi0118), .ZN(new_n7953_));
  INV_X1     g05155(.I(pi0138), .ZN(new_n7954_));
  INV_X1     g05156(.I(pi0139), .ZN(new_n7955_));
  INV_X1     g05157(.I(pi0195), .ZN(new_n7956_));
  INV_X1     g05158(.I(pi0196), .ZN(new_n7957_));
  NOR4_X1    g05159(.A1(new_n7954_), .A2(new_n7955_), .A3(new_n7956_), .A4(new_n7957_), .ZN(new_n7958_));
  INV_X1     g05160(.I(new_n7958_), .ZN(new_n7959_));
  NOR4_X1    g05161(.A1(new_n7959_), .A2(new_n7951_), .A3(new_n7952_), .A4(new_n7953_), .ZN(new_n7960_));
  NOR2_X1    g05162(.A1(new_n7960_), .A2(pi0033), .ZN(new_n7961_));
  NAND2_X1   g05163(.A1(new_n7950_), .A2(new_n7961_), .ZN(new_n7962_));
  NAND2_X1   g05164(.A1(new_n7961_), .A2(pi0954), .ZN(new_n7963_));
  XOR2_X1    g05165(.A1(new_n7962_), .A2(new_n7963_), .Z(new_n7964_));
  NAND2_X1   g05166(.A1(new_n7950_), .A2(pi0954), .ZN(new_n7965_));
  NAND2_X1   g05167(.A1(pi0033), .A2(pi0954), .ZN(new_n7966_));
  XOR2_X1    g05168(.A1(new_n7965_), .A2(new_n7966_), .Z(new_n7967_));
  OAI21_X1   g05169(.A1(new_n7964_), .A2(new_n7967_), .B(new_n7575_), .ZN(po0191));
  INV_X1     g05170(.I(pi0144), .ZN(new_n7969_));
  NOR2_X1    g05171(.A1(new_n7480_), .A2(new_n3089_), .ZN(new_n7970_));
  INV_X1     g05172(.I(pi0140), .ZN(new_n7971_));
  NOR2_X1    g05173(.A1(new_n7971_), .A2(new_n3089_), .ZN(new_n7972_));
  XNOR2_X1   g05174(.A1(new_n7970_), .A2(new_n7972_), .ZN(new_n7973_));
  NOR2_X1    g05175(.A1(new_n7349_), .A2(pi0140), .ZN(new_n7974_));
  NAND2_X1   g05176(.A1(new_n7396_), .A2(new_n7972_), .ZN(new_n7975_));
  OAI21_X1   g05177(.A1(new_n7975_), .A2(new_n7974_), .B(new_n7419_), .ZN(new_n7976_));
  AOI22_X1   g05178(.A1(new_n7976_), .A2(new_n7972_), .B1(pi0144), .B2(new_n5373_), .ZN(new_n7977_));
  OAI22_X1   g05179(.A1(new_n7973_), .A2(new_n7430_), .B1(new_n7969_), .B2(new_n7977_), .ZN(new_n7978_));
  NOR2_X1    g05180(.A1(new_n7374_), .A2(pi0140), .ZN(new_n7979_));
  NOR3_X1    g05181(.A1(new_n7979_), .A2(new_n3089_), .A3(new_n7386_), .ZN(new_n7980_));
  AOI21_X1   g05182(.A1(new_n7980_), .A2(new_n7978_), .B(pi0299), .ZN(new_n7981_));
  NAND2_X1   g05183(.A1(new_n7435_), .A2(pi0181), .ZN(new_n7982_));
  NOR2_X1    g05184(.A1(new_n3211_), .A2(pi0232), .ZN(new_n7983_));
  OAI21_X1   g05185(.A1(new_n7981_), .A2(new_n7982_), .B(new_n7983_), .ZN(new_n7984_));
  OAI21_X1   g05186(.A1(new_n7470_), .A2(new_n4981_), .B(new_n7386_), .ZN(new_n7985_));
  NAND2_X1   g05187(.A1(new_n5373_), .A2(pi0162), .ZN(new_n7986_));
  NOR2_X1    g05188(.A1(new_n7986_), .A2(new_n2847_), .ZN(new_n7987_));
  OAI21_X1   g05189(.A1(new_n7473_), .A2(new_n4981_), .B(new_n7395_), .ZN(new_n7988_));
  AOI21_X1   g05190(.A1(new_n7988_), .A2(pi0146), .B(pi0299), .ZN(new_n7989_));
  NAND3_X1   g05191(.A1(new_n7436_), .A2(new_n5662_), .A3(new_n3098_), .ZN(new_n7990_));
  NAND4_X1   g05192(.A1(new_n7990_), .A2(pi0159), .A3(pi0162), .A4(new_n2827_), .ZN(new_n7991_));
  NOR2_X1    g05193(.A1(new_n7480_), .A2(new_n2847_), .ZN(new_n7992_));
  NOR2_X1    g05194(.A1(new_n2847_), .A2(new_n4981_), .ZN(new_n7993_));
  XOR2_X1    g05195(.A1(new_n7992_), .A2(new_n7993_), .Z(new_n7994_));
  NAND2_X1   g05196(.A1(new_n7994_), .A2(new_n7429_), .ZN(new_n7995_));
  NOR2_X1    g05197(.A1(new_n7418_), .A2(pi0161), .ZN(new_n7996_));
  AOI21_X1   g05198(.A1(new_n7995_), .A2(new_n7996_), .B(new_n2847_), .ZN(new_n7997_));
  OAI22_X1   g05199(.A1(new_n7997_), .A2(pi0162), .B1(new_n7989_), .B2(new_n7991_), .ZN(new_n7998_));
  AOI21_X1   g05200(.A1(new_n7985_), .A2(new_n7987_), .B(new_n7998_), .ZN(new_n7999_));
  INV_X1     g05201(.I(pi0188), .ZN(new_n8000_));
  INV_X1     g05202(.I(new_n7490_), .ZN(new_n8001_));
  NAND2_X1   g05203(.A1(new_n8001_), .A2(pi0188), .ZN(new_n8002_));
  NAND3_X1   g05204(.A1(new_n7494_), .A2(pi0167), .A3(pi0188), .ZN(new_n8003_));
  XOR2_X1    g05205(.A1(new_n8003_), .A2(new_n8002_), .Z(new_n8004_));
  AOI21_X1   g05206(.A1(new_n8004_), .A2(pi0038), .B(pi0167), .ZN(new_n8005_));
  NOR3_X1    g05207(.A1(new_n8005_), .A2(new_n8000_), .A3(new_n7500_), .ZN(new_n8006_));
  OR2_X2     g05208(.A1(new_n8006_), .A2(pi0100), .Z(new_n8007_));
  AOI21_X1   g05209(.A1(new_n7999_), .A2(new_n7984_), .B(new_n8007_), .ZN(new_n8008_));
  INV_X1     g05210(.I(new_n7453_), .ZN(new_n8009_));
  INV_X1     g05211(.I(pi0177), .ZN(new_n8010_));
  NOR2_X1    g05212(.A1(new_n8010_), .A2(pi0299), .ZN(new_n8011_));
  NAND2_X1   g05213(.A1(new_n7454_), .A2(new_n8011_), .ZN(new_n8012_));
  NAND2_X1   g05214(.A1(new_n8011_), .A2(pi0144), .ZN(new_n8013_));
  XOR2_X1    g05215(.A1(new_n8012_), .A2(new_n8013_), .Z(new_n8014_));
  NAND2_X1   g05216(.A1(new_n3259_), .A2(new_n5551_), .ZN(new_n8015_));
  AOI21_X1   g05217(.A1(new_n8014_), .A2(new_n8009_), .B(new_n8015_), .ZN(new_n8016_));
  NAND2_X1   g05218(.A1(new_n8010_), .A2(new_n3098_), .ZN(new_n8017_));
  NAND4_X1   g05219(.A1(new_n7463_), .A2(pi0039), .A3(pi0144), .A4(new_n8017_), .ZN(new_n8018_));
  OAI21_X1   g05220(.A1(new_n8016_), .A2(new_n8018_), .B(new_n3098_), .ZN(new_n8019_));
  INV_X1     g05221(.I(pi0155), .ZN(new_n8020_));
  NAND2_X1   g05222(.A1(new_n7443_), .A2(new_n7439_), .ZN(new_n8021_));
  NAND2_X1   g05223(.A1(new_n7439_), .A2(pi0161), .ZN(new_n8022_));
  XOR2_X1    g05224(.A1(new_n8021_), .A2(new_n8022_), .Z(new_n8023_));
  AOI21_X1   g05225(.A1(new_n8023_), .A2(new_n7446_), .B(new_n8020_), .ZN(new_n8024_));
  NOR2_X1    g05226(.A1(new_n3259_), .A2(new_n8020_), .ZN(new_n8025_));
  XOR2_X1    g05227(.A1(new_n8024_), .A2(new_n8025_), .Z(new_n8026_));
  NOR2_X1    g05228(.A1(new_n7440_), .A2(pi0161), .ZN(new_n8027_));
  NAND4_X1   g05229(.A1(new_n8026_), .A2(new_n7445_), .A3(new_n8019_), .A4(new_n8027_), .ZN(new_n8028_));
  INV_X1     g05230(.I(pi0167), .ZN(new_n8029_));
  NAND2_X1   g05231(.A1(new_n6493_), .A2(new_n8029_), .ZN(new_n8030_));
  XOR2_X1    g05232(.A1(new_n7492_), .A2(new_n8030_), .Z(new_n8031_));
  NOR2_X1    g05233(.A1(new_n8031_), .A2(new_n8000_), .ZN(new_n8032_));
  NOR2_X1    g05234(.A1(new_n8032_), .A2(pi0100), .ZN(new_n8033_));
  XOR2_X1    g05235(.A1(pi0140), .A2(pi0145), .Z(new_n8034_));
  OAI21_X1   g05236(.A1(pi0178), .A2(pi0183), .B(new_n5373_), .ZN(new_n8035_));
  OAI21_X1   g05237(.A1(new_n8034_), .A2(new_n8035_), .B(new_n3098_), .ZN(new_n8036_));
  NOR2_X1    g05238(.A1(pi0178), .A2(pi0183), .ZN(new_n8037_));
  NOR4_X1    g05239(.A1(new_n5386_), .A2(new_n7971_), .A3(new_n5641_), .A4(new_n8037_), .ZN(new_n8038_));
  AOI21_X1   g05240(.A1(new_n8036_), .A2(new_n8038_), .B(pi0232), .ZN(new_n8039_));
  NOR2_X1    g05241(.A1(pi0149), .A2(pi0157), .ZN(new_n8040_));
  XOR2_X1    g05242(.A1(pi0162), .A2(pi0197), .Z(new_n8041_));
  XOR2_X1    g05243(.A1(new_n8041_), .A2(new_n5373_), .Z(new_n8042_));
  NAND3_X1   g05244(.A1(new_n8042_), .A2(pi0299), .A3(new_n8040_), .ZN(new_n8043_));
  NOR2_X1    g05245(.A1(new_n8043_), .A2(new_n8039_), .ZN(new_n8044_));
  NOR2_X1    g05246(.A1(new_n8044_), .A2(new_n3462_), .ZN(new_n8045_));
  NAND2_X1   g05247(.A1(new_n3133_), .A2(new_n3455_), .ZN(new_n8046_));
  OAI21_X1   g05248(.A1(new_n8045_), .A2(new_n8046_), .B(new_n8033_), .ZN(new_n8047_));
  OAI22_X1   g05249(.A1(new_n8008_), .A2(new_n8028_), .B1(new_n3455_), .B2(new_n8047_), .ZN(new_n8048_));
  INV_X1     g05250(.I(new_n8044_), .ZN(new_n8049_));
  NOR3_X1    g05251(.A1(new_n3259_), .A2(new_n8029_), .A3(new_n3098_), .ZN(new_n8050_));
  NOR3_X1    g05252(.A1(new_n3259_), .A2(pi0167), .A3(pi0299), .ZN(new_n8051_));
  NOR2_X1    g05253(.A1(new_n6494_), .A2(new_n8000_), .ZN(new_n8052_));
  OAI21_X1   g05254(.A1(new_n8050_), .A2(new_n8051_), .B(new_n8052_), .ZN(new_n8053_));
  NAND2_X1   g05255(.A1(new_n3140_), .A2(new_n8053_), .ZN(new_n8054_));
  NAND3_X1   g05256(.A1(new_n3211_), .A2(pi0155), .A3(pi0299), .ZN(new_n8055_));
  NAND3_X1   g05257(.A1(new_n3211_), .A2(new_n8020_), .A3(new_n3098_), .ZN(new_n8056_));
  AOI21_X1   g05258(.A1(new_n8055_), .A2(new_n8056_), .B(new_n8010_), .ZN(new_n8057_));
  AOI21_X1   g05259(.A1(new_n8054_), .A2(new_n8057_), .B(new_n3462_), .ZN(new_n8058_));
  XNOR2_X1   g05260(.A1(new_n8058_), .A2(new_n3477_), .ZN(new_n8059_));
  NOR2_X1    g05261(.A1(new_n8044_), .A2(new_n3235_), .ZN(new_n8060_));
  INV_X1     g05262(.I(new_n8060_), .ZN(new_n8061_));
  OAI22_X1   g05263(.A1(new_n8059_), .A2(new_n8049_), .B1(new_n7529_), .B2(new_n8061_), .ZN(new_n8062_));
  NOR2_X1    g05264(.A1(new_n8047_), .A2(new_n3115_), .ZN(new_n8063_));
  AOI21_X1   g05265(.A1(new_n8062_), .A2(new_n8063_), .B(new_n3188_), .ZN(new_n8064_));
  NOR3_X1    g05266(.A1(new_n8064_), .A2(new_n3462_), .A3(new_n8044_), .ZN(new_n8065_));
  NOR2_X1    g05267(.A1(new_n8045_), .A2(new_n8060_), .ZN(new_n8066_));
  NOR2_X1    g05268(.A1(pi0141), .A2(pi0299), .ZN(new_n8067_));
  AOI21_X1   g05269(.A1(new_n4329_), .A2(pi0299), .B(new_n8067_), .ZN(new_n8068_));
  AND2_X2    g05270(.A1(new_n6493_), .A2(new_n8068_), .Z(new_n8069_));
  OAI21_X1   g05271(.A1(new_n7538_), .A2(new_n8069_), .B(new_n8066_), .ZN(new_n8070_));
  NOR3_X1    g05272(.A1(new_n8070_), .A2(pi0055), .A3(new_n3175_), .ZN(new_n8071_));
  AOI21_X1   g05273(.A1(new_n8048_), .A2(new_n8065_), .B(new_n8071_), .ZN(new_n8072_));
  AOI21_X1   g05274(.A1(new_n8066_), .A2(pi0054), .B(new_n8033_), .ZN(new_n8073_));
  NOR2_X1    g05275(.A1(new_n8073_), .A2(new_n3235_), .ZN(new_n8074_));
  NAND4_X1   g05276(.A1(new_n7467_), .A2(pi0092), .A3(pi0162), .A4(new_n7523_), .ZN(new_n8075_));
  NOR3_X1    g05277(.A1(new_n6494_), .A2(new_n3259_), .A3(new_n8029_), .ZN(new_n8076_));
  NAND2_X1   g05278(.A1(new_n8076_), .A2(new_n7537_), .ZN(new_n8077_));
  NAND2_X1   g05279(.A1(new_n8077_), .A2(new_n8075_), .ZN(new_n8078_));
  AOI21_X1   g05280(.A1(new_n5440_), .A2(new_n8078_), .B(new_n3115_), .ZN(new_n8079_));
  NAND3_X1   g05281(.A1(new_n8042_), .A2(pi0232), .A3(new_n8040_), .ZN(new_n8080_));
  NOR2_X1    g05282(.A1(new_n8080_), .A2(new_n7537_), .ZN(new_n8081_));
  NAND2_X1   g05283(.A1(new_n8081_), .A2(pi0054), .ZN(new_n8082_));
  XNOR2_X1   g05284(.A1(new_n8079_), .A2(new_n8082_), .ZN(new_n8083_));
  NAND2_X1   g05285(.A1(new_n7539_), .A2(pi0167), .ZN(new_n8084_));
  INV_X1     g05286(.I(new_n8084_), .ZN(new_n8085_));
  INV_X1     g05287(.I(new_n8080_), .ZN(new_n8086_));
  NOR4_X1    g05288(.A1(new_n6494_), .A2(new_n7538_), .A3(new_n3175_), .A4(new_n4329_), .ZN(new_n8087_));
  OR2_X2     g05289(.A1(new_n8087_), .A2(new_n3258_), .Z(new_n8088_));
  OAI21_X1   g05290(.A1(new_n8088_), .A2(new_n3226_), .B(new_n3175_), .ZN(new_n8089_));
  AND3_X2    g05291(.A1(new_n8083_), .A2(new_n8085_), .A3(new_n8089_), .Z(new_n8090_));
  NOR2_X1    g05292(.A1(new_n8084_), .A2(new_n3259_), .ZN(new_n8091_));
  OAI21_X1   g05293(.A1(new_n8081_), .A2(pi0054), .B(new_n8091_), .ZN(new_n8092_));
  NOR2_X1    g05294(.A1(new_n8081_), .A2(new_n8085_), .ZN(new_n8093_));
  AOI21_X1   g05295(.A1(new_n8093_), .A2(new_n3175_), .B(new_n8087_), .ZN(new_n8094_));
  NAND2_X1   g05296(.A1(new_n8094_), .A2(new_n3225_), .ZN(new_n8095_));
  NAND2_X1   g05297(.A1(new_n8095_), .A2(new_n8092_), .ZN(new_n8096_));
  AOI21_X1   g05298(.A1(new_n8096_), .A2(pi0074), .B(new_n3426_), .ZN(new_n8097_));
  INV_X1     g05299(.I(new_n8097_), .ZN(new_n8098_));
  NAND2_X1   g05300(.A1(new_n8094_), .A2(new_n3426_), .ZN(new_n8099_));
  NOR2_X1    g05301(.A1(new_n8098_), .A2(new_n8099_), .ZN(new_n8100_));
  OAI21_X1   g05302(.A1(new_n8090_), .A2(new_n8100_), .B(new_n8074_), .ZN(new_n8101_));
  NOR2_X1    g05303(.A1(new_n8072_), .A2(new_n8101_), .ZN(new_n8102_));
  NAND2_X1   g05304(.A1(new_n7943_), .A2(new_n3202_), .ZN(new_n8103_));
  AOI21_X1   g05305(.A1(new_n8103_), .A2(new_n3226_), .B(new_n3426_), .ZN(new_n8104_));
  NOR2_X1    g05306(.A1(new_n7827_), .A2(new_n2847_), .ZN(new_n8105_));
  XNOR2_X1   g05307(.A1(new_n8105_), .A2(new_n7993_), .ZN(new_n8106_));
  NOR2_X1    g05308(.A1(new_n8106_), .A2(new_n7778_), .ZN(new_n8107_));
  INV_X1     g05309(.I(pi0162), .ZN(new_n8108_));
  NOR2_X1    g05310(.A1(new_n5662_), .A2(new_n3098_), .ZN(new_n8109_));
  INV_X1     g05311(.I(new_n8109_), .ZN(new_n8110_));
  NAND2_X1   g05312(.A1(new_n8110_), .A2(new_n8108_), .ZN(new_n8111_));
  NAND2_X1   g05313(.A1(new_n7830_), .A2(pi0161), .ZN(new_n8112_));
  XOR2_X1    g05314(.A1(new_n8112_), .A2(new_n7993_), .Z(new_n8113_));
  NOR2_X1    g05315(.A1(new_n8113_), .A2(new_n7781_), .ZN(new_n8114_));
  OAI21_X1   g05316(.A1(new_n8107_), .A2(new_n8111_), .B(new_n8114_), .ZN(new_n8115_));
  NAND2_X1   g05317(.A1(new_n7878_), .A2(pi0146), .ZN(new_n8116_));
  XNOR2_X1   g05318(.A1(new_n8116_), .A2(new_n7993_), .ZN(new_n8117_));
  AOI21_X1   g05319(.A1(new_n8117_), .A2(new_n7868_), .B(pi0162), .ZN(new_n8118_));
  NAND2_X1   g05320(.A1(new_n7870_), .A2(pi0161), .ZN(new_n8119_));
  XNOR2_X1   g05321(.A1(new_n8119_), .A2(new_n7993_), .ZN(new_n8120_));
  NAND2_X1   g05322(.A1(new_n8120_), .A2(new_n7876_), .ZN(new_n8121_));
  AOI21_X1   g05323(.A1(new_n8115_), .A2(new_n8118_), .B(new_n8121_), .ZN(new_n8122_));
  NOR2_X1    g05324(.A1(new_n7892_), .A2(new_n7971_), .ZN(new_n8123_));
  XNOR2_X1   g05325(.A1(new_n8123_), .A2(new_n7972_), .ZN(new_n8124_));
  NAND2_X1   g05326(.A1(new_n7890_), .A2(pi0142), .ZN(new_n8125_));
  XOR2_X1    g05327(.A1(new_n8125_), .A2(new_n7972_), .Z(new_n8126_));
  OAI22_X1   g05328(.A1(new_n8126_), .A2(new_n7742_), .B1(new_n7719_), .B2(new_n8124_), .ZN(new_n8127_));
  NAND2_X1   g05329(.A1(new_n8127_), .A2(pi0181), .ZN(new_n8128_));
  NAND3_X1   g05330(.A1(new_n8128_), .A2(new_n7969_), .A3(new_n3098_), .ZN(new_n8129_));
  NOR3_X1    g05331(.A1(new_n7750_), .A2(pi0140), .A3(pi0142), .ZN(new_n8130_));
  NOR2_X1    g05332(.A1(new_n7853_), .A2(new_n7889_), .ZN(new_n8131_));
  NAND3_X1   g05333(.A1(new_n7675_), .A2(pi0142), .A3(new_n5373_), .ZN(new_n8132_));
  NAND3_X1   g05334(.A1(new_n7676_), .A2(pi0142), .A3(new_n5386_), .ZN(new_n8133_));
  NAND2_X1   g05335(.A1(new_n8133_), .A2(new_n8132_), .ZN(new_n8134_));
  AOI21_X1   g05336(.A1(new_n8134_), .A2(new_n8131_), .B(pi0140), .ZN(new_n8135_));
  OR3_X2     g05337(.A1(new_n7761_), .A2(new_n3089_), .A3(new_n5643_), .Z(new_n8136_));
  OAI22_X1   g05338(.A1(new_n8136_), .A2(new_n8135_), .B1(new_n7807_), .B2(new_n8130_), .ZN(new_n8137_));
  NOR2_X1    g05339(.A1(new_n7897_), .A2(new_n3089_), .ZN(new_n8138_));
  XOR2_X1    g05340(.A1(new_n8138_), .A2(new_n7972_), .Z(new_n8139_));
  AOI22_X1   g05341(.A1(new_n8139_), .A2(new_n7711_), .B1(pi0144), .B2(pi0181), .ZN(new_n8140_));
  OAI21_X1   g05342(.A1(new_n7677_), .A2(new_n7899_), .B(pi0140), .ZN(new_n8141_));
  XNOR2_X1   g05343(.A1(new_n8141_), .A2(new_n7972_), .ZN(new_n8142_));
  NAND4_X1   g05344(.A1(new_n8142_), .A2(new_n3089_), .A3(new_n7686_), .A4(new_n7751_), .ZN(new_n8143_));
  NOR2_X1    g05345(.A1(new_n8140_), .A2(new_n8143_), .ZN(new_n8144_));
  NAND3_X1   g05346(.A1(new_n8129_), .A2(new_n8137_), .A3(new_n8144_), .ZN(new_n8145_));
  NOR2_X1    g05347(.A1(new_n7677_), .A2(new_n7768_), .ZN(new_n8146_));
  NAND2_X1   g05348(.A1(new_n7770_), .A2(pi0142), .ZN(new_n8147_));
  XOR2_X1    g05349(.A1(new_n8147_), .A2(new_n7972_), .Z(new_n8148_));
  NOR4_X1    g05350(.A1(new_n8148_), .A2(new_n7676_), .A3(new_n7820_), .A4(new_n8130_), .ZN(new_n8149_));
  OAI21_X1   g05351(.A1(new_n8149_), .A2(pi0142), .B(new_n8146_), .ZN(new_n8150_));
  AOI21_X1   g05352(.A1(new_n8145_), .A2(new_n5643_), .B(new_n8150_), .ZN(new_n8151_));
  NAND2_X1   g05353(.A1(new_n7788_), .A2(pi0161), .ZN(new_n8152_));
  XOR2_X1    g05354(.A1(new_n8152_), .A2(new_n7993_), .Z(new_n8153_));
  NOR2_X1    g05355(.A1(new_n7835_), .A2(new_n4981_), .ZN(new_n8154_));
  XNOR2_X1   g05356(.A1(new_n8154_), .A2(new_n7993_), .ZN(new_n8155_));
  NOR2_X1    g05357(.A1(new_n7775_), .A2(new_n2847_), .ZN(new_n8156_));
  XOR2_X1    g05358(.A1(new_n8156_), .A2(new_n7993_), .Z(new_n8157_));
  NOR2_X1    g05359(.A1(new_n7861_), .A2(new_n8108_), .ZN(new_n8158_));
  NAND4_X1   g05360(.A1(new_n8157_), .A2(new_n7777_), .A3(new_n7856_), .A4(new_n8158_), .ZN(new_n8159_));
  OAI22_X1   g05361(.A1(new_n8153_), .A2(new_n7821_), .B1(new_n8155_), .B2(new_n8159_), .ZN(new_n8160_));
  NAND2_X1   g05362(.A1(new_n7808_), .A2(pi0146), .ZN(new_n8161_));
  XNOR2_X1   g05363(.A1(new_n8161_), .A2(new_n7993_), .ZN(new_n8162_));
  OAI21_X1   g05364(.A1(new_n7905_), .A2(new_n3212_), .B(new_n5551_), .ZN(new_n8163_));
  OAI21_X1   g05365(.A1(new_n7629_), .A2(new_n3259_), .B(new_n5551_), .ZN(new_n8164_));
  NAND2_X1   g05366(.A1(new_n7600_), .A2(new_n8011_), .ZN(new_n8165_));
  NAND3_X1   g05367(.A1(new_n7601_), .A2(new_n7969_), .A3(new_n7635_), .ZN(new_n8166_));
  NAND4_X1   g05368(.A1(new_n8166_), .A2(new_n8010_), .A3(new_n3098_), .A4(new_n7595_), .ZN(new_n8167_));
  OAI21_X1   g05369(.A1(new_n8167_), .A2(new_n8165_), .B(new_n7969_), .ZN(new_n8168_));
  NAND4_X1   g05370(.A1(new_n8164_), .A2(new_n8168_), .A3(pi0039), .A4(new_n7626_), .ZN(new_n8169_));
  NOR2_X1    g05371(.A1(pi0038), .A2(pi0155), .ZN(new_n8170_));
  INV_X1     g05372(.I(new_n8170_), .ZN(new_n8171_));
  AOI21_X1   g05373(.A1(new_n7604_), .A2(new_n8171_), .B(new_n8022_), .ZN(new_n8172_));
  OAI21_X1   g05374(.A1(new_n7627_), .A2(new_n7614_), .B(new_n8172_), .ZN(new_n8173_));
  NAND2_X1   g05375(.A1(new_n3259_), .A2(pi0155), .ZN(new_n8174_));
  NAND3_X1   g05376(.A1(new_n8173_), .A2(new_n7604_), .A3(new_n8174_), .ZN(new_n8175_));
  NAND2_X1   g05377(.A1(new_n7610_), .A2(new_n7440_), .ZN(new_n8176_));
  NOR2_X1    g05378(.A1(new_n3098_), .A2(pi0159), .ZN(new_n8177_));
  INV_X1     g05379(.I(new_n8177_), .ZN(new_n8178_));
  NOR4_X1    g05380(.A1(new_n7607_), .A2(new_n3455_), .A3(new_n4981_), .A4(new_n8178_), .ZN(new_n8179_));
  NAND4_X1   g05381(.A1(new_n8175_), .A2(new_n8006_), .A3(new_n8176_), .A4(new_n8179_), .ZN(new_n8180_));
  AOI21_X1   g05382(.A1(new_n8169_), .A2(new_n5551_), .B(new_n8180_), .ZN(new_n8181_));
  AND3_X2    g05383(.A1(new_n7786_), .A2(new_n8163_), .A3(new_n8181_), .Z(new_n8182_));
  AND3_X2    g05384(.A1(new_n8160_), .A2(new_n8162_), .A3(new_n8182_), .Z(new_n8183_));
  OAI21_X1   g05385(.A1(new_n8151_), .A2(new_n8122_), .B(new_n8183_), .ZN(new_n8184_));
  NAND2_X1   g05386(.A1(new_n8032_), .A2(pi0038), .ZN(new_n8185_));
  NAND2_X1   g05387(.A1(new_n8185_), .A2(new_n7942_), .ZN(new_n8186_));
  NAND2_X1   g05388(.A1(new_n8186_), .A2(pi0087), .ZN(new_n8187_));
  AOI21_X1   g05389(.A1(new_n8184_), .A2(new_n3462_), .B(new_n8187_), .ZN(new_n8188_));
  OAI21_X1   g05390(.A1(new_n8188_), .A2(new_n8045_), .B(new_n3188_), .ZN(new_n8189_));
  NOR2_X1    g05391(.A1(new_n8060_), .A2(pi0054), .ZN(new_n8190_));
  AOI21_X1   g05392(.A1(new_n7933_), .A2(new_n8186_), .B(new_n6493_), .ZN(new_n8191_));
  NOR3_X1    g05393(.A1(new_n3259_), .A2(new_n8020_), .A3(new_n3098_), .ZN(new_n8192_));
  NOR3_X1    g05394(.A1(new_n3098_), .A2(pi0038), .A3(pi0155), .ZN(new_n8193_));
  OAI21_X1   g05395(.A1(new_n8192_), .A2(new_n8193_), .B(pi0177), .ZN(new_n8194_));
  OAI21_X1   g05396(.A1(new_n8191_), .A2(new_n8194_), .B(new_n7528_), .ZN(new_n8195_));
  NAND2_X1   g05397(.A1(new_n7528_), .A2(pi0100), .ZN(new_n8196_));
  XOR2_X1    g05398(.A1(new_n8195_), .A2(new_n8196_), .Z(new_n8197_));
  NAND2_X1   g05399(.A1(new_n8197_), .A2(new_n8044_), .ZN(new_n8198_));
  AOI21_X1   g05400(.A1(new_n8189_), .A2(new_n8190_), .B(new_n8198_), .ZN(new_n8199_));
  OAI21_X1   g05401(.A1(new_n8199_), .A2(new_n8071_), .B(new_n8074_), .ZN(new_n8200_));
  NOR4_X1    g05402(.A1(new_n7588_), .A2(new_n3192_), .A3(new_n7942_), .A4(new_n7986_), .ZN(new_n8201_));
  OAI21_X1   g05403(.A1(new_n8201_), .A2(pi0232), .B(pi0100), .ZN(new_n8202_));
  AOI21_X1   g05404(.A1(new_n8086_), .A2(new_n8076_), .B(new_n3235_), .ZN(new_n8203_));
  NAND2_X1   g05405(.A1(new_n8202_), .A2(new_n8203_), .ZN(new_n8204_));
  XOR2_X1    g05406(.A1(new_n8204_), .A2(new_n3483_), .Z(new_n8205_));
  NAND3_X1   g05407(.A1(new_n8205_), .A2(new_n5499_), .A3(new_n8086_), .ZN(new_n8206_));
  NAND2_X1   g05408(.A1(new_n7943_), .A2(pi0074), .ZN(new_n8207_));
  AOI21_X1   g05409(.A1(new_n8206_), .A2(new_n8092_), .B(new_n8207_), .ZN(new_n8208_));
  NOR4_X1    g05410(.A1(new_n8099_), .A2(new_n8081_), .A3(new_n8085_), .A4(new_n8088_), .ZN(new_n8209_));
  OAI21_X1   g05411(.A1(new_n8208_), .A2(pi0054), .B(new_n8209_), .ZN(new_n8210_));
  AOI21_X1   g05412(.A1(new_n8200_), .A2(new_n3226_), .B(new_n8210_), .ZN(new_n8211_));
  OAI21_X1   g05413(.A1(new_n8211_), .A2(new_n8104_), .B(new_n8097_), .ZN(new_n8212_));
  NAND2_X1   g05414(.A1(new_n8212_), .A2(pi0034), .ZN(new_n8213_));
  NOR2_X1    g05415(.A1(pi0033), .A2(pi0954), .ZN(new_n8214_));
  NAND2_X1   g05416(.A1(new_n8214_), .A2(pi0034), .ZN(new_n8215_));
  XOR2_X1    g05417(.A1(new_n8213_), .A2(new_n8215_), .Z(new_n8216_));
  NAND2_X1   g05418(.A1(new_n8212_), .A2(new_n8214_), .ZN(new_n8217_));
  NAND2_X1   g05419(.A1(new_n7959_), .A2(new_n7953_), .ZN(new_n8218_));
  INV_X1     g05420(.I(new_n8214_), .ZN(new_n8219_));
  NOR2_X1    g05421(.A1(new_n8219_), .A2(new_n7952_), .ZN(new_n8220_));
  OAI21_X1   g05422(.A1(new_n8218_), .A2(pi0034), .B(new_n8220_), .ZN(new_n8221_));
  XOR2_X1    g05423(.A1(new_n8217_), .A2(new_n8221_), .Z(new_n8222_));
  OAI21_X1   g05424(.A1(new_n8216_), .A2(new_n8222_), .B(new_n8102_), .ZN(po0192));
  NOR3_X1    g05425(.A1(new_n7325_), .A2(new_n3226_), .A3(new_n3292_), .ZN(new_n8224_));
  NAND2_X1   g05426(.A1(new_n8224_), .A2(new_n3258_), .ZN(new_n8225_));
  INV_X1     g05427(.I(new_n5546_), .ZN(new_n8226_));
  NOR2_X1    g05428(.A1(pi0058), .A2(pi0093), .ZN(new_n8227_));
  AOI21_X1   g05429(.A1(new_n2706_), .A2(new_n8227_), .B(new_n2679_), .ZN(new_n8228_));
  OAI21_X1   g05430(.A1(new_n5427_), .A2(new_n8228_), .B(new_n2692_), .ZN(new_n8229_));
  AOI21_X1   g05431(.A1(new_n2916_), .A2(pi0035), .B(new_n7295_), .ZN(new_n8230_));
  NAND2_X1   g05432(.A1(new_n8230_), .A2(new_n8229_), .ZN(new_n8231_));
  OAI21_X1   g05433(.A1(pi1082), .A2(new_n3142_), .B(new_n2502_), .ZN(new_n8232_));
  OAI21_X1   g05434(.A1(new_n8231_), .A2(new_n8232_), .B(new_n3259_), .ZN(new_n8233_));
  INV_X1     g05435(.I(new_n8230_), .ZN(new_n8234_));
  NAND2_X1   g05436(.A1(new_n7303_), .A2(new_n2478_), .ZN(new_n8235_));
  INV_X1     g05437(.I(po0740), .ZN(new_n8236_));
  NOR2_X1    g05438(.A1(new_n5469_), .A2(pi0137), .ZN(new_n8237_));
  INV_X1     g05439(.I(new_n8237_), .ZN(new_n8238_));
  NOR4_X1    g05440(.A1(new_n8236_), .A2(new_n6410_), .A3(new_n6939_), .A4(new_n8238_), .ZN(new_n8239_));
  NOR4_X1    g05441(.A1(new_n6504_), .A2(new_n8237_), .A3(new_n2730_), .A4(new_n6668_), .ZN(new_n8240_));
  NOR2_X1    g05442(.A1(new_n5468_), .A2(new_n7401_), .ZN(new_n8241_));
  OAI21_X1   g05443(.A1(new_n8240_), .A2(new_n8239_), .B(new_n8241_), .ZN(new_n8242_));
  NOR4_X1    g05444(.A1(new_n8234_), .A2(new_n8229_), .A3(new_n8235_), .A4(new_n8242_), .ZN(new_n8243_));
  NAND2_X1   g05445(.A1(new_n5468_), .A2(new_n2436_), .ZN(new_n8244_));
  AOI21_X1   g05446(.A1(new_n8243_), .A2(new_n8233_), .B(new_n8244_), .ZN(new_n8245_));
  NAND2_X1   g05447(.A1(new_n6307_), .A2(pi0038), .ZN(new_n8246_));
  NOR2_X1    g05448(.A1(new_n6403_), .A2(new_n2987_), .ZN(new_n8247_));
  INV_X1     g05449(.I(new_n8247_), .ZN(new_n8248_));
  NOR2_X1    g05450(.A1(new_n8248_), .A2(new_n5528_), .ZN(new_n8249_));
  OAI21_X1   g05451(.A1(po1057), .A2(pi0252), .B(new_n8249_), .ZN(new_n8250_));
  NAND2_X1   g05452(.A1(pi0142), .A2(pi0146), .ZN(new_n8251_));
  AND2_X2    g05453(.A1(new_n8250_), .A2(new_n8251_), .Z(new_n8252_));
  OAI22_X1   g05454(.A1(new_n8252_), .A2(new_n6494_), .B1(new_n6492_), .B2(new_n8251_), .ZN(new_n8253_));
  NAND4_X1   g05455(.A1(new_n8253_), .A2(new_n5508_), .A3(new_n7315_), .A4(new_n8250_), .ZN(new_n8254_));
  AOI21_X1   g05456(.A1(new_n8254_), .A2(new_n3721_), .B(new_n2776_), .ZN(new_n8255_));
  NAND2_X1   g05457(.A1(new_n7314_), .A2(new_n7319_), .ZN(new_n8256_));
  NAND4_X1   g05458(.A1(new_n8256_), .A2(pi0100), .A3(new_n3171_), .A4(new_n3211_), .ZN(new_n8257_));
  OAI22_X1   g05459(.A1(new_n8255_), .A2(new_n8257_), .B1(new_n7325_), .B2(new_n8246_), .ZN(new_n8258_));
  NOR2_X1    g05460(.A1(new_n2471_), .A2(pi0841), .ZN(new_n8259_));
  NAND4_X1   g05461(.A1(new_n8259_), .A2(pi0032), .A3(pi0093), .A4(new_n7273_), .ZN(new_n8260_));
  NAND3_X1   g05462(.A1(new_n8230_), .A2(new_n2794_), .A3(new_n8229_), .ZN(new_n8261_));
  NAND3_X1   g05463(.A1(new_n8258_), .A2(new_n8260_), .A3(new_n8261_), .ZN(new_n8262_));
  INV_X1     g05464(.I(new_n7325_), .ZN(new_n8263_));
  NOR2_X1    g05465(.A1(new_n8263_), .A2(new_n7337_), .ZN(new_n8264_));
  OAI21_X1   g05466(.A1(new_n8262_), .A2(new_n8245_), .B(new_n8264_), .ZN(new_n8265_));
  NOR4_X1    g05467(.A1(new_n6328_), .A2(new_n7272_), .A3(new_n3115_), .A4(new_n3226_), .ZN(new_n8266_));
  OAI21_X1   g05468(.A1(new_n6288_), .A2(new_n6398_), .B(new_n8266_), .ZN(new_n8267_));
  NAND2_X1   g05469(.A1(new_n7294_), .A2(new_n2776_), .ZN(new_n8268_));
  OAI21_X1   g05470(.A1(new_n7326_), .A2(new_n8268_), .B(new_n5527_), .ZN(new_n8269_));
  AOI21_X1   g05471(.A1(new_n8267_), .A2(new_n3303_), .B(new_n8269_), .ZN(new_n8270_));
  AOI21_X1   g05472(.A1(new_n8265_), .A2(new_n8270_), .B(new_n3229_), .ZN(new_n8271_));
  XOR2_X1    g05473(.A1(new_n8271_), .A2(new_n8226_), .Z(new_n8272_));
  NOR2_X1    g05474(.A1(new_n8272_), .A2(new_n8225_), .ZN(po0193));
  NAND3_X1   g05475(.A1(new_n2617_), .A2(new_n2630_), .A3(new_n2534_), .ZN(new_n8274_));
  NOR4_X1    g05476(.A1(new_n7353_), .A2(new_n2449_), .A3(new_n7281_), .A4(new_n2448_), .ZN(new_n8275_));
  INV_X1     g05477(.I(new_n8275_), .ZN(new_n8276_));
  NAND3_X1   g05478(.A1(pi0069), .A2(pi0071), .A3(pi0103), .ZN(new_n8277_));
  NOR4_X1    g05479(.A1(new_n8276_), .A2(new_n2605_), .A3(new_n2606_), .A4(new_n8277_), .ZN(new_n8278_));
  INV_X1     g05480(.I(new_n8278_), .ZN(new_n8279_));
  NOR2_X1    g05481(.A1(new_n8274_), .A2(new_n8279_), .ZN(new_n8280_));
  INV_X1     g05482(.I(new_n8280_), .ZN(new_n8281_));
  NOR2_X1    g05483(.A1(new_n2903_), .A2(new_n2522_), .ZN(new_n8282_));
  INV_X1     g05484(.I(new_n8282_), .ZN(new_n8283_));
  NOR2_X1    g05485(.A1(new_n8281_), .A2(new_n8283_), .ZN(new_n8284_));
  AOI21_X1   g05486(.A1(new_n6422_), .A2(new_n2686_), .B(new_n8284_), .ZN(new_n8285_));
  NOR2_X1    g05487(.A1(po1038), .A2(new_n3203_), .ZN(new_n8286_));
  NOR2_X1    g05488(.A1(new_n3495_), .A2(pi0092), .ZN(new_n8287_));
  NAND2_X1   g05489(.A1(new_n8287_), .A2(new_n8286_), .ZN(new_n8288_));
  NOR2_X1    g05490(.A1(new_n3138_), .A2(new_n2479_), .ZN(new_n8289_));
  NAND2_X1   g05491(.A1(new_n8289_), .A2(new_n5463_), .ZN(new_n8290_));
  NOR2_X1    g05492(.A1(new_n8288_), .A2(new_n8290_), .ZN(new_n8291_));
  INV_X1     g05493(.I(new_n8291_), .ZN(new_n8292_));
  NOR3_X1    g05494(.A1(new_n8285_), .A2(new_n8236_), .A3(new_n8292_), .ZN(po0194));
  NOR3_X1    g05495(.A1(new_n3304_), .A2(new_n7272_), .A3(new_n3183_), .ZN(new_n8294_));
  NAND2_X1   g05496(.A1(new_n2482_), .A2(new_n8294_), .ZN(new_n8295_));
  INV_X1     g05497(.I(new_n8295_), .ZN(new_n8296_));
  NOR2_X1    g05498(.A1(new_n3290_), .A2(po1038), .ZN(new_n8297_));
  NAND3_X1   g05499(.A1(new_n8296_), .A2(pi0038), .A3(new_n8297_), .ZN(new_n8298_));
  NAND3_X1   g05500(.A1(new_n8295_), .A2(new_n3259_), .A3(new_n8297_), .ZN(new_n8299_));
  NOR4_X1    g05501(.A1(new_n3138_), .A2(new_n2671_), .A3(new_n2490_), .A4(new_n7687_), .ZN(new_n8300_));
  INV_X1     g05502(.I(new_n8300_), .ZN(new_n8301_));
  NOR2_X1    g05503(.A1(new_n8301_), .A2(new_n2499_), .ZN(new_n8302_));
  INV_X1     g05504(.I(new_n8302_), .ZN(new_n8303_));
  INV_X1     g05505(.I(new_n2457_), .ZN(new_n8304_));
  NAND4_X1   g05506(.A1(new_n8304_), .A2(pi0039), .A3(pi0064), .A4(pi0841), .ZN(new_n8305_));
  OAI21_X1   g05507(.A1(new_n8303_), .A2(new_n8305_), .B(new_n2955_), .ZN(new_n8306_));
  NOR2_X1    g05508(.A1(new_n2572_), .A2(new_n2574_), .ZN(new_n8307_));
  INV_X1     g05509(.I(new_n8307_), .ZN(new_n8308_));
  NOR2_X1    g05510(.A1(new_n2592_), .A2(new_n8308_), .ZN(new_n8309_));
  INV_X1     g05511(.I(pi0089), .ZN(new_n8310_));
  NOR3_X1    g05512(.A1(new_n8310_), .A2(pi0082), .A3(pi0084), .ZN(new_n8311_));
  NAND4_X1   g05513(.A1(new_n8309_), .A2(pi0048), .A3(new_n8311_), .A4(pi0065), .ZN(new_n8312_));
  NOR4_X1    g05514(.A1(new_n2448_), .A2(new_n2438_), .A3(new_n2450_), .A4(new_n2585_), .ZN(new_n8313_));
  INV_X1     g05515(.I(new_n8313_), .ZN(new_n8314_));
  NOR3_X1    g05516(.A1(new_n8312_), .A2(new_n7364_), .A3(new_n8314_), .ZN(new_n8315_));
  NAND4_X1   g05517(.A1(new_n2651_), .A2(new_n2492_), .A3(new_n8306_), .A4(new_n8315_), .ZN(new_n8316_));
  AOI21_X1   g05518(.A1(new_n8298_), .A2(new_n8299_), .B(new_n8316_), .ZN(po0196));
  NAND2_X1   g05519(.A1(new_n3183_), .A2(new_n2436_), .ZN(new_n8318_));
  INV_X1     g05520(.I(pi0786), .ZN(new_n8319_));
  INV_X1     g05521(.I(pi1082), .ZN(new_n8320_));
  AOI22_X1   g05522(.A1(new_n5461_), .A2(new_n3381_), .B1(new_n5190_), .B2(new_n5400_), .ZN(new_n8321_));
  NOR4_X1    g05523(.A1(new_n8321_), .A2(new_n8319_), .A3(new_n8320_), .A4(new_n8236_), .ZN(new_n8322_));
  NOR2_X1    g05524(.A1(new_n5679_), .A2(new_n5407_), .ZN(new_n8323_));
  OAI21_X1   g05525(.A1(new_n5406_), .A2(new_n5402_), .B(new_n5403_), .ZN(new_n8324_));
  NAND2_X1   g05526(.A1(new_n8324_), .A2(new_n2980_), .ZN(new_n8325_));
  NAND3_X1   g05527(.A1(new_n5434_), .A2(new_n5437_), .A3(new_n8325_), .ZN(new_n8326_));
  NOR2_X1    g05528(.A1(new_n8323_), .A2(new_n8326_), .ZN(new_n8327_));
  INV_X1     g05529(.I(new_n8323_), .ZN(new_n8328_));
  NAND4_X1   g05530(.A1(new_n8328_), .A2(new_n5385_), .A3(new_n5437_), .A4(new_n8325_), .ZN(new_n8329_));
  NAND2_X1   g05531(.A1(new_n8329_), .A2(new_n5398_), .ZN(new_n8330_));
  NAND2_X1   g05532(.A1(new_n5398_), .A2(pi0299), .ZN(new_n8331_));
  XOR2_X1    g05533(.A1(new_n8330_), .A2(new_n8331_), .Z(new_n8332_));
  NAND2_X1   g05534(.A1(new_n8332_), .A2(new_n8327_), .ZN(new_n8333_));
  INV_X1     g05535(.I(new_n8333_), .ZN(new_n8334_));
  NAND4_X1   g05536(.A1(new_n8328_), .A2(pi1093), .A3(new_n5437_), .A4(new_n8325_), .ZN(new_n8335_));
  OAI21_X1   g05537(.A1(pi0223), .A2(new_n8335_), .B(new_n8334_), .ZN(new_n8336_));
  NAND2_X1   g05538(.A1(new_n8329_), .A2(pi0299), .ZN(new_n8337_));
  NAND2_X1   g05539(.A1(new_n5454_), .A2(pi0299), .ZN(new_n8338_));
  XOR2_X1    g05540(.A1(new_n8337_), .A2(new_n8338_), .Z(new_n8339_));
  NAND2_X1   g05541(.A1(new_n8339_), .A2(new_n8327_), .ZN(new_n8340_));
  INV_X1     g05542(.I(new_n8340_), .ZN(new_n8341_));
  OAI21_X1   g05543(.A1(pi0215), .A2(new_n8335_), .B(new_n8341_), .ZN(new_n8342_));
  NAND3_X1   g05544(.A1(pi0039), .A2(pi0786), .A3(pi1082), .ZN(new_n8343_));
  AOI21_X1   g05545(.A1(new_n8336_), .A2(new_n8342_), .B(new_n8343_), .ZN(new_n8344_));
  INV_X1     g05546(.I(new_n8297_), .ZN(new_n8345_));
  NOR2_X1    g05547(.A1(new_n8345_), .A2(pi0038), .ZN(new_n8346_));
  INV_X1     g05548(.I(new_n8346_), .ZN(new_n8347_));
  NOR2_X1    g05549(.A1(new_n8347_), .A2(new_n5681_), .ZN(new_n8348_));
  OAI21_X1   g05550(.A1(new_n8344_), .A2(new_n8322_), .B(new_n8348_), .ZN(new_n8349_));
  NAND2_X1   g05551(.A1(pi0097), .A2(pi0108), .ZN(new_n8350_));
  NOR3_X1    g05552(.A1(new_n2522_), .A2(new_n7266_), .A3(new_n8350_), .ZN(new_n8351_));
  NAND4_X1   g05553(.A1(new_n2514_), .A2(new_n8351_), .A3(pi0102), .A4(new_n2513_), .ZN(new_n8352_));
  NOR2_X1    g05554(.A1(new_n2673_), .A2(pi0841), .ZN(new_n8353_));
  NAND4_X1   g05555(.A1(pi0048), .A2(pi0068), .A3(pi0073), .A4(pi0082), .ZN(new_n8354_));
  NOR4_X1    g05556(.A1(new_n7277_), .A2(new_n8354_), .A3(pi0089), .A4(pi0102), .ZN(new_n8355_));
  NAND4_X1   g05557(.A1(pi0064), .A2(pi0066), .A3(pi0081), .A4(pi0084), .ZN(new_n8356_));
  NOR3_X1    g05558(.A1(new_n8356_), .A2(pi0065), .A3(pi0069), .ZN(new_n8357_));
  NOR4_X1    g05559(.A1(new_n8314_), .A2(new_n7281_), .A3(new_n2607_), .A4(new_n8308_), .ZN(new_n8358_));
  NAND4_X1   g05560(.A1(new_n8358_), .A2(new_n7363_), .A3(new_n8355_), .A4(new_n8357_), .ZN(new_n8359_));
  NOR3_X1    g05561(.A1(new_n8359_), .A2(new_n2459_), .A3(new_n2673_), .ZN(new_n8360_));
  XOR2_X1    g05562(.A1(new_n8360_), .A2(new_n8353_), .Z(new_n8361_));
  OAI21_X1   g05563(.A1(po0740), .A2(pi0986), .B(pi0252), .ZN(new_n8362_));
  NAND4_X1   g05564(.A1(new_n8362_), .A2(new_n2672_), .A3(pi0314), .A4(new_n2468_), .ZN(new_n8363_));
  NOR2_X1    g05565(.A1(new_n8363_), .A2(new_n5422_), .ZN(new_n8364_));
  AOI22_X1   g05566(.A1(new_n8361_), .A2(new_n8364_), .B1(new_n2673_), .B2(new_n8352_), .ZN(new_n8365_));
  INV_X1     g05567(.I(new_n2525_), .ZN(new_n8366_));
  NAND2_X1   g05568(.A1(new_n6381_), .A2(pi0035), .ZN(new_n8367_));
  OAI21_X1   g05569(.A1(new_n2500_), .A2(new_n2751_), .B(pi0035), .ZN(new_n8368_));
  OAI21_X1   g05570(.A1(new_n8367_), .A2(new_n8368_), .B(new_n2479_), .ZN(new_n8369_));
  NAND4_X1   g05571(.A1(new_n2516_), .A2(pi0053), .A3(pi0060), .A4(pi0841), .ZN(new_n8370_));
  NOR3_X1    g05572(.A1(new_n8359_), .A2(new_n2461_), .A3(new_n8370_), .ZN(new_n8371_));
  NAND4_X1   g05573(.A1(new_n8366_), .A2(new_n2900_), .A3(new_n8369_), .A4(new_n8371_), .ZN(new_n8372_));
  NOR2_X1    g05574(.A1(new_n5469_), .A2(pi0032), .ZN(new_n8373_));
  OAI21_X1   g05575(.A1(new_n8365_), .A2(new_n8372_), .B(new_n8373_), .ZN(new_n8374_));
  NAND2_X1   g05576(.A1(new_n8374_), .A2(new_n5557_), .ZN(new_n8375_));
  AOI21_X1   g05577(.A1(new_n8349_), .A2(new_n8318_), .B(new_n8375_), .ZN(po0197));
  NAND4_X1   g05578(.A1(new_n2487_), .A2(new_n2492_), .A3(pi0093), .A4(pi0102), .ZN(new_n8377_));
  NOR2_X1    g05579(.A1(new_n7351_), .A2(new_n8377_), .ZN(new_n8378_));
  NAND4_X1   g05580(.A1(new_n8378_), .A2(new_n2542_), .A3(new_n2491_), .A4(new_n5463_), .ZN(new_n8379_));
  OAI21_X1   g05581(.A1(new_n2750_), .A2(new_n2486_), .B(new_n3142_), .ZN(new_n8380_));
  INV_X1     g05582(.I(new_n8380_), .ZN(new_n8381_));
  NAND2_X1   g05583(.A1(new_n8379_), .A2(new_n2486_), .ZN(new_n8382_));
  AOI21_X1   g05584(.A1(new_n8381_), .A2(new_n8382_), .B(new_n8288_), .ZN(new_n8383_));
  INV_X1     g05585(.I(new_n8288_), .ZN(new_n8384_));
  NAND2_X1   g05586(.A1(new_n8384_), .A2(pi1082), .ZN(new_n8385_));
  XOR2_X1    g05587(.A1(new_n8383_), .A2(new_n8385_), .Z(new_n8386_));
  NOR3_X1    g05588(.A1(new_n8386_), .A2(new_n3138_), .A3(new_n8379_), .ZN(po0198));
  NAND2_X1   g05589(.A1(pi0041), .A2(pi0101), .ZN(new_n8388_));
  INV_X1     g05590(.I(pi0101), .ZN(new_n8389_));
  INV_X1     g05591(.I(pi0044), .ZN(new_n8390_));
  NOR2_X1    g05592(.A1(new_n8390_), .A2(pi0072), .ZN(new_n8391_));
  INV_X1     g05593(.I(new_n8391_), .ZN(new_n8392_));
  INV_X1     g05594(.I(new_n2711_), .ZN(new_n8393_));
  INV_X1     g05595(.I(new_n6364_), .ZN(new_n8394_));
  AOI22_X1   g05596(.A1(new_n6422_), .A2(new_n2487_), .B1(new_n8394_), .B2(new_n2931_), .ZN(new_n8395_));
  OAI21_X1   g05597(.A1(new_n8395_), .A2(new_n2930_), .B(new_n6370_), .ZN(new_n8396_));
  AOI21_X1   g05598(.A1(new_n8396_), .A2(new_n6373_), .B(new_n2702_), .ZN(new_n8397_));
  NAND2_X1   g05599(.A1(pi0051), .A2(pi0096), .ZN(new_n8398_));
  XOR2_X1    g05600(.A1(new_n8397_), .A2(new_n8398_), .Z(new_n8399_));
  NOR2_X1    g05601(.A1(new_n8399_), .A2(new_n8393_), .ZN(new_n8400_));
  NOR2_X1    g05602(.A1(new_n6387_), .A2(new_n6379_), .ZN(new_n8401_));
  INV_X1     g05603(.I(new_n6382_), .ZN(new_n8402_));
  NAND2_X1   g05604(.A1(new_n8402_), .A2(new_n3137_), .ZN(new_n8403_));
  NAND2_X1   g05605(.A1(new_n6379_), .A2(new_n2437_), .ZN(new_n8404_));
  NAND2_X1   g05606(.A1(new_n8403_), .A2(new_n8404_), .ZN(new_n8405_));
  OAI21_X1   g05607(.A1(new_n8401_), .A2(new_n8405_), .B(new_n8400_), .ZN(new_n8406_));
  OAI21_X1   g05608(.A1(new_n2984_), .A2(new_n8404_), .B(new_n8403_), .ZN(new_n8407_));
  NAND2_X1   g05609(.A1(new_n6380_), .A2(new_n2437_), .ZN(new_n8408_));
  AOI21_X1   g05610(.A1(new_n6377_), .A2(new_n8407_), .B(new_n8408_), .ZN(new_n8409_));
  OR3_X2     g05611(.A1(new_n8409_), .A2(new_n2984_), .A3(new_n6387_), .Z(new_n8410_));
  AOI21_X1   g05612(.A1(new_n8406_), .A2(new_n8410_), .B(new_n2437_), .ZN(new_n8411_));
  NAND2_X1   g05613(.A1(new_n8411_), .A2(new_n8390_), .ZN(new_n8412_));
  NAND2_X1   g05614(.A1(new_n8412_), .A2(new_n8392_), .ZN(new_n8413_));
  NOR2_X1    g05615(.A1(new_n8413_), .A2(new_n8389_), .ZN(new_n8414_));
  XOR2_X1    g05616(.A1(new_n8414_), .A2(new_n8388_), .Z(new_n8415_));
  NOR2_X1    g05617(.A1(new_n8415_), .A2(new_n2437_), .ZN(new_n8416_));
  INV_X1     g05618(.I(pi0041), .ZN(new_n8417_));
  NOR3_X1    g05619(.A1(new_n6385_), .A2(pi0044), .A3(pi1093), .ZN(new_n8418_));
  NOR3_X1    g05620(.A1(new_n8418_), .A2(new_n6379_), .A3(new_n6387_), .ZN(new_n8419_));
  OAI21_X1   g05621(.A1(new_n2984_), .A2(new_n8406_), .B(new_n8419_), .ZN(new_n8420_));
  NOR2_X1    g05622(.A1(new_n8420_), .A2(pi0101), .ZN(new_n8421_));
  INV_X1     g05623(.I(new_n8421_), .ZN(new_n8422_));
  NOR2_X1    g05624(.A1(new_n8422_), .A2(new_n8417_), .ZN(new_n8423_));
  OAI21_X1   g05625(.A1(new_n8416_), .A2(new_n2729_), .B(new_n8423_), .ZN(new_n8424_));
  NAND2_X1   g05626(.A1(new_n6387_), .A2(new_n2437_), .ZN(new_n8425_));
  NOR2_X1    g05627(.A1(new_n8425_), .A2(pi0044), .ZN(new_n8426_));
  NOR3_X1    g05628(.A1(new_n8426_), .A2(new_n8389_), .A3(new_n8391_), .ZN(new_n8427_));
  XOR2_X1    g05629(.A1(new_n8427_), .A2(new_n8388_), .Z(new_n8428_));
  NOR2_X1    g05630(.A1(new_n8428_), .A2(new_n2437_), .ZN(new_n8429_));
  INV_X1     g05631(.I(new_n8429_), .ZN(new_n8430_));
  NAND2_X1   g05632(.A1(new_n8430_), .A2(new_n2730_), .ZN(new_n8431_));
  OAI21_X1   g05633(.A1(new_n2984_), .A2(new_n6388_), .B(new_n8419_), .ZN(new_n8432_));
  NOR2_X1    g05634(.A1(new_n8432_), .A2(pi0101), .ZN(new_n8433_));
  INV_X1     g05635(.I(new_n8433_), .ZN(new_n8434_));
  NOR2_X1    g05636(.A1(new_n8434_), .A2(new_n8417_), .ZN(new_n8435_));
  AOI21_X1   g05637(.A1(new_n8431_), .A2(new_n8435_), .B(new_n3005_), .ZN(new_n8436_));
  NAND2_X1   g05638(.A1(new_n8424_), .A2(new_n8436_), .ZN(new_n8437_));
  NOR2_X1    g05639(.A1(new_n5386_), .A2(pi0189), .ZN(new_n8438_));
  INV_X1     g05640(.I(new_n8438_), .ZN(new_n8439_));
  NOR3_X1    g05641(.A1(new_n8439_), .A2(new_n7969_), .A3(pi0174), .ZN(new_n8440_));
  OAI21_X1   g05642(.A1(new_n8440_), .A2(pi0299), .B(new_n5551_), .ZN(new_n8441_));
  NOR2_X1    g05643(.A1(new_n5386_), .A2(pi0166), .ZN(new_n8442_));
  INV_X1     g05644(.I(new_n8442_), .ZN(new_n8443_));
  NOR4_X1    g05645(.A1(new_n8443_), .A2(pi0152), .A3(new_n4981_), .A4(new_n6878_), .ZN(new_n8444_));
  NAND2_X1   g05646(.A1(new_n8441_), .A2(new_n8444_), .ZN(new_n8445_));
  NOR2_X1    g05647(.A1(new_n3145_), .A2(new_n5401_), .ZN(new_n8447_));
  NOR2_X1    g05648(.A1(new_n3132_), .A2(pi0039), .ZN(new_n8449_));
  NAND2_X1   g05649(.A1(new_n2549_), .A2(new_n2902_), .ZN(new_n8450_));
  INV_X1     g05650(.I(new_n8450_), .ZN(new_n8451_));
  NOR2_X1    g05651(.A1(new_n8451_), .A2(new_n2480_), .ZN(new_n8452_));
  NOR3_X1    g05652(.A1(new_n2873_), .A2(pi0046), .A3(pi0109), .ZN(new_n8453_));
  AOI21_X1   g05653(.A1(new_n2549_), .A2(new_n8453_), .B(pi0110), .ZN(new_n8454_));
  NAND2_X1   g05654(.A1(new_n5413_), .A2(new_n2468_), .ZN(new_n8455_));
  AND3_X2    g05655(.A1(pi0901), .A2(pi0949), .A3(pi0959), .Z(new_n8456_));
  NAND4_X1   g05656(.A1(new_n2480_), .A2(pi0047), .A3(pi0480), .A4(new_n8456_), .ZN(new_n8457_));
  NOR4_X1    g05657(.A1(new_n8452_), .A2(new_n8454_), .A3(new_n8455_), .A4(new_n8457_), .ZN(new_n8458_));
  INV_X1     g05658(.I(pi0480), .ZN(new_n8459_));
  INV_X1     g05659(.I(pi0949), .ZN(new_n8460_));
  NOR4_X1    g05660(.A1(new_n2467_), .A2(new_n2673_), .A3(new_n2664_), .A4(new_n5420_), .ZN(new_n8461_));
  INV_X1     g05661(.I(new_n8461_), .ZN(new_n8462_));
  NOR2_X1    g05662(.A1(new_n8462_), .A2(new_n2665_), .ZN(new_n8463_));
  INV_X1     g05663(.I(new_n8463_), .ZN(new_n8464_));
  NOR4_X1    g05664(.A1(new_n8464_), .A2(new_n8459_), .A3(new_n8460_), .A4(new_n2481_), .ZN(new_n8465_));
  INV_X1     g05665(.I(new_n8465_), .ZN(new_n8466_));
  NOR4_X1    g05666(.A1(new_n8466_), .A2(pi0250), .A3(new_n3721_), .A4(new_n3138_), .ZN(new_n8467_));
  OAI21_X1   g05667(.A1(new_n8467_), .A2(pi0901), .B(pi0959), .ZN(new_n8468_));
  NOR2_X1    g05668(.A1(new_n8468_), .A2(new_n8458_), .ZN(new_n8469_));
  NAND2_X1   g05669(.A1(pi0250), .A2(pi0252), .ZN(new_n8470_));
  NOR2_X1    g05670(.A1(new_n8465_), .A2(new_n3137_), .ZN(new_n8471_));
  OAI21_X1   g05671(.A1(new_n8471_), .A2(new_n8470_), .B(new_n2437_), .ZN(new_n8472_));
  NOR2_X1    g05672(.A1(new_n8469_), .A2(new_n8472_), .ZN(new_n8473_));
  AOI21_X1   g05673(.A1(new_n8473_), .A2(new_n8390_), .B(new_n8391_), .ZN(new_n8474_));
  NAND2_X1   g05674(.A1(new_n8474_), .A2(pi0101), .ZN(new_n8475_));
  XOR2_X1    g05675(.A1(new_n8475_), .A2(new_n8388_), .Z(new_n8476_));
  NAND2_X1   g05676(.A1(new_n8476_), .A2(pi0072), .ZN(new_n8477_));
  OAI21_X1   g05677(.A1(new_n8477_), .A2(new_n3005_), .B(new_n8417_), .ZN(new_n8478_));
  NOR2_X1    g05678(.A1(new_n2733_), .A2(new_n3138_), .ZN(new_n8479_));
  INV_X1     g05679(.I(new_n8479_), .ZN(new_n8480_));
  NOR2_X1    g05680(.A1(new_n8480_), .A2(pi0044), .ZN(new_n8481_));
  NOR2_X1    g05681(.A1(new_n8389_), .A2(pi0072), .ZN(new_n8482_));
  NOR2_X1    g05682(.A1(new_n8482_), .A2(pi0041), .ZN(new_n8483_));
  AOI22_X1   g05683(.A1(new_n8481_), .A2(new_n8483_), .B1(new_n8417_), .B2(pi0072), .ZN(new_n8484_));
  AOI21_X1   g05684(.A1(new_n2437_), .A2(new_n6504_), .B(new_n8484_), .ZN(new_n8485_));
  NOR2_X1    g05685(.A1(new_n8485_), .A2(new_n2730_), .ZN(new_n8486_));
  NOR2_X1    g05686(.A1(new_n5519_), .A2(pi0099), .ZN(new_n8487_));
  NAND2_X1   g05687(.A1(new_n8487_), .A2(new_n2729_), .ZN(new_n8488_));
  XOR2_X1    g05688(.A1(new_n8486_), .A2(new_n8488_), .Z(new_n8489_));
  NOR2_X1    g05689(.A1(pi0044), .A2(pi0101), .ZN(new_n8490_));
  NAND2_X1   g05690(.A1(new_n3160_), .A2(new_n8490_), .ZN(new_n8491_));
  NOR2_X1    g05691(.A1(new_n8491_), .A2(new_n6504_), .ZN(new_n8492_));
  NOR3_X1    g05692(.A1(new_n8489_), .A2(pi0041), .A3(new_n2437_), .ZN(new_n8493_));
  INV_X1     g05693(.I(new_n6511_), .ZN(new_n8494_));
  AOI21_X1   g05694(.A1(new_n8445_), .A2(new_n2437_), .B(new_n3183_), .ZN(new_n8495_));
  INV_X1     g05695(.I(new_n8495_), .ZN(new_n8496_));
  OAI21_X1   g05696(.A1(new_n8496_), .A2(new_n5506_), .B(new_n3183_), .ZN(new_n8497_));
  NOR2_X1    g05697(.A1(pi0041), .A2(pi0072), .ZN(new_n8498_));
  NAND4_X1   g05698(.A1(new_n8497_), .A2(new_n2730_), .A3(new_n8494_), .A4(new_n8498_), .ZN(new_n8499_));
  OAI21_X1   g05699(.A1(new_n8493_), .A2(new_n8499_), .B(new_n3455_), .ZN(new_n8500_));
  INV_X1     g05700(.I(new_n8498_), .ZN(new_n8501_));
  AOI21_X1   g05701(.A1(new_n3183_), .A2(new_n8501_), .B(new_n8495_), .ZN(new_n8502_));
  NAND3_X1   g05702(.A1(new_n8500_), .A2(pi0038), .A3(new_n8502_), .ZN(new_n8503_));
  INV_X1     g05703(.I(new_n8492_), .ZN(new_n8504_));
  INV_X1     g05704(.I(new_n8483_), .ZN(new_n8505_));
  NOR2_X1    g05705(.A1(new_n2733_), .A2(pi0024), .ZN(new_n8506_));
  INV_X1     g05706(.I(new_n8506_), .ZN(new_n8507_));
  NOR4_X1    g05707(.A1(new_n8507_), .A2(new_n3721_), .A3(new_n3138_), .A4(new_n6504_), .ZN(new_n8508_));
  INV_X1     g05708(.I(new_n8508_), .ZN(new_n8509_));
  NOR2_X1    g05709(.A1(new_n8509_), .A2(pi0044), .ZN(new_n8510_));
  INV_X1     g05710(.I(new_n8510_), .ZN(new_n8511_));
  NOR2_X1    g05711(.A1(new_n8511_), .A2(new_n8505_), .ZN(new_n8512_));
  OAI21_X1   g05712(.A1(pi0041), .A2(new_n2437_), .B(new_n2730_), .ZN(new_n8513_));
  NAND4_X1   g05713(.A1(new_n8512_), .A2(pi0041), .A3(new_n8487_), .A4(new_n8513_), .ZN(new_n8514_));
  AOI21_X1   g05714(.A1(new_n8514_), .A2(new_n6523_), .B(new_n8504_), .ZN(new_n8515_));
  NOR4_X1    g05715(.A1(new_n6511_), .A2(new_n3183_), .A3(new_n2729_), .A4(new_n8501_), .ZN(new_n8516_));
  OAI21_X1   g05716(.A1(new_n3186_), .A2(new_n8495_), .B(new_n8516_), .ZN(new_n8517_));
  OAI21_X1   g05717(.A1(new_n8515_), .A2(new_n8517_), .B(new_n3235_), .ZN(new_n8518_));
  OAI21_X1   g05718(.A1(new_n3474_), .A2(new_n8498_), .B(new_n3005_), .ZN(new_n8519_));
  NOR2_X1    g05719(.A1(new_n8484_), .A2(new_n8519_), .ZN(new_n8520_));
  NAND2_X1   g05720(.A1(new_n8491_), .A2(pi0041), .ZN(new_n8521_));
  NAND2_X1   g05721(.A1(new_n3133_), .A2(new_n3191_), .ZN(new_n8522_));
  AOI21_X1   g05722(.A1(new_n8522_), .A2(new_n8498_), .B(pi0075), .ZN(new_n8523_));
  OAI21_X1   g05723(.A1(new_n8520_), .A2(new_n8521_), .B(new_n8523_), .ZN(new_n8524_));
  NOR2_X1    g05724(.A1(new_n8496_), .A2(new_n3187_), .ZN(new_n8525_));
  NAND4_X1   g05725(.A1(new_n8518_), .A2(new_n8502_), .A3(new_n8524_), .A4(new_n8525_), .ZN(new_n8526_));
  NAND2_X1   g05726(.A1(new_n8503_), .A2(new_n8526_), .ZN(new_n8527_));
  AOI21_X1   g05727(.A1(new_n8459_), .A2(new_n8460_), .B(new_n8470_), .ZN(new_n8528_));
  INV_X1     g05728(.I(new_n8290_), .ZN(new_n8529_));
  NAND2_X1   g05729(.A1(new_n8463_), .A2(new_n8529_), .ZN(new_n8530_));
  NOR2_X1    g05730(.A1(new_n8530_), .A2(new_n2437_), .ZN(new_n8531_));
  AOI21_X1   g05731(.A1(new_n8469_), .A2(new_n8528_), .B(new_n8531_), .ZN(new_n8532_));
  NAND2_X1   g05732(.A1(new_n8532_), .A2(new_n8390_), .ZN(new_n8533_));
  NOR2_X1    g05733(.A1(new_n8533_), .A2(pi0101), .ZN(new_n8534_));
  INV_X1     g05734(.I(new_n8502_), .ZN(new_n8535_));
  NOR2_X1    g05735(.A1(new_n3183_), .A2(new_n5551_), .ZN(new_n8536_));
  NAND4_X1   g05736(.A1(new_n8442_), .A2(new_n5158_), .A3(pi0161), .A4(new_n8536_), .ZN(new_n8537_));
  NOR2_X1    g05737(.A1(new_n3183_), .A2(new_n8417_), .ZN(new_n8538_));
  NAND4_X1   g05738(.A1(new_n7240_), .A2(pi0072), .A3(new_n8537_), .A4(new_n8538_), .ZN(new_n8539_));
  OAI21_X1   g05739(.A1(new_n8535_), .A2(new_n8539_), .B(new_n6400_), .ZN(new_n8540_));
  NAND4_X1   g05740(.A1(new_n8478_), .A2(new_n8527_), .A3(new_n8534_), .A4(new_n8540_), .ZN(new_n8541_));
  AOI21_X1   g05741(.A1(new_n8437_), .A2(new_n8449_), .B(new_n8541_), .ZN(po0199));
  NOR2_X1    g05742(.A1(new_n5509_), .A2(pi0072), .ZN(new_n8543_));
  NOR2_X1    g05743(.A1(new_n8543_), .A2(pi0039), .ZN(new_n8544_));
  INV_X1     g05744(.I(pi0207), .ZN(new_n8545_));
  INV_X1     g05745(.I(pi0208), .ZN(new_n8546_));
  NOR2_X1    g05746(.A1(new_n8545_), .A2(new_n8546_), .ZN(new_n8547_));
  NOR2_X1    g05747(.A1(new_n8544_), .A2(new_n8547_), .ZN(new_n8548_));
  INV_X1     g05748(.I(pi0199), .ZN(new_n8549_));
  AOI21_X1   g05749(.A1(new_n6216_), .A2(new_n8549_), .B(new_n2437_), .ZN(new_n8550_));
  NAND2_X1   g05750(.A1(new_n8550_), .A2(pi0232), .ZN(new_n8551_));
  NOR2_X1    g05751(.A1(new_n8438_), .A2(pi0072), .ZN(new_n8552_));
  INV_X1     g05752(.I(new_n8552_), .ZN(new_n8553_));
  AOI21_X1   g05753(.A1(new_n8551_), .A2(new_n8553_), .B(new_n8549_), .ZN(new_n8554_));
  INV_X1     g05754(.I(pi0200), .ZN(new_n8555_));
  AOI21_X1   g05755(.A1(new_n6216_), .A2(new_n8555_), .B(new_n2437_), .ZN(new_n8556_));
  INV_X1     g05756(.I(new_n8556_), .ZN(new_n8557_));
  NOR2_X1    g05757(.A1(new_n8557_), .A2(new_n5551_), .ZN(new_n8558_));
  OAI21_X1   g05758(.A1(new_n8558_), .A2(new_n8552_), .B(pi0200), .ZN(new_n8559_));
  INV_X1     g05759(.I(new_n8559_), .ZN(new_n8560_));
  NOR2_X1    g05760(.A1(new_n8560_), .A2(new_n3183_), .ZN(new_n8561_));
  INV_X1     g05761(.I(new_n8561_), .ZN(new_n8562_));
  NOR2_X1    g05762(.A1(new_n8562_), .A2(new_n8554_), .ZN(new_n8563_));
  INV_X1     g05763(.I(new_n8563_), .ZN(new_n8564_));
  AOI21_X1   g05764(.A1(new_n8564_), .A2(new_n8548_), .B(new_n6400_), .ZN(new_n8565_));
  NOR2_X1    g05765(.A1(new_n5515_), .A2(pi0072), .ZN(new_n8566_));
  INV_X1     g05766(.I(new_n8566_), .ZN(new_n8567_));
  NOR3_X1    g05767(.A1(new_n5520_), .A2(pi0072), .A3(new_n5512_), .ZN(new_n8569_));
  INV_X1     g05768(.I(new_n8569_), .ZN(new_n8570_));
  OAI21_X1   g05769(.A1(new_n8570_), .A2(pi0116), .B(new_n8567_), .ZN(new_n8571_));
  NOR2_X1    g05770(.A1(new_n8571_), .A2(new_n5509_), .ZN(new_n8572_));
  NOR2_X1    g05771(.A1(new_n5509_), .A2(new_n5513_), .ZN(new_n8573_));
  XOR2_X1    g05772(.A1(new_n8572_), .A2(new_n8573_), .Z(new_n8574_));
  NOR3_X1    g05773(.A1(new_n5521_), .A2(new_n5512_), .A3(new_n5515_), .ZN(new_n8575_));
  INV_X1     g05774(.I(new_n8575_), .ZN(new_n8576_));
  NOR2_X1    g05775(.A1(new_n8434_), .A2(new_n8576_), .ZN(new_n8577_));
  NOR2_X1    g05776(.A1(new_n8543_), .A2(new_n5513_), .ZN(new_n8578_));
  NAND2_X1   g05777(.A1(new_n2730_), .A2(new_n5514_), .ZN(new_n8579_));
  NAND4_X1   g05778(.A1(new_n8577_), .A2(new_n8574_), .A3(new_n8578_), .A4(new_n8579_), .ZN(new_n8580_));
  NAND2_X1   g05779(.A1(new_n8580_), .A2(new_n3005_), .ZN(new_n8581_));
  NOR3_X1    g05780(.A1(new_n5520_), .A2(pi0072), .A3(new_n5512_), .ZN(new_n8582_));
  NAND2_X1   g05781(.A1(new_n8582_), .A2(new_n5515_), .ZN(new_n8583_));
  NAND2_X1   g05782(.A1(new_n8583_), .A2(new_n8567_), .ZN(new_n8584_));
  NOR2_X1    g05783(.A1(pi0042), .A2(pi0114), .ZN(new_n8585_));
  NOR2_X1    g05784(.A1(pi0113), .A2(pi0116), .ZN(new_n8586_));
  INV_X1     g05785(.I(new_n8586_), .ZN(new_n8587_));
  NOR2_X1    g05786(.A1(new_n8422_), .A2(new_n5521_), .ZN(new_n8588_));
  INV_X1     g05787(.I(new_n8588_), .ZN(new_n8589_));
  NOR2_X1    g05788(.A1(new_n8589_), .A2(new_n8587_), .ZN(new_n8590_));
  NOR2_X1    g05789(.A1(new_n8590_), .A2(pi0042), .ZN(new_n8591_));
  OAI21_X1   g05790(.A1(new_n8591_), .A2(new_n8578_), .B(new_n8585_), .ZN(new_n8592_));
  NAND2_X1   g05791(.A1(new_n8592_), .A2(new_n8584_), .ZN(new_n8593_));
  INV_X1     g05792(.I(new_n8543_), .ZN(new_n8594_));
  NOR2_X1    g05793(.A1(new_n5512_), .A2(pi0072), .ZN(new_n8595_));
  INV_X1     g05794(.I(new_n8595_), .ZN(new_n8596_));
  NAND3_X1   g05795(.A1(new_n8417_), .A2(new_n2437_), .A3(pi0099), .ZN(new_n8597_));
  OAI21_X1   g05796(.A1(new_n8597_), .A2(pi0113), .B(new_n8596_), .ZN(new_n8598_));
  AOI21_X1   g05797(.A1(new_n8598_), .A2(new_n5515_), .B(new_n8566_), .ZN(new_n8599_));
  NAND2_X1   g05798(.A1(new_n8534_), .A2(new_n5520_), .ZN(new_n8600_));
  NOR2_X1    g05799(.A1(new_n8600_), .A2(new_n8587_), .ZN(new_n8601_));
  OAI22_X1   g05800(.A1(new_n8601_), .A2(pi0042), .B1(new_n5513_), .B2(new_n8543_), .ZN(new_n8602_));
  AOI21_X1   g05801(.A1(new_n8602_), .A2(new_n8585_), .B(new_n8599_), .ZN(new_n8603_));
  NOR2_X1    g05802(.A1(new_n8603_), .A2(new_n5514_), .ZN(new_n8604_));
  NAND2_X1   g05803(.A1(pi0115), .A2(pi0228), .ZN(new_n8605_));
  XOR2_X1    g05804(.A1(new_n8604_), .A2(new_n8605_), .Z(new_n8606_));
  OAI21_X1   g05805(.A1(new_n8606_), .A2(new_n8594_), .B(new_n3183_), .ZN(new_n8607_));
  NOR2_X1    g05806(.A1(new_n2730_), .A2(pi0115), .ZN(new_n8608_));
  INV_X1     g05807(.I(new_n8608_), .ZN(new_n8609_));
  NOR3_X1    g05808(.A1(new_n8609_), .A2(new_n5514_), .A3(new_n8594_), .ZN(new_n8610_));
  NAND4_X1   g05809(.A1(new_n8607_), .A2(new_n8581_), .A3(new_n8593_), .A4(new_n8610_), .ZN(new_n8611_));
  INV_X1     g05810(.I(new_n8481_), .ZN(new_n8612_));
  NOR2_X1    g05811(.A1(new_n8612_), .A2(new_n5523_), .ZN(new_n8613_));
  INV_X1     g05812(.I(new_n8613_), .ZN(new_n8614_));
  NOR2_X1    g05813(.A1(new_n8614_), .A2(new_n8587_), .ZN(new_n8615_));
  AOI21_X1   g05814(.A1(new_n8615_), .A2(new_n6486_), .B(pi0072), .ZN(new_n8616_));
  NAND2_X1   g05815(.A1(new_n8616_), .A2(pi0042), .ZN(new_n8617_));
  XOR2_X1    g05816(.A1(new_n8617_), .A2(new_n8573_), .Z(new_n8618_));
  NOR2_X1    g05817(.A1(new_n8491_), .A2(new_n8576_), .ZN(new_n8619_));
  NAND2_X1   g05818(.A1(new_n8619_), .A2(new_n6486_), .ZN(new_n8620_));
  INV_X1     g05819(.I(new_n8620_), .ZN(new_n8621_));
  AOI21_X1   g05820(.A1(new_n8585_), .A2(new_n5511_), .B(new_n5510_), .ZN(new_n8622_));
  NAND2_X1   g05821(.A1(new_n8621_), .A2(new_n8622_), .ZN(new_n8623_));
  AOI21_X1   g05822(.A1(new_n8543_), .A2(new_n8609_), .B(new_n8494_), .ZN(new_n8624_));
  NOR3_X1    g05823(.A1(new_n8624_), .A2(new_n8578_), .A3(new_n8608_), .ZN(new_n8625_));
  NOR4_X1    g05824(.A1(new_n8618_), .A2(new_n3183_), .A3(new_n8623_), .A4(new_n8625_), .ZN(new_n8626_));
  OAI21_X1   g05825(.A1(new_n8626_), .A2(new_n8543_), .B(new_n6511_), .ZN(new_n8627_));
  INV_X1     g05826(.I(new_n8627_), .ZN(new_n8628_));
  AOI21_X1   g05827(.A1(new_n6493_), .A2(new_n4808_), .B(pi0072), .ZN(new_n8629_));
  INV_X1     g05828(.I(new_n8629_), .ZN(new_n8630_));
  NOR2_X1    g05829(.A1(new_n8630_), .A2(new_n3098_), .ZN(new_n8631_));
  NOR2_X1    g05830(.A1(new_n8631_), .A2(new_n3183_), .ZN(new_n8632_));
  INV_X1     g05831(.I(new_n8632_), .ZN(new_n8633_));
  NOR2_X1    g05832(.A1(new_n8633_), .A2(new_n8554_), .ZN(new_n8634_));
  NOR2_X1    g05833(.A1(new_n8634_), .A2(new_n8544_), .ZN(new_n8635_));
  INV_X1     g05834(.I(new_n8635_), .ZN(new_n8636_));
  AOI21_X1   g05835(.A1(new_n8636_), .A2(pi0038), .B(pi0087), .ZN(new_n8637_));
  NAND4_X1   g05836(.A1(new_n8628_), .A2(new_n3259_), .A3(new_n3462_), .A4(new_n8634_), .ZN(new_n8638_));
  INV_X1     g05837(.I(new_n8447_), .ZN(new_n8639_));
  NOR2_X1    g05838(.A1(new_n8639_), .A2(new_n8443_), .ZN(new_n8640_));
  NOR3_X1    g05839(.A1(new_n8640_), .A2(new_n6216_), .A3(new_n8629_), .ZN(new_n8641_));
  INV_X1     g05840(.I(pi0189), .ZN(new_n8642_));
  NOR2_X1    g05841(.A1(new_n5386_), .A2(new_n8642_), .ZN(new_n8643_));
  INV_X1     g05842(.I(new_n8643_), .ZN(new_n8644_));
  NOR3_X1    g05843(.A1(new_n8639_), .A2(new_n2437_), .A3(new_n8644_), .ZN(new_n8645_));
  NOR3_X1    g05844(.A1(new_n8447_), .A2(pi0072), .A3(new_n8644_), .ZN(new_n8646_));
  NOR2_X1    g05845(.A1(new_n8645_), .A2(new_n8646_), .ZN(new_n8647_));
  NOR2_X1    g05846(.A1(pi0232), .A2(pi0299), .ZN(new_n8648_));
  NOR3_X1    g05847(.A1(new_n8647_), .A2(new_n8549_), .A3(new_n8648_), .ZN(new_n8649_));
  OAI21_X1   g05848(.A1(new_n2437_), .A2(new_n5551_), .B(new_n3098_), .ZN(new_n8650_));
  NAND2_X1   g05849(.A1(new_n8650_), .A2(pi0199), .ZN(new_n8651_));
  NAND2_X1   g05850(.A1(new_n8651_), .A2(new_n3183_), .ZN(new_n8652_));
  OAI21_X1   g05851(.A1(new_n8649_), .A2(new_n8652_), .B(new_n8641_), .ZN(new_n8653_));
  AOI21_X1   g05852(.A1(new_n8611_), .A2(new_n8638_), .B(new_n8653_), .ZN(new_n8654_));
  INV_X1     g05853(.I(new_n8634_), .ZN(new_n8655_));
  NOR2_X1    g05854(.A1(new_n8614_), .A2(new_n3005_), .ZN(new_n8656_));
  INV_X1     g05855(.I(new_n8656_), .ZN(new_n8657_));
  OAI21_X1   g05856(.A1(new_n8657_), .A2(new_n5517_), .B(new_n8543_), .ZN(new_n8658_));
  NAND2_X1   g05857(.A1(new_n8619_), .A2(pi0228), .ZN(new_n8659_));
  NOR3_X1    g05858(.A1(new_n8659_), .A2(pi0114), .A3(pi0115), .ZN(new_n8660_));
  NAND2_X1   g05859(.A1(new_n8660_), .A2(pi0042), .ZN(new_n8661_));
  AOI21_X1   g05860(.A1(new_n8658_), .A2(new_n3474_), .B(new_n8661_), .ZN(new_n8662_));
  AOI21_X1   g05861(.A1(new_n8544_), .A2(new_n3133_), .B(new_n3455_), .ZN(new_n8663_));
  INV_X1     g05862(.I(new_n8663_), .ZN(new_n8664_));
  NOR2_X1    g05863(.A1(new_n8662_), .A2(new_n8664_), .ZN(new_n8665_));
  INV_X1     g05864(.I(new_n8665_), .ZN(new_n8666_));
  NOR2_X1    g05865(.A1(new_n8666_), .A2(new_n8655_), .ZN(new_n8667_));
  OAI21_X1   g05866(.A1(new_n8654_), .A2(pi0075), .B(new_n8667_), .ZN(new_n8668_));
  INV_X1     g05867(.I(new_n8625_), .ZN(new_n8669_));
  NOR2_X1    g05868(.A1(new_n8511_), .A2(new_n5523_), .ZN(new_n8670_));
  NAND2_X1   g05869(.A1(new_n8670_), .A2(new_n8586_), .ZN(new_n8671_));
  NAND2_X1   g05870(.A1(new_n8671_), .A2(new_n8543_), .ZN(new_n8672_));
  NOR2_X1    g05871(.A1(new_n8623_), .A2(new_n6523_), .ZN(new_n8673_));
  NAND2_X1   g05872(.A1(new_n8673_), .A2(new_n5509_), .ZN(new_n8674_));
  NAND4_X1   g05873(.A1(new_n8672_), .A2(new_n5513_), .A3(new_n8669_), .A4(new_n8674_), .ZN(new_n8675_));
  NAND2_X1   g05874(.A1(new_n8675_), .A2(new_n3187_), .ZN(new_n8676_));
  NAND3_X1   g05875(.A1(new_n8676_), .A2(new_n6511_), .A3(new_n8543_), .ZN(new_n8677_));
  NAND2_X1   g05876(.A1(new_n3186_), .A2(new_n8543_), .ZN(new_n8678_));
  AOI21_X1   g05877(.A1(new_n8677_), .A2(new_n3183_), .B(new_n8678_), .ZN(new_n8679_));
  NOR2_X1    g05878(.A1(new_n6400_), .A2(new_n3235_), .ZN(new_n8680_));
  NOR2_X1    g05879(.A1(new_n8679_), .A2(new_n8680_), .ZN(new_n8681_));
  NOR2_X1    g05880(.A1(new_n8681_), .A2(new_n8655_), .ZN(new_n8682_));
  INV_X1     g05881(.I(pi0219), .ZN(new_n8683_));
  INV_X1     g05882(.I(pi0211), .ZN(new_n8684_));
  INV_X1     g05883(.I(pi0214), .ZN(new_n8685_));
  NOR2_X1    g05884(.A1(new_n8684_), .A2(new_n8685_), .ZN(new_n8686_));
  NAND2_X1   g05885(.A1(new_n8686_), .A2(pi0212), .ZN(new_n8687_));
  NAND2_X1   g05886(.A1(new_n8687_), .A2(new_n8683_), .ZN(new_n8688_));
  INV_X1     g05887(.I(new_n8688_), .ZN(new_n8689_));
  NOR2_X1    g05888(.A1(new_n8689_), .A2(new_n8547_), .ZN(new_n8690_));
  OAI21_X1   g05889(.A1(new_n8636_), .A2(new_n6399_), .B(new_n8690_), .ZN(new_n8691_));
  AOI21_X1   g05890(.A1(new_n8668_), .A2(new_n8682_), .B(new_n8691_), .ZN(new_n8692_));
  NOR2_X1    g05891(.A1(new_n8655_), .A2(new_n8562_), .ZN(new_n8693_));
  INV_X1     g05892(.I(new_n8693_), .ZN(new_n8694_));
  AOI21_X1   g05893(.A1(new_n8627_), .A2(new_n8694_), .B(new_n5506_), .ZN(new_n8695_));
  INV_X1     g05894(.I(new_n7487_), .ZN(new_n8696_));
  NOR3_X1    g05895(.A1(new_n8696_), .A2(pi0039), .A3(new_n8543_), .ZN(new_n8697_));
  NOR2_X1    g05896(.A1(new_n8637_), .A2(new_n8697_), .ZN(new_n8698_));
  OR3_X2     g05897(.A1(new_n8695_), .A2(new_n3133_), .A3(new_n8698_), .Z(new_n8699_));
  NOR2_X1    g05898(.A1(new_n8681_), .A2(new_n8694_), .ZN(new_n8700_));
  NAND2_X1   g05899(.A1(new_n8694_), .A2(new_n8663_), .ZN(new_n8701_));
  OAI21_X1   g05900(.A1(new_n8662_), .A2(new_n8701_), .B(new_n3235_), .ZN(new_n8702_));
  OAI21_X1   g05901(.A1(new_n8647_), .A2(new_n5551_), .B(new_n8555_), .ZN(new_n8703_));
  NAND2_X1   g05902(.A1(new_n8703_), .A2(pi0199), .ZN(new_n8704_));
  INV_X1     g05903(.I(new_n8641_), .ZN(new_n8705_));
  OAI21_X1   g05904(.A1(new_n8705_), .A2(new_n8651_), .B(new_n8555_), .ZN(new_n8706_));
  NOR2_X1    g05905(.A1(new_n3183_), .A2(new_n2437_), .ZN(new_n8707_));
  NAND2_X1   g05906(.A1(new_n8706_), .A2(new_n8707_), .ZN(new_n8708_));
  AOI21_X1   g05907(.A1(new_n8708_), .A2(new_n8704_), .B(new_n3098_), .ZN(new_n8709_));
  OAI21_X1   g05908(.A1(new_n8700_), .A2(new_n8702_), .B(new_n8709_), .ZN(new_n8710_));
  AOI21_X1   g05909(.A1(new_n8611_), .A2(new_n8699_), .B(new_n8710_), .ZN(new_n8711_));
  OAI21_X1   g05910(.A1(new_n8692_), .A2(new_n8565_), .B(new_n8711_), .ZN(new_n8712_));
  OAI21_X1   g05911(.A1(new_n8630_), .A2(new_n8689_), .B(po1038), .ZN(new_n8713_));
  NOR2_X1    g05912(.A1(new_n7240_), .A2(new_n3183_), .ZN(new_n8714_));
  XNOR2_X1   g05913(.A1(new_n8713_), .A2(new_n8714_), .ZN(new_n8715_));
  AOI21_X1   g05914(.A1(new_n8715_), .A2(new_n8543_), .B(po1038), .ZN(new_n8716_));
  INV_X1     g05915(.I(new_n8554_), .ZN(new_n8717_));
  NAND2_X1   g05916(.A1(new_n8717_), .A2(pi0039), .ZN(new_n8718_));
  AOI21_X1   g05917(.A1(new_n8718_), .A2(new_n8548_), .B(new_n6400_), .ZN(new_n8719_));
  NAND4_X1   g05918(.A1(new_n8628_), .A2(new_n3259_), .A3(new_n3462_), .A4(new_n8563_), .ZN(new_n8720_));
  OAI21_X1   g05919(.A1(new_n8704_), .A2(new_n3183_), .B(new_n8557_), .ZN(new_n8721_));
  NAND2_X1   g05920(.A1(new_n8721_), .A2(new_n8550_), .ZN(new_n8722_));
  AOI21_X1   g05921(.A1(new_n8611_), .A2(new_n8720_), .B(new_n8722_), .ZN(new_n8723_));
  NOR2_X1    g05922(.A1(new_n8666_), .A2(new_n8564_), .ZN(new_n8724_));
  OAI21_X1   g05923(.A1(new_n8723_), .A2(pi0075), .B(new_n8724_), .ZN(new_n8725_));
  NOR2_X1    g05924(.A1(new_n8681_), .A2(new_n8564_), .ZN(new_n8726_));
  NAND2_X1   g05925(.A1(new_n8565_), .A2(new_n8689_), .ZN(new_n8727_));
  AOI21_X1   g05926(.A1(new_n8725_), .A2(new_n8726_), .B(new_n8727_), .ZN(new_n8728_));
  OR2_X2     g05927(.A1(new_n8611_), .A2(new_n3133_), .Z(new_n8729_));
  NAND4_X1   g05928(.A1(new_n8594_), .A2(new_n3183_), .A3(new_n5505_), .A4(new_n7487_), .ZN(new_n8730_));
  AOI21_X1   g05929(.A1(new_n8627_), .A2(new_n8730_), .B(new_n8718_), .ZN(new_n8731_));
  NAND3_X1   g05930(.A1(new_n8717_), .A2(pi0039), .A3(new_n3235_), .ZN(new_n8732_));
  NOR2_X1    g05931(.A1(new_n8681_), .A2(new_n8732_), .ZN(new_n8733_));
  AOI21_X1   g05932(.A1(new_n8549_), .A2(new_n8551_), .B(new_n8647_), .ZN(new_n8734_));
  OAI21_X1   g05933(.A1(new_n8733_), .A2(new_n8731_), .B(new_n8734_), .ZN(new_n8735_));
  AOI21_X1   g05934(.A1(new_n8729_), .A2(new_n3183_), .B(new_n8735_), .ZN(new_n8736_));
  OAI21_X1   g05935(.A1(new_n8728_), .A2(new_n8719_), .B(new_n8736_), .ZN(new_n8737_));
  AOI21_X1   g05936(.A1(new_n8712_), .A2(new_n8716_), .B(new_n8737_), .ZN(po0200));
  INV_X1     g05937(.I(pi0212), .ZN(new_n8739_));
  NOR2_X1    g05938(.A1(new_n8739_), .A2(new_n8685_), .ZN(new_n8740_));
  NOR2_X1    g05939(.A1(new_n8740_), .A2(new_n8684_), .ZN(new_n8741_));
  NOR2_X1    g05940(.A1(pi0211), .A2(pi0219), .ZN(new_n8742_));
  AOI21_X1   g05941(.A1(new_n8740_), .A2(new_n8742_), .B(new_n8741_), .ZN(new_n8743_));
  INV_X1     g05942(.I(new_n8680_), .ZN(new_n8744_));
  NOR2_X1    g05943(.A1(new_n5510_), .A2(pi0072), .ZN(new_n8745_));
  INV_X1     g05944(.I(new_n8745_), .ZN(new_n8746_));
  INV_X1     g05945(.I(new_n8585_), .ZN(new_n8747_));
  NOR2_X1    g05946(.A1(new_n8747_), .A2(pi0115), .ZN(new_n8748_));
  INV_X1     g05947(.I(new_n8748_), .ZN(new_n8749_));
  NOR3_X1    g05948(.A1(new_n8494_), .A2(new_n2730_), .A3(new_n8749_), .ZN(new_n8750_));
  INV_X1     g05949(.I(new_n8750_), .ZN(new_n8751_));
  NOR2_X1    g05950(.A1(new_n8751_), .A2(new_n8746_), .ZN(new_n8752_));
  INV_X1     g05951(.I(new_n8752_), .ZN(new_n8753_));
  AOI21_X1   g05952(.A1(new_n8621_), .A2(new_n6485_), .B(new_n5510_), .ZN(new_n8754_));
  INV_X1     g05953(.I(new_n8754_), .ZN(new_n8755_));
  NOR2_X1    g05954(.A1(new_n5510_), .A2(new_n5511_), .ZN(new_n8756_));
  INV_X1     g05955(.I(new_n8756_), .ZN(new_n8757_));
  INV_X1     g05956(.I(new_n8671_), .ZN(new_n8758_));
  NOR2_X1    g05957(.A1(new_n8758_), .A2(pi0072), .ZN(new_n8759_));
  INV_X1     g05958(.I(new_n8759_), .ZN(new_n8760_));
  NOR2_X1    g05959(.A1(new_n8760_), .A2(new_n8757_), .ZN(new_n8761_));
  NOR2_X1    g05960(.A1(new_n8761_), .A2(new_n8755_), .ZN(new_n8762_));
  NAND2_X1   g05961(.A1(new_n8761_), .A2(new_n8755_), .ZN(new_n8763_));
  NAND2_X1   g05962(.A1(new_n8763_), .A2(new_n8750_), .ZN(new_n8764_));
  NOR2_X1    g05963(.A1(new_n8764_), .A2(new_n8762_), .ZN(new_n8765_));
  NAND2_X1   g05964(.A1(new_n8765_), .A2(new_n8753_), .ZN(new_n8766_));
  OAI21_X1   g05965(.A1(new_n8764_), .A2(new_n8762_), .B(new_n8752_), .ZN(new_n8767_));
  NAND3_X1   g05966(.A1(new_n8766_), .A2(new_n3186_), .A3(new_n8767_), .ZN(new_n8768_));
  NOR2_X1    g05967(.A1(new_n3187_), .A2(new_n3183_), .ZN(new_n8769_));
  XOR2_X1    g05968(.A1(new_n8768_), .A2(new_n8769_), .Z(new_n8770_));
  OAI21_X1   g05969(.A1(new_n8770_), .A2(new_n8746_), .B(new_n8744_), .ZN(new_n8771_));
  NOR2_X1    g05970(.A1(pi0199), .A2(pi0200), .ZN(new_n8772_));
  INV_X1     g05971(.I(new_n8772_), .ZN(new_n8773_));
  NOR2_X1    g05972(.A1(new_n8772_), .A2(pi0299), .ZN(new_n8774_));
  INV_X1     g05973(.I(new_n8774_), .ZN(new_n8775_));
  AOI21_X1   g05974(.A1(new_n8775_), .A2(new_n2437_), .B(pi0232), .ZN(new_n8776_));
  NOR2_X1    g05975(.A1(new_n8776_), .A2(pi0299), .ZN(new_n8777_));
  AOI21_X1   g05976(.A1(new_n8777_), .A2(pi0039), .B(pi0232), .ZN(new_n8778_));
  NOR3_X1    g05977(.A1(new_n8778_), .A2(new_n8553_), .A3(new_n8773_), .ZN(new_n8779_));
  INV_X1     g05978(.I(new_n8779_), .ZN(new_n8780_));
  NOR2_X1    g05979(.A1(new_n8780_), .A2(new_n8631_), .ZN(new_n8781_));
  NOR2_X1    g05980(.A1(new_n8599_), .A2(pi0228), .ZN(new_n8782_));
  NAND2_X1   g05981(.A1(new_n8571_), .A2(new_n2730_), .ZN(new_n8783_));
  NAND2_X1   g05982(.A1(new_n8584_), .A2(new_n2729_), .ZN(new_n8784_));
  AOI21_X1   g05983(.A1(new_n8783_), .A2(new_n8784_), .B(new_n3005_), .ZN(new_n8785_));
  NOR2_X1    g05984(.A1(new_n8785_), .A2(new_n8782_), .ZN(new_n8786_));
  NAND2_X1   g05985(.A1(new_n8589_), .A2(new_n2729_), .ZN(new_n8787_));
  OAI21_X1   g05986(.A1(new_n8434_), .A2(new_n5521_), .B(new_n2730_), .ZN(new_n8788_));
  NAND2_X1   g05987(.A1(new_n8787_), .A2(new_n8788_), .ZN(new_n8789_));
  NOR3_X1    g05988(.A1(new_n8789_), .A2(new_n3005_), .A3(new_n8587_), .ZN(new_n8790_));
  AOI21_X1   g05989(.A1(new_n3005_), .A2(new_n8601_), .B(new_n8790_), .ZN(new_n8791_));
  NOR2_X1    g05990(.A1(new_n8748_), .A2(pi0072), .ZN(new_n8792_));
  OAI22_X1   g05991(.A1(new_n8791_), .A2(new_n8792_), .B1(new_n5510_), .B2(new_n2437_), .ZN(new_n8793_));
  AOI22_X1   g05992(.A1(new_n8793_), .A2(pi0039), .B1(pi0043), .B2(new_n8748_), .ZN(new_n8794_));
  OR2_X2     g05993(.A1(new_n8794_), .A2(new_n8786_), .Z(new_n8795_));
  NOR2_X1    g05994(.A1(new_n8616_), .A2(new_n8757_), .ZN(new_n8796_));
  INV_X1     g05995(.I(new_n8796_), .ZN(new_n8797_));
  NAND3_X1   g05996(.A1(new_n8797_), .A2(pi0043), .A3(new_n8620_), .ZN(new_n8798_));
  OAI21_X1   g05997(.A1(new_n5510_), .A2(new_n8621_), .B(new_n8796_), .ZN(new_n8799_));
  NAND3_X1   g05998(.A1(new_n8798_), .A2(new_n8750_), .A3(new_n8799_), .ZN(new_n8800_));
  NOR2_X1    g05999(.A1(new_n8800_), .A2(new_n8752_), .ZN(new_n8801_));
  AND2_X2    g06000(.A1(new_n8800_), .A2(new_n8752_), .Z(new_n8802_));
  NOR3_X1    g06001(.A1(new_n8802_), .A2(new_n8801_), .A3(pi0039), .ZN(new_n8803_));
  NOR2_X1    g06002(.A1(new_n8745_), .A2(pi0039), .ZN(new_n8804_));
  NAND2_X1   g06003(.A1(new_n8804_), .A2(new_n5505_), .ZN(new_n8805_));
  NOR2_X1    g06004(.A1(new_n8633_), .A2(new_n8560_), .ZN(new_n8806_));
  INV_X1     g06005(.I(new_n8806_), .ZN(new_n8807_));
  AOI21_X1   g06006(.A1(new_n8807_), .A2(new_n8696_), .B(new_n8805_), .ZN(new_n8808_));
  NOR2_X1    g06007(.A1(new_n8807_), .A2(new_n3133_), .ZN(new_n8809_));
  OAI21_X1   g06008(.A1(new_n8803_), .A2(new_n8808_), .B(new_n8809_), .ZN(new_n8810_));
  NAND2_X1   g06009(.A1(new_n8795_), .A2(new_n8810_), .ZN(new_n8811_));
  NAND2_X1   g06010(.A1(new_n8647_), .A2(pi0200), .ZN(new_n8812_));
  NAND3_X1   g06011(.A1(new_n8812_), .A2(pi0232), .A3(new_n3098_), .ZN(new_n8813_));
  AOI21_X1   g06012(.A1(new_n8650_), .A2(pi0200), .B(pi0039), .ZN(new_n8814_));
  AOI21_X1   g06013(.A1(new_n8813_), .A2(new_n8814_), .B(new_n8705_), .ZN(new_n8815_));
  AOI21_X1   g06014(.A1(new_n8811_), .A2(new_n8815_), .B(pi0075), .ZN(new_n8816_));
  INV_X1     g06015(.I(new_n8615_), .ZN(new_n8817_));
  NAND2_X1   g06016(.A1(new_n8817_), .A2(new_n2437_), .ZN(new_n8818_));
  NOR2_X1    g06017(.A1(new_n8749_), .A2(new_n3005_), .ZN(new_n8819_));
  NAND2_X1   g06018(.A1(new_n8818_), .A2(new_n8819_), .ZN(new_n8820_));
  NAND2_X1   g06019(.A1(new_n8819_), .A2(pi0043), .ZN(new_n8821_));
  XOR2_X1    g06020(.A1(new_n8820_), .A2(new_n8821_), .Z(new_n8822_));
  AOI21_X1   g06021(.A1(new_n8822_), .A2(new_n8619_), .B(new_n3134_), .ZN(new_n8823_));
  NAND2_X1   g06022(.A1(new_n8819_), .A2(new_n8745_), .ZN(new_n8824_));
  OAI21_X1   g06023(.A1(new_n8823_), .A2(new_n8824_), .B(new_n3455_), .ZN(new_n8825_));
  NAND4_X1   g06024(.A1(new_n8825_), .A2(new_n3132_), .A3(new_n8804_), .A4(new_n8806_), .ZN(new_n8826_));
  AND2_X2    g06025(.A1(new_n8771_), .A2(new_n8806_), .Z(new_n8827_));
  OAI21_X1   g06026(.A1(new_n8816_), .A2(new_n8826_), .B(new_n8827_), .ZN(new_n8828_));
  INV_X1     g06027(.I(new_n8781_), .ZN(new_n8829_));
  NOR2_X1    g06028(.A1(new_n8804_), .A2(new_n8547_), .ZN(new_n8830_));
  NAND2_X1   g06029(.A1(new_n8807_), .A2(new_n8830_), .ZN(new_n8831_));
  NAND2_X1   g06030(.A1(new_n8831_), .A2(new_n6399_), .ZN(new_n8832_));
  AOI21_X1   g06031(.A1(new_n8829_), .A2(new_n8830_), .B(new_n8832_), .ZN(new_n8833_));
  AOI22_X1   g06032(.A1(new_n8828_), .A2(new_n8833_), .B1(new_n8771_), .B2(new_n8781_), .ZN(new_n8834_));
  NOR3_X1    g06033(.A1(new_n8647_), .A2(new_n8648_), .A3(new_n8773_), .ZN(new_n8835_));
  OR3_X2     g06034(.A1(new_n8835_), .A2(pi0039), .A3(new_n8776_), .Z(new_n8836_));
  NAND2_X1   g06035(.A1(new_n8836_), .A2(new_n8641_), .ZN(new_n8837_));
  AOI21_X1   g06036(.A1(new_n8829_), .A2(new_n8696_), .B(new_n8805_), .ZN(new_n8838_));
  NOR2_X1    g06037(.A1(new_n8829_), .A2(new_n3133_), .ZN(new_n8839_));
  OAI21_X1   g06038(.A1(new_n8803_), .A2(new_n8838_), .B(new_n8839_), .ZN(new_n8840_));
  AOI21_X1   g06039(.A1(new_n8795_), .A2(new_n8840_), .B(new_n8837_), .ZN(new_n8841_));
  NAND3_X1   g06040(.A1(new_n8825_), .A2(new_n3132_), .A3(new_n8804_), .ZN(new_n8842_));
  NOR2_X1    g06041(.A1(new_n8842_), .A2(new_n8829_), .ZN(new_n8843_));
  OAI21_X1   g06042(.A1(new_n8841_), .A2(pi0075), .B(new_n8843_), .ZN(new_n8844_));
  NOR2_X1    g06043(.A1(new_n8834_), .A2(new_n8844_), .ZN(new_n8845_));
  NOR2_X1    g06044(.A1(new_n8845_), .A2(new_n8743_), .ZN(new_n8846_));
  NOR2_X1    g06045(.A1(new_n7240_), .A2(new_n8743_), .ZN(new_n8847_));
  XOR2_X1    g06046(.A1(new_n8846_), .A2(new_n8847_), .Z(new_n8848_));
  NOR2_X1    g06047(.A1(new_n8779_), .A2(new_n8804_), .ZN(new_n8849_));
  NOR3_X1    g06048(.A1(new_n3462_), .A2(pi0038), .A3(pi0087), .ZN(new_n8850_));
  NOR2_X1    g06049(.A1(new_n8780_), .A2(new_n3133_), .ZN(new_n8851_));
  OAI21_X1   g06050(.A1(new_n8803_), .A2(new_n8850_), .B(new_n8851_), .ZN(new_n8852_));
  NAND2_X1   g06051(.A1(new_n8795_), .A2(new_n8852_), .ZN(new_n8853_));
  OAI21_X1   g06052(.A1(new_n8842_), .A2(new_n3235_), .B(new_n3214_), .ZN(new_n8854_));
  NAND2_X1   g06053(.A1(new_n8854_), .A2(new_n8849_), .ZN(new_n8855_));
  NAND2_X1   g06054(.A1(new_n8849_), .A2(new_n6400_), .ZN(new_n8856_));
  NAND4_X1   g06055(.A1(new_n8771_), .A2(new_n8547_), .A3(new_n8779_), .A4(new_n8856_), .ZN(new_n8857_));
  NOR3_X1    g06056(.A1(new_n8645_), .A2(new_n8646_), .A3(new_n8773_), .ZN(new_n8858_));
  OAI21_X1   g06057(.A1(new_n8858_), .A2(new_n5551_), .B(new_n8777_), .ZN(new_n8859_));
  NAND2_X1   g06058(.A1(new_n8562_), .A2(new_n8830_), .ZN(new_n8860_));
  NAND4_X1   g06059(.A1(new_n8859_), .A2(pi0039), .A3(new_n6399_), .A4(new_n8860_), .ZN(new_n8861_));
  AOI21_X1   g06060(.A1(new_n8857_), .A2(new_n8855_), .B(new_n8861_), .ZN(new_n8862_));
  AOI22_X1   g06061(.A1(new_n8853_), .A2(new_n8862_), .B1(new_n8561_), .B2(new_n8771_), .ZN(new_n8863_));
  AOI21_X1   g06062(.A1(new_n8562_), .A2(new_n8696_), .B(new_n8805_), .ZN(new_n8864_));
  NOR2_X1    g06063(.A1(new_n8562_), .A2(new_n3133_), .ZN(new_n8865_));
  OAI21_X1   g06064(.A1(new_n8803_), .A2(new_n8864_), .B(new_n8865_), .ZN(new_n8866_));
  NAND2_X1   g06065(.A1(new_n8795_), .A2(new_n8866_), .ZN(new_n8867_));
  AOI21_X1   g06066(.A1(new_n8556_), .A2(pi0039), .B(pi0232), .ZN(new_n8868_));
  NOR2_X1    g06067(.A1(new_n8812_), .A2(new_n8868_), .ZN(new_n8869_));
  AOI21_X1   g06068(.A1(new_n8867_), .A2(new_n8869_), .B(pi0075), .ZN(new_n8870_));
  NAND3_X1   g06069(.A1(new_n8559_), .A2(pi0039), .A3(po1038), .ZN(new_n8871_));
  NOR4_X1    g06070(.A1(new_n8863_), .A2(new_n8870_), .A3(new_n8842_), .A4(new_n8871_), .ZN(new_n8872_));
  AOI21_X1   g06071(.A1(new_n8848_), .A2(new_n8872_), .B(pi0039), .ZN(new_n8873_));
  NOR3_X1    g06072(.A1(new_n8873_), .A2(new_n8630_), .A3(new_n8743_), .ZN(po0201));
  NAND2_X1   g06073(.A1(new_n8432_), .A2(new_n2730_), .ZN(new_n8875_));
  NOR2_X1    g06074(.A1(new_n8425_), .A2(new_n8390_), .ZN(new_n8876_));
  NAND2_X1   g06075(.A1(new_n8875_), .A2(new_n8876_), .ZN(new_n8877_));
  NAND2_X1   g06076(.A1(new_n8420_), .A2(new_n2730_), .ZN(new_n8878_));
  NAND3_X1   g06077(.A1(new_n8878_), .A2(pi0044), .A3(new_n8411_), .ZN(new_n8879_));
  AOI21_X1   g06078(.A1(new_n8879_), .A2(new_n8877_), .B(new_n3005_), .ZN(new_n8880_));
  NOR2_X1    g06079(.A1(new_n8480_), .A2(new_n5401_), .ZN(new_n8881_));
  NOR2_X1    g06080(.A1(new_n8881_), .A2(pi0072), .ZN(new_n8882_));
  NOR2_X1    g06081(.A1(new_n3132_), .A2(pi0039), .ZN(new_n8883_));
  INV_X1     g06082(.I(new_n8883_), .ZN(new_n8884_));
  OAI21_X1   g06083(.A1(new_n8882_), .A2(new_n8884_), .B(new_n6495_), .ZN(new_n8885_));
  NAND2_X1   g06084(.A1(new_n8885_), .A2(new_n3183_), .ZN(new_n8886_));
  INV_X1     g06085(.I(new_n8473_), .ZN(new_n8887_));
  OR3_X2     g06086(.A1(new_n8532_), .A2(new_n8390_), .A3(new_n3005_), .Z(new_n8888_));
  NAND3_X1   g06087(.A1(new_n8532_), .A2(pi0044), .A3(new_n3005_), .ZN(new_n8889_));
  AOI21_X1   g06088(.A1(new_n8888_), .A2(new_n8889_), .B(new_n8887_), .ZN(new_n8890_));
  OAI21_X1   g06089(.A1(new_n8880_), .A2(new_n8886_), .B(new_n8890_), .ZN(new_n8891_));
  NOR3_X1    g06090(.A1(new_n6531_), .A2(new_n3183_), .A3(new_n2437_), .ZN(new_n8892_));
  NOR3_X1    g06091(.A1(new_n6495_), .A2(new_n3183_), .A3(pi0072), .ZN(new_n8893_));
  OAI21_X1   g06092(.A1(new_n8892_), .A2(new_n8893_), .B(pi0044), .ZN(new_n8894_));
  NAND2_X1   g06093(.A1(new_n8894_), .A2(pi0038), .ZN(new_n8895_));
  NAND2_X1   g06094(.A1(new_n8895_), .A2(new_n3455_), .ZN(new_n8896_));
  NOR2_X1    g06095(.A1(new_n8390_), .A2(new_n2437_), .ZN(new_n8897_));
  OAI21_X1   g06096(.A1(new_n6483_), .A2(pi1091), .B(new_n8897_), .ZN(new_n8898_));
  NOR4_X1    g06097(.A1(new_n6523_), .A2(new_n8390_), .A3(new_n3145_), .A4(new_n6504_), .ZN(new_n8899_));
  INV_X1     g06098(.I(new_n8899_), .ZN(new_n8900_));
  OAI21_X1   g06099(.A1(new_n8898_), .A2(new_n8900_), .B(new_n8390_), .ZN(new_n8901_));
  AOI21_X1   g06100(.A1(new_n2730_), .A2(new_n8391_), .B(new_n8494_), .ZN(new_n8902_));
  NOR3_X1    g06101(.A1(new_n6531_), .A2(new_n3183_), .A3(pi0072), .ZN(new_n8903_));
  AOI21_X1   g06102(.A1(new_n8494_), .A2(new_n8392_), .B(pi0039), .ZN(new_n8904_));
  AOI21_X1   g06103(.A1(new_n8903_), .A2(new_n8904_), .B(new_n8902_), .ZN(new_n8905_));
  NOR2_X1    g06104(.A1(new_n8509_), .A2(new_n8905_), .ZN(new_n8906_));
  AOI21_X1   g06105(.A1(new_n8906_), .A2(new_n8901_), .B(new_n3235_), .ZN(new_n8907_));
  NOR2_X1    g06106(.A1(new_n3187_), .A2(new_n3235_), .ZN(new_n8908_));
  XNOR2_X1   g06107(.A1(new_n8907_), .A2(new_n8908_), .ZN(new_n8909_));
  NOR2_X1    g06108(.A1(new_n8909_), .A2(new_n8894_), .ZN(new_n8910_));
  NAND4_X1   g06109(.A1(new_n3160_), .A2(pi0044), .A3(pi0228), .A4(new_n3132_), .ZN(new_n8911_));
  NAND3_X1   g06110(.A1(new_n8480_), .A2(new_n3005_), .A3(new_n8392_), .ZN(new_n8912_));
  AOI21_X1   g06111(.A1(pi0039), .A2(pi0087), .B(new_n6495_), .ZN(new_n8913_));
  OAI21_X1   g06112(.A1(new_n8913_), .A2(new_n2437_), .B(new_n3183_), .ZN(new_n8914_));
  AOI21_X1   g06113(.A1(new_n8912_), .A2(new_n3132_), .B(new_n8914_), .ZN(new_n8915_));
  OAI21_X1   g06114(.A1(new_n8915_), .A2(new_n8911_), .B(new_n3235_), .ZN(new_n8916_));
  NOR3_X1    g06115(.A1(new_n8479_), .A2(new_n3145_), .A3(new_n6504_), .ZN(new_n8917_));
  NOR3_X1    g06116(.A1(new_n8479_), .A2(new_n8390_), .A3(new_n6486_), .ZN(new_n8918_));
  XNOR2_X1   g06117(.A1(new_n8917_), .A2(new_n8918_), .ZN(new_n8919_));
  NAND3_X1   g06118(.A1(new_n8714_), .A2(new_n7240_), .A3(new_n8391_), .ZN(new_n8921_));
  OAI21_X1   g06119(.A1(new_n8894_), .A2(new_n8921_), .B(new_n6400_), .ZN(new_n8922_));
  NAND2_X1   g06120(.A1(new_n8902_), .A2(new_n8904_), .ZN(new_n8923_));
  NAND2_X1   g06121(.A1(new_n8923_), .A2(new_n8898_), .ZN(new_n8924_));
  NOR2_X1    g06122(.A1(new_n8903_), .A2(new_n5506_), .ZN(new_n8925_));
  NAND3_X1   g06123(.A1(new_n8924_), .A2(new_n8922_), .A3(new_n8925_), .ZN(new_n8926_));
  NOR2_X1    g06124(.A1(new_n8919_), .A2(new_n8926_), .ZN(new_n8927_));
  OAI21_X1   g06125(.A1(new_n8910_), .A2(new_n8916_), .B(new_n8927_), .ZN(new_n8928_));
  AOI21_X1   g06126(.A1(new_n8891_), .A2(new_n8896_), .B(new_n8928_), .ZN(po0202));
  INV_X1     g06127(.I(new_n5679_), .ZN(new_n8930_));
  NOR2_X1    g06128(.A1(new_n3183_), .A2(pi0038), .ZN(new_n8931_));
  INV_X1     g06129(.I(new_n8931_), .ZN(new_n8932_));
  NOR2_X1    g06130(.A1(new_n8345_), .A2(new_n8932_), .ZN(new_n8933_));
  INV_X1     g06131(.I(new_n8933_), .ZN(new_n8934_));
  NOR3_X1    g06132(.A1(new_n8934_), .A2(new_n5405_), .A3(new_n8930_), .ZN(po0203));
  NOR3_X1    g06133(.A1(new_n2448_), .A2(new_n7285_), .A3(new_n2450_), .ZN(new_n8936_));
  NAND4_X1   g06134(.A1(new_n7284_), .A2(new_n6361_), .A3(new_n7288_), .A4(new_n8936_), .ZN(new_n8937_));
  INV_X1     g06135(.I(new_n8937_), .ZN(new_n8938_));
  NAND4_X1   g06136(.A1(pi0049), .A2(pi0068), .A3(pi0073), .A4(pi0076), .ZN(new_n8939_));
  NOR3_X1    g06137(.A1(pi0102), .A2(pi0104), .A3(pi0111), .ZN(new_n8940_));
  INV_X1     g06138(.I(new_n8940_), .ZN(new_n8941_));
  NAND2_X1   g06139(.A1(pi0082), .A2(pi0083), .ZN(new_n8942_));
  NOR4_X1    g06140(.A1(new_n8941_), .A2(new_n8310_), .A3(new_n8939_), .A4(new_n8942_), .ZN(new_n8943_));
  NAND4_X1   g06141(.A1(new_n8938_), .A2(new_n7275_), .A3(new_n8357_), .A4(new_n8943_), .ZN(new_n8944_));
  INV_X1     g06142(.I(new_n2469_), .ZN(new_n8945_));
  NAND2_X1   g06143(.A1(new_n2875_), .A2(new_n8945_), .ZN(new_n8946_));
  NOR2_X1    g06144(.A1(new_n8946_), .A2(new_n8944_), .ZN(new_n8947_));
  NAND2_X1   g06145(.A1(new_n8291_), .A2(new_n7262_), .ZN(new_n8948_));
  NOR2_X1    g06146(.A1(new_n8947_), .A2(new_n8948_), .ZN(po0204));
  NOR2_X1    g06147(.A1(new_n7277_), .A2(new_n6360_), .ZN(new_n8950_));
  INV_X1     g06148(.I(new_n8950_), .ZN(new_n8951_));
  AOI21_X1   g06149(.A1(new_n2544_), .A2(new_n8951_), .B(new_n2558_), .ZN(new_n8952_));
  NOR2_X1    g06150(.A1(new_n8952_), .A2(new_n2681_), .ZN(new_n8953_));
  NAND3_X1   g06151(.A1(new_n8309_), .A2(pi0104), .A3(new_n2599_), .ZN(new_n8954_));
  NAND2_X1   g06152(.A1(new_n2573_), .A2(new_n8310_), .ZN(new_n8955_));
  NAND3_X1   g06153(.A1(new_n8954_), .A2(new_n2605_), .A3(new_n8955_), .ZN(new_n8956_));
  NAND2_X1   g06154(.A1(new_n7286_), .A2(new_n7352_), .ZN(new_n8957_));
  NOR3_X1    g06155(.A1(new_n2448_), .A2(pi0067), .A3(pi0103), .ZN(new_n8958_));
  INV_X1     g06156(.I(new_n8958_), .ZN(new_n8959_));
  NOR4_X1    g06157(.A1(new_n8957_), .A2(new_n7361_), .A3(new_n8959_), .A4(new_n2558_), .ZN(new_n8960_));
  NAND2_X1   g06158(.A1(new_n8956_), .A2(new_n8960_), .ZN(new_n8961_));
  OR3_X2     g06159(.A1(new_n2618_), .A2(new_n6360_), .A3(new_n8961_), .Z(new_n8962_));
  NOR2_X1    g06160(.A1(new_n8962_), .A2(new_n8953_), .ZN(new_n8963_));
  INV_X1     g06161(.I(new_n8963_), .ZN(new_n8964_));
  NAND2_X1   g06162(.A1(new_n6422_), .A2(pi0058), .ZN(new_n8965_));
  NAND2_X1   g06163(.A1(new_n8964_), .A2(new_n8965_), .ZN(new_n8966_));
  AOI21_X1   g06164(.A1(new_n8966_), .A2(pi0091), .B(new_n8290_), .ZN(new_n8967_));
  NOR2_X1    g06165(.A1(new_n8967_), .A2(new_n2983_), .ZN(new_n8968_));
  NOR2_X1    g06166(.A1(new_n8961_), .A2(pi0036), .ZN(new_n8969_));
  OAI21_X1   g06167(.A1(new_n8969_), .A2(pi0088), .B(new_n8952_), .ZN(new_n8970_));
  NOR2_X1    g06168(.A1(new_n8970_), .A2(new_n8303_), .ZN(new_n8971_));
  NAND2_X1   g06169(.A1(new_n2981_), .A2(new_n2721_), .ZN(new_n8972_));
  OAI21_X1   g06170(.A1(new_n8971_), .A2(new_n8972_), .B(new_n5684_), .ZN(new_n8973_));
  AOI21_X1   g06171(.A1(new_n8967_), .A2(new_n2981_), .B(new_n8973_), .ZN(new_n8974_));
  NAND2_X1   g06172(.A1(new_n8974_), .A2(new_n2728_), .ZN(new_n8975_));
  XOR2_X1    g06173(.A1(new_n8975_), .A2(new_n8968_), .Z(new_n8976_));
  NAND2_X1   g06174(.A1(new_n8967_), .A2(new_n6403_), .ZN(new_n8977_));
  INV_X1     g06175(.I(new_n8977_), .ZN(new_n8978_));
  OR2_X2     g06176(.A1(new_n8974_), .A2(pi0829), .Z(new_n8979_));
  OAI21_X1   g06177(.A1(new_n5686_), .A2(new_n6940_), .B(new_n6403_), .ZN(new_n8980_));
  OAI21_X1   g06178(.A1(new_n8529_), .A2(new_n8980_), .B(new_n8285_), .ZN(new_n8981_));
  OR2_X2     g06179(.A1(new_n8978_), .A2(new_n8981_), .Z(new_n8982_));
  AOI22_X1   g06180(.A1(new_n8982_), .A2(new_n8384_), .B1(new_n8978_), .B2(new_n8979_), .ZN(new_n8983_));
  NOR3_X1    g06181(.A1(new_n8983_), .A2(new_n8976_), .A3(new_n2726_), .ZN(po0205));
  NOR3_X1    g06182(.A1(new_n2473_), .A2(pi0072), .A3(new_n2732_), .ZN(new_n8985_));
  NAND2_X1   g06183(.A1(new_n8985_), .A2(new_n2702_), .ZN(new_n8986_));
  NOR4_X1    g06184(.A1(new_n8288_), .A2(new_n8301_), .A3(new_n8359_), .A4(new_n8986_), .ZN(po0206));
  NAND4_X1   g06185(.A1(new_n8263_), .A2(pi0074), .A3(new_n6325_), .A4(new_n7240_), .ZN(new_n8988_));
  NAND4_X1   g06186(.A1(new_n7325_), .A2(new_n3175_), .A3(new_n6325_), .A4(new_n7240_), .ZN(new_n8989_));
  NOR4_X1    g06187(.A1(new_n8955_), .A2(new_n7361_), .A3(new_n8308_), .A4(new_n8941_), .ZN(new_n8990_));
  NOR2_X1    g06188(.A1(new_n7351_), .A2(new_n2448_), .ZN(new_n8991_));
  INV_X1     g06189(.I(new_n8991_), .ZN(new_n8992_));
  NOR3_X1    g06190(.A1(new_n2607_), .A2(new_n8356_), .A3(pi0103), .ZN(new_n8993_));
  NAND4_X1   g06191(.A1(new_n8993_), .A2(new_n7286_), .A3(pi0068), .A4(pi0073), .ZN(new_n8994_));
  NOR2_X1    g06192(.A1(new_n8992_), .A2(new_n8994_), .ZN(new_n8995_));
  NAND2_X1   g06193(.A1(new_n8995_), .A2(new_n8990_), .ZN(new_n8996_));
  NOR3_X1    g06194(.A1(new_n8996_), .A2(new_n2475_), .A3(new_n7408_), .ZN(new_n8997_));
  NAND3_X1   g06195(.A1(new_n8997_), .A2(new_n8289_), .A3(new_n8985_), .ZN(new_n8998_));
  AOI21_X1   g06196(.A1(new_n8988_), .A2(new_n8989_), .B(new_n8998_), .ZN(po0207));
  NAND2_X1   g06197(.A1(new_n5502_), .A2(pi0100), .ZN(new_n9000_));
  AOI21_X1   g06198(.A1(new_n7272_), .A2(new_n2530_), .B(new_n2460_), .ZN(new_n9001_));
  NAND2_X1   g06199(.A1(new_n7264_), .A2(new_n9001_), .ZN(new_n9002_));
  INV_X1     g06200(.I(new_n7315_), .ZN(new_n9003_));
  NAND2_X1   g06201(.A1(po0840), .A2(pi0252), .ZN(new_n9004_));
  OAI21_X1   g06202(.A1(new_n9003_), .A2(pi0252), .B(new_n9004_), .ZN(new_n9005_));
  NAND4_X1   g06203(.A1(new_n8451_), .A2(new_n8529_), .A3(new_n9002_), .A4(new_n9005_), .ZN(new_n9006_));
  AOI21_X1   g06204(.A1(new_n9006_), .A2(new_n7272_), .B(new_n7270_), .ZN(new_n9007_));
  INV_X1     g06205(.I(new_n6386_), .ZN(new_n9008_));
  NOR2_X1    g06206(.A1(new_n9008_), .A2(new_n2796_), .ZN(new_n9009_));
  NOR2_X1    g06207(.A1(new_n7272_), .A2(new_n2679_), .ZN(new_n9010_));
  AND4_X2    g06208(.A1(new_n7271_), .A2(new_n9005_), .A3(new_n9009_), .A4(new_n9010_), .Z(new_n9011_));
  NOR4_X1    g06209(.A1(new_n9007_), .A2(new_n3462_), .A3(new_n5730_), .A4(new_n9011_), .ZN(new_n9012_));
  XOR2_X1    g06210(.A1(new_n9012_), .A2(new_n9000_), .Z(new_n9013_));
  INV_X1     g06211(.I(new_n5527_), .ZN(new_n9014_));
  INV_X1     g06212(.I(new_n7337_), .ZN(new_n9015_));
  NOR4_X1    g06213(.A1(new_n9014_), .A2(new_n7294_), .A3(new_n7331_), .A4(new_n9015_), .ZN(new_n9016_));
  AOI22_X1   g06214(.A1(new_n9016_), .A2(new_n8263_), .B1(new_n3171_), .B2(new_n3211_), .ZN(new_n9017_));
  NOR2_X1    g06215(.A1(new_n9013_), .A2(new_n9017_), .ZN(po0208));
  NOR3_X1    g06216(.A1(new_n8292_), .A2(new_n5420_), .A3(new_n2682_), .ZN(new_n9019_));
  INV_X1     g06217(.I(new_n9019_), .ZN(new_n9020_));
  NOR2_X1    g06218(.A1(new_n8992_), .A2(new_n7355_), .ZN(new_n9021_));
  NAND3_X1   g06219(.A1(new_n9021_), .A2(new_n2623_), .A3(new_n2446_), .ZN(new_n9022_));
  NOR4_X1    g06220(.A1(new_n9020_), .A2(new_n2604_), .A3(new_n2607_), .A4(new_n9022_), .ZN(po0209));
  NOR2_X1    g06221(.A1(new_n5511_), .A2(pi0072), .ZN(new_n9024_));
  INV_X1     g06222(.I(new_n9024_), .ZN(new_n9025_));
  NOR2_X1    g06223(.A1(new_n9025_), .A2(pi0039), .ZN(new_n9026_));
  NOR2_X1    g06224(.A1(new_n8747_), .A2(pi0043), .ZN(new_n9027_));
  NOR2_X1    g06225(.A1(new_n8494_), .A2(new_n8609_), .ZN(new_n9028_));
  NAND2_X1   g06226(.A1(new_n9028_), .A2(new_n9027_), .ZN(new_n9029_));
  NOR2_X1    g06227(.A1(new_n6486_), .A2(new_n9024_), .ZN(new_n9030_));
  AOI21_X1   g06228(.A1(new_n8817_), .A2(new_n9030_), .B(new_n9029_), .ZN(new_n9031_));
  NOR2_X1    g06229(.A1(new_n8609_), .A2(new_n8584_), .ZN(new_n9032_));
  NAND2_X1   g06230(.A1(new_n8608_), .A2(pi0052), .ZN(new_n9033_));
  XNOR2_X1   g06231(.A1(new_n9032_), .A2(new_n9033_), .ZN(new_n9034_));
  AOI21_X1   g06232(.A1(new_n2730_), .A2(new_n5514_), .B(new_n5511_), .ZN(new_n9035_));
  NAND4_X1   g06233(.A1(new_n8590_), .A2(new_n8577_), .A3(new_n9034_), .A4(new_n9035_), .ZN(new_n9036_));
  NAND2_X1   g06234(.A1(new_n9036_), .A2(new_n5511_), .ZN(new_n9037_));
  AND3_X2    g06235(.A1(new_n9037_), .A2(new_n8571_), .A3(new_n9027_), .Z(new_n9038_));
  NAND3_X1   g06236(.A1(new_n9038_), .A2(pi0039), .A3(pi0100), .ZN(new_n9039_));
  INV_X1     g06237(.I(new_n9038_), .ZN(new_n9040_));
  NAND3_X1   g06238(.A1(new_n9040_), .A2(new_n3183_), .A3(pi0100), .ZN(new_n9041_));
  NAND2_X1   g06239(.A1(new_n9041_), .A2(new_n9039_), .ZN(new_n9042_));
  AOI21_X1   g06240(.A1(new_n9042_), .A2(new_n9031_), .B(new_n3259_), .ZN(new_n9043_));
  XOR2_X1    g06241(.A1(new_n9043_), .A2(new_n7487_), .Z(new_n9044_));
  NOR2_X1    g06242(.A1(new_n8932_), .A2(pi0100), .ZN(new_n9045_));
  OAI22_X1   g06243(.A1(new_n3455_), .A2(new_n9045_), .B1(new_n9026_), .B2(new_n3462_), .ZN(new_n9046_));
  AOI21_X1   g06244(.A1(new_n9044_), .A2(new_n9026_), .B(new_n9046_), .ZN(new_n9047_));
  INV_X1     g06245(.I(new_n8573_), .ZN(new_n9048_));
  NOR4_X1    g06246(.A1(new_n9048_), .A2(new_n5510_), .A3(new_n5514_), .A4(new_n3005_), .ZN(new_n9049_));
  OAI21_X1   g06247(.A1(new_n8619_), .A2(pi0052), .B(new_n9049_), .ZN(new_n9050_));
  AOI21_X1   g06248(.A1(new_n8818_), .A2(pi0052), .B(new_n9050_), .ZN(new_n9051_));
  NAND2_X1   g06249(.A1(new_n9049_), .A2(new_n9024_), .ZN(new_n9052_));
  XOR2_X1    g06250(.A1(new_n9051_), .A2(new_n9052_), .Z(new_n9053_));
  NAND2_X1   g06251(.A1(new_n9053_), .A2(pi0038), .ZN(new_n9054_));
  XOR2_X1    g06252(.A1(new_n9054_), .A2(new_n5486_), .Z(new_n9055_));
  NAND2_X1   g06253(.A1(new_n9055_), .A2(new_n9026_), .ZN(new_n9056_));
  OAI21_X1   g06254(.A1(new_n9047_), .A2(new_n9056_), .B(new_n6399_), .ZN(new_n9057_));
  XOR2_X1    g06255(.A1(new_n9057_), .A2(new_n8744_), .Z(new_n9058_));
  INV_X1     g06256(.I(new_n9026_), .ZN(new_n9059_));
  NOR2_X1    g06257(.A1(new_n8671_), .A2(new_n9029_), .ZN(new_n9060_));
  AOI21_X1   g06258(.A1(new_n9060_), .A2(new_n3186_), .B(new_n9059_), .ZN(new_n9061_));
  OAI21_X1   g06259(.A1(new_n9026_), .A2(new_n6399_), .B(new_n8547_), .ZN(new_n9062_));
  NAND2_X1   g06260(.A1(new_n8859_), .A2(pi0039), .ZN(new_n9063_));
  NOR2_X1    g06261(.A1(new_n9031_), .A2(pi0039), .ZN(new_n9064_));
  NOR2_X1    g06262(.A1(new_n9024_), .A2(pi0039), .ZN(new_n9065_));
  NOR2_X1    g06263(.A1(new_n8779_), .A2(new_n9065_), .ZN(new_n9066_));
  NOR3_X1    g06264(.A1(new_n3462_), .A2(pi0038), .A3(pi0087), .ZN(new_n9067_));
  OAI21_X1   g06265(.A1(new_n9064_), .A2(new_n9067_), .B(new_n8851_), .ZN(new_n9068_));
  AOI21_X1   g06266(.A1(new_n9040_), .A2(new_n9068_), .B(new_n9063_), .ZN(new_n9069_));
  NOR2_X1    g06267(.A1(new_n9053_), .A2(pi0039), .ZN(new_n9070_));
  NOR2_X1    g06268(.A1(new_n9070_), .A2(new_n3133_), .ZN(new_n9071_));
  NAND2_X1   g06269(.A1(new_n8851_), .A2(new_n9066_), .ZN(new_n9072_));
  XOR2_X1    g06270(.A1(new_n9071_), .A2(new_n9072_), .Z(new_n9073_));
  INV_X1     g06271(.I(new_n9066_), .ZN(new_n9074_));
  OAI21_X1   g06272(.A1(new_n9074_), .A2(new_n3186_), .B(pi0075), .ZN(new_n9075_));
  NOR2_X1    g06273(.A1(new_n8779_), .A2(new_n3186_), .ZN(new_n9076_));
  NOR2_X1    g06274(.A1(new_n8740_), .A2(pi0211), .ZN(new_n9077_));
  INV_X1     g06275(.I(new_n9077_), .ZN(new_n9078_));
  NOR2_X1    g06276(.A1(new_n9078_), .A2(pi0219), .ZN(new_n9079_));
  NOR2_X1    g06277(.A1(new_n3455_), .A2(pi0039), .ZN(new_n9080_));
  NAND4_X1   g06278(.A1(new_n9079_), .A2(new_n6399_), .A3(new_n8547_), .A4(new_n9080_), .ZN(new_n9081_));
  AOI21_X1   g06279(.A1(new_n9075_), .A2(new_n9076_), .B(new_n9081_), .ZN(new_n9082_));
  OAI21_X1   g06280(.A1(new_n9060_), .A2(new_n9025_), .B(new_n9082_), .ZN(new_n9083_));
  NOR2_X1    g06281(.A1(new_n9073_), .A2(new_n9083_), .ZN(new_n9084_));
  OAI21_X1   g06282(.A1(new_n9069_), .A2(pi0075), .B(new_n9084_), .ZN(new_n9085_));
  NAND2_X1   g06283(.A1(new_n9085_), .A2(new_n9062_), .ZN(new_n9086_));
  NAND3_X1   g06284(.A1(new_n9058_), .A2(new_n9061_), .A3(new_n9086_), .ZN(new_n9087_));
  NAND3_X1   g06285(.A1(new_n9079_), .A2(pi0039), .A3(new_n8629_), .ZN(new_n9088_));
  AOI21_X1   g06286(.A1(new_n7240_), .A2(new_n9059_), .B(new_n9088_), .ZN(new_n9089_));
  INV_X1     g06287(.I(new_n8547_), .ZN(new_n9090_));
  NAND3_X1   g06288(.A1(new_n9074_), .A2(new_n7240_), .A3(new_n9090_), .ZN(new_n9091_));
  AOI21_X1   g06289(.A1(new_n9091_), .A2(new_n6399_), .B(new_n9089_), .ZN(new_n9092_));
  AOI21_X1   g06290(.A1(new_n9038_), .A2(new_n3132_), .B(pi0039), .ZN(new_n9093_));
  NAND3_X1   g06291(.A1(pi0072), .A2(pi0232), .A3(pi0299), .ZN(new_n9094_));
  NOR2_X1    g06292(.A1(new_n9064_), .A2(new_n8632_), .ZN(new_n9095_));
  OAI22_X1   g06293(.A1(new_n9093_), .A2(new_n9094_), .B1(new_n5506_), .B2(new_n9095_), .ZN(new_n9096_));
  INV_X1     g06294(.I(new_n8839_), .ZN(new_n9097_));
  INV_X1     g06295(.I(new_n9064_), .ZN(new_n9098_));
  NOR2_X1    g06296(.A1(new_n8632_), .A2(new_n9065_), .ZN(new_n9099_));
  INV_X1     g06297(.I(new_n9099_), .ZN(new_n9100_));
  NAND4_X1   g06298(.A1(new_n9074_), .A2(pi0038), .A3(new_n5505_), .A4(new_n9100_), .ZN(new_n9101_));
  AOI21_X1   g06299(.A1(new_n9098_), .A2(new_n9101_), .B(new_n9097_), .ZN(new_n9102_));
  AOI21_X1   g06300(.A1(new_n9099_), .A2(new_n3133_), .B(new_n3455_), .ZN(new_n9103_));
  OAI21_X1   g06301(.A1(new_n9074_), .A2(new_n3132_), .B(new_n9103_), .ZN(new_n9104_));
  NAND3_X1   g06302(.A1(new_n9104_), .A2(new_n3133_), .A3(new_n8829_), .ZN(new_n9105_));
  AOI21_X1   g06303(.A1(new_n9070_), .A2(new_n9105_), .B(new_n8547_), .ZN(new_n9106_));
  INV_X1     g06304(.I(new_n9103_), .ZN(new_n9107_));
  NOR3_X1    g06305(.A1(new_n9070_), .A2(new_n3133_), .A3(new_n8632_), .ZN(new_n9108_));
  NOR2_X1    g06306(.A1(new_n9108_), .A2(new_n9107_), .ZN(new_n9109_));
  NAND2_X1   g06307(.A1(new_n8547_), .A2(pi0087), .ZN(new_n9110_));
  NOR4_X1    g06308(.A1(new_n9109_), .A2(new_n8837_), .A3(new_n9106_), .A4(new_n9110_), .ZN(new_n9111_));
  OAI21_X1   g06309(.A1(new_n9038_), .A2(new_n9102_), .B(new_n9111_), .ZN(new_n9112_));
  NAND2_X1   g06310(.A1(new_n9112_), .A2(new_n3455_), .ZN(new_n9113_));
  NOR3_X1    g06311(.A1(new_n8829_), .A2(new_n3235_), .A3(new_n9090_), .ZN(new_n9114_));
  NOR3_X1    g06312(.A1(new_n8781_), .A2(new_n3235_), .A3(new_n8547_), .ZN(new_n9115_));
  NOR2_X1    g06313(.A1(new_n8633_), .A2(new_n6400_), .ZN(new_n9116_));
  OAI21_X1   g06314(.A1(new_n9114_), .A2(new_n9115_), .B(new_n9116_), .ZN(new_n9117_));
  NAND2_X1   g06315(.A1(new_n9117_), .A2(new_n3183_), .ZN(new_n9118_));
  NAND2_X1   g06316(.A1(new_n9100_), .A2(new_n6400_), .ZN(new_n9119_));
  NAND4_X1   g06317(.A1(new_n9061_), .A2(new_n9079_), .A3(new_n9118_), .A4(new_n9119_), .ZN(new_n9120_));
  NAND2_X1   g06318(.A1(new_n9120_), .A2(new_n3235_), .ZN(new_n9121_));
  NOR2_X1    g06319(.A1(new_n9100_), .A2(new_n3259_), .ZN(new_n9122_));
  NAND4_X1   g06320(.A1(new_n9096_), .A2(new_n9113_), .A3(new_n9121_), .A4(new_n9122_), .ZN(new_n9123_));
  AOI21_X1   g06321(.A1(new_n9087_), .A2(new_n9092_), .B(new_n9123_), .ZN(po0210));
  INV_X1     g06322(.I(new_n2860_), .ZN(new_n9125_));
  NOR4_X1    g06323(.A1(new_n9125_), .A2(new_n2518_), .A3(new_n2897_), .A4(new_n2903_), .ZN(new_n9126_));
  NAND3_X1   g06324(.A1(new_n9126_), .A2(pi0024), .A3(new_n8529_), .ZN(new_n9127_));
  NOR2_X1    g06325(.A1(new_n5404_), .A2(pi0979), .ZN(new_n9128_));
  AOI21_X1   g06326(.A1(new_n9128_), .A2(new_n3183_), .B(new_n5401_), .ZN(new_n9129_));
  NOR2_X1    g06327(.A1(new_n8347_), .A2(new_n9129_), .ZN(new_n9130_));
  NAND2_X1   g06328(.A1(new_n9127_), .A2(new_n9130_), .ZN(new_n9131_));
  NAND2_X1   g06329(.A1(new_n9130_), .A2(pi0039), .ZN(new_n9132_));
  XNOR2_X1   g06330(.A1(new_n9131_), .A2(new_n9132_), .ZN(new_n9133_));
  NOR2_X1    g06331(.A1(new_n9133_), .A2(new_n3145_), .ZN(po0211));
  NOR2_X1    g06332(.A1(new_n3187_), .A2(new_n3189_), .ZN(new_n9135_));
  NAND2_X1   g06333(.A1(new_n8296_), .A2(new_n9135_), .ZN(new_n9136_));
  NAND2_X1   g06334(.A1(new_n9136_), .A2(new_n7330_), .ZN(new_n9137_));
  NAND2_X1   g06335(.A1(new_n7330_), .A2(pi0054), .ZN(new_n9138_));
  XNOR2_X1   g06336(.A1(new_n9137_), .A2(new_n9138_), .ZN(new_n9139_));
  NAND3_X1   g06337(.A1(pi0089), .A2(pi0102), .A3(pi0106), .ZN(new_n9140_));
  NAND2_X1   g06338(.A1(new_n2519_), .A2(new_n2575_), .ZN(new_n9141_));
  NOR4_X1    g06339(.A1(new_n2610_), .A2(new_n9141_), .A3(new_n8939_), .A4(new_n9140_), .ZN(new_n9142_));
  NAND4_X1   g06340(.A1(new_n7290_), .A2(new_n8991_), .A3(new_n8993_), .A4(new_n9142_), .ZN(new_n9143_));
  NOR4_X1    g06341(.A1(new_n9143_), .A2(new_n7580_), .A3(pi0053), .A4(new_n7270_), .ZN(new_n9144_));
  NOR3_X1    g06342(.A1(new_n7323_), .A2(pi0841), .A3(new_n2479_), .ZN(new_n9145_));
  NAND4_X1   g06343(.A1(new_n9144_), .A2(new_n2474_), .A3(new_n3195_), .A4(new_n9145_), .ZN(new_n9146_));
  NOR2_X1    g06344(.A1(new_n9139_), .A2(new_n9146_), .ZN(po0212));
  NOR2_X1    g06345(.A1(new_n9136_), .A2(pi0054), .ZN(new_n9148_));
  INV_X1     g06346(.I(new_n9148_), .ZN(new_n9149_));
  NOR4_X1    g06347(.A1(new_n7680_), .A2(new_n2457_), .A3(new_n3292_), .A4(new_n3138_), .ZN(new_n9150_));
  NOR2_X1    g06348(.A1(new_n7329_), .A2(new_n3258_), .ZN(new_n9151_));
  NAND4_X1   g06349(.A1(new_n2440_), .A2(new_n2534_), .A3(new_n2536_), .A4(new_n2539_), .ZN(new_n9152_));
  NOR2_X1    g06350(.A1(new_n8994_), .A2(new_n9152_), .ZN(new_n9153_));
  INV_X1     g06351(.I(new_n9153_), .ZN(new_n9154_));
  NOR2_X1    g06352(.A1(new_n9154_), .A2(new_n3258_), .ZN(new_n9155_));
  OAI21_X1   g06353(.A1(new_n9150_), .A2(new_n9151_), .B(new_n9155_), .ZN(new_n9156_));
  AOI21_X1   g06354(.A1(new_n9149_), .A2(new_n9156_), .B(new_n3175_), .ZN(po0213));
  OAI21_X1   g06355(.A1(new_n3258_), .A2(new_n3201_), .B(new_n3426_), .ZN(new_n9158_));
  AOI21_X1   g06356(.A1(new_n8224_), .A2(pi0056), .B(new_n9158_), .ZN(new_n9159_));
  NOR2_X1    g06357(.A1(new_n3224_), .A2(new_n7401_), .ZN(new_n9160_));
  NAND2_X1   g06358(.A1(new_n5465_), .A2(new_n9160_), .ZN(new_n9161_));
  NOR3_X1    g06359(.A1(new_n9161_), .A2(new_n3219_), .A3(new_n9159_), .ZN(po0214));
  INV_X1     g06360(.I(new_n5785_), .ZN(new_n9163_));
  NAND3_X1   g06361(.A1(new_n9148_), .A2(new_n3175_), .A3(new_n9163_), .ZN(new_n9164_));
  NAND2_X1   g06362(.A1(new_n9164_), .A2(pi0057), .ZN(new_n9165_));
  XOR2_X1    g06363(.A1(new_n9165_), .A2(new_n5546_), .Z(new_n9166_));
  INV_X1     g06364(.I(pi0924), .ZN(new_n9167_));
  NAND2_X1   g06365(.A1(new_n9160_), .A2(new_n5557_), .ZN(new_n9168_));
  NOR2_X1    g06366(.A1(new_n9168_), .A2(pi0062), .ZN(new_n9169_));
  AOI21_X1   g06367(.A1(new_n9160_), .A2(new_n5557_), .B(new_n3201_), .ZN(new_n9170_));
  OAI22_X1   g06368(.A1(new_n9169_), .A2(new_n9170_), .B1(new_n9167_), .B2(new_n3225_), .ZN(new_n9171_));
  NOR2_X1    g06369(.A1(new_n9166_), .A2(new_n9171_), .ZN(po0215));
  INV_X1     g06370(.I(new_n9009_), .ZN(new_n9173_));
  NOR4_X1    g06371(.A1(new_n8288_), .A2(new_n2679_), .A3(pi0093), .A4(new_n9173_), .ZN(new_n9174_));
  AND2_X2    g06372(.A1(new_n8259_), .A2(new_n9174_), .Z(po0216));
  NAND2_X1   g06373(.A1(new_n9164_), .A2(pi0059), .ZN(new_n9176_));
  XOR2_X1    g06374(.A1(new_n9176_), .A2(new_n5546_), .Z(new_n9177_));
  NOR4_X1    g06375(.A1(new_n9177_), .A2(new_n9167_), .A3(new_n3221_), .A4(new_n9168_), .ZN(po0217));
  NOR2_X1    g06376(.A1(new_n3183_), .A2(new_n3721_), .ZN(new_n9179_));
  NAND4_X1   g06377(.A1(new_n5679_), .A2(pi1001), .A3(new_n9128_), .A4(new_n9179_), .ZN(new_n9180_));
  NOR3_X1    g06378(.A1(new_n7270_), .A2(pi0053), .A3(new_n7580_), .ZN(new_n9181_));
  NAND4_X1   g06379(.A1(new_n9181_), .A2(pi0024), .A3(pi0039), .A4(new_n8529_), .ZN(new_n9182_));
  NAND3_X1   g06380(.A1(new_n9182_), .A2(new_n9180_), .A3(new_n2519_), .ZN(new_n9183_));
  AOI21_X1   g06381(.A1(new_n9183_), .A2(new_n2458_), .B(new_n8347_), .ZN(po0218));
  NOR2_X1    g06382(.A1(new_n7272_), .A2(new_n2519_), .ZN(new_n9185_));
  NAND4_X1   g06383(.A1(new_n8291_), .A2(new_n2458_), .A3(new_n9181_), .A4(new_n9185_), .ZN(new_n9186_));
  AOI21_X1   g06384(.A1(new_n9186_), .A2(new_n2732_), .B(new_n8944_), .ZN(po0219));
  NAND2_X1   g06385(.A1(new_n8225_), .A2(pi0057), .ZN(new_n9188_));
  XOR2_X1    g06386(.A1(new_n9188_), .A2(new_n5546_), .Z(new_n9189_));
  NOR4_X1    g06387(.A1(new_n9189_), .A2(pi0056), .A3(new_n3201_), .A4(new_n9161_), .ZN(po0220));
  INV_X1     g06388(.I(pi0063), .ZN(new_n9191_));
  NOR4_X1    g06389(.A1(new_n7578_), .A2(new_n9191_), .A3(new_n2565_), .A4(new_n7408_), .ZN(new_n9192_));
  INV_X1     g06390(.I(new_n9192_), .ZN(new_n9193_));
  NOR2_X1    g06391(.A1(new_n9193_), .A2(new_n8946_), .ZN(new_n9194_));
  NAND2_X1   g06392(.A1(pi0024), .A2(pi0999), .ZN(new_n9195_));
  NAND2_X1   g06393(.A1(new_n8291_), .A2(new_n9195_), .ZN(new_n9196_));
  NOR2_X1    g06394(.A1(new_n9194_), .A2(new_n9196_), .ZN(po0221));
  NAND3_X1   g06395(.A1(new_n2642_), .A2(new_n2644_), .A3(new_n2565_), .ZN(new_n9198_));
  NOR2_X1    g06396(.A1(new_n9191_), .A2(new_n2492_), .ZN(new_n9199_));
  NAND4_X1   g06397(.A1(new_n9198_), .A2(new_n8304_), .A3(new_n2645_), .A4(new_n9199_), .ZN(new_n9200_));
  NAND2_X1   g06398(.A1(new_n9200_), .A2(new_n9019_), .ZN(new_n9201_));
  NAND2_X1   g06399(.A1(new_n9019_), .A2(pi0841), .ZN(new_n9202_));
  XNOR2_X1   g06400(.A1(new_n9201_), .A2(new_n9202_), .ZN(new_n9203_));
  NOR4_X1    g06401(.A1(new_n9203_), .A2(pi0063), .A3(new_n2565_), .A4(new_n7578_), .ZN(po0222));
  NOR3_X1    g06402(.A1(new_n3183_), .A2(new_n8319_), .A3(pi1082), .ZN(new_n9205_));
  INV_X1     g06403(.I(new_n9205_), .ZN(new_n9206_));
  NOR4_X1    g06404(.A1(new_n8333_), .A2(new_n8340_), .A3(new_n8347_), .A4(new_n9206_), .ZN(po0223));
  NOR2_X1    g06405(.A1(pi0199), .A2(pi0299), .ZN(new_n9208_));
  INV_X1     g06406(.I(new_n9208_), .ZN(new_n9209_));
  NAND4_X1   g06407(.A1(new_n7679_), .A2(pi0314), .A3(new_n2456_), .A4(new_n3137_), .ZN(new_n9210_));
  NOR4_X1    g06408(.A1(new_n9210_), .A2(new_n2492_), .A3(new_n2454_), .A4(new_n2453_), .ZN(new_n9211_));
  NAND2_X1   g06409(.A1(new_n9211_), .A2(new_n3291_), .ZN(new_n9212_));
  NOR2_X1    g06410(.A1(new_n7240_), .A2(new_n8683_), .ZN(new_n9213_));
  NOR2_X1    g06411(.A1(new_n8549_), .A2(pi0299), .ZN(new_n9214_));
  NAND4_X1   g06412(.A1(new_n9214_), .A2(pi0219), .A3(new_n3132_), .A4(new_n3191_), .ZN(new_n9215_));
  NOR2_X1    g06413(.A1(new_n3288_), .A2(new_n9215_), .ZN(new_n9216_));
  OAI21_X1   g06414(.A1(new_n9211_), .A2(new_n9213_), .B(new_n9216_), .ZN(new_n9217_));
  AOI21_X1   g06415(.A1(new_n9217_), .A2(new_n9212_), .B(new_n9209_), .ZN(po0224));
  NAND3_X1   g06416(.A1(new_n9021_), .A2(pi0083), .A3(pi0103), .ZN(new_n9219_));
  NOR4_X1    g06417(.A1(new_n2626_), .A2(new_n8288_), .A3(new_n9210_), .A4(new_n9219_), .ZN(po0225));
  INV_X1     g06418(.I(new_n5689_), .ZN(new_n9221_));
  NAND2_X1   g06419(.A1(new_n9221_), .A2(new_n5460_), .ZN(new_n9222_));
  NOR3_X1    g06420(.A1(new_n5293_), .A2(new_n3011_), .A3(pi0221), .ZN(new_n9223_));
  NOR2_X1    g06421(.A1(new_n5689_), .A2(new_n5400_), .ZN(new_n9224_));
  NAND2_X1   g06422(.A1(new_n3386_), .A2(new_n3381_), .ZN(new_n9225_));
  NOR2_X1    g06423(.A1(new_n8934_), .A2(new_n9225_), .ZN(new_n9226_));
  AOI21_X1   g06424(.A1(new_n9224_), .A2(new_n9226_), .B(new_n9223_), .ZN(new_n9227_));
  NOR2_X1    g06425(.A1(new_n9227_), .A2(new_n9222_), .ZN(po0226));
  NAND4_X1   g06426(.A1(new_n8275_), .A2(pi0071), .A3(pi0314), .A4(new_n6361_), .ZN(new_n9229_));
  NOR3_X1    g06427(.A1(new_n2607_), .A2(new_n2623_), .A3(pi0103), .ZN(new_n9230_));
  INV_X1     g06428(.I(pi0314), .ZN(new_n9231_));
  INV_X1     g06429(.I(new_n5579_), .ZN(new_n9232_));
  NOR4_X1    g06430(.A1(new_n9232_), .A2(new_n2450_), .A3(new_n9231_), .A4(new_n2457_), .ZN(new_n9233_));
  NOR2_X1    g06431(.A1(new_n9020_), .A2(new_n8274_), .ZN(new_n9234_));
  OAI21_X1   g06432(.A1(new_n9233_), .A2(new_n9230_), .B(new_n9234_), .ZN(new_n9235_));
  AOI21_X1   g06433(.A1(new_n9235_), .A2(new_n9229_), .B(new_n2569_), .ZN(po0227));
  NOR2_X1    g06434(.A1(new_n2702_), .A2(new_n2707_), .ZN(new_n9237_));
  INV_X1     g06435(.I(new_n9237_), .ZN(new_n9238_));
  NOR3_X1    g06436(.A1(new_n2853_), .A2(new_n2755_), .A3(new_n9238_), .ZN(new_n9239_));
  NAND3_X1   g06437(.A1(new_n9239_), .A2(new_n8294_), .A3(new_n8346_), .ZN(new_n9240_));
  NOR2_X1    g06438(.A1(new_n4822_), .A2(new_n5293_), .ZN(new_n9241_));
  NAND2_X1   g06439(.A1(new_n5461_), .A2(new_n9241_), .ZN(new_n9242_));
  INV_X1     g06440(.I(pi0589), .ZN(new_n9243_));
  NOR2_X1    g06441(.A1(new_n3072_), .A2(new_n9243_), .ZN(new_n9244_));
  NAND3_X1   g06442(.A1(new_n5400_), .A2(new_n3383_), .A3(new_n9244_), .ZN(new_n9245_));
  NOR2_X1    g06443(.A1(pi0210), .A2(pi0589), .ZN(new_n9246_));
  AOI21_X1   g06444(.A1(new_n9245_), .A2(new_n9246_), .B(new_n9242_), .ZN(new_n9247_));
  NAND3_X1   g06445(.A1(new_n5407_), .A2(pi0593), .A3(pi0835), .ZN(new_n9248_));
  OAI22_X1   g06446(.A1(new_n5694_), .A2(new_n9248_), .B1(new_n3183_), .B2(new_n5401_), .ZN(new_n9249_));
  NAND2_X1   g06447(.A1(new_n9247_), .A2(new_n9249_), .ZN(new_n9250_));
  AOI21_X1   g06448(.A1(new_n3145_), .A2(new_n9240_), .B(new_n9250_), .ZN(po0228));
  NOR2_X1    g06449(.A1(new_n7408_), .A2(pi0050), .ZN(new_n9252_));
  INV_X1     g06450(.I(new_n9252_), .ZN(new_n9253_));
  NOR2_X1    g06451(.A1(new_n5585_), .A2(new_n9253_), .ZN(new_n9254_));
  NOR2_X1    g06452(.A1(new_n2610_), .A2(new_n2441_), .ZN(new_n9255_));
  NAND3_X1   g06453(.A1(new_n5564_), .A2(new_n9255_), .A3(new_n2445_), .ZN(new_n9256_));
  NOR2_X1    g06454(.A1(new_n9256_), .A2(new_n8959_), .ZN(new_n9257_));
  NOR2_X1    g06455(.A1(new_n9209_), .A2(new_n8555_), .ZN(new_n9258_));
  NOR2_X1    g06456(.A1(new_n8684_), .A2(pi0219), .ZN(new_n9259_));
  INV_X1     g06457(.I(new_n9259_), .ZN(new_n9260_));
  NOR2_X1    g06458(.A1(new_n9260_), .A2(new_n3098_), .ZN(new_n9261_));
  NOR2_X1    g06459(.A1(new_n9261_), .A2(new_n9258_), .ZN(new_n9262_));
  INV_X1     g06460(.I(new_n9262_), .ZN(new_n9263_));
  NOR4_X1    g06461(.A1(new_n9210_), .A2(new_n8288_), .A3(new_n8957_), .A4(new_n9263_), .ZN(new_n9264_));
  AOI21_X1   g06462(.A1(new_n9257_), .A2(new_n9264_), .B(new_n9254_), .ZN(new_n9265_));
  NAND2_X1   g06463(.A1(new_n7287_), .A2(new_n2492_), .ZN(new_n9266_));
  NOR4_X1    g06464(.A1(new_n8290_), .A2(new_n2644_), .A3(new_n9263_), .A4(new_n9231_), .ZN(new_n9267_));
  OAI21_X1   g06465(.A1(new_n9257_), .A2(new_n9266_), .B(new_n9267_), .ZN(new_n9268_));
  NOR2_X1    g06466(.A1(new_n9265_), .A2(new_n9268_), .ZN(po0229));
  NOR3_X1    g06467(.A1(new_n9224_), .A2(pi0039), .A3(new_n6545_), .ZN(new_n9270_));
  NOR3_X1    g06468(.A1(new_n9270_), .A2(new_n3100_), .A3(new_n8347_), .ZN(new_n9271_));
  NOR2_X1    g06469(.A1(new_n9222_), .A2(new_n3183_), .ZN(new_n9272_));
  OAI21_X1   g06470(.A1(new_n9271_), .A2(new_n6541_), .B(new_n9272_), .ZN(new_n9273_));
  NAND2_X1   g06471(.A1(pi0024), .A2(pi0072), .ZN(new_n9274_));
  NOR3_X1    g06472(.A1(new_n5693_), .A2(new_n6360_), .A3(new_n7422_), .ZN(new_n9275_));
  NAND4_X1   g06473(.A1(new_n9275_), .A2(new_n2557_), .A3(new_n2558_), .A4(new_n8282_), .ZN(new_n9276_));
  OAI21_X1   g06474(.A1(new_n2733_), .A2(new_n9274_), .B(new_n9276_), .ZN(new_n9277_));
  AOI21_X1   g06475(.A1(new_n9273_), .A2(new_n3138_), .B(new_n9277_), .ZN(po0230));
  INV_X1     g06476(.I(pi1050), .ZN(new_n9279_));
  OAI21_X1   g06477(.A1(new_n9222_), .A2(new_n7440_), .B(pi0299), .ZN(new_n9280_));
  NAND2_X1   g06478(.A1(new_n9224_), .A2(new_n7450_), .ZN(new_n9281_));
  NAND2_X1   g06479(.A1(new_n9281_), .A2(new_n3098_), .ZN(new_n9282_));
  NAND2_X1   g06480(.A1(new_n9280_), .A2(new_n9282_), .ZN(new_n9283_));
  NAND2_X1   g06481(.A1(new_n9283_), .A2(new_n8346_), .ZN(new_n9284_));
  NAND2_X1   g06482(.A1(new_n8346_), .A2(pi0039), .ZN(new_n9285_));
  XNOR2_X1   g06483(.A1(new_n9284_), .A2(new_n9285_), .ZN(new_n9286_));
  NAND2_X1   g06484(.A1(new_n7411_), .A2(new_n8529_), .ZN(new_n9287_));
  NOR4_X1    g06485(.A1(new_n9286_), .A2(pi0314), .A3(new_n9279_), .A4(new_n9287_), .ZN(po0231));
  NAND2_X1   g06486(.A1(new_n6424_), .A2(new_n2801_), .ZN(new_n9289_));
  NAND2_X1   g06487(.A1(new_n9289_), .A2(new_n2755_), .ZN(new_n9290_));
  INV_X1     g06488(.I(new_n9290_), .ZN(new_n9291_));
  AOI21_X1   g06489(.A1(po0840), .A2(pi0479), .B(pi0096), .ZN(new_n9292_));
  NAND3_X1   g06490(.A1(new_n6402_), .A2(new_n2755_), .A3(new_n2984_), .ZN(new_n9293_));
  NOR2_X1    g06491(.A1(new_n6400_), .A2(new_n5468_), .ZN(new_n9294_));
  NAND4_X1   g06492(.A1(new_n9293_), .A2(new_n3437_), .A3(new_n9294_), .A4(po1038), .ZN(new_n9295_));
  NOR3_X1    g06493(.A1(new_n6384_), .A2(new_n9292_), .A3(new_n9295_), .ZN(new_n9296_));
  AOI21_X1   g06494(.A1(new_n9291_), .A2(new_n9296_), .B(pi0074), .ZN(new_n9297_));
  NOR2_X1    g06495(.A1(new_n9149_), .A2(new_n9297_), .ZN(po0232));
  INV_X1     g06496(.I(new_n6428_), .ZN(new_n9299_));
  NOR4_X1    g06497(.A1(new_n9291_), .A2(new_n2728_), .A3(new_n2986_), .A4(new_n3194_), .ZN(new_n9300_));
  OAI21_X1   g06498(.A1(new_n9300_), .A2(pi0096), .B(pi1093), .ZN(new_n9301_));
  NOR2_X1    g06499(.A1(new_n7331_), .A2(new_n3235_), .ZN(new_n9302_));
  OAI21_X1   g06500(.A1(new_n8296_), .A2(new_n9302_), .B(new_n8908_), .ZN(new_n9303_));
  AOI21_X1   g06501(.A1(new_n9301_), .A2(new_n9303_), .B(new_n9299_), .ZN(po0233));
  NOR2_X1    g06502(.A1(new_n8303_), .A2(new_n7291_), .ZN(new_n9305_));
  INV_X1     g06503(.I(new_n9305_), .ZN(new_n9306_));
  AOI21_X1   g06504(.A1(new_n7302_), .A2(new_n2530_), .B(new_n8290_), .ZN(new_n9307_));
  OAI21_X1   g06505(.A1(new_n8451_), .A2(new_n7269_), .B(new_n9307_), .ZN(new_n9308_));
  INV_X1     g06506(.I(new_n9308_), .ZN(new_n9309_));
  NAND3_X1   g06507(.A1(new_n9309_), .A2(pi0252), .A3(new_n2982_), .ZN(new_n9310_));
  NAND3_X1   g06508(.A1(new_n9308_), .A2(new_n3721_), .A3(new_n2982_), .ZN(new_n9311_));
  AOI21_X1   g06509(.A1(new_n9310_), .A2(new_n9311_), .B(new_n9306_), .ZN(new_n9312_));
  NOR2_X1    g06510(.A1(new_n9309_), .A2(new_n2982_), .ZN(new_n9313_));
  NOR2_X1    g06511(.A1(new_n9312_), .A2(new_n9313_), .ZN(new_n9314_));
  INV_X1     g06512(.I(new_n9314_), .ZN(new_n9315_));
  NAND2_X1   g06513(.A1(new_n9315_), .A2(new_n2984_), .ZN(new_n9316_));
  NAND2_X1   g06514(.A1(new_n9316_), .A2(pi0137), .ZN(new_n9317_));
  NOR2_X1    g06515(.A1(new_n6427_), .A2(pi0252), .ZN(new_n9318_));
  NOR2_X1    g06516(.A1(new_n2481_), .A2(new_n3304_), .ZN(new_n9319_));
  NAND2_X1   g06517(.A1(new_n8451_), .A2(new_n9319_), .ZN(new_n9320_));
  INV_X1     g06518(.I(new_n9320_), .ZN(new_n9321_));
  NAND3_X1   g06519(.A1(new_n9309_), .A2(new_n9321_), .A3(new_n2982_), .ZN(new_n9322_));
  XOR2_X1    g06520(.A1(new_n9322_), .A2(new_n9318_), .Z(new_n9323_));
  NAND2_X1   g06521(.A1(new_n9323_), .A2(pi0122), .ZN(new_n9324_));
  NAND2_X1   g06522(.A1(new_n9314_), .A2(new_n6472_), .ZN(new_n9325_));
  XNOR2_X1   g06523(.A1(new_n9324_), .A2(new_n9325_), .ZN(new_n9326_));
  NOR3_X1    g06524(.A1(new_n9326_), .A2(new_n2776_), .A3(new_n9323_), .ZN(new_n9327_));
  XOR2_X1    g06525(.A1(new_n9327_), .A2(new_n9317_), .Z(new_n9328_));
  INV_X1     g06526(.I(new_n9328_), .ZN(new_n9329_));
  NAND2_X1   g06527(.A1(new_n9323_), .A2(pi1093), .ZN(new_n9330_));
  NAND3_X1   g06528(.A1(new_n9309_), .A2(pi0137), .A3(pi1093), .ZN(new_n9331_));
  XOR2_X1    g06529(.A1(new_n9330_), .A2(new_n9331_), .Z(new_n9332_));
  OAI21_X1   g06530(.A1(new_n2776_), .A2(new_n9316_), .B(new_n9332_), .ZN(new_n9333_));
  NAND2_X1   g06531(.A1(new_n9333_), .A2(new_n2730_), .ZN(new_n9334_));
  OAI21_X1   g06532(.A1(new_n9329_), .A2(new_n2730_), .B(new_n9334_), .ZN(new_n9335_));
  NAND2_X1   g06533(.A1(new_n9326_), .A2(new_n2729_), .ZN(new_n9336_));
  NOR2_X1    g06534(.A1(new_n9316_), .A2(new_n2730_), .ZN(new_n9337_));
  XNOR2_X1   g06535(.A1(new_n9336_), .A2(new_n9337_), .ZN(new_n9338_));
  NAND3_X1   g06536(.A1(new_n9338_), .A2(pi1093), .A3(new_n9308_), .ZN(new_n9339_));
  INV_X1     g06537(.I(new_n9339_), .ZN(new_n9340_));
  NOR2_X1    g06538(.A1(new_n9340_), .A2(new_n3072_), .ZN(new_n9341_));
  AOI21_X1   g06539(.A1(new_n3072_), .A2(new_n9335_), .B(new_n9341_), .ZN(new_n9342_));
  NOR2_X1    g06540(.A1(new_n3080_), .A2(new_n5386_), .ZN(new_n9343_));
  NAND2_X1   g06541(.A1(new_n9343_), .A2(pi0299), .ZN(new_n9344_));
  NOR2_X1    g06542(.A1(new_n7293_), .A2(new_n2729_), .ZN(new_n9345_));
  AOI21_X1   g06543(.A1(new_n5526_), .A2(new_n9345_), .B(new_n2776_), .ZN(new_n9346_));
  NAND2_X1   g06544(.A1(new_n9333_), .A2(new_n9346_), .ZN(new_n9347_));
  NAND2_X1   g06545(.A1(po1057), .A2(pi0137), .ZN(new_n9348_));
  XOR2_X1    g06546(.A1(new_n9347_), .A2(new_n9348_), .Z(new_n9349_));
  AOI21_X1   g06547(.A1(po1057), .A2(new_n2729_), .B(new_n9305_), .ZN(new_n9350_));
  NOR2_X1    g06548(.A1(new_n6404_), .A2(new_n2776_), .ZN(new_n9351_));
  NOR4_X1    g06549(.A1(new_n9350_), .A2(new_n6427_), .A3(new_n9306_), .A4(new_n9351_), .ZN(new_n9352_));
  NAND2_X1   g06550(.A1(new_n9349_), .A2(new_n9352_), .ZN(new_n9353_));
  NAND2_X1   g06551(.A1(new_n9353_), .A2(new_n5526_), .ZN(new_n9354_));
  NAND2_X1   g06552(.A1(new_n9354_), .A2(new_n9329_), .ZN(new_n9355_));
  NOR2_X1    g06553(.A1(new_n9355_), .A2(pi0198), .ZN(new_n9356_));
  AOI21_X1   g06554(.A1(new_n2729_), .A2(new_n6486_), .B(new_n5526_), .ZN(new_n9357_));
  NOR2_X1    g06555(.A1(new_n9306_), .A2(new_n5526_), .ZN(new_n9358_));
  INV_X1     g06556(.I(new_n9358_), .ZN(new_n9359_));
  NOR2_X1    g06557(.A1(new_n9339_), .A2(new_n9359_), .ZN(new_n9360_));
  XOR2_X1    g06558(.A1(new_n9360_), .A2(new_n9357_), .Z(new_n9361_));
  AOI21_X1   g06559(.A1(new_n9361_), .A2(pi0198), .B(new_n9356_), .ZN(new_n9362_));
  NAND2_X1   g06560(.A1(new_n9362_), .A2(new_n9343_), .ZN(new_n9363_));
  XNOR2_X1   g06561(.A1(new_n9363_), .A2(new_n9344_), .ZN(new_n9364_));
  NOR2_X1    g06562(.A1(new_n8443_), .A2(new_n2786_), .ZN(new_n9365_));
  INV_X1     g06563(.I(new_n9365_), .ZN(new_n9366_));
  NOR2_X1    g06564(.A1(new_n9335_), .A2(new_n9366_), .ZN(new_n9367_));
  NOR2_X1    g06565(.A1(new_n9366_), .A2(new_n2777_), .ZN(new_n9368_));
  XOR2_X1    g06566(.A1(new_n9367_), .A2(new_n9368_), .Z(new_n9369_));
  AOI21_X1   g06567(.A1(new_n9369_), .A2(new_n9340_), .B(pi0299), .ZN(new_n9370_));
  OAI21_X1   g06568(.A1(new_n9364_), .A2(new_n9342_), .B(new_n9370_), .ZN(new_n9371_));
  NOR2_X1    g06569(.A1(new_n9355_), .A2(pi0210), .ZN(new_n9372_));
  AOI21_X1   g06570(.A1(new_n9361_), .A2(pi0210), .B(new_n9372_), .ZN(new_n9373_));
  NAND2_X1   g06571(.A1(new_n9373_), .A2(pi0299), .ZN(new_n9374_));
  XOR2_X1    g06572(.A1(new_n9374_), .A2(new_n5912_), .Z(new_n9375_));
  OR2_X2     g06573(.A1(new_n9375_), .A2(new_n9362_), .Z(new_n9376_));
  NAND4_X1   g06574(.A1(new_n9373_), .A2(pi0232), .A3(new_n8384_), .A4(new_n9366_), .ZN(new_n9377_));
  AOI21_X1   g06575(.A1(new_n9376_), .A2(new_n6939_), .B(new_n9377_), .ZN(new_n9378_));
  AOI21_X1   g06576(.A1(new_n9378_), .A2(new_n9371_), .B(new_n6668_), .ZN(new_n9379_));
  NOR3_X1    g06577(.A1(new_n3721_), .A2(new_n2979_), .A3(pi1093), .ZN(new_n9380_));
  NAND2_X1   g06578(.A1(new_n2776_), .A2(new_n2721_), .ZN(new_n9381_));
  OAI21_X1   g06579(.A1(pi0950), .A2(new_n9381_), .B(new_n9380_), .ZN(new_n9382_));
  NOR2_X1    g06580(.A1(new_n9314_), .A2(new_n6410_), .ZN(new_n9383_));
  XNOR2_X1   g06581(.A1(new_n9383_), .A2(new_n6472_), .ZN(new_n9384_));
  AOI21_X1   g06582(.A1(new_n6402_), .A2(new_n9313_), .B(new_n9312_), .ZN(new_n9385_));
  NOR2_X1    g06583(.A1(new_n9320_), .A2(new_n5533_), .ZN(new_n9386_));
  INV_X1     g06584(.I(new_n9386_), .ZN(new_n9387_));
  NOR2_X1    g06585(.A1(new_n9385_), .A2(new_n9387_), .ZN(new_n9388_));
  INV_X1     g06586(.I(new_n9388_), .ZN(new_n9389_));
  NOR2_X1    g06587(.A1(new_n9384_), .A2(new_n9389_), .ZN(new_n9390_));
  NOR2_X1    g06588(.A1(new_n6427_), .A2(new_n3721_), .ZN(new_n9391_));
  NOR2_X1    g06589(.A1(new_n9314_), .A2(new_n2984_), .ZN(new_n9392_));
  XNOR2_X1   g06590(.A1(new_n9392_), .A2(new_n6472_), .ZN(new_n9393_));
  NOR3_X1    g06591(.A1(new_n9393_), .A2(new_n9391_), .A3(new_n9320_), .ZN(new_n9394_));
  OAI21_X1   g06592(.A1(new_n9394_), .A2(new_n9390_), .B(new_n2729_), .ZN(new_n9395_));
  NAND2_X1   g06593(.A1(new_n9320_), .A2(pi1093), .ZN(new_n9396_));
  XOR2_X1    g06594(.A1(new_n9396_), .A2(new_n6472_), .Z(new_n9397_));
  NOR2_X1    g06595(.A1(new_n9397_), .A2(new_n9308_), .ZN(new_n9398_));
  OAI21_X1   g06596(.A1(new_n9390_), .A2(new_n9398_), .B(new_n2730_), .ZN(new_n9399_));
  NOR2_X1    g06597(.A1(new_n9320_), .A2(new_n9391_), .ZN(new_n9400_));
  NOR3_X1    g06598(.A1(new_n9400_), .A2(new_n2776_), .A3(new_n2729_), .ZN(new_n9401_));
  NAND3_X1   g06599(.A1(new_n9395_), .A2(new_n9399_), .A3(new_n9401_), .ZN(new_n9402_));
  AOI21_X1   g06600(.A1(new_n9402_), .A2(new_n9382_), .B(new_n9320_), .ZN(new_n9403_));
  NAND2_X1   g06601(.A1(new_n9403_), .A2(new_n2777_), .ZN(new_n9404_));
  NAND2_X1   g06602(.A1(new_n9395_), .A2(new_n9399_), .ZN(new_n9405_));
  OAI21_X1   g06603(.A1(new_n2777_), .A2(new_n9405_), .B(new_n9404_), .ZN(new_n9406_));
  AOI21_X1   g06604(.A1(new_n9359_), .A2(new_n6410_), .B(new_n8236_), .ZN(new_n9407_));
  AND3_X2    g06605(.A1(new_n9403_), .A2(po1057), .A3(new_n9407_), .Z(new_n9408_));
  NOR3_X1    g06606(.A1(new_n9403_), .A2(new_n5526_), .A3(new_n9407_), .ZN(new_n9409_));
  OAI21_X1   g06607(.A1(new_n9408_), .A2(new_n9409_), .B(pi0137), .ZN(new_n9410_));
  AOI21_X1   g06608(.A1(new_n9405_), .A2(new_n5526_), .B(new_n9407_), .ZN(new_n9411_));
  AOI21_X1   g06609(.A1(new_n9411_), .A2(pi0210), .B(new_n3098_), .ZN(new_n9412_));
  OAI21_X1   g06610(.A1(new_n9410_), .A2(pi0210), .B(new_n9412_), .ZN(new_n9413_));
  NAND2_X1   g06611(.A1(new_n9365_), .A2(pi0299), .ZN(new_n9414_));
  XOR2_X1    g06612(.A1(new_n9413_), .A2(new_n9414_), .Z(new_n9415_));
  XOR2_X1    g06613(.A1(new_n9413_), .A2(new_n6216_), .Z(new_n9416_));
  NAND2_X1   g06614(.A1(new_n9411_), .A2(pi0198), .ZN(new_n9417_));
  OAI21_X1   g06615(.A1(new_n9410_), .A2(pi0198), .B(new_n9417_), .ZN(new_n9418_));
  AND2_X2    g06616(.A1(new_n9418_), .A2(pi0232), .Z(new_n9419_));
  AOI22_X1   g06617(.A1(new_n9406_), .A2(new_n9415_), .B1(new_n9416_), .B2(new_n9419_), .ZN(new_n9420_));
  NOR2_X1    g06618(.A1(new_n9405_), .A2(new_n3072_), .ZN(new_n9421_));
  AOI21_X1   g06619(.A1(new_n9403_), .A2(new_n3072_), .B(new_n9421_), .ZN(new_n9422_));
  INV_X1     g06620(.I(new_n9343_), .ZN(new_n9423_));
  NOR2_X1    g06621(.A1(new_n9418_), .A2(new_n9423_), .ZN(new_n9424_));
  XOR2_X1    g06622(.A1(new_n9424_), .A2(new_n9344_), .Z(new_n9425_));
  NOR4_X1    g06623(.A1(new_n9379_), .A2(new_n9420_), .A3(new_n9422_), .A4(new_n9425_), .ZN(po0234));
  INV_X1     g06624(.I(pi0086), .ZN(new_n9427_));
  NOR3_X1    g06625(.A1(new_n2548_), .A2(new_n9427_), .A3(new_n7270_), .ZN(new_n9428_));
  INV_X1     g06626(.I(new_n9428_), .ZN(new_n9429_));
  INV_X1     g06627(.I(new_n2554_), .ZN(new_n9430_));
  NOR2_X1    g06628(.A1(new_n9430_), .A2(new_n2520_), .ZN(new_n9431_));
  NOR2_X1    g06629(.A1(new_n9431_), .A2(pi0086), .ZN(new_n9432_));
  NOR2_X1    g06630(.A1(new_n5599_), .A2(new_n9432_), .ZN(new_n9433_));
  NAND2_X1   g06631(.A1(new_n9433_), .A2(new_n8945_), .ZN(new_n9434_));
  NAND2_X1   g06632(.A1(new_n9434_), .A2(new_n8291_), .ZN(new_n9435_));
  NAND2_X1   g06633(.A1(new_n8291_), .A2(pi0314), .ZN(new_n9436_));
  XNOR2_X1   g06634(.A1(new_n9435_), .A2(new_n9436_), .ZN(new_n9437_));
  NOR2_X1    g06635(.A1(new_n9437_), .A2(new_n9429_), .ZN(po0235));
  INV_X1     g06636(.I(pi0468), .ZN(new_n9439_));
  AND3_X2    g06637(.A1(new_n9439_), .A2(pi0119), .A3(pi0232), .Z(po0236));
  OAI21_X1   g06638(.A1(new_n7470_), .A2(new_n8443_), .B(new_n2837_), .ZN(new_n9441_));
  NOR2_X1    g06639(.A1(new_n5386_), .A2(new_n4808_), .ZN(new_n9442_));
  INV_X1     g06640(.I(new_n9442_), .ZN(new_n9443_));
  OAI21_X1   g06641(.A1(new_n7473_), .A2(new_n9443_), .B(new_n2837_), .ZN(new_n9444_));
  NAND4_X1   g06642(.A1(new_n9444_), .A2(pi0040), .A3(pi0163), .A4(new_n7396_), .ZN(new_n9445_));
  NOR2_X1    g06643(.A1(new_n7386_), .A2(new_n9445_), .ZN(new_n9446_));
  AOI21_X1   g06644(.A1(new_n9441_), .A2(new_n9446_), .B(new_n5664_), .ZN(new_n9447_));
  NOR3_X1    g06645(.A1(new_n2501_), .A2(new_n2890_), .A3(new_n2774_), .ZN(new_n9448_));
  NOR2_X1    g06646(.A1(new_n9448_), .A2(pi0040), .ZN(new_n9449_));
  INV_X1     g06647(.I(new_n9449_), .ZN(new_n9450_));
  NOR2_X1    g06648(.A1(new_n7387_), .A2(new_n9450_), .ZN(new_n9451_));
  AOI21_X1   g06649(.A1(new_n9451_), .A2(new_n8442_), .B(pi0210), .ZN(new_n9452_));
  NAND3_X1   g06650(.A1(new_n7472_), .A2(new_n5657_), .A3(new_n9449_), .ZN(new_n9453_));
  AND2_X2    g06651(.A1(new_n9453_), .A2(new_n9442_), .Z(new_n9454_));
  NOR4_X1    g06652(.A1(new_n9452_), .A2(pi0153), .A3(new_n7390_), .A4(new_n9454_), .ZN(new_n9455_));
  INV_X1     g06653(.I(pi0163), .ZN(new_n9456_));
  NOR2_X1    g06654(.A1(new_n7470_), .A2(new_n9450_), .ZN(new_n9457_));
  OAI21_X1   g06655(.A1(new_n2837_), .A2(new_n9443_), .B(new_n9453_), .ZN(new_n9458_));
  NAND3_X1   g06656(.A1(new_n9458_), .A2(new_n7396_), .A3(new_n8442_), .ZN(new_n9459_));
  OAI21_X1   g06657(.A1(new_n9457_), .A2(new_n9459_), .B(new_n9456_), .ZN(new_n9460_));
  OAI21_X1   g06658(.A1(pi0040), .A2(pi0163), .B(new_n8442_), .ZN(new_n9461_));
  NOR2_X1    g06659(.A1(new_n7402_), .A2(pi0153), .ZN(new_n9462_));
  OAI21_X1   g06660(.A1(new_n7426_), .A2(new_n9461_), .B(new_n9462_), .ZN(new_n9463_));
  NAND2_X1   g06661(.A1(new_n9463_), .A2(new_n7416_), .ZN(new_n9464_));
  NOR4_X1    g06662(.A1(new_n9464_), .A2(new_n2486_), .A3(new_n5664_), .A4(new_n5386_), .ZN(new_n9465_));
  OAI21_X1   g06663(.A1(new_n9455_), .A2(new_n9460_), .B(new_n9465_), .ZN(new_n9466_));
  XNOR2_X1   g06664(.A1(new_n9466_), .A2(new_n9447_), .ZN(new_n9467_));
  NAND3_X1   g06665(.A1(new_n7374_), .A2(pi0184), .A3(pi0189), .ZN(new_n9468_));
  NAND3_X1   g06666(.A1(new_n7379_), .A2(pi0184), .A3(new_n8642_), .ZN(new_n9469_));
  AOI21_X1   g06667(.A1(new_n9469_), .A2(new_n9468_), .B(new_n7426_), .ZN(new_n9470_));
  INV_X1     g06668(.I(pi0184), .ZN(new_n9471_));
  NOR3_X1    g06669(.A1(new_n7349_), .A2(new_n9471_), .A3(new_n8642_), .ZN(new_n9472_));
  INV_X1     g06670(.I(new_n9448_), .ZN(new_n9473_));
  NOR2_X1    g06671(.A1(pi0175), .A2(pi0299), .ZN(new_n9474_));
  AOI21_X1   g06672(.A1(pi0040), .A2(new_n9474_), .B(new_n5373_), .ZN(new_n9475_));
  NOR3_X1    g06673(.A1(new_n9473_), .A2(new_n5644_), .A3(new_n9475_), .ZN(new_n9476_));
  OAI21_X1   g06674(.A1(new_n9470_), .A2(new_n9472_), .B(new_n9476_), .ZN(new_n9477_));
  NOR2_X1    g06675(.A1(pi0182), .A2(pi0184), .ZN(new_n9478_));
  NOR3_X1    g06676(.A1(new_n7397_), .A2(new_n8642_), .A3(new_n9478_), .ZN(new_n9479_));
  OAI21_X1   g06677(.A1(new_n7393_), .A2(new_n8439_), .B(new_n9479_), .ZN(new_n9480_));
  NAND2_X1   g06678(.A1(new_n9450_), .A2(new_n8644_), .ZN(new_n9481_));
  OAI21_X1   g06679(.A1(new_n7396_), .A2(new_n9481_), .B(new_n5559_), .ZN(new_n9482_));
  OR3_X2     g06680(.A1(new_n5386_), .A2(new_n2486_), .A3(new_n9478_), .Z(new_n9483_));
  AOI21_X1   g06681(.A1(new_n9482_), .A2(new_n9483_), .B(new_n8439_), .ZN(new_n9484_));
  NAND2_X1   g06682(.A1(new_n9451_), .A2(new_n9484_), .ZN(new_n9485_));
  INV_X1     g06683(.I(pi0175), .ZN(new_n9486_));
  NOR2_X1    g06684(.A1(new_n9486_), .A2(pi0299), .ZN(new_n9487_));
  INV_X1     g06685(.I(new_n9487_), .ZN(new_n9488_));
  OAI21_X1   g06686(.A1(new_n7392_), .A2(new_n9485_), .B(new_n9488_), .ZN(new_n9489_));
  NAND3_X1   g06687(.A1(new_n7413_), .A2(pi0189), .A3(new_n3142_), .ZN(new_n9490_));
  NAND3_X1   g06688(.A1(new_n7414_), .A2(new_n8642_), .A3(new_n3142_), .ZN(new_n9491_));
  NAND2_X1   g06689(.A1(new_n7416_), .A2(new_n5373_), .ZN(new_n9492_));
  AOI21_X1   g06690(.A1(new_n9491_), .A2(new_n9490_), .B(new_n9492_), .ZN(new_n9493_));
  OAI21_X1   g06691(.A1(new_n9493_), .A2(pi0182), .B(new_n9448_), .ZN(new_n9494_));
  NAND2_X1   g06692(.A1(new_n9494_), .A2(new_n9471_), .ZN(new_n9495_));
  NAND4_X1   g06693(.A1(new_n9480_), .A2(pi0040), .A3(new_n9489_), .A4(new_n9495_), .ZN(new_n9496_));
  OAI21_X1   g06694(.A1(new_n9464_), .A2(new_n3098_), .B(new_n5386_), .ZN(new_n9497_));
  NAND2_X1   g06695(.A1(new_n2486_), .A2(new_n3098_), .ZN(new_n9498_));
  NOR2_X1    g06696(.A1(new_n2501_), .A2(new_n7403_), .ZN(new_n9499_));
  INV_X1     g06697(.I(new_n7589_), .ZN(new_n9500_));
  AOI22_X1   g06698(.A1(new_n9500_), .A2(new_n5411_), .B1(pi0179), .B2(pi0189), .ZN(new_n9501_));
  NOR2_X1    g06699(.A1(new_n9498_), .A2(pi0039), .ZN(new_n9502_));
  NOR4_X1    g06700(.A1(new_n9501_), .A2(new_n5397_), .A3(new_n7451_), .A4(new_n9502_), .ZN(new_n9503_));
  AOI21_X1   g06701(.A1(new_n9503_), .A2(new_n9499_), .B(new_n9498_), .ZN(new_n9504_));
  INV_X1     g06702(.I(pi0156), .ZN(new_n9505_));
  OAI22_X1   g06703(.A1(new_n7597_), .A2(new_n7589_), .B1(new_n9505_), .B2(new_n4808_), .ZN(new_n9506_));
  NAND4_X1   g06704(.A1(new_n9506_), .A2(new_n5454_), .A3(new_n7439_), .A4(new_n9499_), .ZN(new_n9507_));
  OAI21_X1   g06705(.A1(new_n9504_), .A2(new_n9507_), .B(new_n5551_), .ZN(new_n9508_));
  NAND4_X1   g06706(.A1(new_n9497_), .A2(pi0039), .A3(new_n9448_), .A4(new_n9508_), .ZN(new_n9509_));
  AOI21_X1   g06707(.A1(new_n9496_), .A2(new_n9477_), .B(new_n9509_), .ZN(new_n9510_));
  AOI21_X1   g06708(.A1(new_n9510_), .A2(new_n9467_), .B(pi0038), .ZN(new_n9511_));
  NAND2_X1   g06709(.A1(pi0040), .A2(pi0232), .ZN(new_n9512_));
  NOR2_X1    g06710(.A1(new_n5373_), .A2(new_n8040_), .ZN(new_n9513_));
  NOR4_X1    g06711(.A1(new_n9513_), .A2(new_n8108_), .A3(new_n9456_), .A4(new_n5665_), .ZN(new_n9514_));
  INV_X1     g06712(.I(new_n9514_), .ZN(new_n9515_));
  NOR4_X1    g06713(.A1(new_n7986_), .A2(pi0149), .A3(pi0157), .A4(new_n5665_), .ZN(new_n9516_));
  OAI21_X1   g06714(.A1(new_n9515_), .A2(new_n9516_), .B(new_n5386_), .ZN(new_n9517_));
  XOR2_X1    g06715(.A1(new_n9517_), .A2(new_n9515_), .Z(new_n9518_));
  NOR2_X1    g06716(.A1(pi0140), .A2(pi0145), .ZN(new_n9519_));
  NOR3_X1    g06717(.A1(new_n8037_), .A2(new_n7971_), .A3(new_n5641_), .ZN(new_n9520_));
  NOR3_X1    g06718(.A1(new_n9520_), .A2(new_n5386_), .A3(new_n9519_), .ZN(new_n9521_));
  INV_X1     g06719(.I(new_n9521_), .ZN(new_n9522_));
  NOR2_X1    g06720(.A1(new_n9471_), .A2(pi0299), .ZN(new_n9523_));
  NOR3_X1    g06721(.A1(new_n9522_), .A2(new_n5386_), .A3(new_n9523_), .ZN(new_n9524_));
  OAI21_X1   g06722(.A1(new_n9524_), .A2(pi0232), .B(pi0299), .ZN(new_n9525_));
  NOR2_X1    g06723(.A1(new_n9518_), .A2(new_n9525_), .ZN(new_n9526_));
  NOR2_X1    g06724(.A1(new_n9526_), .A2(new_n3462_), .ZN(new_n9527_));
  INV_X1     g06725(.I(pi0187), .ZN(new_n9528_));
  NAND3_X1   g06726(.A1(new_n6493_), .A2(pi0147), .A3(pi0299), .ZN(new_n9529_));
  INV_X1     g06727(.I(pi0147), .ZN(new_n9530_));
  NAND3_X1   g06728(.A1(new_n6493_), .A2(new_n9530_), .A3(new_n3098_), .ZN(new_n9531_));
  AOI21_X1   g06729(.A1(new_n9529_), .A2(new_n9531_), .B(new_n9528_), .ZN(new_n9532_));
  OAI21_X1   g06730(.A1(new_n9532_), .A2(new_n3259_), .B(new_n3462_), .ZN(new_n9533_));
  INV_X1     g06731(.I(new_n9533_), .ZN(new_n9534_));
  NOR3_X1    g06732(.A1(new_n9527_), .A2(pi0087), .A3(new_n9534_), .ZN(new_n9535_));
  NOR2_X1    g06733(.A1(pi0038), .A2(pi0040), .ZN(new_n9536_));
  NAND2_X1   g06734(.A1(new_n3184_), .A2(new_n9536_), .ZN(new_n9537_));
  OAI22_X1   g06735(.A1(new_n9511_), .A2(new_n9512_), .B1(new_n9535_), .B2(new_n9537_), .ZN(new_n9538_));
  NOR2_X1    g06736(.A1(new_n7494_), .A2(new_n9530_), .ZN(new_n9539_));
  NOR2_X1    g06737(.A1(new_n9530_), .A2(new_n9528_), .ZN(new_n9540_));
  XOR2_X1    g06738(.A1(new_n9539_), .A2(new_n9540_), .Z(new_n9541_));
  NAND2_X1   g06739(.A1(new_n7500_), .A2(new_n9528_), .ZN(new_n9542_));
  AOI21_X1   g06740(.A1(new_n9541_), .A2(new_n7490_), .B(new_n9542_), .ZN(new_n9543_));
  NOR2_X1    g06741(.A1(new_n9543_), .A2(new_n9530_), .ZN(new_n9544_));
  INV_X1     g06742(.I(pi0179), .ZN(new_n9545_));
  NAND3_X1   g06743(.A1(new_n6493_), .A2(pi0156), .A3(pi0299), .ZN(new_n9546_));
  NAND3_X1   g06744(.A1(new_n6493_), .A2(new_n9505_), .A3(new_n3098_), .ZN(new_n9547_));
  AOI21_X1   g06745(.A1(new_n9547_), .A2(new_n9546_), .B(new_n9545_), .ZN(new_n9548_));
  NAND4_X1   g06746(.A1(new_n2750_), .A2(new_n9548_), .A3(new_n3142_), .A4(new_n3191_), .ZN(new_n9549_));
  NAND2_X1   g06747(.A1(new_n9549_), .A2(new_n9536_), .ZN(new_n9550_));
  NOR3_X1    g06748(.A1(new_n9526_), .A2(new_n3235_), .A3(new_n7529_), .ZN(new_n9551_));
  AOI21_X1   g06749(.A1(new_n9534_), .A2(new_n9550_), .B(new_n9551_), .ZN(new_n9552_));
  NOR4_X1    g06750(.A1(new_n9552_), .A2(new_n3115_), .A3(new_n3462_), .A4(new_n9526_), .ZN(new_n9553_));
  OAI21_X1   g06751(.A1(new_n9553_), .A2(new_n3188_), .B(pi0038), .ZN(new_n9554_));
  NOR2_X1    g06752(.A1(new_n9544_), .A2(new_n9554_), .ZN(new_n9555_));
  INV_X1     g06753(.I(new_n9526_), .ZN(new_n9556_));
  AOI21_X1   g06754(.A1(new_n9556_), .A2(new_n6328_), .B(new_n7538_), .ZN(new_n9557_));
  AOI22_X1   g06755(.A1(new_n9538_), .A2(new_n9555_), .B1(pi0074), .B2(new_n9557_), .ZN(new_n9558_));
  NOR2_X1    g06756(.A1(new_n9526_), .A2(new_n3115_), .ZN(new_n9559_));
  NAND2_X1   g06757(.A1(new_n7537_), .A2(pi0054), .ZN(new_n9560_));
  XNOR2_X1   g06758(.A1(new_n9559_), .A2(new_n9560_), .ZN(new_n9561_));
  AND2_X2    g06759(.A1(new_n9561_), .A2(new_n9532_), .Z(new_n9562_));
  NOR2_X1    g06760(.A1(new_n9518_), .A2(new_n5551_), .ZN(new_n9563_));
  INV_X1     g06761(.I(new_n9563_), .ZN(new_n9564_));
  OAI21_X1   g06762(.A1(new_n9564_), .A2(new_n7537_), .B(pi0074), .ZN(new_n9565_));
  NAND3_X1   g06763(.A1(new_n9564_), .A2(new_n9530_), .A3(new_n7538_), .ZN(new_n9566_));
  NAND2_X1   g06764(.A1(new_n9566_), .A2(new_n6493_), .ZN(new_n9567_));
  INV_X1     g06765(.I(new_n9567_), .ZN(new_n9568_));
  NOR2_X1    g06766(.A1(new_n3115_), .A2(new_n3175_), .ZN(new_n9569_));
  NAND4_X1   g06767(.A1(new_n3191_), .A2(pi0092), .A3(pi0163), .A4(pi0232), .ZN(new_n9570_));
  NOR3_X1    g06768(.A1(new_n2501_), .A2(new_n7403_), .A3(new_n9570_), .ZN(new_n9571_));
  AOI21_X1   g06769(.A1(new_n9530_), .A2(new_n5486_), .B(new_n6494_), .ZN(new_n9572_));
  INV_X1     g06770(.I(new_n9572_), .ZN(new_n9573_));
  NAND4_X1   g06771(.A1(new_n9564_), .A2(new_n3235_), .A3(pi0100), .A4(new_n9573_), .ZN(new_n9574_));
  NAND2_X1   g06772(.A1(new_n9574_), .A2(new_n9536_), .ZN(new_n9575_));
  OAI21_X1   g06773(.A1(new_n9575_), .A2(new_n9571_), .B(pi0054), .ZN(new_n9576_));
  XNOR2_X1   g06774(.A1(new_n9576_), .A2(new_n9569_), .ZN(new_n9577_));
  NAND2_X1   g06775(.A1(new_n9577_), .A2(new_n9568_), .ZN(new_n9578_));
  AOI21_X1   g06776(.A1(new_n9578_), .A2(new_n5975_), .B(new_n9565_), .ZN(new_n9579_));
  OAI22_X1   g06777(.A1(new_n9568_), .A2(new_n3115_), .B1(new_n3175_), .B2(new_n9565_), .ZN(new_n9580_));
  OAI22_X1   g06778(.A1(new_n9563_), .A2(new_n3462_), .B1(new_n9536_), .B2(new_n9573_), .ZN(new_n9581_));
  NAND2_X1   g06779(.A1(new_n9581_), .A2(pi0075), .ZN(new_n9582_));
  XOR2_X1    g06780(.A1(new_n9582_), .A2(new_n7928_), .Z(new_n9583_));
  NOR2_X1    g06781(.A1(new_n9583_), .A2(new_n9564_), .ZN(new_n9584_));
  AOI21_X1   g06782(.A1(new_n9584_), .A2(new_n9580_), .B(new_n3225_), .ZN(new_n9585_));
  NAND3_X1   g06783(.A1(new_n9568_), .A2(new_n3426_), .A3(new_n9565_), .ZN(new_n9586_));
  NOR3_X1    g06784(.A1(new_n9585_), .A2(new_n3426_), .A3(new_n9586_), .ZN(new_n9587_));
  OAI21_X1   g06785(.A1(new_n9579_), .A2(new_n9587_), .B(new_n9562_), .ZN(new_n9588_));
  OR2_X2     g06786(.A1(new_n9558_), .A2(new_n9588_), .Z(new_n9589_));
  INV_X1     g06787(.I(new_n7695_), .ZN(new_n9590_));
  NOR2_X1    g06788(.A1(new_n5398_), .A2(new_n8642_), .ZN(new_n9591_));
  AOI21_X1   g06789(.A1(new_n2486_), .A2(new_n5373_), .B(new_n2539_), .ZN(new_n9592_));
  NOR2_X1    g06790(.A1(new_n7591_), .A2(new_n9592_), .ZN(new_n9593_));
  NOR2_X1    g06791(.A1(new_n7599_), .A2(pi0040), .ZN(new_n9594_));
  NAND3_X1   g06792(.A1(new_n9594_), .A2(pi0189), .A3(new_n9593_), .ZN(new_n9595_));
  OAI21_X1   g06793(.A1(new_n9595_), .A2(new_n9591_), .B(pi0179), .ZN(new_n9596_));
  AOI21_X1   g06794(.A1(new_n9591_), .A2(new_n9595_), .B(new_n9596_), .ZN(new_n9597_));
  NOR2_X1    g06795(.A1(new_n2448_), .A2(new_n2486_), .ZN(new_n9598_));
  OAI21_X1   g06796(.A1(new_n7598_), .A2(new_n9598_), .B(new_n5434_), .ZN(new_n9599_));
  NOR2_X1    g06797(.A1(new_n7633_), .A2(new_n9592_), .ZN(new_n9600_));
  NOR3_X1    g06798(.A1(new_n9600_), .A2(pi0179), .A3(new_n5398_), .ZN(new_n9601_));
  NAND3_X1   g06799(.A1(new_n5397_), .A2(new_n9545_), .A3(pi0189), .ZN(new_n9602_));
  XOR2_X1    g06800(.A1(new_n9601_), .A2(new_n9602_), .Z(new_n9603_));
  OAI22_X1   g06801(.A1(new_n9603_), .A2(new_n9599_), .B1(new_n5397_), .B2(new_n9594_), .ZN(new_n9604_));
  OAI21_X1   g06802(.A1(new_n9604_), .A2(new_n9597_), .B(new_n7450_), .ZN(new_n9605_));
  NOR2_X1    g06803(.A1(new_n7451_), .A2(new_n3098_), .ZN(new_n9606_));
  XOR2_X1    g06804(.A1(new_n9605_), .A2(new_n9606_), .Z(new_n9607_));
  NOR2_X1    g06805(.A1(new_n9607_), .A2(new_n9590_), .ZN(new_n9608_));
  INV_X1     g06806(.I(new_n9594_), .ZN(new_n9609_));
  NOR2_X1    g06807(.A1(new_n9593_), .A2(new_n7440_), .ZN(new_n9610_));
  NAND3_X1   g06808(.A1(new_n5455_), .A2(pi0166), .A3(new_n7439_), .ZN(new_n9611_));
  XOR2_X1    g06809(.A1(new_n9610_), .A2(new_n9611_), .Z(new_n9612_));
  OAI21_X1   g06810(.A1(new_n9612_), .A2(new_n9609_), .B(new_n3098_), .ZN(new_n9613_));
  NAND2_X1   g06811(.A1(new_n9599_), .A2(new_n5455_), .ZN(new_n9614_));
  OAI21_X1   g06812(.A1(new_n9609_), .A2(new_n5455_), .B(new_n9614_), .ZN(new_n9615_));
  NOR2_X1    g06813(.A1(pi0156), .A2(pi0232), .ZN(new_n9616_));
  NOR4_X1    g06814(.A1(new_n7440_), .A2(new_n3183_), .A3(new_n9590_), .A4(new_n9616_), .ZN(new_n9617_));
  NAND4_X1   g06815(.A1(new_n9613_), .A2(new_n7605_), .A3(new_n9615_), .A4(new_n9617_), .ZN(new_n9618_));
  NOR2_X1    g06816(.A1(new_n9600_), .A2(new_n7440_), .ZN(new_n9619_));
  NOR3_X1    g06817(.A1(new_n5454_), .A2(new_n7440_), .A3(pi0166), .ZN(new_n9620_));
  XOR2_X1    g06818(.A1(new_n9619_), .A2(new_n9620_), .Z(new_n9621_));
  AOI21_X1   g06819(.A1(new_n9621_), .A2(new_n9615_), .B(pi0299), .ZN(new_n9622_));
  AOI21_X1   g06820(.A1(new_n9599_), .A2(new_n5397_), .B(new_n7451_), .ZN(new_n9623_));
  OAI21_X1   g06821(.A1(new_n9609_), .A2(new_n5397_), .B(new_n9623_), .ZN(new_n9624_));
  XNOR2_X1   g06822(.A1(new_n9624_), .A2(new_n9606_), .ZN(new_n9625_));
  AOI21_X1   g06823(.A1(new_n9625_), .A2(new_n7695_), .B(pi0232), .ZN(new_n9626_));
  NOR3_X1    g06824(.A1(new_n9626_), .A2(new_n9618_), .A3(new_n9622_), .ZN(new_n9627_));
  AOI21_X1   g06825(.A1(new_n9608_), .A2(new_n9627_), .B(new_n3259_), .ZN(new_n9628_));
  AOI21_X1   g06826(.A1(new_n7803_), .A2(new_n2486_), .B(pi0095), .ZN(new_n9629_));
  NAND3_X1   g06827(.A1(new_n7817_), .A2(new_n2486_), .A3(pi0166), .ZN(new_n9630_));
  NAND2_X1   g06828(.A1(new_n9630_), .A2(new_n9629_), .ZN(new_n9631_));
  AOI21_X1   g06829(.A1(new_n7665_), .A2(new_n7706_), .B(new_n7662_), .ZN(new_n9632_));
  INV_X1     g06830(.I(new_n9632_), .ZN(new_n9633_));
  AOI21_X1   g06831(.A1(new_n7682_), .A2(new_n2486_), .B(pi0095), .ZN(new_n9634_));
  NAND2_X1   g06832(.A1(new_n9634_), .A2(pi0153), .ZN(new_n9635_));
  NAND2_X1   g06833(.A1(new_n9635_), .A2(new_n9287_), .ZN(new_n9636_));
  NOR2_X1    g06834(.A1(new_n5664_), .A2(new_n9456_), .ZN(new_n9637_));
  NAND4_X1   g06835(.A1(new_n9633_), .A2(new_n9442_), .A3(new_n9636_), .A4(new_n9637_), .ZN(new_n9638_));
  AOI21_X1   g06836(.A1(new_n9631_), .A2(new_n9638_), .B(new_n2837_), .ZN(new_n9639_));
  NOR2_X1    g06837(.A1(new_n7735_), .A2(new_n9443_), .ZN(new_n9640_));
  AOI21_X1   g06838(.A1(new_n9634_), .A2(new_n9640_), .B(pi0153), .ZN(new_n9641_));
  NAND2_X1   g06839(.A1(new_n8442_), .A2(new_n7695_), .ZN(new_n9642_));
  OAI21_X1   g06840(.A1(new_n9641_), .A2(new_n9642_), .B(new_n5664_), .ZN(new_n9643_));
  NOR2_X1    g06841(.A1(new_n5373_), .A2(pi0153), .ZN(new_n9644_));
  AOI21_X1   g06842(.A1(new_n9631_), .A2(new_n9644_), .B(new_n7735_), .ZN(new_n9645_));
  OAI21_X1   g06843(.A1(new_n9639_), .A2(new_n9643_), .B(new_n9645_), .ZN(new_n9646_));
  NOR2_X1    g06844(.A1(new_n7896_), .A2(pi0040), .ZN(new_n9647_));
  NOR2_X1    g06845(.A1(new_n9647_), .A2(pi0095), .ZN(new_n9648_));
  NOR2_X1    g06846(.A1(new_n9648_), .A2(new_n9633_), .ZN(new_n9649_));
  NOR2_X1    g06847(.A1(new_n7696_), .A2(pi0095), .ZN(new_n9650_));
  NOR2_X1    g06848(.A1(new_n9590_), .A2(new_n2436_), .ZN(new_n9651_));
  NOR2_X1    g06849(.A1(new_n9650_), .A2(new_n9651_), .ZN(new_n9652_));
  NOR2_X1    g06850(.A1(new_n7707_), .A2(new_n8644_), .ZN(new_n9653_));
  NAND2_X1   g06851(.A1(new_n8643_), .A2(pi0198), .ZN(new_n9654_));
  XOR2_X1    g06852(.A1(new_n9653_), .A2(new_n9654_), .Z(new_n9655_));
  OAI21_X1   g06853(.A1(new_n9655_), .A2(new_n9652_), .B(pi0182), .ZN(new_n9656_));
  NAND2_X1   g06854(.A1(new_n7696_), .A2(new_n2436_), .ZN(new_n9657_));
  NAND2_X1   g06855(.A1(new_n9657_), .A2(new_n9632_), .ZN(new_n9658_));
  NAND2_X1   g06856(.A1(new_n9658_), .A2(new_n8643_), .ZN(new_n9659_));
  XNOR2_X1   g06857(.A1(new_n9659_), .A2(new_n9654_), .ZN(new_n9660_));
  OAI21_X1   g06858(.A1(new_n7693_), .A2(new_n7704_), .B(new_n9632_), .ZN(new_n9661_));
  NAND2_X1   g06859(.A1(new_n8438_), .A2(pi0182), .ZN(new_n9662_));
  NOR4_X1    g06860(.A1(new_n9660_), .A2(new_n7740_), .A3(new_n9661_), .A4(new_n9662_), .ZN(new_n9663_));
  NOR2_X1    g06861(.A1(new_n9663_), .A2(new_n9656_), .ZN(new_n9664_));
  NAND2_X1   g06862(.A1(new_n9663_), .A2(new_n9656_), .ZN(new_n9665_));
  NAND3_X1   g06863(.A1(new_n9665_), .A2(new_n8439_), .A3(new_n9632_), .ZN(new_n9666_));
  NAND2_X1   g06864(.A1(new_n5373_), .A2(pi0184), .ZN(new_n9667_));
  NOR2_X1    g06865(.A1(new_n9632_), .A2(pi0182), .ZN(new_n9668_));
  AND3_X2    g06866(.A1(new_n7682_), .A2(new_n2486_), .A3(pi0182), .Z(new_n9669_));
  NOR3_X1    g06867(.A1(new_n2436_), .A2(pi0063), .A3(pi0107), .ZN(new_n9670_));
  NOR4_X1    g06868(.A1(new_n9668_), .A2(new_n9669_), .A3(new_n9670_), .A4(new_n9667_), .ZN(new_n9671_));
  NOR2_X1    g06869(.A1(new_n9671_), .A2(new_n9487_), .ZN(new_n9672_));
  NOR2_X1    g06870(.A1(new_n2436_), .A2(pi0182), .ZN(new_n9673_));
  NOR4_X1    g06871(.A1(new_n7741_), .A2(new_n9667_), .A3(new_n9672_), .A4(new_n9673_), .ZN(new_n9674_));
  OAI21_X1   g06872(.A1(new_n9666_), .A2(new_n9664_), .B(new_n9674_), .ZN(new_n9675_));
  NAND2_X1   g06873(.A1(new_n9647_), .A2(new_n8643_), .ZN(new_n9676_));
  OAI21_X1   g06874(.A1(new_n7845_), .A2(pi0040), .B(new_n2794_), .ZN(new_n9677_));
  OAI21_X1   g06875(.A1(new_n9677_), .A2(new_n2436_), .B(new_n2794_), .ZN(new_n9678_));
  AOI21_X1   g06876(.A1(new_n9678_), .A2(new_n7695_), .B(new_n7706_), .ZN(new_n9679_));
  NAND2_X1   g06877(.A1(new_n8438_), .A2(pi0198), .ZN(new_n9680_));
  NAND2_X1   g06878(.A1(new_n9677_), .A2(new_n7702_), .ZN(new_n9681_));
  NAND2_X1   g06879(.A1(new_n9681_), .A2(new_n2436_), .ZN(new_n9682_));
  NAND2_X1   g06880(.A1(new_n9682_), .A2(new_n7735_), .ZN(new_n9683_));
  NAND2_X1   g06881(.A1(new_n9683_), .A2(new_n8438_), .ZN(new_n9684_));
  XOR2_X1    g06882(.A1(new_n9684_), .A2(new_n9680_), .Z(new_n9685_));
  NAND3_X1   g06883(.A1(new_n9474_), .A2(pi0182), .A3(new_n9471_), .ZN(new_n9686_));
  AOI21_X1   g06884(.A1(new_n9685_), .A2(new_n9679_), .B(new_n9686_), .ZN(new_n9687_));
  AOI21_X1   g06885(.A1(new_n9676_), .A2(new_n9687_), .B(pi0184), .ZN(new_n9688_));
  INV_X1     g06886(.I(new_n9629_), .ZN(new_n9689_));
  NAND2_X1   g06887(.A1(new_n5373_), .A2(pi0182), .ZN(new_n9690_));
  AOI21_X1   g06888(.A1(new_n9632_), .A2(new_n5373_), .B(new_n9690_), .ZN(new_n9691_));
  NOR3_X1    g06889(.A1(new_n9633_), .A2(pi0182), .A3(new_n5386_), .ZN(new_n9692_));
  OAI21_X1   g06890(.A1(new_n9692_), .A2(new_n9691_), .B(new_n7706_), .ZN(new_n9693_));
  OAI21_X1   g06891(.A1(new_n9689_), .A2(new_n9693_), .B(new_n8642_), .ZN(new_n9694_));
  NAND4_X1   g06892(.A1(new_n9649_), .A2(new_n2486_), .A3(new_n7817_), .A4(new_n9694_), .ZN(new_n9695_));
  OAI21_X1   g06893(.A1(new_n9695_), .A2(new_n9688_), .B(new_n9675_), .ZN(new_n9696_));
  NAND2_X1   g06894(.A1(new_n9678_), .A2(new_n7695_), .ZN(new_n9697_));
  NAND2_X1   g06895(.A1(new_n9697_), .A2(new_n9632_), .ZN(new_n9698_));
  NAND2_X1   g06896(.A1(new_n9698_), .A2(new_n8438_), .ZN(new_n9699_));
  XNOR2_X1   g06897(.A1(new_n9699_), .A2(new_n9680_), .ZN(new_n9700_));
  AOI21_X1   g06898(.A1(new_n9681_), .A2(new_n2436_), .B(new_n9633_), .ZN(new_n9701_));
  NAND4_X1   g06899(.A1(new_n9701_), .A2(pi0182), .A3(pi0184), .A4(new_n9474_), .ZN(new_n9702_));
  NOR2_X1    g06900(.A1(new_n9700_), .A2(new_n9702_), .ZN(new_n9703_));
  AOI21_X1   g06901(.A1(new_n9696_), .A2(new_n9703_), .B(new_n9649_), .ZN(new_n9704_));
  NAND2_X1   g06902(.A1(new_n7875_), .A2(new_n2486_), .ZN(new_n9705_));
  AOI21_X1   g06903(.A1(new_n9705_), .A2(new_n2436_), .B(new_n9633_), .ZN(new_n9706_));
  NAND3_X1   g06904(.A1(new_n5373_), .A2(new_n8642_), .A3(pi0299), .ZN(new_n9707_));
  OAI21_X1   g06905(.A1(new_n9704_), .A2(new_n9707_), .B(new_n9646_), .ZN(new_n9708_));
  NOR2_X1    g06906(.A1(new_n9706_), .A2(new_n3098_), .ZN(new_n9709_));
  XOR2_X1    g06907(.A1(new_n9709_), .A2(new_n5912_), .Z(new_n9710_));
  NAND2_X1   g06908(.A1(new_n9710_), .A2(new_n9649_), .ZN(new_n9711_));
  NAND2_X1   g06909(.A1(new_n9683_), .A2(new_n8442_), .ZN(new_n9712_));
  NAND2_X1   g06910(.A1(new_n8442_), .A2(pi0210), .ZN(new_n9713_));
  XOR2_X1    g06911(.A1(new_n9712_), .A2(new_n9713_), .Z(new_n9714_));
  NAND2_X1   g06912(.A1(new_n9714_), .A2(new_n9679_), .ZN(new_n9715_));
  INV_X1     g06913(.I(new_n9652_), .ZN(new_n9716_));
  NOR2_X1    g06914(.A1(new_n7707_), .A2(new_n9443_), .ZN(new_n9717_));
  NAND2_X1   g06915(.A1(new_n9442_), .A2(pi0210), .ZN(new_n9718_));
  XNOR2_X1   g06916(.A1(new_n9717_), .A2(new_n9718_), .ZN(new_n9719_));
  NAND2_X1   g06917(.A1(new_n2837_), .A2(new_n5664_), .ZN(new_n9720_));
  AOI21_X1   g06918(.A1(new_n9719_), .A2(new_n9716_), .B(new_n9720_), .ZN(new_n9721_));
  NAND2_X1   g06919(.A1(new_n7738_), .A2(new_n8442_), .ZN(new_n9722_));
  XNOR2_X1   g06920(.A1(new_n9722_), .A2(new_n9713_), .ZN(new_n9723_));
  NOR4_X1    g06921(.A1(new_n9721_), .A2(pi0153), .A3(new_n7733_), .A4(new_n9723_), .ZN(new_n9724_));
  AOI21_X1   g06922(.A1(new_n9715_), .A2(new_n9724_), .B(new_n9442_), .ZN(new_n9725_));
  OAI21_X1   g06923(.A1(new_n9705_), .A2(new_n9725_), .B(new_n9456_), .ZN(new_n9726_));
  NAND2_X1   g06924(.A1(new_n9698_), .A2(new_n8442_), .ZN(new_n9727_));
  XOR2_X1    g06925(.A1(new_n9727_), .A2(new_n9713_), .Z(new_n9728_));
  AOI21_X1   g06926(.A1(new_n9728_), .A2(new_n9701_), .B(pi0153), .ZN(new_n9729_));
  NAND2_X1   g06927(.A1(new_n9658_), .A2(new_n9442_), .ZN(new_n9730_));
  XNOR2_X1   g06928(.A1(new_n9730_), .A2(new_n9718_), .ZN(new_n9731_));
  NOR2_X1    g06929(.A1(new_n9731_), .A2(new_n9661_), .ZN(new_n9732_));
  NAND2_X1   g06930(.A1(new_n7737_), .A2(new_n9713_), .ZN(new_n9733_));
  NAND3_X1   g06931(.A1(new_n9733_), .A2(pi0210), .A3(new_n9633_), .ZN(new_n9734_));
  NOR2_X1    g06932(.A1(new_n3259_), .A2(new_n4808_), .ZN(new_n9735_));
  NAND4_X1   g06933(.A1(new_n7731_), .A2(pi0232), .A3(new_n9544_), .A4(new_n9735_), .ZN(new_n9736_));
  AOI21_X1   g06934(.A1(new_n9734_), .A2(new_n9632_), .B(new_n9736_), .ZN(new_n9737_));
  OAI21_X1   g06935(.A1(new_n9732_), .A2(new_n9720_), .B(new_n9737_), .ZN(new_n9738_));
  NOR2_X1    g06936(.A1(new_n9738_), .A2(new_n9729_), .ZN(new_n9739_));
  NAND3_X1   g06937(.A1(new_n9726_), .A2(new_n9739_), .A3(new_n9706_), .ZN(new_n9740_));
  AOI21_X1   g06938(.A1(new_n9711_), .A2(new_n3183_), .B(new_n9740_), .ZN(new_n9741_));
  NAND2_X1   g06939(.A1(new_n9741_), .A2(new_n9708_), .ZN(new_n9742_));
  XOR2_X1    g06940(.A1(new_n9742_), .A2(new_n9628_), .Z(new_n9743_));
  NOR2_X1    g06941(.A1(new_n9563_), .A2(new_n3462_), .ZN(new_n9744_));
  OAI21_X1   g06942(.A1(new_n7695_), .A2(new_n3183_), .B(new_n7523_), .ZN(new_n9745_));
  AOI21_X1   g06943(.A1(new_n7587_), .A2(new_n5386_), .B(new_n7577_), .ZN(new_n9746_));
  AOI21_X1   g06944(.A1(new_n7588_), .A2(new_n2539_), .B(pi0040), .ZN(new_n9747_));
  NAND2_X1   g06945(.A1(new_n9456_), .A2(new_n5551_), .ZN(new_n9748_));
  OAI21_X1   g06946(.A1(new_n9747_), .A2(new_n9748_), .B(new_n9746_), .ZN(new_n9749_));
  AOI21_X1   g06947(.A1(new_n9749_), .A2(new_n3183_), .B(new_n9745_), .ZN(new_n9750_));
  NAND3_X1   g06948(.A1(new_n2448_), .A2(pi0087), .A3(new_n9536_), .ZN(new_n9751_));
  NAND2_X1   g06949(.A1(new_n9572_), .A2(new_n9751_), .ZN(new_n9752_));
  OAI21_X1   g06950(.A1(new_n9581_), .A2(new_n7938_), .B(pi0075), .ZN(new_n9753_));
  NOR2_X1    g06951(.A1(new_n9564_), .A2(new_n3483_), .ZN(new_n9754_));
  XOR2_X1    g06952(.A1(new_n9753_), .A2(new_n9754_), .Z(new_n9755_));
  OAI22_X1   g06953(.A1(new_n9750_), .A2(new_n9752_), .B1(new_n3189_), .B2(new_n9755_), .ZN(new_n9756_));
  AOI21_X1   g06954(.A1(new_n9756_), .A2(new_n9744_), .B(new_n3115_), .ZN(new_n9757_));
  XNOR2_X1   g06955(.A1(new_n9757_), .A2(new_n9569_), .ZN(new_n9758_));
  OAI21_X1   g06956(.A1(new_n9758_), .A2(new_n9567_), .B(new_n5975_), .ZN(new_n9759_));
  INV_X1     g06957(.I(new_n9557_), .ZN(new_n9760_));
  NOR2_X1    g06958(.A1(new_n9760_), .A2(new_n9565_), .ZN(new_n9761_));
  AOI21_X1   g06959(.A1(new_n9759_), .A2(new_n9761_), .B(pi0074), .ZN(new_n9762_));
  NOR2_X1    g06960(.A1(new_n9585_), .A2(new_n3426_), .ZN(new_n9763_));
  NAND2_X1   g06961(.A1(new_n9586_), .A2(new_n7944_), .ZN(new_n9764_));
  NAND2_X1   g06962(.A1(new_n9534_), .A2(new_n9751_), .ZN(new_n9765_));
  NOR2_X1    g06963(.A1(new_n9765_), .A2(new_n3455_), .ZN(new_n9766_));
  OR3_X2     g06964(.A1(new_n9527_), .A2(new_n3189_), .A3(new_n9766_), .Z(new_n9767_));
  NAND2_X1   g06965(.A1(new_n9548_), .A2(new_n2539_), .ZN(new_n9768_));
  OAI21_X1   g06966(.A1(new_n9765_), .A2(new_n9745_), .B(new_n3183_), .ZN(new_n9769_));
  AND3_X2    g06967(.A1(new_n9747_), .A2(new_n9768_), .A3(new_n9769_), .Z(new_n9770_));
  OAI21_X1   g06968(.A1(new_n9770_), .A2(new_n9551_), .B(new_n9527_), .ZN(new_n9771_));
  NAND2_X1   g06969(.A1(new_n9562_), .A2(pi0054), .ZN(new_n9772_));
  AOI22_X1   g06970(.A1(new_n9771_), .A2(new_n9772_), .B1(new_n3185_), .B2(new_n9767_), .ZN(new_n9773_));
  OAI21_X1   g06971(.A1(new_n9763_), .A2(new_n9764_), .B(new_n9773_), .ZN(new_n9774_));
  OR3_X2     g06972(.A1(new_n9743_), .A2(new_n9762_), .A3(new_n9774_), .Z(new_n9775_));
  NAND2_X1   g06973(.A1(new_n9775_), .A2(pi0079), .ZN(new_n9776_));
  NOR2_X1    g06974(.A1(new_n8219_), .A2(pi0034), .ZN(new_n9777_));
  INV_X1     g06975(.I(new_n9777_), .ZN(new_n9778_));
  NOR2_X1    g06976(.A1(new_n9778_), .A2(new_n7952_), .ZN(new_n9779_));
  XOR2_X1    g06977(.A1(new_n9776_), .A2(new_n9779_), .Z(new_n9780_));
  NAND2_X1   g06978(.A1(new_n9775_), .A2(new_n9777_), .ZN(new_n9781_));
  NOR2_X1    g06979(.A1(new_n9778_), .A2(pi0079), .ZN(new_n9782_));
  INV_X1     g06980(.I(new_n9782_), .ZN(new_n9783_));
  AOI21_X1   g06981(.A1(new_n7953_), .A2(new_n7958_), .B(new_n9783_), .ZN(new_n9784_));
  XOR2_X1    g06982(.A1(new_n9781_), .A2(new_n9784_), .Z(new_n9785_));
  AOI21_X1   g06983(.A1(new_n9780_), .A2(new_n9785_), .B(new_n9589_), .ZN(po0237));
  INV_X1     g06984(.I(pi0588), .ZN(new_n9787_));
  NOR2_X1    g06985(.A1(new_n2558_), .A2(new_n2979_), .ZN(new_n9788_));
  INV_X1     g06986(.I(new_n9788_), .ZN(new_n9789_));
  NOR2_X1    g06987(.A1(new_n9789_), .A2(new_n2984_), .ZN(new_n9790_));
  NOR2_X1    g06988(.A1(new_n2723_), .A2(pi0567), .ZN(new_n9791_));
  NOR2_X1    g06989(.A1(new_n9790_), .A2(new_n9791_), .ZN(new_n9792_));
  AOI21_X1   g06990(.A1(new_n9792_), .A2(new_n7129_), .B(new_n9787_), .ZN(new_n9793_));
  INV_X1     g06991(.I(new_n9792_), .ZN(new_n9796_));
  NAND2_X1   g06992(.A1(new_n9792_), .A2(pi0592), .ZN(new_n9798_));
  INV_X1     g06993(.I(new_n9790_), .ZN(new_n9799_));
  NOR2_X1    g06994(.A1(new_n9799_), .A2(new_n3474_), .ZN(new_n9800_));
  NOR2_X1    g06995(.A1(new_n5420_), .A2(new_n2512_), .ZN(new_n9801_));
  INV_X1     g06996(.I(new_n9801_), .ZN(new_n9802_));
  NAND3_X1   g06997(.A1(new_n8453_), .A2(new_n6360_), .A3(new_n2667_), .ZN(new_n9803_));
  NOR3_X1    g06998(.A1(new_n6362_), .A2(new_n9802_), .A3(new_n9803_), .ZN(new_n9804_));
  XOR2_X1    g06999(.A1(new_n2795_), .A2(new_n2509_), .Z(new_n9805_));
  NOR3_X1    g07000(.A1(new_n9805_), .A2(new_n2679_), .A3(new_n2732_), .ZN(new_n9806_));
  AOI21_X1   g07001(.A1(new_n9804_), .A2(new_n9806_), .B(pi0051), .ZN(new_n9807_));
  NOR4_X1    g07002(.A1(new_n3304_), .A2(new_n2755_), .A3(new_n5683_), .A4(new_n2722_), .ZN(new_n9808_));
  OAI21_X1   g07003(.A1(new_n9808_), .A2(new_n9788_), .B(new_n6369_), .ZN(new_n9809_));
  NOR2_X1    g07004(.A1(new_n9807_), .A2(new_n9809_), .ZN(new_n9810_));
  INV_X1     g07005(.I(new_n9810_), .ZN(new_n9811_));
  NOR2_X1    g07006(.A1(new_n9799_), .A2(new_n2726_), .ZN(new_n9812_));
  AOI21_X1   g07007(.A1(new_n9812_), .A2(new_n3193_), .B(new_n6940_), .ZN(new_n9813_));
  NAND4_X1   g07008(.A1(new_n6369_), .A2(pi0824), .A3(pi0950), .A4(new_n3144_), .ZN(new_n9814_));
  INV_X1     g07009(.I(new_n9814_), .ZN(new_n9815_));
  AOI21_X1   g07010(.A1(new_n9804_), .A2(new_n9815_), .B(pi0098), .ZN(new_n9816_));
  NOR2_X1    g07011(.A1(new_n9816_), .A2(new_n2979_), .ZN(new_n9817_));
  INV_X1     g07012(.I(new_n9812_), .ZN(new_n9818_));
  OAI21_X1   g07013(.A1(new_n9818_), .A2(new_n6989_), .B(new_n6941_), .ZN(new_n9819_));
  NAND2_X1   g07014(.A1(new_n9817_), .A2(new_n9819_), .ZN(new_n9820_));
  OAI21_X1   g07015(.A1(pi0567), .A2(new_n2723_), .B(new_n6399_), .ZN(new_n9825_));
  NAND2_X1   g07016(.A1(new_n9825_), .A2(new_n6358_), .ZN(new_n9826_));
  NAND2_X1   g07017(.A1(new_n9798_), .A2(new_n9826_), .ZN(new_n9827_));
  XOR2_X1    g07018(.A1(pi0426), .A2(pi0430), .Z(new_n9859_));
  NAND3_X1   g07019(.A1(new_n7124_), .A2(pi0448), .A3(new_n9859_), .ZN(new_n9861_));
  NAND2_X1   g07020(.A1(new_n9793_), .A2(new_n9861_), .ZN(new_n9862_));
  INV_X1     g07021(.I(new_n6407_), .ZN(new_n9863_));
  NOR2_X1    g07022(.A1(new_n9863_), .A2(new_n9790_), .ZN(new_n9864_));
  NAND2_X1   g07023(.A1(new_n6940_), .A2(pi0122), .ZN(new_n9865_));
  NOR2_X1    g07024(.A1(new_n9812_), .A2(new_n3474_), .ZN(new_n9866_));
  INV_X1     g07025(.I(new_n9866_), .ZN(new_n9867_));
  NOR2_X1    g07026(.A1(new_n9810_), .A2(new_n9867_), .ZN(new_n9868_));
  NAND2_X1   g07027(.A1(new_n9866_), .A2(pi0087), .ZN(new_n9869_));
  XNOR2_X1   g07028(.A1(new_n9868_), .A2(new_n9869_), .ZN(new_n9870_));
  NAND3_X1   g07029(.A1(new_n9870_), .A2(new_n9817_), .A3(new_n9866_), .ZN(new_n9871_));
  NOR2_X1    g07030(.A1(new_n6400_), .A2(new_n6514_), .ZN(new_n9872_));
  INV_X1     g07031(.I(new_n9872_), .ZN(new_n9873_));
  AOI21_X1   g07032(.A1(new_n9864_), .A2(new_n6394_), .B(new_n9873_), .ZN(new_n9875_));
  NOR2_X1    g07033(.A1(new_n9875_), .A2(pi0075), .ZN(new_n9876_));
  AOI21_X1   g07034(.A1(new_n9871_), .A2(new_n9865_), .B(new_n9876_), .ZN(new_n9877_));
  XOR2_X1    g07035(.A1(pi0426), .A2(pi0430), .Z(new_n9903_));
  NAND3_X1   g07036(.A1(new_n7124_), .A2(pi0448), .A3(new_n9903_), .ZN(new_n9905_));
  NAND2_X1   g07037(.A1(new_n9793_), .A2(new_n9905_), .ZN(new_n9906_));
  NOR2_X1    g07038(.A1(pi0590), .A2(pi0591), .ZN(new_n9907_));
  INV_X1     g07039(.I(new_n9907_), .ZN(new_n9908_));
  NOR2_X1    g07040(.A1(new_n6354_), .A2(new_n6352_), .ZN(new_n9935_));
  NOR2_X1    g07041(.A1(new_n9935_), .A2(pi0356), .ZN(new_n9936_));
  NOR2_X1    g07042(.A1(new_n9935_), .A2(new_n6650_), .ZN(new_n9937_));
  NOR2_X1    g07043(.A1(new_n9936_), .A2(new_n9937_), .ZN(new_n9938_));
  NOR3_X1    g07044(.A1(new_n6657_), .A2(new_n6653_), .A3(new_n9938_), .ZN(new_n9939_));
  NOR2_X1    g07045(.A1(new_n9939_), .A2(new_n9908_), .ZN(new_n9940_));
  OR3_X2     g07046(.A1(new_n6657_), .A2(new_n6653_), .A3(new_n9938_), .Z(new_n9941_));
  OAI21_X1   g07047(.A1(new_n9940_), .A2(new_n9941_), .B(new_n6669_), .ZN(new_n9942_));
  INV_X1     g07048(.I(new_n6657_), .ZN(new_n9943_));
  INV_X1     g07049(.I(new_n6352_), .ZN(new_n9944_));
  NAND2_X1   g07050(.A1(new_n9944_), .A2(new_n6353_), .ZN(new_n9964_));
  NAND2_X1   g07051(.A1(new_n9964_), .A2(new_n6650_), .ZN(new_n9965_));
  NAND2_X1   g07052(.A1(new_n9964_), .A2(pi0356), .ZN(new_n9966_));
  NAND2_X1   g07053(.A1(new_n9965_), .A2(new_n9966_), .ZN(new_n9967_));
  NAND3_X1   g07054(.A1(new_n9943_), .A2(pi0354), .A3(new_n9967_), .ZN(new_n9968_));
  NAND3_X1   g07055(.A1(new_n9943_), .A2(pi0354), .A3(new_n9967_), .ZN(new_n9969_));
  AOI21_X1   g07056(.A1(new_n9907_), .A2(new_n9968_), .B(new_n9969_), .ZN(new_n9970_));
  NOR2_X1    g07057(.A1(new_n6983_), .A2(new_n6728_), .ZN(new_n9971_));
  INV_X1     g07058(.I(new_n9971_), .ZN(new_n9972_));
  NOR2_X1    g07059(.A1(new_n6400_), .A2(new_n9791_), .ZN(new_n9973_));
  AOI21_X1   g07060(.A1(new_n6410_), .A2(new_n9789_), .B(new_n6403_), .ZN(new_n9974_));
  AOI22_X1   g07061(.A1(new_n6833_), .A2(new_n9974_), .B1(new_n6941_), .B2(new_n9818_), .ZN(new_n9975_));
  INV_X1     g07062(.I(new_n9975_), .ZN(new_n9976_));
  INV_X1     g07063(.I(new_n9817_), .ZN(new_n9978_));
  NOR2_X1    g07064(.A1(new_n6833_), .A2(new_n9788_), .ZN(new_n9979_));
  AOI21_X1   g07065(.A1(new_n6833_), .A2(new_n9978_), .B(new_n9979_), .ZN(new_n9980_));
  AOI21_X1   g07066(.A1(new_n6833_), .A2(new_n9811_), .B(new_n9979_), .ZN(new_n9981_));
  NOR2_X1    g07067(.A1(new_n6403_), .A2(pi0122), .ZN(new_n9986_));
  INV_X1     g07068(.I(new_n9986_), .ZN(new_n9987_));
  AOI21_X1   g07069(.A1(new_n9789_), .A2(new_n9987_), .B(new_n9976_), .ZN(new_n9988_));
  INV_X1     g07070(.I(new_n9988_), .ZN(new_n9989_));
  INV_X1     g07071(.I(new_n2723_), .ZN(new_n9992_));
  NOR2_X1    g07072(.A1(new_n9992_), .A2(pi0567), .ZN(new_n9993_));
  AOI21_X1   g07073(.A1(new_n9989_), .A2(pi0567), .B(new_n9993_), .ZN(new_n9994_));
  XNOR2_X1   g07074(.A1(pi0404), .A2(pi0411), .ZN(new_n9997_));
  NOR2_X1    g07075(.A1(pi0404), .A2(pi0411), .ZN(new_n9998_));
  INV_X1     g07076(.I(pi0411), .ZN(new_n9999_));
  NOR2_X1    g07077(.A1(new_n6773_), .A2(new_n9999_), .ZN(new_n10000_));
  OAI21_X1   g07078(.A1(new_n10000_), .A2(new_n9998_), .B(pi0397), .ZN(new_n10001_));
  OAI21_X1   g07079(.A1(pi0397), .A2(new_n9997_), .B(new_n10001_), .ZN(new_n10002_));
  NAND2_X1   g07080(.A1(new_n10002_), .A2(new_n6788_), .ZN(new_n10003_));
  OAI21_X1   g07081(.A1(new_n6789_), .A2(new_n10002_), .B(new_n10003_), .ZN(new_n10004_));
  AOI21_X1   g07082(.A1(new_n10004_), .A2(new_n6402_), .B(new_n9788_), .ZN(new_n10005_));
  AND2_X2    g07083(.A1(new_n6783_), .A2(pi0412), .Z(new_n10006_));
  OAI21_X1   g07084(.A1(new_n10004_), .A2(new_n6403_), .B(new_n9789_), .ZN(new_n10007_));
  NAND2_X1   g07085(.A1(new_n10007_), .A2(pi0412), .ZN(new_n10008_));
  XNOR2_X1   g07086(.A1(new_n10008_), .A2(new_n10006_), .ZN(new_n10009_));
  NAND2_X1   g07087(.A1(new_n10009_), .A2(new_n10005_), .ZN(new_n10010_));
  NAND2_X1   g07088(.A1(new_n10007_), .A2(new_n6783_), .ZN(new_n10011_));
  XNOR2_X1   g07089(.A1(new_n10011_), .A2(new_n10006_), .ZN(new_n10012_));
  NAND2_X1   g07090(.A1(new_n10012_), .A2(new_n10005_), .ZN(new_n10013_));
  NAND3_X1   g07091(.A1(new_n10010_), .A2(new_n10013_), .A3(new_n6410_), .ZN(new_n10014_));
  AOI21_X1   g07092(.A1(new_n10014_), .A2(new_n9789_), .B(new_n6941_), .ZN(new_n10015_));
  NOR2_X1    g07093(.A1(new_n10015_), .A2(new_n9812_), .ZN(new_n10016_));
  INV_X1     g07094(.I(new_n10016_), .ZN(new_n10017_));
  AOI21_X1   g07095(.A1(pi0567), .A2(new_n10017_), .B(new_n9994_), .ZN(new_n10018_));
  NAND2_X1   g07096(.A1(new_n6845_), .A2(new_n9788_), .ZN(new_n10021_));
  NAND2_X1   g07097(.A1(new_n6845_), .A2(new_n9978_), .ZN(new_n10022_));
  XNOR2_X1   g07098(.A1(new_n10021_), .A2(new_n10022_), .ZN(new_n10023_));
  AOI21_X1   g07099(.A1(new_n10016_), .A2(pi0567), .B(new_n9993_), .ZN(new_n10040_));
  NOR2_X1    g07100(.A1(new_n6792_), .A2(new_n9810_), .ZN(new_n10046_));
  XOR2_X1    g07101(.A1(new_n10021_), .A2(new_n10046_), .Z(new_n10047_));
  XNOR2_X1   g07102(.A1(pi0333), .A2(pi0391), .ZN(new_n10057_));
  XNOR2_X1   g07103(.A1(pi0392), .A2(pi0393), .ZN(new_n10062_));
  NOR3_X1    g07104(.A1(new_n6931_), .A2(new_n6350_), .A3(new_n10062_), .ZN(new_n10063_));
  NOR3_X1    g07105(.A1(new_n10063_), .A2(pi0588), .A3(pi0590), .ZN(new_n10064_));
  NAND2_X1   g07106(.A1(new_n9792_), .A2(new_n6358_), .ZN(new_n10065_));
  NAND2_X1   g07107(.A1(new_n9877_), .A2(pi0592), .ZN(new_n10066_));
  NAND2_X1   g07108(.A1(new_n10066_), .A2(new_n10065_), .ZN(new_n10067_));
  NOR2_X1    g07109(.A1(new_n10067_), .A2(new_n7188_), .ZN(new_n10068_));
  AOI21_X1   g07110(.A1(new_n7188_), .A2(new_n9796_), .B(new_n10068_), .ZN(new_n10069_));
  NAND2_X1   g07111(.A1(new_n10069_), .A2(pi1198), .ZN(new_n10070_));
  NAND3_X1   g07112(.A1(new_n10067_), .A2(pi1198), .A3(pi1199), .ZN(new_n10071_));
  XOR2_X1    g07113(.A1(new_n10070_), .A2(new_n10071_), .Z(new_n10072_));
  NOR2_X1    g07114(.A1(new_n10067_), .A2(new_n6731_), .ZN(new_n10073_));
  NOR2_X1    g07115(.A1(new_n9796_), .A2(new_n6731_), .ZN(new_n10074_));
  XNOR2_X1   g07116(.A1(new_n10073_), .A2(new_n10074_), .ZN(new_n10075_));
  AOI21_X1   g07117(.A1(new_n6728_), .A2(new_n9796_), .B(new_n6719_), .ZN(new_n10076_));
  OR3_X2     g07118(.A1(new_n10075_), .A2(new_n6720_), .A3(new_n6725_), .Z(new_n10078_));
  NAND2_X1   g07119(.A1(new_n10067_), .A2(new_n6719_), .ZN(new_n10079_));
  AOI21_X1   g07120(.A1(new_n10078_), .A2(new_n6356_), .B(new_n10079_), .ZN(new_n10080_));
  INV_X1     g07121(.I(new_n10080_), .ZN(new_n10081_));
  OAI21_X1   g07122(.A1(new_n10081_), .A2(pi1198), .B(new_n10072_), .ZN(new_n10082_));
  NOR2_X1    g07123(.A1(new_n10082_), .A2(pi0374), .ZN(new_n10083_));
  OAI21_X1   g07124(.A1(new_n6356_), .A2(new_n10069_), .B(new_n10081_), .ZN(new_n10084_));
  NOR2_X1    g07125(.A1(new_n10084_), .A2(new_n7178_), .ZN(new_n10085_));
  NOR2_X1    g07126(.A1(new_n10085_), .A2(new_n10083_), .ZN(new_n10086_));
  XOR2_X1    g07127(.A1(pi0370), .A2(pi0371), .Z(new_n10087_));
  INV_X1     g07128(.I(new_n10087_), .ZN(new_n10088_));
  XNOR2_X1   g07129(.A1(pi0370), .A2(pi0371), .ZN(new_n10089_));
  NOR2_X1    g07130(.A1(new_n6756_), .A2(new_n10089_), .ZN(new_n10090_));
  AOI21_X1   g07131(.A1(new_n6756_), .A2(new_n10088_), .B(new_n10090_), .ZN(new_n10091_));
  INV_X1     g07132(.I(new_n10091_), .ZN(new_n10092_));
  NAND2_X1   g07133(.A1(new_n10092_), .A2(pi0369), .ZN(new_n10093_));
  NOR2_X1    g07134(.A1(new_n10084_), .A2(pi0374), .ZN(new_n10094_));
  NOR2_X1    g07135(.A1(new_n10082_), .A2(new_n7178_), .ZN(new_n10095_));
  NOR2_X1    g07136(.A1(new_n10094_), .A2(new_n10095_), .ZN(new_n10096_));
  NAND2_X1   g07137(.A1(new_n10096_), .A2(pi0369), .ZN(new_n10097_));
  XNOR2_X1   g07138(.A1(new_n10097_), .A2(new_n10093_), .ZN(new_n10098_));
  NOR2_X1    g07139(.A1(new_n10098_), .A2(new_n10086_), .ZN(new_n10099_));
  NAND2_X1   g07140(.A1(new_n10096_), .A2(new_n10092_), .ZN(new_n10100_));
  XNOR2_X1   g07141(.A1(new_n10100_), .A2(new_n10093_), .ZN(new_n10101_));
  OAI21_X1   g07142(.A1(new_n10101_), .A2(new_n10086_), .B(new_n6350_), .ZN(new_n10102_));
  NOR4_X1    g07143(.A1(new_n10102_), .A2(new_n10099_), .A3(new_n9970_), .A4(new_n10064_), .ZN(new_n10103_));
  INV_X1     g07144(.I(new_n6931_), .ZN(new_n10104_));
  AOI21_X1   g07145(.A1(new_n9792_), .A2(new_n6400_), .B(new_n6816_), .ZN(new_n10105_));
  NOR2_X1    g07146(.A1(new_n9811_), .A2(new_n9813_), .ZN(new_n10106_));
  NAND2_X1   g07147(.A1(new_n9981_), .A2(new_n10106_), .ZN(new_n10107_));
  INV_X1     g07148(.I(new_n10107_), .ZN(new_n10108_));
  AOI21_X1   g07149(.A1(new_n9812_), .A2(new_n6554_), .B(new_n6940_), .ZN(new_n10109_));
  OAI22_X1   g07150(.A1(new_n10023_), .A2(new_n10109_), .B1(new_n10047_), .B2(new_n9813_), .ZN(new_n10110_));
  AND2_X2    g07151(.A1(new_n10110_), .A2(new_n9800_), .Z(new_n10111_));
  NOR2_X1    g07152(.A1(new_n6832_), .A2(new_n9820_), .ZN(new_n10112_));
  OAI21_X1   g07153(.A1(new_n10111_), .A2(new_n10108_), .B(new_n10112_), .ZN(new_n10113_));
  NAND2_X1   g07154(.A1(new_n10113_), .A2(new_n10105_), .ZN(new_n10114_));
  OAI22_X1   g07155(.A1(new_n9980_), .A2(new_n9799_), .B1(new_n3474_), .B2(new_n9820_), .ZN(new_n10115_));
  NAND2_X1   g07156(.A1(new_n10115_), .A2(new_n10107_), .ZN(new_n10116_));
  OAI21_X1   g07157(.A1(pi0592), .A2(pi1196), .B(new_n6399_), .ZN(new_n10117_));
  NOR2_X1    g07158(.A1(new_n9796_), .A2(new_n10117_), .ZN(new_n10118_));
  NOR2_X1    g07159(.A1(new_n9796_), .A2(new_n6356_), .ZN(new_n10119_));
  OAI21_X1   g07160(.A1(new_n10119_), .A2(new_n6991_), .B(new_n9973_), .ZN(new_n10120_));
  NOR2_X1    g07161(.A1(pi0075), .A2(pi0567), .ZN(new_n10121_));
  AOI22_X1   g07162(.A1(new_n10116_), .A2(new_n10118_), .B1(new_n10120_), .B2(new_n10121_), .ZN(new_n10122_));
  AOI21_X1   g07163(.A1(new_n10114_), .A2(new_n10122_), .B(new_n6770_), .ZN(new_n10123_));
  NOR2_X1    g07164(.A1(new_n9790_), .A2(new_n3235_), .ZN(new_n10124_));
  AOI21_X1   g07165(.A1(new_n10111_), .A2(new_n3235_), .B(new_n10124_), .ZN(new_n10125_));
  AOI21_X1   g07166(.A1(new_n10105_), .A2(new_n9973_), .B(pi0567), .ZN(new_n10126_));
  OAI21_X1   g07167(.A1(new_n10119_), .A2(pi1196), .B(pi0592), .ZN(new_n10127_));
  NOR4_X1    g07168(.A1(new_n10123_), .A2(new_n10125_), .A3(new_n10126_), .A4(new_n10127_), .ZN(new_n10128_));
  NOR4_X1    g07169(.A1(new_n10128_), .A2(new_n6728_), .A3(new_n6770_), .A4(new_n9827_), .ZN(new_n10129_));
  NOR2_X1    g07170(.A1(new_n10129_), .A2(new_n10057_), .ZN(new_n10130_));
  NOR2_X1    g07171(.A1(new_n6983_), .A2(new_n9827_), .ZN(new_n10131_));
  NOR3_X1    g07172(.A1(new_n10128_), .A2(new_n10057_), .A3(new_n10131_), .ZN(new_n10132_));
  XNOR2_X1   g07173(.A1(new_n10130_), .A2(new_n10132_), .ZN(new_n10133_));
  NOR2_X1    g07174(.A1(new_n10133_), .A2(pi0392), .ZN(new_n10134_));
  INV_X1     g07175(.I(pi0392), .ZN(new_n10135_));
  NOR2_X1    g07176(.A1(new_n10133_), .A2(new_n10135_), .ZN(new_n10136_));
  NOR2_X1    g07177(.A1(new_n10134_), .A2(new_n10136_), .ZN(new_n10137_));
  INV_X1     g07178(.I(new_n10137_), .ZN(new_n10138_));
  AND3_X2    g07179(.A1(new_n10138_), .A2(pi0393), .A3(new_n10104_), .Z(new_n10139_));
  INV_X1     g07180(.I(pi0369), .ZN(new_n10140_));
  NAND2_X1   g07181(.A1(new_n9825_), .A2(pi0592), .ZN(new_n10141_));
  NAND2_X1   g07182(.A1(new_n10065_), .A2(new_n10141_), .ZN(new_n10142_));
  NOR2_X1    g07183(.A1(new_n10142_), .A2(new_n6675_), .ZN(new_n10143_));
  NOR2_X1    g07184(.A1(new_n10142_), .A2(new_n6356_), .ZN(new_n10144_));
  NOR2_X1    g07185(.A1(new_n7187_), .A2(new_n6356_), .ZN(new_n10145_));
  XNOR2_X1   g07186(.A1(new_n10145_), .A2(new_n10144_), .ZN(new_n10146_));
  AOI21_X1   g07187(.A1(new_n10065_), .A2(new_n10141_), .B(new_n6718_), .ZN(new_n10147_));
  NOR4_X1    g07188(.A1(new_n10146_), .A2(pi1199), .A3(new_n9796_), .A4(new_n10147_), .ZN(new_n10148_));
  NOR2_X1    g07189(.A1(new_n10148_), .A2(new_n10076_), .ZN(new_n10149_));
  NOR2_X1    g07190(.A1(new_n10142_), .A2(new_n6728_), .ZN(new_n10150_));
  XOR2_X1    g07191(.A1(new_n6730_), .A2(pi0367), .Z(new_n10151_));
  NOR2_X1    g07192(.A1(new_n6727_), .A2(new_n10151_), .ZN(new_n10152_));
  NOR2_X1    g07193(.A1(new_n6726_), .A2(new_n6731_), .ZN(new_n10153_));
  OAI21_X1   g07194(.A1(new_n10152_), .A2(new_n10153_), .B(pi1197), .ZN(new_n10154_));
  XOR2_X1    g07195(.A1(new_n10154_), .A2(new_n10150_), .Z(new_n10155_));
  NOR4_X1    g07196(.A1(new_n10149_), .A2(new_n6675_), .A3(new_n9796_), .A4(new_n10155_), .ZN(new_n10156_));
  XNOR2_X1   g07197(.A1(new_n10156_), .A2(new_n10143_), .ZN(new_n10157_));
  NOR3_X1    g07198(.A1(new_n10157_), .A2(new_n10140_), .A3(new_n10091_), .ZN(new_n10158_));
  NOR2_X1    g07199(.A1(new_n10158_), .A2(new_n7129_), .ZN(new_n10159_));
  OR3_X2     g07200(.A1(new_n10157_), .A2(new_n10140_), .A3(new_n10091_), .Z(new_n10160_));
  OAI21_X1   g07201(.A1(new_n10159_), .A2(new_n10160_), .B(new_n6350_), .ZN(new_n10161_));
  NOR2_X1    g07202(.A1(new_n10139_), .A2(new_n10161_), .ZN(new_n10162_));
  INV_X1     g07203(.I(pi0080), .ZN(new_n10163_));
  NOR3_X1    g07204(.A1(new_n7240_), .A2(new_n10163_), .A3(new_n6668_), .ZN(new_n10164_));
  NAND4_X1   g07205(.A1(new_n10138_), .A2(pi0393), .A3(new_n10104_), .A4(new_n10164_), .ZN(new_n10165_));
  NOR3_X1    g07206(.A1(new_n10162_), .A2(new_n10103_), .A3(new_n10165_), .ZN(new_n10166_));
  NAND4_X1   g07207(.A1(new_n10166_), .A2(new_n9862_), .A3(new_n9906_), .A4(new_n9942_), .ZN(new_n10167_));
  INV_X1     g07208(.I(pi0217), .ZN(new_n10168_));
  INV_X1     g07209(.I(new_n7250_), .ZN(new_n10169_));
  OAI21_X1   g07210(.A1(new_n10168_), .A2(new_n10169_), .B(new_n9796_), .ZN(new_n10170_));
  AOI21_X1   g07211(.A1(new_n10170_), .A2(pi0080), .B(pi0217), .ZN(new_n10171_));
  NOR2_X1    g07212(.A1(new_n6358_), .A2(new_n6595_), .ZN(new_n10172_));
  NAND2_X1   g07213(.A1(new_n10040_), .A2(new_n10172_), .ZN(new_n10173_));
  NAND2_X1   g07214(.A1(new_n9792_), .A2(new_n10172_), .ZN(new_n10174_));
  XNOR2_X1   g07215(.A1(new_n10173_), .A2(new_n10174_), .ZN(new_n10175_));
  NAND2_X1   g07216(.A1(new_n9994_), .A2(pi0592), .ZN(new_n10176_));
  XNOR2_X1   g07217(.A1(new_n10176_), .A2(new_n10174_), .ZN(new_n10177_));
  OAI21_X1   g07218(.A1(new_n10018_), .A2(new_n6816_), .B(pi1199), .ZN(new_n10178_));
  OAI22_X1   g07219(.A1(new_n10177_), .A2(new_n10178_), .B1(pi1199), .B2(new_n10175_), .ZN(new_n10179_));
  NOR2_X1    g07220(.A1(new_n10179_), .A2(new_n9972_), .ZN(new_n10180_));
  NOR2_X1    g07221(.A1(new_n7191_), .A2(new_n9796_), .ZN(new_n10181_));
  NAND2_X1   g07222(.A1(new_n9971_), .A2(new_n10181_), .ZN(new_n10182_));
  XNOR2_X1   g07223(.A1(new_n10180_), .A2(new_n10182_), .ZN(new_n10183_));
  NOR3_X1    g07224(.A1(new_n6983_), .A2(new_n7191_), .A3(new_n9796_), .ZN(new_n10184_));
  AOI21_X1   g07225(.A1(new_n10179_), .A2(new_n6983_), .B(new_n10184_), .ZN(new_n10185_));
  NOR2_X1    g07226(.A1(new_n10185_), .A2(new_n6757_), .ZN(new_n10186_));
  AOI21_X1   g07227(.A1(new_n10183_), .A2(new_n6757_), .B(new_n10186_), .ZN(new_n10187_));
  XOR2_X1    g07228(.A1(new_n6932_), .A2(new_n10135_), .Z(new_n10188_));
  NAND2_X1   g07229(.A1(new_n10188_), .A2(pi0391), .ZN(new_n10189_));
  NOR2_X1    g07230(.A1(new_n10185_), .A2(pi0333), .ZN(new_n10190_));
  AOI21_X1   g07231(.A1(new_n10183_), .A2(pi0333), .B(new_n10190_), .ZN(new_n10191_));
  NAND2_X1   g07232(.A1(new_n10191_), .A2(pi0391), .ZN(new_n10192_));
  XNOR2_X1   g07233(.A1(new_n10192_), .A2(new_n10189_), .ZN(new_n10193_));
  OAI22_X1   g07234(.A1(new_n7185_), .A2(new_n6577_), .B1(pi0592), .B2(new_n7153_), .ZN(new_n10194_));
  NOR2_X1    g07235(.A1(new_n7190_), .A2(new_n7153_), .ZN(new_n10195_));
  NAND2_X1   g07236(.A1(new_n7152_), .A2(pi1198), .ZN(new_n10196_));
  XOR2_X1    g07237(.A1(new_n10195_), .A2(new_n10196_), .Z(new_n10197_));
  OAI21_X1   g07238(.A1(new_n9792_), .A2(new_n6934_), .B(pi0592), .ZN(new_n10198_));
  NOR2_X1    g07239(.A1(new_n10197_), .A2(new_n10198_), .ZN(new_n10199_));
  AOI21_X1   g07240(.A1(new_n10199_), .A2(new_n10194_), .B(pi0591), .ZN(new_n10200_));
  OAI21_X1   g07241(.A1(new_n10193_), .A2(new_n10187_), .B(new_n10200_), .ZN(new_n10201_));
  NAND2_X1   g07242(.A1(new_n10191_), .A2(new_n10188_), .ZN(new_n10202_));
  XNOR2_X1   g07243(.A1(new_n10202_), .A2(new_n10189_), .ZN(new_n10203_));
  NOR2_X1    g07244(.A1(new_n10203_), .A2(new_n10187_), .ZN(new_n10204_));
  NOR2_X1    g07245(.A1(new_n6354_), .A2(new_n6352_), .ZN(new_n10207_));
  NOR2_X1    g07246(.A1(new_n10207_), .A2(pi0356), .ZN(new_n10208_));
  NOR2_X1    g07247(.A1(new_n10207_), .A2(new_n6650_), .ZN(new_n10209_));
  NOR2_X1    g07248(.A1(new_n10208_), .A2(new_n10209_), .ZN(new_n10210_));
  NOR3_X1    g07249(.A1(new_n6657_), .A2(new_n6653_), .A3(new_n10210_), .ZN(new_n10211_));
  NOR2_X1    g07250(.A1(new_n10211_), .A2(new_n9908_), .ZN(new_n10212_));
  OR3_X2     g07251(.A1(new_n6657_), .A2(new_n6653_), .A3(new_n10210_), .Z(new_n10213_));
  OAI21_X1   g07252(.A1(new_n10212_), .A2(new_n10213_), .B(new_n9787_), .ZN(new_n10214_));
  AOI21_X1   g07253(.A1(new_n10201_), .A2(new_n10204_), .B(new_n10214_), .ZN(new_n10215_));
  NOR3_X1    g07254(.A1(new_n6667_), .A2(new_n6662_), .A3(new_n6663_), .ZN(new_n10217_));
  INV_X1     g07255(.I(new_n9793_), .ZN(new_n10218_));
  XOR2_X1    g07256(.A1(pi0426), .A2(pi0430), .Z(new_n10223_));
  AND3_X2    g07257(.A1(new_n7124_), .A2(pi0448), .A3(new_n10223_), .Z(new_n10226_));
  NOR2_X1    g07258(.A1(new_n10218_), .A2(new_n10226_), .ZN(new_n10227_));
  OAI21_X1   g07259(.A1(new_n10215_), .A2(new_n10217_), .B(new_n10227_), .ZN(new_n10228_));
  AOI21_X1   g07260(.A1(new_n10167_), .A2(new_n10171_), .B(new_n10228_), .ZN(po0238));
  NOR2_X1    g07261(.A1(new_n2644_), .A2(new_n2492_), .ZN(new_n10230_));
  INV_X1     g07262(.I(new_n10230_), .ZN(new_n10231_));
  NOR4_X1    g07263(.A1(new_n10231_), .A2(new_n2605_), .A3(new_n2611_), .A4(new_n2610_), .ZN(new_n10232_));
  NAND4_X1   g07264(.A1(new_n2603_), .A2(new_n7286_), .A3(new_n8958_), .A4(new_n10232_), .ZN(new_n10233_));
  NAND3_X1   g07265(.A1(new_n10233_), .A2(new_n2492_), .A3(new_n2453_), .ZN(new_n10234_));
  NAND2_X1   g07266(.A1(new_n9150_), .A2(new_n7240_), .ZN(new_n10235_));
  AOI21_X1   g07267(.A1(pi0314), .A2(new_n10234_), .B(new_n10235_), .ZN(po0239));
  NAND2_X1   g07268(.A1(pi0067), .A2(pi0069), .ZN(new_n10237_));
  NOR3_X1    g07269(.A1(new_n2620_), .A2(new_n9231_), .A3(new_n10237_), .ZN(new_n10238_));
  NOR4_X1    g07270(.A1(new_n2567_), .A2(new_n2571_), .A3(pi0073), .A4(new_n2624_), .ZN(new_n10239_));
  NAND2_X1   g07271(.A1(new_n9021_), .A2(new_n2446_), .ZN(new_n10240_));
  NOR4_X1    g07272(.A1(new_n9020_), .A2(new_n10238_), .A3(new_n10239_), .A4(new_n10240_), .ZN(po0240));
  INV_X1     g07273(.I(new_n9021_), .ZN(new_n10242_));
  NOR2_X1    g07274(.A1(new_n10242_), .A2(new_n7408_), .ZN(new_n10243_));
  INV_X1     g07275(.I(new_n10243_), .ZN(new_n10244_));
  NAND3_X1   g07276(.A1(new_n2609_), .A2(new_n2605_), .A3(new_n2534_), .ZN(new_n10245_));
  NOR4_X1    g07277(.A1(new_n10245_), .A2(new_n2611_), .A3(new_n2598_), .A4(new_n2624_), .ZN(new_n10246_));
  INV_X1     g07278(.I(new_n10246_), .ZN(new_n10247_));
  NOR2_X1    g07279(.A1(new_n2627_), .A2(new_n10243_), .ZN(new_n10248_));
  NAND2_X1   g07280(.A1(new_n10246_), .A2(pi0083), .ZN(new_n10249_));
  OAI21_X1   g07281(.A1(new_n10248_), .A2(new_n10249_), .B(new_n8291_), .ZN(new_n10250_));
  XNOR2_X1   g07282(.A1(new_n10250_), .A2(new_n9436_), .ZN(new_n10251_));
  NOR4_X1    g07283(.A1(new_n10251_), .A2(new_n7362_), .A3(new_n10244_), .A4(new_n10247_), .ZN(po0241));
  NOR2_X1    g07284(.A1(new_n3098_), .A2(pi0211), .ZN(new_n10253_));
  NOR2_X1    g07285(.A1(new_n8683_), .A2(new_n3098_), .ZN(new_n10254_));
  NAND2_X1   g07286(.A1(new_n10254_), .A2(new_n8772_), .ZN(new_n10255_));
  XOR2_X1    g07287(.A1(new_n10255_), .A2(new_n10253_), .Z(new_n10256_));
  NOR3_X1    g07288(.A1(new_n9212_), .A2(po1038), .A3(new_n10256_), .ZN(po0242));
  NOR2_X1    g07289(.A1(new_n9022_), .A2(new_n2607_), .ZN(new_n10258_));
  INV_X1     g07290(.I(new_n9256_), .ZN(new_n10259_));
  NAND4_X1   g07291(.A1(new_n10259_), .A2(new_n9231_), .A3(new_n9019_), .A4(new_n10258_), .ZN(new_n10260_));
  AOI21_X1   g07292(.A1(new_n10260_), .A2(new_n2634_), .B(new_n9022_), .ZN(po0243));
  AOI21_X1   g07293(.A1(new_n6542_), .A2(new_n9226_), .B(new_n9223_), .ZN(new_n10262_));
  NOR2_X1    g07294(.A1(new_n10262_), .A2(new_n6539_), .ZN(po0244));
  NOR3_X1    g07295(.A1(new_n2636_), .A2(new_n2465_), .A3(new_n10242_), .ZN(new_n10264_));
  INV_X1     g07296(.I(new_n10264_), .ZN(new_n10265_));
  NOR4_X1    g07297(.A1(new_n10265_), .A2(new_n8292_), .A3(new_n9231_), .A4(new_n2469_), .ZN(po0245));
  INV_X1     g07298(.I(new_n9803_), .ZN(new_n10267_));
  NAND4_X1   g07299(.A1(new_n8969_), .A2(pi0094), .A3(new_n6361_), .A4(new_n10267_), .ZN(new_n10268_));
  NOR4_X1    g07300(.A1(new_n10268_), .A2(new_n6403_), .A3(new_n8290_), .A4(new_n9802_), .ZN(new_n10269_));
  INV_X1     g07301(.I(new_n10269_), .ZN(new_n10270_));
  OAI21_X1   g07302(.A1(new_n3291_), .A2(new_n2987_), .B(pi1093), .ZN(new_n10271_));
  OAI22_X1   g07303(.A1(new_n10270_), .A2(new_n10271_), .B1(new_n8303_), .B2(new_n8970_), .ZN(new_n10272_));
  AOI21_X1   g07304(.A1(new_n10272_), .A2(new_n6402_), .B(new_n6939_), .ZN(new_n10273_));
  XOR2_X1    g07305(.A1(new_n10273_), .A2(new_n7253_), .Z(new_n10274_));
  INV_X1     g07306(.I(new_n3304_), .ZN(new_n10275_));
  NAND3_X1   g07307(.A1(new_n10275_), .A2(pi0088), .A3(pi1093), .ZN(new_n10276_));
  NOR4_X1    g07308(.A1(new_n3292_), .A2(new_n10276_), .A3(new_n2481_), .A4(new_n6403_), .ZN(new_n10277_));
  NAND4_X1   g07309(.A1(new_n10277_), .A2(new_n2558_), .A3(new_n2557_), .A4(new_n8282_), .ZN(new_n10278_));
  NOR2_X1    g07310(.A1(new_n10274_), .A2(new_n10278_), .ZN(po0246));
  NAND4_X1   g07311(.A1(new_n8315_), .A2(new_n8304_), .A3(new_n7275_), .A4(new_n10230_), .ZN(new_n10280_));
  INV_X1     g07312(.I(new_n10280_), .ZN(new_n10281_));
  NOR3_X1    g07313(.A1(new_n10281_), .A2(pi0070), .A3(pi0841), .ZN(new_n10282_));
  NOR3_X1    g07314(.A1(new_n8288_), .A2(new_n2707_), .A3(new_n3143_), .ZN(new_n10283_));
  OAI21_X1   g07315(.A1(new_n10282_), .A2(new_n6368_), .B(new_n10283_), .ZN(new_n10284_));
  AOI21_X1   g07316(.A1(new_n10284_), .A2(new_n2853_), .B(new_n7272_), .ZN(po0247));
  NOR2_X1    g07317(.A1(new_n2679_), .A2(new_n9279_), .ZN(new_n10286_));
  OAI21_X1   g07318(.A1(new_n7411_), .A2(new_n9174_), .B(new_n10286_), .ZN(new_n10287_));
  AOI21_X1   g07319(.A1(new_n10287_), .A2(new_n2732_), .B(new_n2471_), .ZN(po0248));
  OAI22_X1   g07320(.A1(new_n8281_), .A2(new_n8283_), .B1(pi0058), .B2(new_n2868_), .ZN(new_n10289_));
  NOR2_X1    g07321(.A1(new_n9009_), .A2(pi0039), .ZN(new_n10290_));
  NAND2_X1   g07322(.A1(new_n2868_), .A2(new_n10290_), .ZN(new_n10291_));
  NOR3_X1    g07323(.A1(new_n2731_), .A2(new_n7272_), .A3(new_n2798_), .ZN(new_n10292_));
  NAND2_X1   g07324(.A1(new_n8290_), .A2(new_n2745_), .ZN(new_n10293_));
  AOI21_X1   g07325(.A1(new_n10291_), .A2(new_n10292_), .B(new_n10293_), .ZN(new_n10294_));
  OAI21_X1   g07326(.A1(new_n10289_), .A2(new_n10294_), .B(new_n8297_), .ZN(new_n10295_));
  NOR2_X1    g07327(.A1(new_n6551_), .A2(new_n10295_), .ZN(po0249));
  NOR3_X1    g07328(.A1(new_n3382_), .A2(new_n3099_), .A3(new_n3100_), .ZN(new_n10297_));
  AOI22_X1   g07329(.A1(new_n6538_), .A2(new_n10297_), .B1(new_n6542_), .B2(new_n9241_), .ZN(new_n10298_));
  INV_X1     g07330(.I(new_n8286_), .ZN(new_n10299_));
  NAND4_X1   g07331(.A1(new_n3437_), .A2(pi0092), .A3(new_n9231_), .A4(pi1050), .ZN(new_n10300_));
  NOR2_X1    g07332(.A1(new_n10300_), .A2(new_n10299_), .ZN(new_n10301_));
  AOI22_X1   g07333(.A1(new_n10301_), .A2(new_n3160_), .B1(new_n3205_), .B2(new_n9045_), .ZN(new_n10302_));
  NOR2_X1    g07334(.A1(new_n10298_), .A2(new_n10302_), .ZN(po0250));
  NOR2_X1    g07335(.A1(new_n8286_), .A2(new_n3437_), .ZN(new_n10304_));
  NOR4_X1    g07336(.A1(new_n10304_), .A2(new_n9173_), .A3(new_n3303_), .A4(new_n2732_), .ZN(new_n10305_));
  NAND2_X1   g07337(.A1(new_n2879_), .A2(new_n10305_), .ZN(new_n10306_));
  AOI21_X1   g07338(.A1(new_n10306_), .A2(new_n3145_), .B(new_n9279_), .ZN(po0251));
  NAND2_X1   g07339(.A1(new_n8997_), .A2(new_n9145_), .ZN(new_n10308_));
  NAND2_X1   g07340(.A1(new_n2982_), .A2(pi1093), .ZN(new_n10309_));
  AOI21_X1   g07341(.A1(new_n10308_), .A2(new_n10309_), .B(new_n2730_), .ZN(new_n10310_));
  OAI21_X1   g07342(.A1(new_n8290_), .A2(new_n2903_), .B(new_n3721_), .ZN(new_n10311_));
  NOR2_X1    g07343(.A1(new_n8996_), .A2(new_n8370_), .ZN(new_n10312_));
  NOR2_X1    g07344(.A1(new_n2549_), .A2(new_n10312_), .ZN(new_n10313_));
  OAI21_X1   g07345(.A1(new_n10310_), .A2(new_n10311_), .B(new_n10313_), .ZN(new_n10314_));
  NAND2_X1   g07346(.A1(new_n10314_), .A2(new_n3721_), .ZN(new_n10315_));
  OAI21_X1   g07347(.A1(new_n10308_), .A2(new_n3721_), .B(new_n8384_), .ZN(new_n10316_));
  AOI21_X1   g07348(.A1(new_n10315_), .A2(po0840), .B(new_n10316_), .ZN(new_n10317_));
  NOR2_X1    g07349(.A1(new_n9003_), .A2(new_n8288_), .ZN(new_n10318_));
  XNOR2_X1   g07350(.A1(new_n10317_), .A2(new_n10318_), .ZN(new_n10319_));
  NOR2_X1    g07351(.A1(new_n10319_), .A2(new_n10308_), .ZN(po0252));
  NOR3_X1    g07352(.A1(new_n5400_), .A2(new_n3384_), .A3(new_n9244_), .ZN(new_n10321_));
  NAND3_X1   g07353(.A1(new_n2734_), .A2(new_n2794_), .A3(pi0095), .ZN(new_n10322_));
  NOR3_X1    g07354(.A1(new_n2733_), .A2(new_n7272_), .A3(new_n10322_), .ZN(new_n10323_));
  NOR3_X1    g07355(.A1(new_n10323_), .A2(pi0039), .A3(new_n8346_), .ZN(new_n10324_));
  NOR4_X1    g07356(.A1(new_n8290_), .A2(new_n2955_), .A3(pi0841), .A4(new_n2479_), .ZN(new_n10325_));
  NAND2_X1   g07357(.A1(new_n10281_), .A2(new_n10325_), .ZN(new_n10326_));
  OAI21_X1   g07358(.A1(new_n10324_), .A2(new_n10326_), .B(new_n3183_), .ZN(new_n10327_));
  AOI21_X1   g07359(.A1(new_n5698_), .A2(new_n10321_), .B(new_n10327_), .ZN(new_n10328_));
  AOI21_X1   g07360(.A1(new_n5461_), .A2(new_n9241_), .B(new_n5699_), .ZN(new_n10329_));
  NOR4_X1    g07361(.A1(new_n10328_), .A2(new_n2777_), .A3(new_n9243_), .A4(new_n10329_), .ZN(po0253));
  NOR2_X1    g07362(.A1(po0840), .A2(new_n2890_), .ZN(new_n10331_));
  INV_X1     g07363(.I(new_n10331_), .ZN(new_n10332_));
  NOR4_X1    g07364(.A1(new_n2816_), .A2(new_n2436_), .A3(new_n2755_), .A4(new_n5431_), .ZN(new_n10333_));
  AND3_X2    g07365(.A1(new_n2917_), .A2(new_n10332_), .A3(new_n10333_), .Z(new_n10334_));
  NOR4_X1    g07366(.A1(new_n2817_), .A2(pi0072), .A3(new_n2816_), .A4(new_n8288_), .ZN(new_n10335_));
  OAI21_X1   g07367(.A1(new_n10334_), .A2(new_n10331_), .B(new_n10335_), .ZN(new_n10336_));
  AOI21_X1   g07368(.A1(new_n10336_), .A2(new_n10322_), .B(new_n8507_), .ZN(po0254));
  NOR4_X1    g07369(.A1(new_n8236_), .A2(pi0039), .A3(pi0096), .A4(new_n3304_), .ZN(new_n10338_));
  OAI21_X1   g07370(.A1(new_n10338_), .A2(new_n5469_), .B(new_n10331_), .ZN(new_n10339_));
  AND2_X2    g07371(.A1(pi0039), .A2(pi0593), .Z(new_n10340_));
  NAND4_X1   g07372(.A1(new_n5699_), .A2(new_n8346_), .A3(new_n9247_), .A4(new_n10340_), .ZN(new_n10341_));
  AOI21_X1   g07373(.A1(new_n10341_), .A2(new_n10339_), .B(new_n9289_), .ZN(po0255));
  NOR4_X1    g07374(.A1(new_n10299_), .A2(new_n9231_), .A3(new_n3495_), .A4(new_n9279_), .ZN(new_n10343_));
  NAND3_X1   g07375(.A1(new_n10343_), .A2(pi0092), .A3(new_n3160_), .ZN(new_n10344_));
  NAND3_X1   g07376(.A1(new_n10343_), .A2(new_n3303_), .A3(new_n3145_), .ZN(new_n10345_));
  AOI21_X1   g07377(.A1(new_n10344_), .A2(new_n10345_), .B(new_n9287_), .ZN(po0256));
  INV_X1     g07378(.I(pi0099), .ZN(new_n10347_));
  AOI21_X1   g07379(.A1(pi0041), .A2(pi0072), .B(new_n10347_), .ZN(new_n10348_));
  NAND2_X1   g07380(.A1(new_n8430_), .A2(new_n10348_), .ZN(new_n10349_));
  NOR2_X1    g07381(.A1(new_n8787_), .A2(new_n8788_), .ZN(new_n10350_));
  AOI21_X1   g07382(.A1(new_n10350_), .A2(new_n10349_), .B(new_n10348_), .ZN(new_n10351_));
  INV_X1     g07383(.I(new_n8600_), .ZN(new_n10352_));
  OAI21_X1   g07384(.A1(new_n10352_), .A2(pi0228), .B(new_n10348_), .ZN(new_n10353_));
  OAI21_X1   g07385(.A1(new_n8477_), .A2(new_n10353_), .B(new_n3183_), .ZN(new_n10354_));
  NAND2_X1   g07386(.A1(new_n8899_), .A2(new_n5522_), .ZN(new_n10355_));
  NOR2_X1    g07387(.A1(new_n10347_), .A2(pi0072), .ZN(new_n10356_));
  OAI21_X1   g07388(.A1(new_n8511_), .A2(new_n8505_), .B(new_n10356_), .ZN(new_n10357_));
  INV_X1     g07389(.I(new_n8487_), .ZN(new_n10358_));
  NAND2_X1   g07390(.A1(new_n10358_), .A2(new_n2729_), .ZN(new_n10359_));
  AOI21_X1   g07391(.A1(new_n10357_), .A2(new_n10355_), .B(new_n10359_), .ZN(new_n10360_));
  AOI21_X1   g07392(.A1(new_n8438_), .A2(pi0144), .B(new_n3098_), .ZN(new_n10361_));
  NAND4_X1   g07393(.A1(new_n8442_), .A2(pi0072), .A3(pi0152), .A4(pi0161), .ZN(new_n10362_));
  NOR4_X1    g07394(.A1(new_n10362_), .A2(pi0072), .A3(new_n7378_), .A4(new_n3098_), .ZN(new_n10363_));
  XOR2_X1    g07395(.A1(new_n10363_), .A2(new_n10361_), .Z(new_n10364_));
  OAI21_X1   g07396(.A1(new_n10364_), .A2(new_n5551_), .B(pi0039), .ZN(new_n10365_));
  INV_X1     g07397(.I(new_n10365_), .ZN(new_n10366_));
  INV_X1     g07398(.I(new_n10356_), .ZN(new_n10367_));
  NOR4_X1    g07399(.A1(new_n6511_), .A2(new_n3183_), .A3(new_n2729_), .A4(new_n10367_), .ZN(new_n10368_));
  OAI21_X1   g07400(.A1(new_n10366_), .A2(new_n3186_), .B(new_n10368_), .ZN(new_n10369_));
  OAI21_X1   g07401(.A1(new_n10360_), .A2(new_n10369_), .B(new_n3235_), .ZN(new_n10370_));
  AOI21_X1   g07402(.A1(new_n3183_), .A2(new_n10367_), .B(new_n10366_), .ZN(new_n10371_));
  INV_X1     g07403(.I(new_n10371_), .ZN(new_n10372_));
  NOR2_X1    g07404(.A1(new_n10372_), .A2(new_n3187_), .ZN(new_n10373_));
  NOR3_X1    g07405(.A1(new_n8491_), .A2(new_n3005_), .A3(new_n5521_), .ZN(new_n10374_));
  AOI21_X1   g07406(.A1(new_n3213_), .A2(new_n10356_), .B(pi0228), .ZN(new_n10375_));
  NOR4_X1    g07407(.A1(new_n8612_), .A2(new_n8505_), .A3(new_n10374_), .A4(new_n10375_), .ZN(new_n10376_));
  OAI21_X1   g07408(.A1(new_n10371_), .A2(new_n3213_), .B(pi0087), .ZN(new_n10377_));
  OAI21_X1   g07409(.A1(new_n10376_), .A2(new_n10377_), .B(new_n3235_), .ZN(new_n10378_));
  AOI21_X1   g07410(.A1(new_n10370_), .A2(new_n10373_), .B(new_n10378_), .ZN(new_n10379_));
  AOI21_X1   g07411(.A1(new_n5520_), .A2(new_n10356_), .B(new_n2730_), .ZN(new_n10380_));
  NAND2_X1   g07412(.A1(new_n10358_), .A2(new_n10380_), .ZN(new_n10381_));
  AOI21_X1   g07413(.A1(new_n8485_), .A2(new_n8492_), .B(new_n10381_), .ZN(new_n10382_));
  OAI21_X1   g07414(.A1(new_n10365_), .A2(new_n5506_), .B(new_n3183_), .ZN(new_n10383_));
  NAND4_X1   g07415(.A1(new_n10383_), .A2(new_n2730_), .A3(new_n8494_), .A4(new_n10356_), .ZN(new_n10384_));
  OAI21_X1   g07416(.A1(new_n10382_), .A2(new_n10384_), .B(new_n3455_), .ZN(new_n10385_));
  NOR2_X1    g07417(.A1(new_n10372_), .A2(new_n3259_), .ZN(new_n10386_));
  OAI21_X1   g07418(.A1(new_n8536_), .A2(new_n10364_), .B(new_n8881_), .ZN(new_n10387_));
  NAND2_X1   g07419(.A1(new_n10387_), .A2(new_n3133_), .ZN(new_n10388_));
  AOI21_X1   g07420(.A1(new_n10385_), .A2(new_n10386_), .B(new_n10388_), .ZN(new_n10389_));
  NAND3_X1   g07421(.A1(new_n8714_), .A2(new_n7240_), .A3(new_n10356_), .ZN(new_n10391_));
  OAI21_X1   g07422(.A1(new_n10372_), .A2(new_n10391_), .B(new_n6400_), .ZN(new_n10392_));
  NAND2_X1   g07423(.A1(new_n10392_), .A2(pi0228), .ZN(new_n10393_));
  NOR3_X1    g07424(.A1(new_n10379_), .A2(new_n10389_), .A3(new_n10393_), .ZN(new_n10394_));
  NAND3_X1   g07425(.A1(new_n8416_), .A2(new_n10354_), .A3(new_n10394_), .ZN(new_n10395_));
  NOR2_X1    g07426(.A1(new_n10395_), .A2(new_n10351_), .ZN(po0257));
  NOR2_X1    g07427(.A1(new_n7332_), .A2(new_n3160_), .ZN(new_n10397_));
  OAI21_X1   g07428(.A1(new_n7318_), .A2(new_n6492_), .B(new_n8250_), .ZN(new_n10398_));
  NAND2_X1   g07429(.A1(new_n8250_), .A2(pi0129), .ZN(new_n10399_));
  AOI22_X1   g07430(.A1(new_n10398_), .A2(new_n6493_), .B1(new_n8251_), .B2(new_n10399_), .ZN(new_n10400_));
  NAND4_X1   g07431(.A1(new_n5505_), .A2(pi0024), .A3(pi0075), .A4(new_n3191_), .ZN(new_n10401_));
  NOR4_X1    g07432(.A1(new_n5502_), .A2(new_n7294_), .A3(new_n9015_), .A4(new_n10401_), .ZN(new_n10402_));
  NAND2_X1   g07433(.A1(new_n5538_), .A2(new_n10402_), .ZN(new_n10403_));
  NOR4_X1    g07434(.A1(new_n10400_), .A2(new_n7327_), .A3(new_n10397_), .A4(new_n10403_), .ZN(po0258));
  NAND2_X1   g07435(.A1(new_n2729_), .A2(pi0101), .ZN(new_n10405_));
  XOR2_X1    g07436(.A1(new_n8427_), .A2(new_n10405_), .Z(new_n10406_));
  NOR2_X1    g07437(.A1(new_n8413_), .A2(new_n2730_), .ZN(new_n10407_));
  XOR2_X1    g07438(.A1(new_n10407_), .A2(new_n10405_), .Z(new_n10408_));
  OAI22_X1   g07439(.A1(new_n10408_), .A2(new_n8420_), .B1(new_n8432_), .B2(new_n10406_), .ZN(new_n10409_));
  NAND2_X1   g07440(.A1(new_n10409_), .A2(pi0228), .ZN(new_n10410_));
  AOI21_X1   g07441(.A1(pi0299), .A2(new_n8536_), .B(new_n8882_), .ZN(new_n10411_));
  NOR3_X1    g07442(.A1(new_n8439_), .A2(pi0144), .A3(new_n7378_), .ZN(new_n10412_));
  NAND2_X1   g07443(.A1(new_n10412_), .A2(new_n3132_), .ZN(new_n10413_));
  OAI21_X1   g07444(.A1(new_n10411_), .A2(new_n10413_), .B(new_n3098_), .ZN(new_n10414_));
  NOR4_X1    g07445(.A1(new_n8881_), .A2(pi0072), .A3(new_n3397_), .A4(new_n5386_), .ZN(new_n10415_));
  AOI21_X1   g07446(.A1(new_n10414_), .A2(new_n10415_), .B(pi0039), .ZN(new_n10416_));
  NOR3_X1    g07447(.A1(new_n8533_), .A2(new_n8389_), .A3(new_n3005_), .ZN(new_n10417_));
  AND3_X2    g07448(.A1(new_n8533_), .A2(pi0101), .A3(new_n3005_), .Z(new_n10418_));
  NOR3_X1    g07449(.A1(new_n8479_), .A2(new_n6486_), .A3(new_n8482_), .ZN(new_n10419_));
  NAND2_X1   g07450(.A1(new_n5525_), .A2(new_n2730_), .ZN(new_n10420_));
  NAND3_X1   g07451(.A1(new_n10420_), .A2(new_n8492_), .A3(pi0044), .ZN(new_n10421_));
  INV_X1     g07452(.I(new_n8482_), .ZN(new_n10422_));
  NAND4_X1   g07453(.A1(new_n3394_), .A2(new_n5373_), .A3(new_n2437_), .A4(pi0152), .ZN(new_n10423_));
  OAI21_X1   g07454(.A1(new_n10412_), .A2(new_n5912_), .B(new_n8707_), .ZN(new_n10424_));
  AOI21_X1   g07455(.A1(new_n10424_), .A2(new_n3098_), .B(new_n10423_), .ZN(new_n10425_));
  AOI21_X1   g07456(.A1(new_n10425_), .A2(new_n5505_), .B(pi0039), .ZN(new_n10426_));
  OAI21_X1   g07457(.A1(new_n8494_), .A2(new_n10422_), .B(new_n2730_), .ZN(new_n10427_));
  NOR3_X1    g07458(.A1(new_n10427_), .A2(new_n10422_), .A3(new_n10426_), .ZN(new_n10428_));
  OAI21_X1   g07459(.A1(new_n10419_), .A2(new_n10421_), .B(new_n10428_), .ZN(new_n10429_));
  AOI21_X1   g07460(.A1(new_n3183_), .A2(new_n10422_), .B(new_n10425_), .ZN(new_n10430_));
  NAND2_X1   g07461(.A1(new_n10430_), .A2(pi0038), .ZN(new_n10431_));
  AOI21_X1   g07462(.A1(new_n10429_), .A2(new_n3455_), .B(new_n10431_), .ZN(new_n10432_));
  NOR2_X1    g07463(.A1(new_n8511_), .A2(new_n8504_), .ZN(new_n10433_));
  NOR2_X1    g07464(.A1(new_n5524_), .A2(new_n2730_), .ZN(new_n10434_));
  OAI21_X1   g07465(.A1(new_n6523_), .A2(new_n10422_), .B(new_n10434_), .ZN(new_n10435_));
  NOR2_X1    g07466(.A1(new_n10425_), .A2(new_n3186_), .ZN(new_n10436_));
  NOR4_X1    g07467(.A1(new_n10427_), .A2(new_n3183_), .A3(new_n10422_), .A4(new_n10436_), .ZN(new_n10437_));
  OAI21_X1   g07468(.A1(new_n10433_), .A2(new_n10435_), .B(new_n10437_), .ZN(new_n10438_));
  NAND2_X1   g07469(.A1(new_n10438_), .A2(new_n3235_), .ZN(new_n10439_));
  NOR2_X1    g07470(.A1(new_n8482_), .A2(pi0228), .ZN(new_n10440_));
  AOI21_X1   g07471(.A1(new_n8612_), .A2(new_n10440_), .B(new_n3133_), .ZN(new_n10441_));
  NOR2_X1    g07472(.A1(new_n8911_), .A2(new_n8389_), .ZN(new_n10442_));
  OAI21_X1   g07473(.A1(new_n10441_), .A2(pi0039), .B(new_n10442_), .ZN(new_n10443_));
  NAND3_X1   g07474(.A1(new_n10430_), .A2(new_n3186_), .A3(new_n10425_), .ZN(new_n10444_));
  AOI21_X1   g07475(.A1(new_n10443_), .A2(new_n3171_), .B(new_n10444_), .ZN(new_n10445_));
  AOI21_X1   g07476(.A1(new_n10439_), .A2(new_n10445_), .B(new_n10432_), .ZN(new_n10446_));
  INV_X1     g07477(.I(new_n8714_), .ZN(new_n10447_));
  NOR3_X1    g07478(.A1(new_n10447_), .A2(po1038), .A3(new_n10422_), .ZN(new_n10449_));
  AOI21_X1   g07479(.A1(new_n10430_), .A2(new_n10449_), .B(new_n6399_), .ZN(new_n10450_));
  NOR3_X1    g07480(.A1(new_n10446_), .A2(new_n8474_), .A3(new_n10450_), .ZN(new_n10451_));
  OAI21_X1   g07481(.A1(new_n10418_), .A2(new_n10417_), .B(new_n10451_), .ZN(new_n10452_));
  AOI21_X1   g07482(.A1(new_n10410_), .A2(new_n10416_), .B(new_n10452_), .ZN(po0259));
  NOR3_X1    g07483(.A1(new_n2652_), .A2(new_n2448_), .A3(new_n10231_), .ZN(new_n10454_));
  INV_X1     g07484(.I(new_n10454_), .ZN(new_n10455_));
  NOR2_X1    g07485(.A1(new_n10235_), .A2(new_n10455_), .ZN(po0260));
  AOI21_X1   g07486(.A1(new_n5617_), .A2(pi0314), .B(pi0109), .ZN(new_n10457_));
  NOR3_X1    g07487(.A1(new_n2466_), .A2(pi0109), .A3(pi0314), .ZN(new_n10458_));
  NAND2_X1   g07488(.A1(new_n8291_), .A2(new_n9801_), .ZN(new_n10459_));
  NOR4_X1    g07489(.A1(new_n10265_), .A2(new_n10457_), .A3(new_n10458_), .A4(new_n10459_), .ZN(po0261));
  INV_X1     g07490(.I(new_n2987_), .ZN(new_n10461_));
  NAND4_X1   g07491(.A1(new_n10269_), .A2(new_n10461_), .A3(po1057), .A4(new_n6495_), .ZN(new_n10462_));
  NOR2_X1    g07492(.A1(new_n6531_), .A2(new_n2987_), .ZN(new_n10463_));
  NOR2_X1    g07493(.A1(new_n6403_), .A2(pi0047), .ZN(new_n10464_));
  AOI22_X1   g07494(.A1(new_n5413_), .A2(new_n2468_), .B1(new_n8529_), .B2(new_n10464_), .ZN(new_n10465_));
  NOR3_X1    g07495(.A1(new_n10465_), .A2(new_n2665_), .A3(new_n10268_), .ZN(new_n10466_));
  OAI21_X1   g07496(.A1(new_n10466_), .A2(new_n10463_), .B(po1057), .ZN(new_n10467_));
  NOR2_X1    g07497(.A1(new_n8530_), .A2(new_n8248_), .ZN(new_n10468_));
  AOI21_X1   g07498(.A1(new_n10468_), .A2(new_n10318_), .B(new_n6668_), .ZN(new_n10469_));
  AOI21_X1   g07499(.A1(new_n10467_), .A2(new_n10462_), .B(new_n10469_), .ZN(po0262));
  NOR2_X1    g07500(.A1(new_n2732_), .A2(pi0024), .ZN(new_n10471_));
  AOI21_X1   g07501(.A1(new_n2518_), .A2(new_n9143_), .B(new_n2899_), .ZN(new_n10472_));
  NOR2_X1    g07502(.A1(new_n10472_), .A2(new_n7272_), .ZN(new_n10473_));
  NAND3_X1   g07503(.A1(new_n9144_), .A2(pi0024), .A3(new_n2902_), .ZN(new_n10474_));
  XNOR2_X1   g07504(.A1(new_n10473_), .A2(new_n10474_), .ZN(new_n10475_));
  NAND3_X1   g07505(.A1(new_n10475_), .A2(pi0841), .A3(new_n9126_), .ZN(new_n10476_));
  OAI21_X1   g07506(.A1(new_n10476_), .A2(new_n10471_), .B(new_n8291_), .ZN(new_n10477_));
  AOI21_X1   g07507(.A1(new_n10471_), .A2(new_n10476_), .B(new_n10477_), .ZN(po0264));
  NOR3_X1    g07508(.A1(new_n9193_), .A2(pi0999), .A3(new_n8292_), .ZN(po0265));
  NAND2_X1   g07509(.A1(new_n6363_), .A2(new_n2461_), .ZN(new_n10480_));
  NAND4_X1   g07510(.A1(new_n10480_), .A2(pi0047), .A3(new_n2462_), .A4(new_n2468_), .ZN(new_n10481_));
  NOR3_X1    g07511(.A1(new_n10481_), .A2(new_n2525_), .A3(new_n7266_), .ZN(new_n10482_));
  NAND2_X1   g07512(.A1(new_n8362_), .A2(new_n6369_), .ZN(new_n10483_));
  NOR2_X1    g07513(.A1(new_n10482_), .A2(new_n10483_), .ZN(new_n10484_));
  NOR2_X1    g07514(.A1(new_n10483_), .A2(new_n9231_), .ZN(new_n10485_));
  XNOR2_X1   g07515(.A1(new_n10484_), .A2(new_n10485_), .ZN(new_n10486_));
  NOR3_X1    g07516(.A1(new_n10482_), .A2(pi0051), .A3(new_n6369_), .ZN(new_n10487_));
  NOR2_X1    g07517(.A1(new_n6411_), .A2(new_n3134_), .ZN(new_n10488_));
  NOR4_X1    g07518(.A1(new_n6366_), .A2(new_n3455_), .A3(new_n10488_), .A4(new_n8362_), .ZN(new_n10489_));
  OAI21_X1   g07519(.A1(new_n5498_), .A2(new_n7332_), .B(new_n10489_), .ZN(new_n10490_));
  NOR3_X1    g07520(.A1(new_n10486_), .A2(new_n10487_), .A3(new_n10490_), .ZN(po0266));
  NOR3_X1    g07521(.A1(new_n9436_), .A2(new_n9430_), .A3(new_n9253_), .ZN(po0267));
  NOR4_X1    g07522(.A1(new_n2465_), .A2(new_n9802_), .A3(new_n2664_), .A4(new_n2612_), .ZN(new_n10493_));
  NAND3_X1   g07523(.A1(new_n10258_), .A2(new_n2617_), .A3(new_n10493_), .ZN(new_n10494_));
  NOR2_X1    g07524(.A1(new_n9003_), .A2(new_n8248_), .ZN(new_n10495_));
  INV_X1     g07525(.I(new_n10495_), .ZN(new_n10496_));
  OAI21_X1   g07526(.A1(new_n10496_), .A2(new_n10494_), .B(new_n8291_), .ZN(new_n10497_));
  AOI21_X1   g07527(.A1(pi0314), .A2(new_n8463_), .B(new_n10497_), .ZN(po0268));
  NOR2_X1    g07528(.A1(new_n10494_), .A2(pi0314), .ZN(new_n10499_));
  INV_X1     g07529(.I(new_n10499_), .ZN(new_n10500_));
  NOR2_X1    g07530(.A1(new_n8507_), .A2(new_n10500_), .ZN(new_n10501_));
  NOR2_X1    g07531(.A1(new_n7422_), .A2(new_n2437_), .ZN(new_n10502_));
  NOR4_X1    g07532(.A1(new_n10501_), .A2(new_n3138_), .A3(new_n8288_), .A4(new_n10502_), .ZN(po0269));
  NAND2_X1   g07533(.A1(new_n9439_), .A2(pi0124), .ZN(po0270));
  NOR2_X1    g07534(.A1(new_n8494_), .A2(new_n2730_), .ZN(new_n10505_));
  INV_X1     g07535(.I(new_n10505_), .ZN(new_n10506_));
  NOR2_X1    g07536(.A1(new_n10506_), .A2(new_n5518_), .ZN(new_n10507_));
  NAND4_X1   g07537(.A1(new_n10507_), .A2(new_n8492_), .A3(pi0113), .A4(new_n5520_), .ZN(new_n10508_));
  AOI21_X1   g07538(.A1(new_n10505_), .A2(new_n8595_), .B(new_n5518_), .ZN(new_n10509_));
  NOR2_X1    g07539(.A1(new_n10509_), .A2(new_n3194_), .ZN(new_n10510_));
  AOI21_X1   g07540(.A1(new_n8670_), .A2(new_n10510_), .B(new_n6485_), .ZN(new_n10511_));
  OAI21_X1   g07541(.A1(new_n10511_), .A2(new_n10508_), .B(new_n3235_), .ZN(new_n10512_));
  NAND2_X1   g07542(.A1(new_n8595_), .A2(new_n3183_), .ZN(new_n10513_));
  NOR2_X1    g07543(.A1(new_n3187_), .A2(new_n10513_), .ZN(new_n10514_));
  AOI21_X1   g07544(.A1(new_n10512_), .A2(new_n10514_), .B(new_n7331_), .ZN(new_n10515_));
  NOR2_X1    g07545(.A1(new_n8416_), .A2(new_n2730_), .ZN(new_n10516_));
  NOR2_X1    g07546(.A1(new_n2730_), .A2(new_n10347_), .ZN(new_n10517_));
  XOR2_X1    g07547(.A1(new_n10516_), .A2(new_n10517_), .Z(new_n10518_));
  AOI21_X1   g07548(.A1(new_n10518_), .A2(new_n8429_), .B(pi0113), .ZN(new_n10519_));
  NOR3_X1    g07549(.A1(new_n10519_), .A2(new_n2437_), .A3(new_n5521_), .ZN(new_n10520_));
  NOR2_X1    g07550(.A1(new_n8789_), .A2(new_n5512_), .ZN(new_n10521_));
  OAI21_X1   g07551(.A1(new_n10520_), .A2(pi0228), .B(new_n10521_), .ZN(new_n10522_));
  NAND2_X1   g07552(.A1(new_n8597_), .A2(pi0113), .ZN(new_n10523_));
  NAND2_X1   g07553(.A1(pi0113), .A2(pi0228), .ZN(new_n10524_));
  XOR2_X1    g07554(.A1(new_n10523_), .A2(new_n10524_), .Z(new_n10525_));
  NAND2_X1   g07555(.A1(new_n10352_), .A2(new_n10525_), .ZN(new_n10526_));
  AOI21_X1   g07556(.A1(new_n10522_), .A2(new_n8883_), .B(new_n10526_), .ZN(new_n10527_));
  OR3_X2     g07557(.A1(new_n8614_), .A2(new_n6504_), .A3(new_n10509_), .Z(new_n10528_));
  NAND2_X1   g07558(.A1(new_n5505_), .A2(pi0039), .ZN(new_n10529_));
  AOI21_X1   g07559(.A1(new_n10528_), .A2(new_n10529_), .B(new_n10508_), .ZN(new_n10530_));
  NOR2_X1    g07560(.A1(new_n3214_), .A2(pi0113), .ZN(new_n10531_));
  AOI21_X1   g07561(.A1(new_n10374_), .A2(new_n10531_), .B(new_n8595_), .ZN(new_n10532_));
  NOR2_X1    g07562(.A1(new_n8657_), .A2(new_n10532_), .ZN(new_n10533_));
  NOR3_X1    g07563(.A1(new_n10513_), .A2(new_n3235_), .A3(new_n3133_), .ZN(new_n10534_));
  AOI21_X1   g07564(.A1(new_n10533_), .A2(new_n10534_), .B(pi0087), .ZN(new_n10535_));
  NOR4_X1    g07565(.A1(new_n10535_), .A2(new_n3259_), .A3(new_n7331_), .A4(new_n10513_), .ZN(new_n10536_));
  OAI21_X1   g07566(.A1(new_n10527_), .A2(new_n10530_), .B(new_n10536_), .ZN(new_n10537_));
  XNOR2_X1   g07567(.A1(new_n10537_), .A2(new_n10515_), .ZN(po0271));
  OAI21_X1   g07568(.A1(new_n8673_), .A2(new_n9028_), .B(pi0114), .ZN(new_n10539_));
  OAI21_X1   g07569(.A1(new_n8760_), .A2(new_n10539_), .B(new_n3194_), .ZN(new_n10540_));
  INV_X1     g07570(.I(new_n9028_), .ZN(new_n10541_));
  NOR2_X1    g07571(.A1(new_n5513_), .A2(pi0072), .ZN(new_n10542_));
  INV_X1     g07572(.I(new_n10542_), .ZN(new_n10543_));
  NOR2_X1    g07573(.A1(new_n10541_), .A2(new_n10543_), .ZN(new_n10544_));
  AOI21_X1   g07574(.A1(new_n10540_), .A2(new_n10544_), .B(pi0075), .ZN(new_n10545_));
  NOR2_X1    g07575(.A1(new_n10543_), .A2(pi0039), .ZN(new_n10546_));
  NAND2_X1   g07576(.A1(new_n10546_), .A2(new_n3186_), .ZN(new_n10547_));
  OAI21_X1   g07577(.A1(new_n10545_), .A2(new_n10547_), .B(new_n7332_), .ZN(new_n10548_));
  NOR2_X1    g07578(.A1(new_n8786_), .A2(new_n5513_), .ZN(new_n10549_));
  OAI21_X1   g07579(.A1(new_n8791_), .A2(pi0114), .B(pi0115), .ZN(new_n10550_));
  NOR2_X1    g07580(.A1(new_n10550_), .A2(new_n10549_), .ZN(new_n10551_));
  NAND2_X1   g07581(.A1(pi0039), .A2(pi0115), .ZN(new_n10552_));
  XNOR2_X1   g07582(.A1(new_n10551_), .A2(new_n10552_), .ZN(new_n10553_));
  INV_X1     g07583(.I(new_n8616_), .ZN(new_n10554_));
  AOI22_X1   g07584(.A1(new_n8615_), .A2(pi0228), .B1(new_n3132_), .B2(new_n10542_), .ZN(new_n10555_));
  NOR2_X1    g07585(.A1(new_n10546_), .A2(new_n3132_), .ZN(new_n10556_));
  NOR2_X1    g07586(.A1(new_n9045_), .A2(new_n3455_), .ZN(new_n10557_));
  NAND2_X1   g07587(.A1(new_n10557_), .A2(pi0075), .ZN(new_n10558_));
  OAI22_X1   g07588(.A1(new_n10555_), .A2(new_n5514_), .B1(new_n10556_), .B2(new_n10558_), .ZN(new_n10559_));
  OAI21_X1   g07589(.A1(new_n9028_), .A2(new_n10542_), .B(new_n3183_), .ZN(new_n10560_));
  NAND3_X1   g07590(.A1(new_n3259_), .A2(new_n3455_), .A3(pi0100), .ZN(new_n10561_));
  NAND2_X1   g07591(.A1(new_n10560_), .A2(new_n10561_), .ZN(new_n10562_));
  NAND3_X1   g07592(.A1(new_n10562_), .A2(pi0114), .A3(new_n8660_), .ZN(new_n10563_));
  AOI21_X1   g07593(.A1(new_n8623_), .A2(new_n10541_), .B(new_n10563_), .ZN(new_n10564_));
  NAND3_X1   g07594(.A1(new_n10559_), .A2(new_n10554_), .A3(new_n10564_), .ZN(new_n10565_));
  NAND2_X1   g07595(.A1(new_n10565_), .A2(new_n3133_), .ZN(new_n10566_));
  NOR2_X1    g07596(.A1(new_n10543_), .A2(pi0039), .ZN(new_n10567_));
  NAND4_X1   g07597(.A1(new_n10553_), .A2(new_n7332_), .A3(new_n10566_), .A4(new_n10567_), .ZN(new_n10568_));
  XOR2_X1    g07598(.A1(new_n10568_), .A2(new_n10548_), .Z(po0272));
  OAI21_X1   g07599(.A1(pi0072), .A2(new_n5514_), .B(new_n10506_), .ZN(new_n10570_));
  NAND2_X1   g07600(.A1(new_n8759_), .A2(pi0115), .ZN(new_n10571_));
  NAND2_X1   g07601(.A1(new_n9027_), .A2(pi0052), .ZN(new_n10572_));
  AOI21_X1   g07602(.A1(new_n8620_), .A2(new_n5514_), .B(new_n10572_), .ZN(new_n10573_));
  AOI21_X1   g07603(.A1(new_n10573_), .A2(new_n6485_), .B(new_n10506_), .ZN(new_n10574_));
  NOR4_X1    g07604(.A1(new_n3186_), .A2(pi0039), .A3(pi0072), .A4(new_n5514_), .ZN(new_n10575_));
  OAI21_X1   g07605(.A1(new_n10575_), .A2(new_n3235_), .B(new_n3194_), .ZN(new_n10576_));
  AOI21_X1   g07606(.A1(new_n10571_), .A2(new_n10574_), .B(new_n10576_), .ZN(new_n10577_));
  OAI21_X1   g07607(.A1(new_n10577_), .A2(new_n10570_), .B(new_n7332_), .ZN(new_n10578_));
  NAND2_X1   g07608(.A1(new_n8786_), .A2(pi0115), .ZN(new_n10579_));
  XNOR2_X1   g07609(.A1(new_n10579_), .A2(new_n10552_), .ZN(new_n10580_));
  NAND4_X1   g07610(.A1(new_n3132_), .A2(new_n3183_), .A3(new_n2437_), .A4(pi0115), .ZN(new_n10581_));
  NOR4_X1    g07611(.A1(new_n8791_), .A2(new_n7331_), .A3(new_n10580_), .A4(new_n10581_), .ZN(new_n10582_));
  XNOR2_X1   g07612(.A1(new_n10582_), .A2(new_n10578_), .ZN(po0273));
  NAND2_X1   g07613(.A1(new_n8670_), .A2(new_n5512_), .ZN(new_n10584_));
  AOI22_X1   g07614(.A1(new_n10584_), .A2(new_n8566_), .B1(new_n6485_), .B2(new_n8621_), .ZN(new_n10585_));
  NAND2_X1   g07615(.A1(new_n10507_), .A2(new_n3193_), .ZN(new_n10586_));
  OAI21_X1   g07616(.A1(new_n10585_), .A2(new_n10586_), .B(new_n8567_), .ZN(new_n10587_));
  AOI21_X1   g07617(.A1(new_n10587_), .A2(new_n10505_), .B(pi0075), .ZN(new_n10588_));
  NOR2_X1    g07618(.A1(new_n8567_), .A2(pi0039), .ZN(new_n10589_));
  NAND2_X1   g07619(.A1(new_n10589_), .A2(new_n3186_), .ZN(new_n10590_));
  OAI21_X1   g07620(.A1(new_n10588_), .A2(new_n10590_), .B(new_n7332_), .ZN(new_n10591_));
  INV_X1     g07621(.I(new_n8598_), .ZN(new_n10592_));
  AOI21_X1   g07622(.A1(new_n2729_), .A2(new_n8582_), .B(pi0116), .ZN(new_n10593_));
  OAI21_X1   g07623(.A1(new_n10593_), .A2(new_n8570_), .B(new_n3005_), .ZN(new_n10594_));
  NOR3_X1    g07624(.A1(new_n8434_), .A2(new_n2730_), .A3(new_n8576_), .ZN(new_n10595_));
  AOI21_X1   g07625(.A1(new_n10595_), .A2(new_n10594_), .B(new_n8884_), .ZN(new_n10596_));
  NAND2_X1   g07626(.A1(new_n8659_), .A2(pi0038), .ZN(new_n10597_));
  NOR2_X1    g07627(.A1(new_n8657_), .A2(pi0113), .ZN(new_n10598_));
  NOR4_X1    g07628(.A1(new_n10598_), .A2(new_n3259_), .A3(pi0039), .A4(new_n8567_), .ZN(new_n10599_));
  OR2_X2     g07629(.A1(new_n10599_), .A2(new_n10597_), .Z(new_n10600_));
  NAND2_X1   g07630(.A1(new_n10599_), .A2(new_n10597_), .ZN(new_n10601_));
  NAND3_X1   g07631(.A1(new_n10600_), .A2(new_n10601_), .A3(new_n10557_), .ZN(new_n10602_));
  NAND2_X1   g07632(.A1(pi0087), .A2(pi0100), .ZN(new_n10603_));
  XOR2_X1    g07633(.A1(new_n10602_), .A2(new_n10603_), .Z(new_n10604_));
  AOI21_X1   g07634(.A1(new_n10604_), .A2(new_n10589_), .B(pi0075), .ZN(new_n10605_));
  OAI22_X1   g07635(.A1(new_n8614_), .A2(new_n6504_), .B1(new_n8567_), .B2(new_n8620_), .ZN(new_n10606_));
  NAND4_X1   g07636(.A1(new_n10606_), .A2(pi0113), .A3(new_n8566_), .A4(new_n10505_), .ZN(new_n10607_));
  XOR2_X1    g07637(.A1(new_n10607_), .A2(new_n10507_), .Z(new_n10608_));
  NAND3_X1   g07638(.A1(new_n3259_), .A2(new_n3455_), .A3(pi0100), .ZN(new_n10609_));
  NAND2_X1   g07639(.A1(new_n10609_), .A2(new_n3183_), .ZN(new_n10610_));
  NAND4_X1   g07640(.A1(new_n7332_), .A2(pi0116), .A3(new_n10589_), .A4(new_n10610_), .ZN(new_n10611_));
  NOR2_X1    g07641(.A1(new_n10608_), .A2(new_n10611_), .ZN(new_n10612_));
  OAI21_X1   g07642(.A1(new_n8601_), .A2(pi0228), .B(new_n10612_), .ZN(new_n10613_));
  NOR4_X1    g07643(.A1(new_n10605_), .A2(new_n10592_), .A3(new_n10596_), .A4(new_n10613_), .ZN(new_n10614_));
  XNOR2_X1   g07644(.A1(new_n10614_), .A2(new_n10591_), .ZN(po0274));
  NOR2_X1    g07645(.A1(new_n5488_), .A2(new_n3258_), .ZN(new_n10616_));
  NAND3_X1   g07646(.A1(new_n3461_), .A2(pi0100), .A3(new_n6306_), .ZN(new_n10617_));
  AND2_X2    g07647(.A1(new_n10617_), .A2(new_n3617_), .Z(new_n10618_));
  INV_X1     g07648(.I(new_n5498_), .ZN(new_n10619_));
  OAI22_X1   g07649(.A1(new_n10617_), .A2(new_n3617_), .B1(new_n3455_), .B2(new_n10619_), .ZN(new_n10620_));
  NOR2_X1    g07650(.A1(new_n6289_), .A2(pi0054), .ZN(new_n10621_));
  INV_X1     g07651(.I(new_n10621_), .ZN(new_n10622_));
  NAND4_X1   g07652(.A1(new_n3207_), .A2(pi0038), .A3(pi0055), .A4(pi0092), .ZN(new_n10623_));
  AOI21_X1   g07653(.A1(new_n10622_), .A2(new_n3175_), .B(new_n10623_), .ZN(new_n10624_));
  OAI21_X1   g07654(.A1(new_n10618_), .A2(new_n10620_), .B(new_n10624_), .ZN(new_n10625_));
  XOR2_X1    g07655(.A1(new_n10625_), .A2(new_n10616_), .Z(new_n10626_));
  NOR4_X1    g07656(.A1(new_n10626_), .A2(new_n5497_), .A3(new_n5544_), .A4(new_n8226_), .ZN(po0275));
  NOR3_X1    g07657(.A1(new_n9513_), .A2(new_n8108_), .A3(new_n5665_), .ZN(new_n10628_));
  INV_X1     g07658(.I(pi0150), .ZN(new_n10629_));
  NOR3_X1    g07659(.A1(new_n10628_), .A2(new_n9456_), .A3(new_n5386_), .ZN(new_n10631_));
  NOR2_X1    g07660(.A1(new_n10631_), .A2(new_n5551_), .ZN(new_n10632_));
  NOR3_X1    g07661(.A1(new_n3230_), .A2(new_n7537_), .A3(pi0165), .ZN(new_n10633_));
  NOR2_X1    g07662(.A1(new_n6494_), .A2(new_n10633_), .ZN(new_n10634_));
  NAND3_X1   g07663(.A1(new_n10632_), .A2(new_n7537_), .A3(new_n10634_), .ZN(new_n10635_));
  INV_X1     g07664(.I(new_n10632_), .ZN(new_n10636_));
  NAND3_X1   g07665(.A1(new_n10636_), .A2(new_n7538_), .A3(new_n10634_), .ZN(new_n10637_));
  AOI21_X1   g07666(.A1(new_n10637_), .A2(new_n10635_), .B(new_n3175_), .ZN(new_n10638_));
  INV_X1     g07667(.I(new_n10638_), .ZN(new_n10639_));
  INV_X1     g07668(.I(pi0165), .ZN(new_n10640_));
  OAI22_X1   g07669(.A1(new_n6494_), .A2(new_n3259_), .B1(new_n3115_), .B2(new_n10640_), .ZN(new_n10641_));
  NAND3_X1   g07670(.A1(new_n10632_), .A2(pi0074), .A3(new_n7537_), .ZN(new_n10642_));
  NAND3_X1   g07671(.A1(new_n10636_), .A2(new_n3175_), .A3(new_n7537_), .ZN(new_n10643_));
  NAND2_X1   g07672(.A1(new_n10643_), .A2(new_n10642_), .ZN(new_n10644_));
  NAND2_X1   g07673(.A1(new_n10644_), .A2(new_n10641_), .ZN(new_n10645_));
  INV_X1     g07674(.I(new_n10645_), .ZN(new_n10646_));
  NOR2_X1    g07675(.A1(new_n10636_), .A2(new_n7537_), .ZN(new_n10647_));
  NOR2_X1    g07676(.A1(new_n10647_), .A2(new_n3175_), .ZN(new_n10648_));
  OAI21_X1   g07677(.A1(new_n7328_), .A2(new_n10648_), .B(new_n10646_), .ZN(new_n10649_));
  INV_X1     g07678(.I(new_n10649_), .ZN(new_n10650_));
  NAND3_X1   g07679(.A1(new_n5699_), .A2(new_n5400_), .A3(new_n9606_), .ZN(new_n10651_));
  NOR2_X1    g07680(.A1(new_n9241_), .A2(pi0232), .ZN(new_n10652_));
  AOI21_X1   g07681(.A1(new_n5698_), .A2(new_n10652_), .B(new_n5460_), .ZN(new_n10653_));
  AOI21_X1   g07682(.A1(new_n10651_), .A2(new_n10653_), .B(new_n3183_), .ZN(new_n10654_));
  AOI21_X1   g07683(.A1(pi0190), .A2(new_n7374_), .B(new_n7387_), .ZN(new_n10655_));
  INV_X1     g07684(.I(pi0190), .ZN(new_n10656_));
  NAND2_X1   g07685(.A1(new_n7349_), .A2(pi0173), .ZN(new_n10657_));
  AOI21_X1   g07686(.A1(new_n7397_), .A2(new_n10656_), .B(new_n10657_), .ZN(new_n10658_));
  INV_X1     g07687(.I(pi0185), .ZN(new_n10659_));
  NAND3_X1   g07688(.A1(new_n7419_), .A2(new_n10659_), .A3(new_n10656_), .ZN(new_n10660_));
  NAND2_X1   g07689(.A1(new_n5386_), .A2(new_n10656_), .ZN(new_n10661_));
  AOI21_X1   g07690(.A1(new_n10660_), .A2(pi0173), .B(new_n10661_), .ZN(new_n10662_));
  NAND3_X1   g07691(.A1(new_n7413_), .A2(pi0173), .A3(new_n3137_), .ZN(new_n10663_));
  INV_X1     g07692(.I(pi0173), .ZN(new_n10664_));
  NAND3_X1   g07693(.A1(new_n7414_), .A2(new_n10664_), .A3(new_n3137_), .ZN(new_n10665_));
  NAND2_X1   g07694(.A1(new_n10665_), .A2(new_n10663_), .ZN(new_n10666_));
  NAND2_X1   g07695(.A1(new_n10666_), .A2(new_n7423_), .ZN(new_n10667_));
  OAI21_X1   g07696(.A1(new_n10662_), .A2(new_n10667_), .B(new_n10659_), .ZN(new_n10668_));
  OAI21_X1   g07697(.A1(new_n10668_), .A2(new_n10658_), .B(pi0173), .ZN(new_n10669_));
  OAI21_X1   g07698(.A1(new_n10655_), .A2(new_n10669_), .B(new_n3098_), .ZN(new_n10670_));
  NOR3_X1    g07699(.A1(new_n7392_), .A2(new_n5386_), .A3(new_n7387_), .ZN(new_n10671_));
  AOI21_X1   g07700(.A1(new_n7387_), .A2(new_n5373_), .B(pi0210), .ZN(new_n10672_));
  OAI21_X1   g07701(.A1(new_n10672_), .A2(new_n7390_), .B(new_n3098_), .ZN(new_n10673_));
  AOI21_X1   g07702(.A1(new_n10671_), .A2(new_n10670_), .B(new_n10673_), .ZN(new_n10674_));
  OAI21_X1   g07703(.A1(new_n7470_), .A2(new_n4635_), .B(new_n7386_), .ZN(new_n10675_));
  AOI21_X1   g07704(.A1(new_n10675_), .A2(pi0151), .B(new_n10629_), .ZN(new_n10676_));
  NOR4_X1    g07705(.A1(new_n7407_), .A2(new_n3538_), .A3(new_n4635_), .A4(new_n5423_), .ZN(new_n10677_));
  NAND2_X1   g07706(.A1(new_n7424_), .A2(new_n3538_), .ZN(new_n10678_));
  OAI21_X1   g07707(.A1(new_n10677_), .A2(new_n10678_), .B(pi0168), .ZN(new_n10679_));
  NOR2_X1    g07708(.A1(new_n5386_), .A2(new_n4635_), .ZN(new_n10680_));
  INV_X1     g07709(.I(new_n10680_), .ZN(new_n10681_));
  OAI21_X1   g07710(.A1(new_n7473_), .A2(new_n10681_), .B(new_n7395_), .ZN(new_n10682_));
  NOR4_X1    g07711(.A1(new_n7403_), .A2(pi0040), .A3(new_n10629_), .A4(new_n3538_), .ZN(new_n10683_));
  NAND3_X1   g07712(.A1(new_n10682_), .A2(new_n10679_), .A3(new_n10683_), .ZN(new_n10684_));
  XOR2_X1    g07713(.A1(new_n10676_), .A2(new_n10684_), .Z(new_n10685_));
  NOR2_X1    g07714(.A1(new_n7387_), .A2(pi0232), .ZN(new_n10686_));
  NAND2_X1   g07715(.A1(new_n7391_), .A2(new_n5469_), .ZN(new_n10687_));
  OAI21_X1   g07716(.A1(new_n10687_), .A2(new_n10686_), .B(new_n3183_), .ZN(new_n10688_));
  NAND3_X1   g07717(.A1(new_n10688_), .A2(pi0038), .A3(pi0232), .ZN(new_n10689_));
  NOR3_X1    g07718(.A1(new_n10674_), .A2(new_n10689_), .A3(new_n10685_), .ZN(new_n10690_));
  NOR2_X1    g07719(.A1(new_n5699_), .A2(new_n6448_), .ZN(new_n10691_));
  INV_X1     g07720(.I(pi0157), .ZN(new_n10692_));
  NOR2_X1    g07721(.A1(new_n7446_), .A2(new_n10692_), .ZN(new_n10693_));
  INV_X1     g07722(.I(new_n7445_), .ZN(new_n10694_));
  NOR3_X1    g07723(.A1(new_n10694_), .A2(new_n10692_), .A3(new_n4635_), .ZN(new_n10695_));
  XOR2_X1    g07724(.A1(new_n10693_), .A2(new_n10695_), .Z(new_n10696_));
  NAND2_X1   g07725(.A1(new_n10696_), .A2(pi0168), .ZN(new_n10697_));
  AOI21_X1   g07726(.A1(new_n10697_), .A2(new_n7443_), .B(new_n10692_), .ZN(new_n10698_));
  OAI21_X1   g07727(.A1(new_n10698_), .A2(new_n10691_), .B(new_n9241_), .ZN(new_n10699_));
  XOR2_X1    g07728(.A1(new_n10632_), .A2(new_n5912_), .Z(new_n10700_));
  NAND2_X1   g07729(.A1(new_n5373_), .A2(pi0185), .ZN(new_n10701_));
  XOR2_X1    g07730(.A1(new_n10701_), .A2(pi0184), .Z(new_n10702_));
  NOR2_X1    g07731(.A1(new_n10702_), .A2(new_n9522_), .ZN(new_n10703_));
  NAND2_X1   g07732(.A1(new_n10700_), .A2(new_n10703_), .ZN(new_n10704_));
  NAND2_X1   g07733(.A1(new_n10704_), .A2(pi0054), .ZN(new_n10705_));
  XNOR2_X1   g07734(.A1(new_n10705_), .A2(new_n9560_), .ZN(new_n10706_));
  NAND3_X1   g07735(.A1(new_n6493_), .A2(pi0143), .A3(pi0299), .ZN(new_n10707_));
  INV_X1     g07736(.I(pi0143), .ZN(new_n10708_));
  NAND3_X1   g07737(.A1(new_n6493_), .A2(new_n10708_), .A3(new_n3098_), .ZN(new_n10709_));
  AOI21_X1   g07738(.A1(new_n10709_), .A2(new_n10707_), .B(new_n10640_), .ZN(new_n10710_));
  NAND2_X1   g07739(.A1(new_n10710_), .A2(pi0074), .ZN(new_n10711_));
  OAI21_X1   g07740(.A1(new_n10706_), .A2(new_n10711_), .B(new_n3115_), .ZN(new_n10712_));
  INV_X1     g07741(.I(new_n10704_), .ZN(new_n10713_));
  NOR2_X1    g07742(.A1(new_n10713_), .A2(new_n3235_), .ZN(new_n10714_));
  OAI21_X1   g07743(.A1(new_n10710_), .A2(new_n3259_), .B(new_n3462_), .ZN(new_n10715_));
  NOR2_X1    g07744(.A1(new_n10713_), .A2(new_n3462_), .ZN(new_n10716_));
  INV_X1     g07745(.I(new_n10716_), .ZN(new_n10717_));
  OAI21_X1   g07746(.A1(new_n10717_), .A2(new_n7529_), .B(new_n10715_), .ZN(new_n10718_));
  NAND3_X1   g07747(.A1(new_n6493_), .A2(pi0157), .A3(pi0299), .ZN(new_n10719_));
  NAND3_X1   g07748(.A1(new_n6493_), .A2(new_n10692_), .A3(new_n3098_), .ZN(new_n10720_));
  AOI21_X1   g07749(.A1(new_n10719_), .A2(new_n10720_), .B(new_n7510_), .ZN(new_n10721_));
  NOR3_X1    g07750(.A1(new_n3145_), .A2(new_n7334_), .A3(new_n10721_), .ZN(new_n10722_));
  AOI21_X1   g07751(.A1(new_n10718_), .A2(new_n10722_), .B(new_n10714_), .ZN(new_n10723_));
  NAND3_X1   g07752(.A1(new_n7494_), .A2(pi0143), .A3(pi0165), .ZN(new_n10724_));
  OR3_X2     g07753(.A1(new_n7494_), .A2(pi0143), .A3(new_n10640_), .Z(new_n10725_));
  AOI21_X1   g07754(.A1(new_n10725_), .A2(new_n10724_), .B(new_n8001_), .ZN(new_n10726_));
  NAND3_X1   g07755(.A1(new_n7500_), .A2(new_n3259_), .A3(new_n10708_), .ZN(new_n10727_));
  NAND2_X1   g07756(.A1(new_n10727_), .A2(pi0165), .ZN(new_n10728_));
  OAI21_X1   g07757(.A1(new_n10726_), .A2(new_n10728_), .B(new_n3184_), .ZN(new_n10729_));
  NOR2_X1    g07758(.A1(new_n10729_), .A2(new_n10723_), .ZN(new_n10730_));
  NAND4_X1   g07759(.A1(new_n7441_), .A2(pi0178), .A3(new_n5373_), .A4(new_n5398_), .ZN(new_n10731_));
  OAI21_X1   g07760(.A1(new_n5689_), .A2(new_n7449_), .B(pi0178), .ZN(new_n10732_));
  NOR2_X1    g07761(.A1(new_n10691_), .A2(new_n10732_), .ZN(new_n10733_));
  OAI21_X1   g07762(.A1(new_n7510_), .A2(new_n10656_), .B(new_n5698_), .ZN(new_n10734_));
  NAND3_X1   g07763(.A1(new_n10734_), .A2(pi0190), .A3(new_n5400_), .ZN(new_n10735_));
  OAI21_X1   g07764(.A1(new_n10733_), .A2(new_n10735_), .B(new_n10731_), .ZN(new_n10736_));
  NOR2_X1    g07765(.A1(new_n6494_), .A2(new_n10629_), .ZN(new_n10737_));
  NAND4_X1   g07766(.A1(new_n10737_), .A2(new_n7333_), .A3(pi0092), .A4(new_n7537_), .ZN(new_n10738_));
  NAND3_X1   g07767(.A1(new_n10738_), .A2(new_n3115_), .A3(new_n10640_), .ZN(new_n10739_));
  NAND3_X1   g07768(.A1(new_n10739_), .A2(new_n3160_), .A3(new_n6493_), .ZN(new_n10740_));
  NAND2_X1   g07769(.A1(new_n10646_), .A2(new_n10740_), .ZN(new_n10741_));
  NOR2_X1    g07770(.A1(new_n10648_), .A2(new_n3258_), .ZN(new_n10742_));
  AOI21_X1   g07771(.A1(new_n10741_), .A2(new_n10742_), .B(new_n3225_), .ZN(new_n10743_));
  NAND3_X1   g07772(.A1(new_n10710_), .A2(pi0038), .A3(new_n3185_), .ZN(new_n10744_));
  NAND2_X1   g07773(.A1(new_n10717_), .A2(new_n10744_), .ZN(new_n10745_));
  AOI21_X1   g07774(.A1(new_n10704_), .A2(new_n6328_), .B(new_n7538_), .ZN(new_n10746_));
  NAND4_X1   g07775(.A1(new_n10745_), .A2(new_n3188_), .A3(new_n10297_), .A4(new_n10746_), .ZN(new_n10747_));
  NOR4_X1    g07776(.A1(new_n5699_), .A2(new_n10747_), .A3(new_n6448_), .A4(new_n10743_), .ZN(new_n10748_));
  NAND4_X1   g07777(.A1(new_n10736_), .A2(new_n10712_), .A3(new_n10730_), .A4(new_n10748_), .ZN(new_n10749_));
  AOI21_X1   g07778(.A1(new_n10699_), .A2(new_n5551_), .B(new_n10749_), .ZN(new_n10750_));
  OAI21_X1   g07779(.A1(new_n10690_), .A2(new_n10654_), .B(new_n10750_), .ZN(new_n10751_));
  NAND2_X1   g07780(.A1(new_n10751_), .A2(new_n10650_), .ZN(new_n10752_));
  NAND2_X1   g07781(.A1(new_n10752_), .A2(new_n10639_), .ZN(new_n10753_));
  INV_X1     g07782(.I(new_n8104_), .ZN(new_n10754_));
  NAND2_X1   g07783(.A1(new_n3538_), .A2(new_n4635_), .ZN(new_n10755_));
  NOR3_X1    g07784(.A1(new_n7676_), .A2(new_n10664_), .A3(new_n5386_), .ZN(new_n10756_));
  NOR3_X1    g07785(.A1(new_n7675_), .A2(new_n10664_), .A3(new_n5373_), .ZN(new_n10757_));
  OAI21_X1   g07786(.A1(new_n10756_), .A2(new_n10757_), .B(new_n7748_), .ZN(new_n10758_));
  NOR2_X1    g07787(.A1(new_n7577_), .A2(new_n5386_), .ZN(new_n10759_));
  INV_X1     g07788(.I(new_n7748_), .ZN(new_n10760_));
  NOR2_X1    g07789(.A1(new_n10760_), .A2(new_n5373_), .ZN(new_n10761_));
  OAI21_X1   g07790(.A1(new_n10761_), .A2(new_n10759_), .B(new_n10664_), .ZN(new_n10762_));
  NOR2_X1    g07791(.A1(new_n5386_), .A2(new_n10664_), .ZN(new_n10763_));
  NOR2_X1    g07792(.A1(new_n7760_), .A2(new_n5386_), .ZN(new_n10764_));
  XOR2_X1    g07793(.A1(new_n10764_), .A2(new_n10763_), .Z(new_n10765_));
  NAND2_X1   g07794(.A1(new_n10765_), .A2(new_n8131_), .ZN(new_n10766_));
  NOR2_X1    g07795(.A1(new_n10761_), .A2(new_n10659_), .ZN(new_n10767_));
  NOR2_X1    g07796(.A1(pi0190), .A2(pi0299), .ZN(new_n10768_));
  INV_X1     g07797(.I(new_n10768_), .ZN(new_n10769_));
  AOI21_X1   g07798(.A1(new_n10766_), .A2(new_n10767_), .B(new_n10769_), .ZN(new_n10770_));
  NOR2_X1    g07799(.A1(new_n7748_), .A2(new_n5373_), .ZN(new_n10771_));
  NOR2_X1    g07800(.A1(new_n7806_), .A2(new_n10771_), .ZN(new_n10772_));
  NOR2_X1    g07801(.A1(new_n10772_), .A2(new_n10664_), .ZN(new_n10773_));
  NOR2_X1    g07802(.A1(new_n10664_), .A2(new_n10659_), .ZN(new_n10774_));
  XOR2_X1    g07803(.A1(new_n10773_), .A2(new_n10774_), .Z(new_n10775_));
  NAND2_X1   g07804(.A1(new_n10775_), .A2(new_n7748_), .ZN(new_n10776_));
  NOR2_X1    g07805(.A1(new_n7819_), .A2(new_n10771_), .ZN(new_n10777_));
  OAI21_X1   g07806(.A1(new_n10761_), .A2(new_n7768_), .B(pi0173), .ZN(new_n10778_));
  XNOR2_X1   g07807(.A1(new_n10778_), .A2(new_n10774_), .ZN(new_n10779_));
  AOI21_X1   g07808(.A1(new_n10779_), .A2(new_n10777_), .B(pi0190), .ZN(new_n10780_));
  OAI21_X1   g07809(.A1(new_n10770_), .A2(new_n10776_), .B(new_n10780_), .ZN(new_n10781_));
  NAND4_X1   g07810(.A1(new_n10781_), .A2(pi0185), .A3(new_n10758_), .A4(new_n10762_), .ZN(new_n10782_));
  NAND2_X1   g07811(.A1(new_n10782_), .A2(new_n5551_), .ZN(new_n10783_));
  NOR2_X1    g07812(.A1(new_n7776_), .A2(new_n5386_), .ZN(new_n10784_));
  NOR2_X1    g07813(.A1(new_n3538_), .A2(new_n4635_), .ZN(new_n10785_));
  OAI21_X1   g07814(.A1(new_n10760_), .A2(new_n5373_), .B(new_n10785_), .ZN(new_n10786_));
  OAI21_X1   g07815(.A1(new_n10784_), .A2(new_n10786_), .B(new_n10629_), .ZN(new_n10787_));
  NOR2_X1    g07816(.A1(new_n10772_), .A2(new_n3538_), .ZN(new_n10788_));
  XOR2_X1    g07817(.A1(new_n10788_), .A2(new_n10785_), .Z(new_n10789_));
  NAND2_X1   g07818(.A1(new_n10629_), .A2(new_n3098_), .ZN(new_n10790_));
  AOI21_X1   g07819(.A1(new_n10789_), .A2(new_n10777_), .B(new_n10790_), .ZN(new_n10791_));
  NOR2_X1    g07820(.A1(new_n7767_), .A2(new_n4635_), .ZN(new_n10792_));
  NAND4_X1   g07821(.A1(new_n7748_), .A2(new_n3538_), .A3(new_n5386_), .A4(new_n10680_), .ZN(new_n10793_));
  NOR4_X1    g07822(.A1(new_n7857_), .A2(new_n10791_), .A3(new_n10792_), .A4(new_n10793_), .ZN(new_n10794_));
  NAND4_X1   g07823(.A1(new_n10783_), .A2(new_n10755_), .A3(new_n10787_), .A4(new_n10794_), .ZN(new_n10795_));
  NAND2_X1   g07824(.A1(new_n10795_), .A2(new_n3183_), .ZN(new_n10796_));
  NAND3_X1   g07825(.A1(new_n10796_), .A2(pi0232), .A3(new_n7748_), .ZN(new_n10797_));
  NAND3_X1   g07826(.A1(new_n10797_), .A2(new_n3259_), .A3(new_n10729_), .ZN(new_n10798_));
  OAI22_X1   g07827(.A1(new_n7591_), .A2(new_n7633_), .B1(new_n10692_), .B2(new_n4635_), .ZN(new_n10799_));
  NOR3_X1    g07828(.A1(new_n5455_), .A2(new_n5386_), .A3(new_n7440_), .ZN(new_n10800_));
  AOI21_X1   g07829(.A1(new_n10799_), .A2(new_n10800_), .B(new_n7577_), .ZN(new_n10801_));
  NOR2_X1    g07830(.A1(new_n7577_), .A2(new_n3098_), .ZN(new_n10802_));
  XOR2_X1    g07831(.A1(new_n10801_), .A2(new_n10802_), .Z(new_n10803_));
  AOI21_X1   g07832(.A1(new_n5398_), .A2(new_n7577_), .B(new_n7451_), .ZN(new_n10804_));
  NOR2_X1    g07833(.A1(new_n7596_), .A2(pi0299), .ZN(new_n10805_));
  NAND2_X1   g07834(.A1(new_n10805_), .A2(pi0190), .ZN(new_n10806_));
  NOR2_X1    g07835(.A1(new_n10804_), .A2(pi0178), .ZN(new_n10807_));
  AOI21_X1   g07836(.A1(new_n10807_), .A2(new_n10806_), .B(new_n5551_), .ZN(new_n10808_));
  AOI22_X1   g07837(.A1(new_n7623_), .A2(new_n10808_), .B1(new_n7510_), .B2(new_n10804_), .ZN(new_n10809_));
  OAI21_X1   g07838(.A1(new_n7577_), .A2(pi0232), .B(pi0039), .ZN(new_n10810_));
  NOR4_X1    g07839(.A1(new_n10809_), .A2(new_n7591_), .A3(new_n7592_), .A4(new_n10810_), .ZN(new_n10811_));
  AOI21_X1   g07840(.A1(new_n10803_), .A2(pi0178), .B(new_n10811_), .ZN(new_n10812_));
  INV_X1     g07841(.I(new_n10647_), .ZN(new_n10813_));
  NOR3_X1    g07842(.A1(new_n7577_), .A2(pi0038), .A3(pi0054), .ZN(new_n10814_));
  OR3_X2     g07843(.A1(new_n7933_), .A2(new_n10737_), .A3(new_n10814_), .Z(new_n10815_));
  AOI21_X1   g07844(.A1(new_n10815_), .A2(pi0092), .B(new_n10641_), .ZN(new_n10816_));
  OAI22_X1   g07845(.A1(new_n10816_), .A2(new_n7538_), .B1(new_n3258_), .B2(new_n10813_), .ZN(new_n10817_));
  AOI21_X1   g07846(.A1(new_n10817_), .A2(pi0074), .B(new_n3225_), .ZN(new_n10818_));
  NOR2_X1    g07847(.A1(new_n10744_), .A2(new_n7941_), .ZN(new_n10819_));
  NOR2_X1    g07848(.A1(new_n10715_), .A2(new_n7942_), .ZN(new_n10820_));
  OR2_X2     g07849(.A1(new_n10820_), .A2(new_n10721_), .Z(new_n10821_));
  AOI22_X1   g07850(.A1(new_n7933_), .A2(new_n10821_), .B1(new_n7528_), .B2(new_n10714_), .ZN(new_n10822_));
  NAND2_X1   g07851(.A1(new_n10716_), .A2(new_n3188_), .ZN(new_n10823_));
  OAI22_X1   g07852(.A1(new_n10822_), .A2(new_n10823_), .B1(new_n10716_), .B2(new_n10819_), .ZN(new_n10824_));
  OAI21_X1   g07853(.A1(new_n10656_), .A2(new_n3098_), .B(new_n7510_), .ZN(new_n10825_));
  NAND2_X1   g07854(.A1(new_n10638_), .A2(new_n10825_), .ZN(new_n10826_));
  NOR2_X1    g07855(.A1(new_n7635_), .A2(new_n10826_), .ZN(new_n10827_));
  NAND4_X1   g07856(.A1(new_n10827_), .A2(new_n10712_), .A3(new_n10746_), .A4(new_n10824_), .ZN(new_n10828_));
  NOR3_X1    g07857(.A1(new_n10812_), .A2(new_n10818_), .A3(new_n10828_), .ZN(new_n10829_));
  NAND2_X1   g07858(.A1(new_n10798_), .A2(new_n10829_), .ZN(new_n10830_));
  AOI21_X1   g07859(.A1(new_n10830_), .A2(new_n10754_), .B(new_n10649_), .ZN(new_n10831_));
  NOR2_X1    g07860(.A1(new_n10831_), .A2(new_n7953_), .ZN(new_n10832_));
  NAND2_X1   g07861(.A1(new_n9782_), .A2(pi0118), .ZN(new_n10833_));
  XOR2_X1    g07862(.A1(new_n10832_), .A2(new_n10833_), .Z(new_n10834_));
  NOR2_X1    g07863(.A1(new_n10831_), .A2(new_n9783_), .ZN(new_n10835_));
  NOR2_X1    g07864(.A1(new_n9783_), .A2(new_n8218_), .ZN(new_n10836_));
  XNOR2_X1   g07865(.A1(new_n10835_), .A2(new_n10836_), .ZN(new_n10837_));
  AOI21_X1   g07866(.A1(new_n10837_), .A2(new_n10834_), .B(new_n10753_), .ZN(po0276));
  INV_X1     g07867(.I(pi0128), .ZN(new_n10839_));
  NOR2_X1    g07868(.A1(new_n10839_), .A2(new_n3005_), .ZN(new_n10840_));
  INV_X1     g07869(.I(new_n10840_), .ZN(new_n10841_));
  NAND2_X1   g07870(.A1(new_n10841_), .A2(pi0092), .ZN(new_n10842_));
  OAI21_X1   g07871(.A1(new_n6312_), .A2(new_n10842_), .B(new_n8286_), .ZN(new_n10843_));
  NAND4_X1   g07872(.A1(new_n2524_), .A2(pi0046), .A3(pi0108), .A4(new_n2731_), .ZN(new_n10844_));
  NAND4_X1   g07873(.A1(new_n6493_), .A2(pi0299), .A3(new_n5663_), .A4(new_n5666_), .ZN(new_n10845_));
  NAND3_X1   g07874(.A1(new_n5667_), .A2(new_n6493_), .A3(new_n3098_), .ZN(new_n10846_));
  AOI21_X1   g07875(.A1(new_n10845_), .A2(new_n10846_), .B(new_n5646_), .ZN(new_n10847_));
  AOI22_X1   g07876(.A1(new_n9433_), .A2(new_n10847_), .B1(pi0109), .B2(new_n2731_), .ZN(new_n10848_));
  NOR2_X1    g07877(.A1(new_n5618_), .A2(new_n10847_), .ZN(new_n10849_));
  AOI21_X1   g07878(.A1(new_n5562_), .A2(new_n10847_), .B(new_n10849_), .ZN(new_n10850_));
  OR2_X2     g07879(.A1(new_n10848_), .A2(new_n10850_), .Z(new_n10851_));
  OAI22_X1   g07880(.A1(new_n5589_), .A2(new_n2461_), .B1(pi0086), .B2(new_n9431_), .ZN(new_n10852_));
  NAND3_X1   g07881(.A1(new_n10852_), .A2(new_n2521_), .A3(new_n8280_), .ZN(new_n10853_));
  AOI21_X1   g07882(.A1(new_n10851_), .A2(new_n10844_), .B(new_n10853_), .ZN(new_n10854_));
  NOR2_X1    g07883(.A1(new_n10854_), .A2(new_n2798_), .ZN(new_n10855_));
  XOR2_X1    g07884(.A1(new_n10855_), .A2(new_n2799_), .Z(new_n10856_));
  NOR4_X1    g07885(.A1(new_n2880_), .A2(new_n2684_), .A3(new_n3259_), .A4(new_n10290_), .ZN(new_n10857_));
  NAND2_X1   g07886(.A1(new_n10856_), .A2(new_n10857_), .ZN(new_n10858_));
  NOR3_X1    g07887(.A1(new_n6543_), .A2(new_n3091_), .A3(new_n3382_), .ZN(new_n10859_));
  NAND2_X1   g07888(.A1(new_n6539_), .A2(new_n5293_), .ZN(new_n10860_));
  OAI21_X1   g07889(.A1(new_n10859_), .A2(new_n10860_), .B(new_n3312_), .ZN(new_n10861_));
  AOI21_X1   g07890(.A1(new_n10858_), .A2(new_n3183_), .B(new_n10861_), .ZN(new_n10862_));
  AOI21_X1   g07891(.A1(new_n10839_), .A2(pi0228), .B(new_n3462_), .ZN(new_n10863_));
  OAI21_X1   g07892(.A1(new_n10862_), .A2(pi0228), .B(new_n10863_), .ZN(new_n10864_));
  XOR2_X1    g07893(.A1(new_n10864_), .A2(new_n3477_), .Z(new_n10865_));
  OAI21_X1   g07894(.A1(new_n3412_), .A2(new_n3212_), .B(new_n10841_), .ZN(new_n10866_));
  AOI21_X1   g07895(.A1(new_n10841_), .A2(pi0087), .B(pi0075), .ZN(new_n10867_));
  OAI21_X1   g07896(.A1(new_n10865_), .A2(new_n10866_), .B(new_n10867_), .ZN(new_n10868_));
  NAND3_X1   g07897(.A1(new_n3411_), .A2(new_n3462_), .A3(new_n7333_), .ZN(new_n10869_));
  NAND2_X1   g07898(.A1(new_n10869_), .A2(new_n3483_), .ZN(new_n10870_));
  NAND4_X1   g07899(.A1(new_n10868_), .A2(new_n8286_), .A3(new_n10840_), .A4(new_n10870_), .ZN(new_n10871_));
  XOR2_X1    g07900(.A1(new_n10871_), .A2(new_n10843_), .Z(po0277));
  OAI21_X1   g07901(.A1(new_n6403_), .A2(new_n6941_), .B(new_n6410_), .ZN(new_n10873_));
  AOI21_X1   g07902(.A1(new_n3160_), .A2(new_n10873_), .B(new_n3474_), .ZN(new_n10874_));
  AOI21_X1   g07903(.A1(new_n6943_), .A2(new_n10874_), .B(pi0087), .ZN(new_n10875_));
  NOR3_X1    g07904(.A1(new_n10875_), .A2(new_n3474_), .A3(new_n6407_), .ZN(new_n10876_));
  NOR2_X1    g07905(.A1(new_n6390_), .A2(pi1093), .ZN(new_n10877_));
  INV_X1     g07906(.I(new_n10877_), .ZN(new_n10878_));
  AOI21_X1   g07907(.A1(pi0122), .A2(new_n2728_), .B(new_n6388_), .ZN(new_n10879_));
  NAND3_X1   g07908(.A1(new_n6387_), .A2(new_n6410_), .A3(new_n6403_), .ZN(new_n10880_));
  NAND3_X1   g07909(.A1(new_n10880_), .A2(pi0829), .A3(new_n5532_), .ZN(new_n10881_));
  OAI21_X1   g07910(.A1(new_n10881_), .A2(new_n10879_), .B(new_n9299_), .ZN(new_n10882_));
  AOI21_X1   g07911(.A1(new_n10882_), .A2(new_n8400_), .B(new_n2986_), .ZN(new_n10883_));
  AOI21_X1   g07912(.A1(new_n6388_), .A2(new_n6402_), .B(new_n6941_), .ZN(new_n10884_));
  AOI21_X1   g07913(.A1(new_n9987_), .A2(new_n10884_), .B(new_n10883_), .ZN(new_n10885_));
  NAND2_X1   g07914(.A1(new_n10885_), .A2(new_n10878_), .ZN(new_n10886_));
  NAND2_X1   g07915(.A1(new_n10886_), .A2(pi0039), .ZN(new_n10887_));
  XOR2_X1    g07916(.A1(new_n10887_), .A2(new_n3262_), .Z(new_n10888_));
  NAND2_X1   g07917(.A1(new_n6406_), .A2(new_n6443_), .ZN(new_n10889_));
  XOR2_X1    g07918(.A1(new_n6440_), .A2(new_n10889_), .Z(new_n10890_));
  NOR2_X1    g07919(.A1(new_n7611_), .A2(new_n6407_), .ZN(new_n10891_));
  AOI21_X1   g07920(.A1(new_n10890_), .A2(new_n7611_), .B(new_n10891_), .ZN(new_n10892_));
  INV_X1     g07921(.I(new_n10892_), .ZN(new_n10893_));
  NOR2_X1    g07922(.A1(new_n6407_), .A2(new_n5385_), .ZN(new_n10894_));
  AOI21_X1   g07923(.A1(new_n10890_), .A2(new_n5385_), .B(new_n10894_), .ZN(new_n10895_));
  NAND2_X1   g07924(.A1(new_n10895_), .A2(new_n6459_), .ZN(new_n10896_));
  XNOR2_X1   g07925(.A1(new_n10896_), .A2(new_n6462_), .ZN(new_n10897_));
  AOI21_X1   g07926(.A1(new_n10897_), .A2(new_n10893_), .B(pi0299), .ZN(new_n10898_));
  NOR3_X1    g07927(.A1(new_n10898_), .A2(new_n6407_), .A3(new_n6461_), .ZN(new_n10899_));
  NAND2_X1   g07928(.A1(new_n9863_), .A2(new_n6453_), .ZN(new_n10900_));
  NAND2_X1   g07929(.A1(new_n10900_), .A2(new_n3098_), .ZN(new_n10901_));
  NAND2_X1   g07930(.A1(new_n10895_), .A2(new_n6451_), .ZN(new_n10902_));
  XOR2_X1    g07931(.A1(new_n10902_), .A2(new_n6454_), .Z(new_n10903_));
  NOR2_X1    g07932(.A1(new_n10903_), .A2(new_n10892_), .ZN(new_n10904_));
  OAI21_X1   g07933(.A1(new_n10899_), .A2(new_n10901_), .B(new_n10904_), .ZN(new_n10905_));
  OAI21_X1   g07934(.A1(new_n10888_), .A2(new_n10905_), .B(new_n3462_), .ZN(new_n10906_));
  NAND3_X1   g07935(.A1(new_n10906_), .A2(new_n9863_), .A3(new_n7487_), .ZN(new_n10907_));
  AOI21_X1   g07936(.A1(new_n10907_), .A2(new_n6534_), .B(new_n6407_), .ZN(new_n10908_));
  NOR2_X1    g07937(.A1(new_n6497_), .A2(new_n3235_), .ZN(new_n10909_));
  OAI21_X1   g07938(.A1(pi1091), .A2(new_n6406_), .B(new_n6894_), .ZN(new_n10910_));
  NAND2_X1   g07939(.A1(new_n10910_), .A2(pi0075), .ZN(new_n10911_));
  XOR2_X1    g07940(.A1(new_n10911_), .A2(new_n10909_), .Z(new_n10912_));
  NOR3_X1    g07941(.A1(new_n10912_), .A2(new_n3235_), .A3(new_n6407_), .ZN(new_n10913_));
  OAI21_X1   g07942(.A1(new_n10908_), .A2(new_n10913_), .B(new_n10876_), .ZN(new_n10914_));
  NAND3_X1   g07943(.A1(new_n6349_), .A2(new_n10163_), .A3(pi0818), .ZN(new_n10915_));
  INV_X1     g07944(.I(new_n10915_), .ZN(new_n10916_));
  INV_X1     g07945(.I(new_n6529_), .ZN(new_n10917_));
  NOR2_X1    g07946(.A1(new_n10883_), .A2(new_n10884_), .ZN(new_n10918_));
  OAI21_X1   g07947(.A1(new_n6551_), .A2(new_n3462_), .B(new_n3183_), .ZN(new_n10919_));
  NAND3_X1   g07948(.A1(new_n10878_), .A2(new_n10918_), .A3(new_n10919_), .ZN(new_n10920_));
  NAND2_X1   g07949(.A1(new_n6946_), .A2(pi0087), .ZN(new_n10921_));
  AOI21_X1   g07950(.A1(new_n10920_), .A2(new_n10921_), .B(new_n6534_), .ZN(new_n10922_));
  OAI21_X1   g07951(.A1(new_n10922_), .A2(pi0075), .B(new_n10917_), .ZN(new_n10923_));
  NAND2_X1   g07952(.A1(new_n10923_), .A2(new_n6939_), .ZN(new_n10924_));
  INV_X1     g07953(.I(pi0120), .ZN(new_n10925_));
  NOR2_X1    g07954(.A1(new_n6400_), .A2(new_n10925_), .ZN(new_n10926_));
  NOR2_X1    g07955(.A1(pi0120), .A2(pi1093), .ZN(new_n10927_));
  NOR3_X1    g07956(.A1(new_n9987_), .A2(new_n2726_), .A3(new_n10927_), .ZN(new_n10928_));
  NOR2_X1    g07957(.A1(new_n9863_), .A2(new_n10925_), .ZN(new_n10929_));
  NOR2_X1    g07958(.A1(new_n10929_), .A2(new_n10928_), .ZN(new_n10930_));
  INV_X1     g07959(.I(new_n10930_), .ZN(new_n10931_));
  NOR2_X1    g07960(.A1(new_n10931_), .A2(new_n6668_), .ZN(new_n10932_));
  INV_X1     g07961(.I(new_n10932_), .ZN(new_n10933_));
  INV_X1     g07962(.I(new_n10927_), .ZN(new_n10934_));
  NAND2_X1   g07963(.A1(new_n10915_), .A2(new_n10934_), .ZN(new_n10935_));
  OAI21_X1   g07964(.A1(po1038), .A2(new_n10935_), .B(new_n7250_), .ZN(new_n10936_));
  OAI21_X1   g07965(.A1(new_n10933_), .A2(new_n10936_), .B(new_n10925_), .ZN(new_n10937_));
  NAND2_X1   g07966(.A1(new_n10937_), .A2(new_n10932_), .ZN(new_n10938_));
  NAND2_X1   g07967(.A1(new_n10938_), .A2(new_n10925_), .ZN(new_n10939_));
  AOI21_X1   g07968(.A1(new_n9863_), .A2(new_n6400_), .B(new_n6668_), .ZN(new_n10940_));
  NAND2_X1   g07969(.A1(new_n10933_), .A2(new_n6400_), .ZN(new_n10941_));
  NAND3_X1   g07970(.A1(new_n10939_), .A2(new_n10940_), .A3(new_n10941_), .ZN(new_n10942_));
  AOI21_X1   g07971(.A1(new_n10924_), .A2(new_n10926_), .B(new_n10942_), .ZN(new_n10943_));
  NAND3_X1   g07972(.A1(pi0951), .A2(pi0982), .A3(pi1092), .ZN(new_n10944_));
  NOR2_X1    g07973(.A1(new_n10944_), .A2(new_n2984_), .ZN(new_n10945_));
  NOR2_X1    g07974(.A1(new_n10945_), .A2(pi0120), .ZN(new_n10946_));
  INV_X1     g07975(.I(new_n10946_), .ZN(new_n10947_));
  AOI21_X1   g07976(.A1(new_n10936_), .A2(new_n10947_), .B(new_n10933_), .ZN(new_n10948_));
  INV_X1     g07977(.I(new_n10948_), .ZN(new_n10949_));
  AOI21_X1   g07978(.A1(new_n10877_), .A2(pi0120), .B(pi0039), .ZN(new_n10958_));
  OAI21_X1   g07979(.A1(pi0120), .A2(pi1093), .B(new_n3462_), .ZN(new_n10961_));
  NOR2_X1    g07980(.A1(new_n6947_), .A2(new_n10927_), .ZN(new_n10962_));
  AOI21_X1   g07981(.A1(new_n10962_), .A2(pi0075), .B(pi0087), .ZN(new_n10963_));
  NOR2_X1    g07982(.A1(new_n6525_), .A2(new_n3145_), .ZN(new_n10964_));
  NOR3_X1    g07983(.A1(new_n6532_), .A2(new_n10925_), .A3(new_n6512_), .ZN(new_n10965_));
  NOR3_X1    g07984(.A1(new_n6507_), .A2(pi0120), .A3(new_n6512_), .ZN(new_n10966_));
  OAI21_X1   g07985(.A1(new_n10965_), .A2(new_n10966_), .B(new_n10964_), .ZN(new_n10967_));
  NOR2_X1    g07986(.A1(new_n10967_), .A2(new_n10963_), .ZN(new_n10968_));
  AOI21_X1   g07987(.A1(new_n10968_), .A2(new_n10961_), .B(new_n6399_), .ZN(new_n10969_));
  AOI21_X1   g07988(.A1(new_n6939_), .A2(new_n10927_), .B(new_n6400_), .ZN(new_n10970_));
  INV_X1     g07989(.I(new_n10885_), .ZN(new_n10971_));
  NAND2_X1   g07990(.A1(new_n2726_), .A2(new_n2979_), .ZN(new_n10972_));
  NAND2_X1   g07991(.A1(new_n6407_), .A2(new_n10925_), .ZN(new_n10973_));
  AOI21_X1   g07992(.A1(new_n6439_), .A2(new_n10972_), .B(new_n10973_), .ZN(new_n10974_));
  NOR2_X1    g07993(.A1(new_n10974_), .A2(new_n6537_), .ZN(new_n10975_));
  NOR2_X1    g07994(.A1(new_n10931_), .A2(new_n7611_), .ZN(new_n10976_));
  AOI21_X1   g07995(.A1(new_n10975_), .A2(new_n7611_), .B(new_n10976_), .ZN(new_n10977_));
  NOR2_X1    g07996(.A1(new_n10975_), .A2(new_n6448_), .ZN(new_n10978_));
  AOI21_X1   g07997(.A1(new_n6448_), .A2(new_n10931_), .B(new_n10978_), .ZN(new_n10979_));
  NAND2_X1   g07998(.A1(new_n10979_), .A2(new_n6459_), .ZN(new_n10980_));
  XOR2_X1    g07999(.A1(new_n10980_), .A2(new_n6462_), .Z(new_n10981_));
  OAI21_X1   g08000(.A1(new_n10981_), .A2(new_n10977_), .B(new_n3098_), .ZN(new_n10982_));
  NAND3_X1   g08001(.A1(new_n10982_), .A2(new_n6459_), .A3(new_n10930_), .ZN(new_n10983_));
  NAND2_X1   g08002(.A1(new_n10979_), .A2(new_n6451_), .ZN(new_n10984_));
  XOR2_X1    g08003(.A1(new_n10984_), .A2(new_n6454_), .Z(new_n10985_));
  OAI21_X1   g08004(.A1(new_n10985_), .A2(new_n10977_), .B(new_n3098_), .ZN(new_n10986_));
  NAND3_X1   g08005(.A1(new_n10986_), .A2(new_n6451_), .A3(new_n10930_), .ZN(new_n10987_));
  NAND3_X1   g08006(.A1(new_n10983_), .A2(new_n10987_), .A3(new_n3262_), .ZN(new_n10988_));
  OAI21_X1   g08007(.A1(new_n9863_), .A2(new_n5485_), .B(new_n10927_), .ZN(new_n10989_));
  NOR2_X1    g08008(.A1(new_n10964_), .A2(new_n10973_), .ZN(new_n10990_));
  OAI21_X1   g08009(.A1(new_n10990_), .A2(new_n6532_), .B(new_n2984_), .ZN(new_n10991_));
  NOR2_X1    g08010(.A1(new_n10930_), .A2(pi0100), .ZN(new_n10992_));
  NOR4_X1    g08011(.A1(new_n10992_), .A2(new_n3455_), .A3(new_n10925_), .A4(new_n6512_), .ZN(new_n10993_));
  NAND2_X1   g08012(.A1(new_n10991_), .A2(new_n10993_), .ZN(new_n10994_));
  AOI21_X1   g08013(.A1(new_n10994_), .A2(new_n10989_), .B(new_n3235_), .ZN(new_n10995_));
  NAND2_X1   g08014(.A1(new_n10958_), .A2(new_n10995_), .ZN(new_n10996_));
  AOI21_X1   g08015(.A1(new_n10988_), .A2(new_n10971_), .B(new_n10996_), .ZN(new_n10997_));
  OAI21_X1   g08016(.A1(new_n10997_), .A2(new_n10876_), .B(new_n10962_), .ZN(new_n10998_));
  NAND2_X1   g08017(.A1(new_n5499_), .A2(new_n3175_), .ZN(new_n10999_));
  NAND2_X1   g08018(.A1(new_n3193_), .A2(pi0075), .ZN(new_n11000_));
  AOI21_X1   g08019(.A1(new_n10910_), .A2(pi0120), .B(new_n6495_), .ZN(new_n11001_));
  NAND2_X1   g08020(.A1(new_n6527_), .A2(new_n10928_), .ZN(new_n11002_));
  AOI22_X1   g08021(.A1(new_n11002_), .A2(new_n11001_), .B1(new_n6495_), .B2(new_n10930_), .ZN(new_n11003_));
  NOR2_X1    g08022(.A1(new_n11003_), .A2(new_n3235_), .ZN(new_n11004_));
  XNOR2_X1   g08023(.A1(new_n11004_), .A2(new_n11000_), .ZN(new_n11005_));
  NAND3_X1   g08024(.A1(new_n11005_), .A2(new_n10930_), .A3(new_n10916_), .ZN(new_n11006_));
  AOI21_X1   g08025(.A1(new_n10998_), .A2(new_n10999_), .B(new_n11006_), .ZN(new_n11007_));
  NOR3_X1    g08026(.A1(new_n10917_), .A2(new_n10934_), .A3(new_n10938_), .ZN(new_n11008_));
  OAI21_X1   g08027(.A1(new_n11007_), .A2(new_n10970_), .B(new_n11008_), .ZN(new_n11009_));
  OAI22_X1   g08028(.A1(new_n11009_), .A2(new_n10969_), .B1(new_n7240_), .B2(new_n10949_), .ZN(new_n11010_));
  AOI22_X1   g08029(.A1(new_n10914_), .A2(new_n10943_), .B1(new_n10916_), .B2(new_n11010_), .ZN(new_n11011_));
  NOR2_X1    g08030(.A1(new_n10930_), .A2(new_n10946_), .ZN(new_n11012_));
  INV_X1     g08031(.I(new_n11012_), .ZN(new_n11013_));
  NAND2_X1   g08032(.A1(new_n6537_), .A2(pi0120), .ZN(new_n11014_));
  INV_X1     g08033(.I(new_n10945_), .ZN(new_n11015_));
  NOR2_X1    g08034(.A1(new_n11015_), .A2(pi1091), .ZN(new_n11016_));
  INV_X1     g08035(.I(new_n11016_), .ZN(new_n11017_));
  NOR2_X1    g08036(.A1(new_n9986_), .A2(new_n11017_), .ZN(new_n11018_));
  NOR3_X1    g08037(.A1(new_n11018_), .A2(new_n6407_), .A3(new_n10925_), .ZN(new_n11019_));
  NOR2_X1    g08038(.A1(new_n2986_), .A2(new_n10944_), .ZN(new_n11020_));
  INV_X1     g08039(.I(new_n11020_), .ZN(new_n11021_));
  OAI21_X1   g08040(.A1(new_n6439_), .A2(new_n11021_), .B(new_n11019_), .ZN(new_n11022_));
  XOR2_X1    g08041(.A1(new_n11014_), .A2(new_n11022_), .Z(new_n11023_));
  NAND2_X1   g08042(.A1(new_n11023_), .A2(new_n7611_), .ZN(new_n11024_));
  OAI21_X1   g08043(.A1(new_n7611_), .A2(new_n11012_), .B(new_n11024_), .ZN(new_n11025_));
  NOR2_X1    g08044(.A1(new_n11012_), .A2(new_n5385_), .ZN(new_n11026_));
  AOI21_X1   g08045(.A1(new_n11023_), .A2(new_n5385_), .B(new_n11026_), .ZN(new_n11027_));
  NAND2_X1   g08046(.A1(new_n11027_), .A2(new_n6459_), .ZN(new_n11028_));
  XNOR2_X1   g08047(.A1(new_n11028_), .A2(new_n6462_), .ZN(new_n11029_));
  NAND2_X1   g08048(.A1(new_n11029_), .A2(new_n11025_), .ZN(new_n11030_));
  NAND2_X1   g08049(.A1(new_n6459_), .A2(pi0299), .ZN(new_n11031_));
  AOI21_X1   g08050(.A1(new_n10931_), .A2(new_n11031_), .B(new_n10947_), .ZN(new_n11032_));
  AOI21_X1   g08051(.A1(new_n11030_), .A2(new_n11032_), .B(new_n3183_), .ZN(new_n11033_));
  INV_X1     g08052(.I(new_n6374_), .ZN(new_n11034_));
  NOR2_X1    g08053(.A1(new_n6411_), .A2(pi0950), .ZN(new_n11035_));
  NOR4_X1    g08054(.A1(new_n2544_), .A2(new_n6360_), .A3(new_n2558_), .A4(new_n2522_), .ZN(new_n11036_));
  NAND4_X1   g08055(.A1(new_n6373_), .A2(pi0090), .A3(new_n2902_), .A4(new_n11036_), .ZN(new_n11037_));
  NOR3_X1    g08056(.A1(new_n11034_), .A2(new_n11035_), .A3(new_n11037_), .ZN(new_n11038_));
  NOR4_X1    g08057(.A1(new_n11034_), .A2(new_n5683_), .A3(new_n11035_), .A4(new_n11037_), .ZN(new_n11039_));
  NOR2_X1    g08058(.A1(new_n11039_), .A2(new_n10944_), .ZN(new_n11040_));
  NAND2_X1   g08059(.A1(new_n11040_), .A2(new_n11038_), .ZN(new_n11041_));
  NAND2_X1   g08060(.A1(pi0122), .A2(pi0829), .ZN(new_n11042_));
  OAI21_X1   g08061(.A1(new_n10944_), .A2(new_n11042_), .B(new_n11041_), .ZN(new_n11043_));
  NOR2_X1    g08062(.A1(new_n2929_), .A2(new_n2931_), .ZN(new_n11044_));
  NAND2_X1   g08063(.A1(new_n11036_), .A2(pi0097), .ZN(new_n11045_));
  OAI22_X1   g08064(.A1(new_n6371_), .A2(new_n2678_), .B1(new_n11044_), .B2(new_n11045_), .ZN(new_n11046_));
  NAND2_X1   g08065(.A1(new_n11046_), .A2(new_n6422_), .ZN(new_n11047_));
  NAND2_X1   g08066(.A1(new_n11047_), .A2(pi0051), .ZN(new_n11048_));
  NOR3_X1    g08067(.A1(new_n6372_), .A2(new_n2702_), .A3(new_n8393_), .ZN(new_n11049_));
  NOR2_X1    g08068(.A1(new_n11048_), .A2(new_n11049_), .ZN(new_n11050_));
  NOR4_X1    g08069(.A1(new_n11047_), .A2(new_n2702_), .A3(new_n8393_), .A4(new_n6372_), .ZN(new_n11051_));
  NOR3_X1    g08070(.A1(new_n11050_), .A2(new_n11051_), .A3(pi0096), .ZN(new_n11052_));
  NAND4_X1   g08071(.A1(new_n8402_), .A2(new_n2437_), .A3(pi0950), .A4(new_n3137_), .ZN(new_n11053_));
  NOR2_X1    g08072(.A1(new_n6378_), .A2(new_n10944_), .ZN(new_n11054_));
  OAI21_X1   g08073(.A1(new_n11052_), .A2(new_n11053_), .B(new_n11054_), .ZN(new_n11055_));
  NAND2_X1   g08074(.A1(new_n6431_), .A2(pi1091), .ZN(new_n11056_));
  AOI21_X1   g08075(.A1(new_n11043_), .A2(new_n11055_), .B(new_n11056_), .ZN(new_n11057_));
  OAI21_X1   g08076(.A1(new_n11057_), .A2(new_n2728_), .B(new_n10945_), .ZN(new_n11058_));
  NAND2_X1   g08077(.A1(new_n11058_), .A2(pi0120), .ZN(new_n11059_));
  NAND4_X1   g08078(.A1(new_n11040_), .A2(pi0120), .A3(new_n6940_), .A4(new_n9987_), .ZN(new_n11060_));
  NOR2_X1    g08079(.A1(new_n10886_), .A2(new_n11060_), .ZN(new_n11061_));
  XNOR2_X1   g08080(.A1(new_n11061_), .A2(new_n11059_), .ZN(new_n11062_));
  NAND2_X1   g08081(.A1(new_n11027_), .A2(new_n6451_), .ZN(new_n11063_));
  XNOR2_X1   g08082(.A1(new_n11063_), .A2(new_n6454_), .ZN(new_n11064_));
  AOI21_X1   g08083(.A1(new_n6453_), .A2(new_n10946_), .B(new_n3098_), .ZN(new_n11065_));
  NAND3_X1   g08084(.A1(new_n10900_), .A2(pi0039), .A3(new_n11065_), .ZN(new_n11066_));
  AOI21_X1   g08085(.A1(new_n11064_), .A2(new_n11025_), .B(new_n11066_), .ZN(new_n11067_));
  NAND2_X1   g08086(.A1(new_n11062_), .A2(new_n11067_), .ZN(new_n11068_));
  OAI21_X1   g08087(.A1(new_n11068_), .A2(new_n11033_), .B(pi0038), .ZN(new_n11069_));
  AOI21_X1   g08088(.A1(new_n11033_), .A2(new_n11068_), .B(new_n11069_), .ZN(new_n11070_));
  XOR2_X1    g08089(.A1(new_n11070_), .A2(new_n5486_), .Z(new_n11071_));
  NOR2_X1    g08090(.A1(new_n11071_), .A2(new_n11013_), .ZN(new_n11072_));
  NOR2_X1    g08091(.A1(new_n2728_), .A2(new_n5531_), .ZN(new_n11073_));
  NOR3_X1    g08092(.A1(new_n11020_), .A2(pi0950), .A3(new_n11073_), .ZN(new_n11074_));
  NOR2_X1    g08093(.A1(new_n3145_), .A2(new_n11074_), .ZN(new_n11075_));
  INV_X1     g08094(.I(new_n11075_), .ZN(new_n11076_));
  NAND2_X1   g08095(.A1(new_n5683_), .A2(new_n2722_), .ZN(new_n11077_));
  OAI21_X1   g08096(.A1(new_n11016_), .A2(new_n11077_), .B(new_n3160_), .ZN(new_n11078_));
  AOI21_X1   g08097(.A1(new_n11076_), .A2(new_n11078_), .B(pi0120), .ZN(new_n11079_));
  NOR2_X1    g08098(.A1(new_n11075_), .A2(new_n11018_), .ZN(new_n11080_));
  AOI21_X1   g08099(.A1(new_n3474_), .A2(new_n10946_), .B(new_n3455_), .ZN(new_n11081_));
  OAI21_X1   g08100(.A1(new_n6407_), .A2(new_n3134_), .B(new_n11081_), .ZN(new_n11082_));
  NOR2_X1    g08101(.A1(new_n11080_), .A2(new_n11082_), .ZN(new_n11083_));
  AOI22_X1   g08102(.A1(new_n11079_), .A2(new_n11083_), .B1(new_n6943_), .B2(new_n10874_), .ZN(new_n11084_));
  AOI21_X1   g08103(.A1(pi0120), .A2(new_n3134_), .B(new_n6944_), .ZN(new_n11085_));
  NOR4_X1    g08104(.A1(new_n11084_), .A2(new_n3455_), .A3(new_n6943_), .A4(new_n11085_), .ZN(new_n11086_));
  OAI21_X1   g08105(.A1(new_n10940_), .A2(new_n10934_), .B(new_n6399_), .ZN(new_n11087_));
  NAND2_X1   g08106(.A1(new_n11039_), .A2(new_n11016_), .ZN(new_n11088_));
  AOI21_X1   g08107(.A1(new_n11058_), .A2(new_n10925_), .B(new_n11088_), .ZN(new_n11089_));
  NOR4_X1    g08108(.A1(new_n10877_), .A2(new_n10925_), .A3(new_n10883_), .A4(new_n10884_), .ZN(new_n11090_));
  OAI21_X1   g08109(.A1(pi0039), .A2(new_n11089_), .B(new_n11090_), .ZN(new_n11091_));
  NOR2_X1    g08110(.A1(new_n6512_), .A2(new_n3259_), .ZN(new_n11092_));
  NAND3_X1   g08111(.A1(new_n3145_), .A2(new_n2722_), .A3(new_n11021_), .ZN(new_n11093_));
  NAND3_X1   g08112(.A1(new_n6483_), .A2(new_n6359_), .A3(new_n11093_), .ZN(new_n11094_));
  NAND2_X1   g08113(.A1(new_n11094_), .A2(pi0120), .ZN(new_n11095_));
  NOR2_X1    g08114(.A1(new_n11017_), .A2(new_n10925_), .ZN(new_n11096_));
  INV_X1     g08115(.I(new_n11096_), .ZN(new_n11097_));
  NOR2_X1    g08116(.A1(new_n6532_), .A2(new_n11097_), .ZN(new_n11098_));
  OR2_X2     g08117(.A1(new_n11098_), .A2(new_n11095_), .Z(new_n11099_));
  NAND2_X1   g08118(.A1(new_n8494_), .A2(new_n3462_), .ZN(new_n11100_));
  AOI21_X1   g08119(.A1(new_n11098_), .A2(new_n11095_), .B(new_n11100_), .ZN(new_n11101_));
  NAND2_X1   g08120(.A1(new_n10946_), .A2(pi0039), .ZN(new_n11102_));
  AOI21_X1   g08121(.A1(new_n11099_), .A2(new_n11101_), .B(new_n11102_), .ZN(new_n11103_));
  OAI21_X1   g08122(.A1(new_n11103_), .A2(new_n11092_), .B(new_n3132_), .ZN(new_n11104_));
  NOR2_X1    g08123(.A1(new_n6797_), .A2(new_n10946_), .ZN(new_n11105_));
  NOR2_X1    g08124(.A1(new_n11105_), .A2(new_n6461_), .ZN(new_n11106_));
  XOR2_X1    g08125(.A1(new_n11106_), .A2(new_n6462_), .Z(new_n11107_));
  NAND3_X1   g08126(.A1(new_n11107_), .A2(new_n6803_), .A3(new_n10947_), .ZN(new_n11108_));
  NAND3_X1   g08127(.A1(new_n6459_), .A2(new_n10946_), .A3(pi0039), .ZN(new_n11109_));
  AOI21_X1   g08128(.A1(new_n11108_), .A2(new_n3098_), .B(new_n11109_), .ZN(new_n11110_));
  NOR2_X1    g08129(.A1(new_n11105_), .A2(new_n6453_), .ZN(new_n11111_));
  XNOR2_X1   g08130(.A1(new_n11111_), .A2(new_n6454_), .ZN(new_n11112_));
  INV_X1     g08131(.I(new_n11081_), .ZN(new_n11113_));
  NOR3_X1    g08132(.A1(new_n11085_), .A2(new_n6943_), .A3(new_n11079_), .ZN(new_n11114_));
  OAI21_X1   g08133(.A1(new_n11114_), .A2(new_n11113_), .B(new_n3235_), .ZN(new_n11115_));
  NAND4_X1   g08134(.A1(new_n6803_), .A2(pi0087), .A3(new_n11115_), .A4(new_n10947_), .ZN(new_n11116_));
  NOR2_X1    g08135(.A1(new_n11112_), .A2(new_n11116_), .ZN(new_n11117_));
  OAI21_X1   g08136(.A1(new_n11110_), .A2(new_n11065_), .B(new_n11117_), .ZN(new_n11118_));
  AOI21_X1   g08137(.A1(new_n11091_), .A2(new_n11104_), .B(new_n11118_), .ZN(new_n11119_));
  NOR2_X1    g08138(.A1(new_n6939_), .A2(new_n6400_), .ZN(new_n11120_));
  NAND4_X1   g08139(.A1(new_n9010_), .A2(pi0093), .A3(pi0122), .A4(new_n2497_), .ZN(new_n11121_));
  NOR2_X1    g08140(.A1(new_n3721_), .A2(new_n2721_), .ZN(new_n11122_));
  NAND4_X1   g08141(.A1(new_n2795_), .A2(new_n3137_), .A3(pi0950), .A4(new_n11122_), .ZN(new_n11123_));
  OAI21_X1   g08142(.A1(new_n11123_), .A2(new_n11121_), .B(new_n11021_), .ZN(new_n11124_));
  OAI21_X1   g08143(.A1(new_n2470_), .A2(new_n11124_), .B(new_n6483_), .ZN(new_n11125_));
  NAND2_X1   g08144(.A1(new_n11125_), .A2(pi0120), .ZN(new_n11126_));
  NOR3_X1    g08145(.A1(new_n6527_), .A2(new_n2984_), .A3(new_n11097_), .ZN(new_n11127_));
  AOI21_X1   g08146(.A1(new_n11127_), .A2(new_n11126_), .B(new_n3194_), .ZN(new_n11128_));
  OAI21_X1   g08147(.A1(new_n11126_), .A2(new_n11127_), .B(new_n11128_), .ZN(new_n11129_));
  NAND2_X1   g08148(.A1(new_n6495_), .A2(new_n3193_), .ZN(new_n11130_));
  XOR2_X1    g08149(.A1(new_n11129_), .A2(new_n11130_), .Z(new_n11131_));
  NAND2_X1   g08150(.A1(new_n11131_), .A2(new_n10946_), .ZN(new_n11132_));
  NAND4_X1   g08151(.A1(new_n10948_), .A2(new_n3193_), .A3(new_n6399_), .A4(new_n10946_), .ZN(new_n11133_));
  AOI21_X1   g08152(.A1(new_n11132_), .A2(new_n3235_), .B(new_n11133_), .ZN(new_n11134_));
  OAI21_X1   g08153(.A1(new_n11119_), .A2(new_n11120_), .B(new_n11134_), .ZN(new_n11135_));
  INV_X1     g08154(.I(new_n11125_), .ZN(new_n11136_));
  NOR3_X1    g08155(.A1(new_n10910_), .A2(new_n10925_), .A3(new_n6495_), .ZN(new_n11137_));
  OAI21_X1   g08156(.A1(new_n11137_), .A2(new_n11018_), .B(new_n11136_), .ZN(new_n11138_));
  NAND2_X1   g08157(.A1(new_n11013_), .A2(new_n6495_), .ZN(new_n11139_));
  AOI21_X1   g08158(.A1(new_n11138_), .A2(new_n11139_), .B(new_n3235_), .ZN(new_n11140_));
  XOR2_X1    g08159(.A1(new_n11140_), .A2(new_n11000_), .Z(new_n11141_));
  OAI21_X1   g08160(.A1(new_n11141_), .A2(new_n11013_), .B(new_n6400_), .ZN(new_n11142_));
  NOR2_X1    g08161(.A1(new_n6507_), .A2(new_n10925_), .ZN(new_n11143_));
  NAND2_X1   g08162(.A1(new_n11094_), .A2(new_n11019_), .ZN(new_n11144_));
  OAI21_X1   g08163(.A1(new_n11143_), .A2(new_n11144_), .B(new_n3211_), .ZN(new_n11145_));
  AOI21_X1   g08164(.A1(new_n11143_), .A2(new_n11144_), .B(new_n11145_), .ZN(new_n11146_));
  XNOR2_X1   g08165(.A1(new_n11146_), .A2(new_n6512_), .ZN(new_n11147_));
  AOI21_X1   g08166(.A1(new_n11147_), .A2(new_n11012_), .B(pi0100), .ZN(new_n11148_));
  NOR4_X1    g08167(.A1(new_n11148_), .A2(new_n3235_), .A3(new_n3212_), .A4(new_n11013_), .ZN(new_n11149_));
  NAND2_X1   g08168(.A1(new_n11149_), .A2(new_n11142_), .ZN(new_n11150_));
  AOI21_X1   g08169(.A1(new_n11135_), .A2(new_n11087_), .B(new_n11150_), .ZN(new_n11151_));
  OAI21_X1   g08170(.A1(new_n11072_), .A2(new_n11086_), .B(new_n11151_), .ZN(new_n11152_));
  NOR2_X1    g08171(.A1(new_n11152_), .A2(new_n11011_), .ZN(po0278));
  NOR4_X1    g08172(.A1(new_n10245_), .A2(new_n2623_), .A3(new_n7362_), .A4(new_n8276_), .ZN(new_n11154_));
  NAND4_X1   g08173(.A1(new_n11154_), .A2(pi0050), .A3(pi0077), .A4(new_n2667_), .ZN(new_n11155_));
  NOR2_X1    g08174(.A1(new_n6368_), .A2(new_n2473_), .ZN(new_n11156_));
  INV_X1     g08175(.I(new_n11156_), .ZN(new_n11157_));
  NOR3_X1    g08176(.A1(new_n11157_), .A2(pi0024), .A3(new_n9231_), .ZN(new_n11158_));
  NAND2_X1   g08177(.A1(new_n11158_), .A2(new_n7269_), .ZN(new_n11159_));
  NOR2_X1    g08178(.A1(new_n11155_), .A2(new_n11159_), .ZN(new_n11160_));
  NAND2_X1   g08179(.A1(new_n11160_), .A2(new_n10275_), .ZN(new_n11161_));
  INV_X1     g08180(.I(new_n11161_), .ZN(new_n11162_));
  NAND2_X1   g08181(.A1(new_n11154_), .A2(new_n2521_), .ZN(new_n11163_));
  OAI21_X1   g08182(.A1(new_n9427_), .A2(new_n11163_), .B(new_n11155_), .ZN(new_n11164_));
  NAND3_X1   g08183(.A1(new_n11164_), .A2(pi0024), .A3(new_n7269_), .ZN(new_n11165_));
  NOR4_X1    g08184(.A1(new_n2606_), .A2(new_n2611_), .A3(new_n2450_), .A4(new_n2598_), .ZN(new_n11166_));
  INV_X1     g08185(.I(new_n11166_), .ZN(new_n11167_));
  NOR4_X1    g08186(.A1(new_n11163_), .A2(new_n7272_), .A3(new_n9427_), .A4(new_n7270_), .ZN(new_n11168_));
  NOR2_X1    g08187(.A1(new_n11168_), .A2(new_n11167_), .ZN(new_n11169_));
  NAND2_X1   g08188(.A1(new_n11165_), .A2(new_n11169_), .ZN(new_n11170_));
  AOI21_X1   g08189(.A1(new_n11157_), .A2(new_n11166_), .B(pi0051), .ZN(new_n11171_));
  NAND2_X1   g08190(.A1(new_n11170_), .A2(new_n11171_), .ZN(new_n11172_));
  NOR2_X1    g08191(.A1(new_n11172_), .A2(new_n3304_), .ZN(new_n11173_));
  INV_X1     g08192(.I(new_n11173_), .ZN(new_n11174_));
  NOR2_X1    g08193(.A1(new_n11167_), .A2(pi0051), .ZN(new_n11175_));
  INV_X1     g08194(.I(new_n11175_), .ZN(new_n11176_));
  INV_X1     g08195(.I(new_n11163_), .ZN(new_n11177_));
  NAND4_X1   g08196(.A1(new_n11177_), .A2(pi0058), .A3(new_n7579_), .A4(new_n11156_), .ZN(new_n11178_));
  NOR3_X1    g08197(.A1(new_n11178_), .A2(new_n2437_), .A3(new_n3138_), .ZN(new_n11179_));
  NOR2_X1    g08198(.A1(new_n11179_), .A2(new_n11176_), .ZN(new_n11180_));
  NAND2_X1   g08199(.A1(new_n11174_), .A2(new_n11180_), .ZN(new_n11181_));
  NOR2_X1    g08200(.A1(new_n11181_), .A2(new_n11162_), .ZN(new_n11182_));
  NOR2_X1    g08201(.A1(new_n11182_), .A2(new_n5373_), .ZN(new_n11183_));
  INV_X1     g08202(.I(new_n11183_), .ZN(new_n11184_));
  NAND3_X1   g08203(.A1(new_n9429_), .A2(pi0024), .A3(pi0314), .ZN(new_n11185_));
  NOR3_X1    g08204(.A1(new_n9434_), .A2(new_n7272_), .A3(new_n9231_), .ZN(new_n11186_));
  XOR2_X1    g08205(.A1(new_n11186_), .A2(new_n11185_), .Z(new_n11187_));
  NOR2_X1    g08206(.A1(new_n11187_), .A2(new_n2481_), .ZN(new_n11188_));
  INV_X1     g08207(.I(new_n11188_), .ZN(new_n11189_));
  AOI21_X1   g08208(.A1(new_n11189_), .A2(new_n2437_), .B(new_n5625_), .ZN(new_n11190_));
  INV_X1     g08209(.I(new_n11190_), .ZN(new_n11191_));
  NOR2_X1    g08210(.A1(new_n11191_), .A2(new_n5386_), .ZN(new_n11192_));
  INV_X1     g08211(.I(new_n11192_), .ZN(new_n11193_));
  NAND2_X1   g08212(.A1(new_n11193_), .A2(new_n11184_), .ZN(new_n11194_));
  INV_X1     g08213(.I(new_n11182_), .ZN(new_n11195_));
  NOR2_X1    g08214(.A1(new_n8480_), .A2(new_n2437_), .ZN(new_n11196_));
  NAND3_X1   g08215(.A1(new_n11187_), .A2(new_n2702_), .A3(new_n6368_), .ZN(new_n11197_));
  NAND2_X1   g08216(.A1(new_n11197_), .A2(new_n7322_), .ZN(new_n11198_));
  NOR2_X1    g08217(.A1(new_n11198_), .A2(new_n11196_), .ZN(new_n11199_));
  NAND2_X1   g08218(.A1(new_n11199_), .A2(new_n5373_), .ZN(new_n11200_));
  OAI21_X1   g08219(.A1(new_n5373_), .A2(new_n11195_), .B(new_n11200_), .ZN(new_n11201_));
  NOR2_X1    g08220(.A1(new_n11201_), .A2(new_n7793_), .ZN(new_n11202_));
  NOR2_X1    g08221(.A1(new_n7793_), .A2(new_n2847_), .ZN(new_n11203_));
  XOR2_X1    g08222(.A1(new_n11202_), .A2(new_n11203_), .Z(new_n11204_));
  NOR2_X1    g08223(.A1(new_n11175_), .A2(new_n5386_), .ZN(new_n11205_));
  NOR2_X1    g08224(.A1(new_n11162_), .A2(new_n11176_), .ZN(new_n11206_));
  INV_X1     g08225(.I(new_n11206_), .ZN(new_n11207_));
  NOR2_X1    g08226(.A1(new_n11173_), .A2(new_n11207_), .ZN(new_n11208_));
  NOR2_X1    g08227(.A1(new_n11208_), .A2(new_n5373_), .ZN(new_n11209_));
  NOR2_X1    g08228(.A1(new_n11209_), .A2(new_n11205_), .ZN(new_n11210_));
  INV_X1     g08229(.I(new_n11210_), .ZN(new_n11211_));
  AOI21_X1   g08230(.A1(new_n11174_), .A2(new_n11175_), .B(new_n5386_), .ZN(new_n11212_));
  INV_X1     g08231(.I(new_n11212_), .ZN(new_n11213_));
  NOR2_X1    g08232(.A1(new_n11213_), .A2(pi0146), .ZN(new_n11214_));
  NOR2_X1    g08233(.A1(new_n11166_), .A2(pi0051), .ZN(new_n11215_));
  NOR2_X1    g08234(.A1(new_n3304_), .A2(new_n5386_), .ZN(new_n11216_));
  INV_X1     g08235(.I(new_n11216_), .ZN(new_n11217_));
  NAND2_X1   g08236(.A1(new_n11172_), .A2(new_n5373_), .ZN(new_n11218_));
  XOR2_X1    g08237(.A1(new_n11218_), .A2(new_n11217_), .Z(new_n11219_));
  NAND2_X1   g08238(.A1(new_n11219_), .A2(new_n11215_), .ZN(new_n11220_));
  INV_X1     g08239(.I(new_n11220_), .ZN(new_n11221_));
  AOI21_X1   g08240(.A1(new_n11221_), .A2(pi0146), .B(new_n11214_), .ZN(new_n11222_));
  INV_X1     g08241(.I(new_n11181_), .ZN(new_n11223_));
  NOR3_X1    g08242(.A1(new_n11223_), .A2(pi0051), .A3(new_n5386_), .ZN(new_n11224_));
  NOR2_X1    g08243(.A1(new_n11183_), .A2(new_n11224_), .ZN(new_n11225_));
  NAND2_X1   g08244(.A1(new_n11225_), .A2(new_n7811_), .ZN(new_n11226_));
  AOI21_X1   g08245(.A1(new_n11226_), .A2(new_n11222_), .B(new_n11211_), .ZN(new_n11227_));
  NOR3_X1    g08246(.A1(new_n11227_), .A2(pi0156), .A3(pi0161), .ZN(new_n11228_));
  NOR2_X1    g08247(.A1(new_n5386_), .A2(new_n2702_), .ZN(new_n11229_));
  INV_X1     g08248(.I(new_n11229_), .ZN(new_n11230_));
  NOR2_X1    g08249(.A1(new_n11230_), .A2(pi0146), .ZN(new_n11231_));
  INV_X1     g08250(.I(new_n11231_), .ZN(new_n11232_));
  NAND3_X1   g08251(.A1(new_n11195_), .A2(new_n7792_), .A3(new_n11232_), .ZN(new_n11233_));
  OAI21_X1   g08252(.A1(new_n11228_), .A2(new_n11233_), .B(new_n4981_), .ZN(new_n11234_));
  AOI21_X1   g08253(.A1(new_n11204_), .A2(new_n11194_), .B(new_n11234_), .ZN(new_n11235_));
  NAND2_X1   g08254(.A1(new_n9434_), .A2(new_n2480_), .ZN(new_n11236_));
  NAND2_X1   g08255(.A1(new_n2480_), .A2(pi0024), .ZN(new_n11237_));
  XOR2_X1    g08256(.A1(new_n11236_), .A2(new_n11237_), .Z(new_n11238_));
  NAND2_X1   g08257(.A1(new_n11238_), .A2(new_n9428_), .ZN(new_n11239_));
  AOI21_X1   g08258(.A1(new_n11239_), .A2(new_n2437_), .B(new_n5625_), .ZN(new_n11240_));
  INV_X1     g08259(.I(new_n11240_), .ZN(new_n11241_));
  NOR2_X1    g08260(.A1(new_n11241_), .A2(new_n5386_), .ZN(new_n11242_));
  NOR2_X1    g08261(.A1(new_n11242_), .A2(new_n11183_), .ZN(new_n11243_));
  INV_X1     g08262(.I(new_n11196_), .ZN(new_n11244_));
  NOR2_X1    g08263(.A1(new_n11239_), .A2(new_n11217_), .ZN(new_n11245_));
  NAND2_X1   g08264(.A1(new_n11245_), .A2(new_n5373_), .ZN(new_n11246_));
  AOI21_X1   g08265(.A1(new_n11246_), .A2(new_n2702_), .B(new_n11244_), .ZN(new_n11247_));
  NAND2_X1   g08266(.A1(new_n11247_), .A2(new_n11184_), .ZN(new_n11248_));
  NAND2_X1   g08267(.A1(new_n11248_), .A2(new_n7811_), .ZN(new_n11249_));
  NOR2_X1    g08268(.A1(new_n7812_), .A2(new_n2847_), .ZN(new_n11250_));
  XOR2_X1    g08269(.A1(new_n11249_), .A2(new_n11250_), .Z(new_n11251_));
  NOR3_X1    g08270(.A1(new_n11235_), .A2(new_n11243_), .A3(new_n11251_), .ZN(new_n11252_));
  NAND2_X1   g08271(.A1(pi0142), .A2(pi0144), .ZN(new_n11253_));
  NAND2_X1   g08272(.A1(new_n11248_), .A2(pi0142), .ZN(new_n11254_));
  XNOR2_X1   g08273(.A1(new_n11254_), .A2(new_n11253_), .ZN(new_n11255_));
  NOR2_X1    g08274(.A1(new_n11255_), .A2(new_n11243_), .ZN(new_n11256_));
  NAND2_X1   g08275(.A1(new_n9545_), .A2(new_n5642_), .ZN(new_n11257_));
  NOR2_X1    g08276(.A1(new_n11213_), .A2(pi0142), .ZN(new_n11258_));
  AOI21_X1   g08277(.A1(new_n11221_), .A2(pi0142), .B(new_n11258_), .ZN(new_n11259_));
  NAND2_X1   g08278(.A1(new_n11225_), .A2(pi0144), .ZN(new_n11260_));
  AOI21_X1   g08279(.A1(new_n11260_), .A2(new_n11259_), .B(new_n11211_), .ZN(new_n11261_));
  OAI21_X1   g08280(.A1(new_n11256_), .A2(new_n11257_), .B(new_n11261_), .ZN(new_n11262_));
  NOR2_X1    g08281(.A1(new_n11196_), .A2(new_n5386_), .ZN(new_n11263_));
  NAND2_X1   g08282(.A1(new_n11182_), .A2(new_n11229_), .ZN(new_n11264_));
  XOR2_X1    g08283(.A1(new_n11264_), .A2(new_n11263_), .Z(new_n11265_));
  NOR2_X1    g08284(.A1(new_n11265_), .A2(pi0144), .ZN(new_n11266_));
  INV_X1     g08285(.I(new_n11179_), .ZN(new_n11267_));
  NAND2_X1   g08286(.A1(new_n11210_), .A2(new_n11267_), .ZN(new_n11268_));
  NOR2_X1    g08287(.A1(new_n11268_), .A2(new_n7969_), .ZN(new_n11269_));
  OAI21_X1   g08288(.A1(new_n11266_), .A2(new_n11269_), .B(pi0180), .ZN(new_n11270_));
  AOI21_X1   g08289(.A1(new_n11270_), .A2(new_n11230_), .B(new_n3089_), .ZN(new_n11271_));
  INV_X1     g08290(.I(new_n11265_), .ZN(new_n11272_));
  NAND4_X1   g08291(.A1(new_n2554_), .A2(new_n2702_), .A3(new_n9252_), .A4(new_n11158_), .ZN(new_n11273_));
  NOR2_X1    g08292(.A1(new_n11273_), .A2(new_n11217_), .ZN(new_n11274_));
  INV_X1     g08293(.I(new_n11274_), .ZN(new_n11275_));
  NAND2_X1   g08294(.A1(new_n11272_), .A2(new_n11275_), .ZN(new_n11276_));
  NAND2_X1   g08295(.A1(new_n11276_), .A2(pi0142), .ZN(new_n11277_));
  XNOR2_X1   g08296(.A1(new_n11277_), .A2(new_n11253_), .ZN(new_n11278_));
  OAI21_X1   g08297(.A1(new_n11230_), .A2(pi0142), .B(pi0144), .ZN(new_n11279_));
  OAI21_X1   g08298(.A1(new_n5642_), .A2(new_n11279_), .B(new_n11268_), .ZN(new_n11280_));
  NAND2_X1   g08299(.A1(new_n11273_), .A2(new_n2437_), .ZN(new_n11281_));
  NAND2_X1   g08300(.A1(new_n5561_), .A2(new_n11281_), .ZN(new_n11282_));
  OAI21_X1   g08301(.A1(new_n5386_), .A2(new_n11282_), .B(new_n11184_), .ZN(new_n11283_));
  NAND4_X1   g08302(.A1(new_n11283_), .A2(new_n11280_), .A3(pi0299), .A4(new_n11162_), .ZN(new_n11284_));
  NOR2_X1    g08303(.A1(new_n11278_), .A2(new_n11284_), .ZN(new_n11285_));
  OAI21_X1   g08304(.A1(pi0179), .A2(new_n11271_), .B(new_n11285_), .ZN(new_n11286_));
  NAND2_X1   g08305(.A1(new_n11286_), .A2(new_n11262_), .ZN(new_n11287_));
  NOR2_X1    g08306(.A1(new_n11201_), .A2(new_n3089_), .ZN(new_n11288_));
  XNOR2_X1   g08307(.A1(new_n11288_), .A2(new_n11253_), .ZN(new_n11289_));
  AOI21_X1   g08308(.A1(new_n11289_), .A2(new_n11194_), .B(pi0180), .ZN(new_n11290_));
  NOR3_X1    g08309(.A1(new_n11290_), .A2(new_n11195_), .A3(new_n11279_), .ZN(new_n11291_));
  AOI21_X1   g08310(.A1(new_n11287_), .A2(new_n11291_), .B(new_n11252_), .ZN(new_n11292_));
  INV_X1     g08311(.I(new_n11205_), .ZN(new_n11293_));
  NOR2_X1    g08312(.A1(new_n2702_), .A2(new_n3089_), .ZN(new_n11294_));
  NOR2_X1    g08313(.A1(new_n11293_), .A2(new_n11294_), .ZN(new_n11295_));
  NAND2_X1   g08314(.A1(new_n11295_), .A2(new_n11279_), .ZN(new_n11296_));
  NOR2_X1    g08315(.A1(new_n11231_), .A2(new_n4981_), .ZN(new_n11297_));
  NOR2_X1    g08316(.A1(new_n2702_), .A2(new_n2847_), .ZN(new_n11298_));
  OAI21_X1   g08317(.A1(new_n11297_), .A2(new_n11205_), .B(new_n11298_), .ZN(new_n11299_));
  INV_X1     g08318(.I(new_n11299_), .ZN(new_n11300_));
  NAND3_X1   g08319(.A1(new_n11300_), .A2(pi0232), .A3(pi0299), .ZN(new_n11301_));
  NOR2_X1    g08320(.A1(new_n11300_), .A2(new_n5551_), .ZN(new_n11302_));
  NAND2_X1   g08321(.A1(new_n11302_), .A2(new_n6216_), .ZN(new_n11303_));
  AOI21_X1   g08322(.A1(new_n11303_), .A2(new_n11301_), .B(new_n11296_), .ZN(new_n11304_));
  INV_X1     g08323(.I(pi0133), .ZN(new_n11305_));
  INV_X1     g08324(.I(pi0121), .ZN(new_n11306_));
  INV_X1     g08325(.I(pi0126), .ZN(new_n11307_));
  INV_X1     g08326(.I(pi0132), .ZN(new_n11308_));
  INV_X1     g08327(.I(pi0130), .ZN(new_n11309_));
  INV_X1     g08328(.I(pi0134), .ZN(new_n11310_));
  INV_X1     g08329(.I(pi0135), .ZN(new_n11311_));
  INV_X1     g08330(.I(pi0136), .ZN(new_n11312_));
  NOR4_X1    g08331(.A1(new_n11309_), .A2(new_n11310_), .A3(new_n11311_), .A4(new_n11312_), .ZN(new_n11313_));
  INV_X1     g08332(.I(new_n11313_), .ZN(new_n11314_));
  NOR4_X1    g08333(.A1(new_n11314_), .A2(new_n11306_), .A3(new_n11307_), .A4(new_n11308_), .ZN(new_n11315_));
  NAND2_X1   g08334(.A1(new_n11315_), .A2(pi0121), .ZN(new_n11316_));
  XOR2_X1    g08335(.A1(new_n11316_), .A2(new_n11305_), .Z(new_n11317_));
  NOR2_X1    g08336(.A1(new_n9456_), .A2(new_n3098_), .ZN(new_n11318_));
  OAI21_X1   g08337(.A1(new_n9523_), .A2(new_n11318_), .B(new_n6493_), .ZN(new_n11319_));
  AOI22_X1   g08338(.A1(new_n11317_), .A2(pi0125), .B1(pi0087), .B2(new_n11319_), .ZN(new_n11320_));
  NOR2_X1    g08339(.A1(new_n3287_), .A2(pi0087), .ZN(new_n11321_));
  NAND2_X1   g08340(.A1(new_n11176_), .A2(new_n11321_), .ZN(new_n11322_));
  NOR2_X1    g08341(.A1(new_n11320_), .A2(new_n11322_), .ZN(new_n11323_));
  INV_X1     g08342(.I(new_n5827_), .ZN(new_n11324_));
  AND2_X2    g08343(.A1(new_n11259_), .A2(new_n7969_), .Z(new_n11325_));
  NAND2_X1   g08344(.A1(new_n5642_), .A2(pi0179), .ZN(new_n11326_));
  OAI21_X1   g08345(.A1(new_n11325_), .A2(new_n11326_), .B(new_n11279_), .ZN(new_n11327_));
  INV_X1     g08346(.I(new_n11215_), .ZN(new_n11328_));
  NOR2_X1    g08347(.A1(new_n11160_), .A2(new_n11167_), .ZN(new_n11329_));
  NOR2_X1    g08348(.A1(new_n11171_), .A2(new_n11156_), .ZN(new_n11330_));
  NAND2_X1   g08349(.A1(new_n11170_), .A2(new_n11330_), .ZN(new_n11331_));
  AOI21_X1   g08350(.A1(new_n11331_), .A2(new_n11329_), .B(new_n5386_), .ZN(new_n11332_));
  XOR2_X1    g08351(.A1(new_n11332_), .A2(new_n11217_), .Z(new_n11333_));
  NOR2_X1    g08352(.A1(new_n11333_), .A2(new_n11328_), .ZN(new_n11334_));
  INV_X1     g08353(.I(new_n11334_), .ZN(new_n11335_));
  INV_X1     g08354(.I(new_n11208_), .ZN(new_n11336_));
  NAND2_X1   g08355(.A1(new_n11336_), .A2(new_n5373_), .ZN(new_n11337_));
  NAND2_X1   g08356(.A1(new_n11337_), .A2(pi0142), .ZN(new_n11338_));
  XNOR2_X1   g08357(.A1(new_n11338_), .A2(new_n11253_), .ZN(new_n11339_));
  OAI21_X1   g08358(.A1(new_n11339_), .A2(new_n11335_), .B(new_n5642_), .ZN(new_n11340_));
  AOI21_X1   g08359(.A1(new_n11327_), .A2(new_n11245_), .B(new_n11340_), .ZN(new_n11341_));
  NAND2_X1   g08360(.A1(new_n11198_), .A2(new_n5373_), .ZN(new_n11342_));
  OAI21_X1   g08361(.A1(new_n11342_), .A2(new_n7969_), .B(new_n3089_), .ZN(new_n11343_));
  NAND2_X1   g08362(.A1(new_n11343_), .A2(pi0051), .ZN(new_n11344_));
  OAI21_X1   g08363(.A1(new_n11341_), .A2(new_n11344_), .B(new_n11324_), .ZN(new_n11345_));
  NOR2_X1    g08364(.A1(new_n11178_), .A2(new_n3304_), .ZN(new_n11346_));
  NOR4_X1    g08365(.A1(new_n11166_), .A2(pi0051), .A3(new_n5401_), .A4(new_n5386_), .ZN(new_n11347_));
  INV_X1     g08366(.I(new_n11295_), .ZN(new_n11348_));
  AOI21_X1   g08367(.A1(new_n11348_), .A2(new_n7969_), .B(new_n7451_), .ZN(new_n11349_));
  AOI21_X1   g08368(.A1(new_n11349_), .A2(new_n11347_), .B(pi0181), .ZN(new_n11350_));
  NOR2_X1    g08369(.A1(new_n5386_), .A2(pi0287), .ZN(new_n11351_));
  INV_X1     g08370(.I(new_n11351_), .ZN(new_n11352_));
  NOR2_X1    g08371(.A1(new_n7451_), .A2(new_n11352_), .ZN(new_n11353_));
  INV_X1     g08372(.I(new_n11353_), .ZN(new_n11354_));
  NOR3_X1    g08373(.A1(new_n11354_), .A2(new_n3145_), .A3(new_n3089_), .ZN(new_n11355_));
  NOR3_X1    g08374(.A1(new_n11354_), .A2(new_n3160_), .A3(pi0142), .ZN(new_n11356_));
  NOR3_X1    g08375(.A1(new_n8393_), .A2(new_n9008_), .A3(new_n11279_), .ZN(new_n11357_));
  OAI21_X1   g08376(.A1(new_n11355_), .A2(new_n11356_), .B(new_n11357_), .ZN(new_n11358_));
  OAI21_X1   g08377(.A1(new_n11350_), .A2(new_n11358_), .B(new_n3098_), .ZN(new_n11359_));
  NOR2_X1    g08378(.A1(new_n11296_), .A2(new_n5643_), .ZN(new_n11360_));
  INV_X1     g08379(.I(new_n8536_), .ZN(new_n11361_));
  NOR3_X1    g08380(.A1(new_n11300_), .A2(pi0159), .A3(new_n3098_), .ZN(new_n11362_));
  OAI21_X1   g08381(.A1(new_n11362_), .A2(new_n11361_), .B(new_n3259_), .ZN(new_n11363_));
  AOI21_X1   g08382(.A1(new_n11359_), .A2(new_n11360_), .B(new_n11363_), .ZN(new_n11364_));
  NOR2_X1    g08383(.A1(new_n11206_), .A2(new_n5386_), .ZN(new_n11365_));
  INV_X1     g08384(.I(new_n11365_), .ZN(new_n11366_));
  OAI21_X1   g08385(.A1(new_n11329_), .A2(pi0051), .B(new_n5373_), .ZN(new_n11367_));
  XOR2_X1    g08386(.A1(new_n11367_), .A2(new_n11217_), .Z(new_n11368_));
  NAND2_X1   g08387(.A1(new_n11368_), .A2(new_n11215_), .ZN(new_n11369_));
  NAND2_X1   g08388(.A1(new_n11369_), .A2(pi0142), .ZN(new_n11370_));
  XNOR2_X1   g08389(.A1(new_n11370_), .A2(new_n11253_), .ZN(new_n11371_));
  OAI21_X1   g08390(.A1(new_n11371_), .A2(new_n11366_), .B(new_n5642_), .ZN(new_n11372_));
  NOR2_X1    g08391(.A1(new_n11275_), .A2(new_n11279_), .ZN(new_n11373_));
  AOI21_X1   g08392(.A1(new_n11372_), .A2(new_n11373_), .B(pi0179), .ZN(new_n11374_));
  NOR2_X1    g08393(.A1(new_n11231_), .A2(pi0161), .ZN(new_n11375_));
  INV_X1     g08394(.I(new_n11375_), .ZN(new_n11376_));
  OAI21_X1   g08395(.A1(new_n11376_), .A2(new_n11347_), .B(new_n7440_), .ZN(new_n11377_));
  NOR2_X1    g08396(.A1(new_n8930_), .A2(new_n5386_), .ZN(new_n11378_));
  AND3_X2    g08397(.A1(new_n11378_), .A2(new_n11297_), .A3(new_n11377_), .Z(new_n11379_));
  NOR4_X1    g08398(.A1(new_n11296_), .A2(new_n5642_), .A3(new_n7440_), .A4(new_n11299_), .ZN(new_n11380_));
  OAI21_X1   g08399(.A1(new_n11379_), .A2(new_n8109_), .B(new_n11380_), .ZN(new_n11381_));
  NOR3_X1    g08400(.A1(new_n11374_), .A2(new_n11364_), .A3(new_n11381_), .ZN(new_n11382_));
  AOI21_X1   g08401(.A1(new_n11345_), .A2(new_n11382_), .B(pi0156), .ZN(new_n11383_));
  NAND2_X1   g08402(.A1(new_n11337_), .A2(pi0146), .ZN(new_n11384_));
  XNOR2_X1   g08403(.A1(new_n11384_), .A2(new_n7993_), .ZN(new_n11385_));
  NOR2_X1    g08404(.A1(new_n11335_), .A2(new_n7812_), .ZN(new_n11386_));
  AOI21_X1   g08405(.A1(new_n11385_), .A2(new_n11386_), .B(pi0161), .ZN(new_n11387_));
  INV_X1     g08406(.I(new_n11342_), .ZN(new_n11388_));
  OAI21_X1   g08407(.A1(new_n2702_), .A2(new_n2847_), .B(new_n11388_), .ZN(new_n11389_));
  OAI21_X1   g08408(.A1(new_n11389_), .A2(new_n11387_), .B(new_n5551_), .ZN(new_n11390_));
  NOR2_X1    g08409(.A1(new_n11245_), .A2(new_n4981_), .ZN(new_n11391_));
  NOR3_X1    g08410(.A1(new_n11222_), .A2(new_n4981_), .A3(new_n11232_), .ZN(new_n11392_));
  XOR2_X1    g08411(.A1(new_n11392_), .A2(new_n11391_), .Z(new_n11393_));
  NAND2_X1   g08412(.A1(new_n11369_), .A2(pi0146), .ZN(new_n11394_));
  XOR2_X1    g08413(.A1(new_n11394_), .A2(new_n7993_), .Z(new_n11395_));
  NOR3_X1    g08414(.A1(new_n11395_), .A2(new_n7812_), .A3(new_n11366_), .ZN(new_n11396_));
  OAI21_X1   g08415(.A1(new_n11396_), .A2(new_n11297_), .B(new_n11274_), .ZN(new_n11397_));
  OAI21_X1   g08416(.A1(new_n11304_), .A2(new_n3259_), .B(new_n3462_), .ZN(new_n11398_));
  NAND3_X1   g08417(.A1(new_n11398_), .A2(new_n9505_), .A3(new_n3212_), .ZN(new_n11399_));
  INV_X1     g08418(.I(new_n11304_), .ZN(new_n11400_));
  NOR2_X1    g08419(.A1(new_n11400_), .A2(new_n3462_), .ZN(new_n11401_));
  NOR2_X1    g08420(.A1(new_n11401_), .A2(new_n3207_), .ZN(new_n11402_));
  NAND2_X1   g08421(.A1(new_n7792_), .A2(pi0158), .ZN(new_n11403_));
  NOR4_X1    g08422(.A1(new_n11402_), .A2(new_n3098_), .A3(new_n11300_), .A4(new_n11403_), .ZN(new_n11404_));
  NAND2_X1   g08423(.A1(new_n11404_), .A2(new_n11399_), .ZN(new_n11405_));
  AOI21_X1   g08424(.A1(new_n11397_), .A2(new_n5551_), .B(new_n11405_), .ZN(new_n11406_));
  NAND3_X1   g08425(.A1(new_n11390_), .A2(new_n11406_), .A3(new_n11393_), .ZN(new_n11407_));
  INV_X1     g08426(.I(new_n11321_), .ZN(new_n11408_));
  NOR3_X1    g08427(.A1(new_n11400_), .A2(new_n11320_), .A3(new_n11408_), .ZN(new_n11409_));
  OAI21_X1   g08428(.A1(new_n11383_), .A2(new_n11407_), .B(new_n11409_), .ZN(new_n11410_));
  NAND2_X1   g08429(.A1(new_n11317_), .A2(pi0125), .ZN(new_n11411_));
  NOR2_X1    g08430(.A1(new_n5386_), .A2(new_n9456_), .ZN(new_n11412_));
  NOR2_X1    g08431(.A1(new_n3455_), .A2(new_n5551_), .ZN(new_n11413_));
  XOR2_X1    g08432(.A1(new_n11302_), .A2(new_n11413_), .Z(new_n11414_));
  NAND2_X1   g08433(.A1(new_n11414_), .A2(new_n11412_), .ZN(new_n11415_));
  NOR2_X1    g08434(.A1(new_n11176_), .A2(pi0087), .ZN(new_n11416_));
  INV_X1     g08435(.I(new_n11416_), .ZN(new_n11417_));
  NOR4_X1    g08436(.A1(new_n11415_), .A2(po1038), .A3(new_n11411_), .A4(new_n11417_), .ZN(new_n11418_));
  AOI22_X1   g08437(.A1(new_n11410_), .A2(new_n11418_), .B1(new_n11304_), .B2(new_n11323_), .ZN(new_n11419_));
  NAND2_X1   g08438(.A1(new_n3183_), .A2(new_n5551_), .ZN(new_n11420_));
  AOI21_X1   g08439(.A1(new_n11299_), .A2(new_n11176_), .B(new_n3361_), .ZN(new_n11421_));
  NOR2_X1    g08440(.A1(new_n11346_), .A2(new_n11176_), .ZN(new_n11422_));
  INV_X1     g08441(.I(new_n11422_), .ZN(new_n11423_));
  AOI21_X1   g08442(.A1(new_n11423_), .A2(new_n11232_), .B(new_n4981_), .ZN(new_n11424_));
  NOR2_X1    g08443(.A1(new_n11423_), .A2(new_n5373_), .ZN(new_n11425_));
  NOR2_X1    g08444(.A1(new_n8393_), .A2(new_n9008_), .ZN(new_n11426_));
  NOR2_X1    g08445(.A1(new_n11426_), .A2(pi0051), .ZN(new_n11427_));
  INV_X1     g08446(.I(new_n11427_), .ZN(new_n11428_));
  NOR2_X1    g08447(.A1(new_n11428_), .A2(new_n5386_), .ZN(new_n11429_));
  NOR2_X1    g08448(.A1(new_n11425_), .A2(new_n11429_), .ZN(new_n11430_));
  NOR2_X1    g08449(.A1(new_n11425_), .A2(new_n5949_), .ZN(new_n11431_));
  NAND2_X1   g08450(.A1(new_n11431_), .A2(pi0146), .ZN(new_n11432_));
  XOR2_X1    g08451(.A1(new_n11432_), .A2(new_n7993_), .Z(new_n11433_));
  NOR2_X1    g08452(.A1(new_n11433_), .A2(new_n11430_), .ZN(new_n11434_));
  OAI21_X1   g08453(.A1(new_n11434_), .A2(new_n11424_), .B(new_n3361_), .ZN(new_n11435_));
  NAND3_X1   g08454(.A1(new_n11435_), .A2(new_n5551_), .A3(new_n8178_), .ZN(new_n11436_));
  NAND2_X1   g08455(.A1(new_n11436_), .A2(new_n11421_), .ZN(new_n11437_));
  INV_X1     g08456(.I(new_n11346_), .ZN(new_n11438_));
  OAI22_X1   g08457(.A1(new_n11175_), .A2(new_n11420_), .B1(new_n5825_), .B2(new_n6545_), .ZN(new_n11439_));
  NOR2_X1    g08458(.A1(new_n11438_), .A2(new_n11439_), .ZN(new_n11440_));
  INV_X1     g08459(.I(new_n11430_), .ZN(new_n11441_));
  NOR3_X1    g08460(.A1(new_n11431_), .A2(new_n3089_), .A3(new_n6544_), .ZN(new_n11442_));
  INV_X1     g08461(.I(new_n11431_), .ZN(new_n11443_));
  NOR3_X1    g08462(.A1(new_n11443_), .A2(pi0142), .A3(new_n6544_), .ZN(new_n11444_));
  OAI21_X1   g08463(.A1(new_n11444_), .A2(new_n11442_), .B(new_n11441_), .ZN(new_n11445_));
  AOI21_X1   g08464(.A1(new_n11422_), .A2(new_n2702_), .B(new_n11229_), .ZN(new_n11446_));
  AOI21_X1   g08465(.A1(new_n11229_), .A2(new_n3089_), .B(new_n11175_), .ZN(new_n11447_));
  NOR4_X1    g08466(.A1(new_n11446_), .A2(new_n7969_), .A3(new_n6544_), .A4(new_n11294_), .ZN(new_n11448_));
  NOR2_X1    g08467(.A1(new_n11328_), .A2(new_n5386_), .ZN(new_n11449_));
  NOR2_X1    g08468(.A1(new_n6544_), .A2(new_n7969_), .ZN(new_n11450_));
  OAI21_X1   g08469(.A1(new_n11447_), .A2(new_n11450_), .B(new_n11449_), .ZN(new_n11451_));
  INV_X1     g08470(.I(new_n11451_), .ZN(new_n11452_));
  OAI21_X1   g08471(.A1(new_n11448_), .A2(pi0181), .B(new_n11452_), .ZN(new_n11453_));
  OAI21_X1   g08472(.A1(new_n11445_), .A2(new_n11453_), .B(new_n3098_), .ZN(new_n11454_));
  INV_X1     g08473(.I(new_n11448_), .ZN(new_n11455_));
  INV_X1     g08474(.I(new_n11347_), .ZN(new_n11456_));
  NOR2_X1    g08475(.A1(new_n7450_), .A2(new_n11166_), .ZN(new_n11457_));
  NOR3_X1    g08476(.A1(new_n11348_), .A2(new_n11456_), .A3(new_n11457_), .ZN(new_n11458_));
  NOR2_X1    g08477(.A1(new_n11455_), .A2(new_n11458_), .ZN(new_n11459_));
  NOR2_X1    g08478(.A1(new_n11352_), .A2(pi0051), .ZN(new_n11460_));
  NOR2_X1    g08479(.A1(new_n11441_), .A2(new_n11460_), .ZN(new_n11461_));
  INV_X1     g08480(.I(new_n11461_), .ZN(new_n11462_));
  NAND2_X1   g08481(.A1(new_n11462_), .A2(new_n3100_), .ZN(new_n11463_));
  NOR3_X1    g08482(.A1(new_n11451_), .A2(new_n3089_), .A3(new_n11230_), .ZN(new_n11464_));
  AOI21_X1   g08483(.A1(new_n11463_), .A2(new_n11464_), .B(new_n7450_), .ZN(new_n11465_));
  NOR4_X1    g08484(.A1(new_n11465_), .A2(new_n11445_), .A3(new_n5643_), .A4(new_n11459_), .ZN(new_n11466_));
  AOI21_X1   g08485(.A1(new_n11466_), .A2(new_n11454_), .B(new_n11440_), .ZN(new_n11467_));
  NAND2_X1   g08486(.A1(new_n11437_), .A2(new_n11467_), .ZN(new_n11468_));
  NAND3_X1   g08487(.A1(new_n11461_), .A2(pi0161), .A3(new_n11231_), .ZN(new_n11469_));
  NAND3_X1   g08488(.A1(new_n11462_), .A2(pi0161), .A3(new_n11232_), .ZN(new_n11470_));
  NAND2_X1   g08489(.A1(new_n11470_), .A2(new_n11469_), .ZN(new_n11471_));
  AOI21_X1   g08490(.A1(new_n11346_), .A2(new_n11352_), .B(new_n11176_), .ZN(new_n11472_));
  INV_X1     g08491(.I(new_n11472_), .ZN(new_n11473_));
  NOR2_X1    g08492(.A1(new_n11473_), .A2(new_n3011_), .ZN(new_n11474_));
  NAND2_X1   g08493(.A1(new_n3362_), .A2(pi0216), .ZN(new_n11475_));
  AOI21_X1   g08494(.A1(new_n11471_), .A2(new_n11474_), .B(new_n11475_), .ZN(new_n11476_));
  OR2_X2     g08495(.A1(new_n11421_), .A2(new_n8110_), .Z(new_n11477_));
  AOI21_X1   g08496(.A1(new_n11476_), .A2(new_n11435_), .B(new_n11477_), .ZN(new_n11478_));
  AOI21_X1   g08497(.A1(new_n11468_), .A2(new_n11478_), .B(new_n11420_), .ZN(new_n11479_));
  NAND2_X1   g08498(.A1(new_n11182_), .A2(pi0038), .ZN(new_n11480_));
  OAI21_X1   g08499(.A1(new_n11479_), .A2(new_n11480_), .B(new_n7468_), .ZN(new_n11481_));
  NOR2_X1    g08500(.A1(new_n11267_), .A2(new_n11167_), .ZN(new_n11482_));
  INV_X1     g08501(.I(new_n11482_), .ZN(new_n11483_));
  NOR2_X1    g08502(.A1(new_n11483_), .A2(new_n11230_), .ZN(new_n11484_));
  INV_X1     g08503(.I(new_n11484_), .ZN(new_n11485_));
  NOR2_X1    g08504(.A1(new_n11485_), .A2(new_n11162_), .ZN(new_n11486_));
  OAI21_X1   g08505(.A1(new_n11176_), .A2(new_n11230_), .B(new_n4981_), .ZN(new_n11487_));
  AOI21_X1   g08506(.A1(new_n11486_), .A2(pi0146), .B(new_n11487_), .ZN(new_n11488_));
  NOR3_X1    g08507(.A1(new_n11488_), .A2(new_n5386_), .A3(new_n11195_), .ZN(new_n11489_));
  NAND2_X1   g08508(.A1(new_n11276_), .A2(pi0146), .ZN(new_n11490_));
  XNOR2_X1   g08509(.A1(new_n11490_), .A2(new_n7993_), .ZN(new_n11491_));
  AOI21_X1   g08510(.A1(new_n11491_), .A2(new_n11283_), .B(new_n11489_), .ZN(new_n11492_));
  NAND2_X1   g08511(.A1(new_n7811_), .A2(new_n7792_), .ZN(new_n11493_));
  OAI22_X1   g08512(.A1(new_n11492_), .A2(new_n11493_), .B1(new_n11272_), .B2(new_n11376_), .ZN(new_n11494_));
  NOR2_X1    g08513(.A1(new_n11195_), .A2(new_n5386_), .ZN(new_n11495_));
  AOI21_X1   g08514(.A1(new_n2702_), .A2(new_n5386_), .B(new_n11483_), .ZN(new_n11496_));
  OR2_X2     g08515(.A1(new_n11496_), .A2(pi0146), .Z(new_n11497_));
  AOI21_X1   g08516(.A1(new_n11495_), .A2(new_n11497_), .B(pi0161), .ZN(new_n11498_));
  NAND2_X1   g08517(.A1(new_n11175_), .A2(pi0100), .ZN(new_n11499_));
  NAND2_X1   g08518(.A1(new_n11499_), .A2(new_n3207_), .ZN(new_n11500_));
  INV_X1     g08519(.I(new_n11500_), .ZN(new_n11501_));
  NOR2_X1    g08520(.A1(new_n11401_), .A2(new_n11501_), .ZN(new_n11502_));
  NAND2_X1   g08521(.A1(new_n11400_), .A2(new_n3132_), .ZN(new_n11503_));
  NAND4_X1   g08522(.A1(new_n11503_), .A2(pi0146), .A3(pi0156), .A4(new_n11175_), .ZN(new_n11504_));
  NOR4_X1    g08523(.A1(new_n11498_), .A2(new_n11268_), .A3(new_n11502_), .A4(new_n11504_), .ZN(new_n11505_));
  NAND3_X1   g08524(.A1(new_n11494_), .A2(new_n11481_), .A3(new_n11505_), .ZN(new_n11506_));
  NOR3_X1    g08525(.A1(new_n11292_), .A2(new_n11419_), .A3(new_n11506_), .ZN(po0279));
  OR2_X2     g08526(.A1(new_n10914_), .A2(new_n6400_), .Z(new_n11509_));
  NOR2_X1    g08527(.A1(new_n9863_), .A2(po1038), .ZN(new_n11510_));
  AOI21_X1   g08528(.A1(new_n11509_), .A2(new_n11510_), .B(new_n6939_), .ZN(po0280));
  NOR4_X1    g08529(.A1(new_n5460_), .A2(new_n2665_), .A3(new_n3362_), .A4(new_n7589_), .ZN(new_n11512_));
  INV_X1     g08530(.I(new_n11512_), .ZN(new_n11513_));
  NAND3_X1   g08531(.A1(new_n9500_), .A2(pi0110), .A3(new_n6545_), .ZN(new_n11514_));
  OAI21_X1   g08532(.A1(new_n11514_), .A2(new_n6272_), .B(new_n3183_), .ZN(new_n11515_));
  NAND3_X1   g08533(.A1(new_n11515_), .A2(pi0299), .A3(new_n11512_), .ZN(new_n11516_));
  INV_X1     g08534(.I(pi0111), .ZN(new_n11517_));
  OAI21_X1   g08535(.A1(new_n2617_), .A2(new_n11517_), .B(new_n7361_), .ZN(new_n11518_));
  AOI21_X1   g08536(.A1(new_n11518_), .A2(new_n2605_), .B(new_n11517_), .ZN(new_n11519_));
  NAND2_X1   g08537(.A1(new_n5573_), .A2(new_n11519_), .ZN(new_n11520_));
  NOR2_X1    g08538(.A1(new_n11520_), .A2(new_n2606_), .ZN(new_n11521_));
  INV_X1     g08539(.I(new_n11521_), .ZN(new_n11522_));
  XOR2_X1    g08540(.A1(new_n11520_), .A2(new_n10237_), .Z(new_n11523_));
  NAND2_X1   g08541(.A1(new_n11523_), .A2(new_n2619_), .ZN(new_n11524_));
  INV_X1     g08542(.I(new_n11524_), .ZN(new_n11525_));
  AOI21_X1   g08543(.A1(new_n11525_), .A2(new_n11522_), .B(pi0083), .ZN(new_n11526_));
  OAI21_X1   g08544(.A1(new_n11522_), .A2(new_n11525_), .B(new_n11526_), .ZN(new_n11527_));
  AOI21_X1   g08545(.A1(pi0090), .A2(new_n2476_), .B(new_n9254_), .ZN(new_n11528_));
  NOR3_X1    g08546(.A1(new_n5580_), .A2(new_n11528_), .A3(new_n2628_), .ZN(new_n11529_));
  AND2_X2    g08547(.A1(new_n11527_), .A2(new_n11529_), .Z(new_n11530_));
  NOR2_X1    g08548(.A1(new_n8462_), .A2(new_n2679_), .ZN(new_n11531_));
  OAI21_X1   g08549(.A1(new_n11530_), .A2(new_n7406_), .B(new_n11531_), .ZN(new_n11532_));
  NOR2_X1    g08550(.A1(new_n2480_), .A2(pi0072), .ZN(new_n11533_));
  OAI21_X1   g08551(.A1(new_n10496_), .A2(new_n2665_), .B(new_n3138_), .ZN(new_n11534_));
  NAND2_X1   g08552(.A1(new_n11534_), .A2(new_n8461_), .ZN(new_n11535_));
  AOI21_X1   g08553(.A1(new_n11532_), .A2(new_n11533_), .B(new_n11535_), .ZN(new_n11536_));
  INV_X1     g08554(.I(new_n2680_), .ZN(new_n11537_));
  INV_X1     g08555(.I(new_n11530_), .ZN(new_n11538_));
  AOI21_X1   g08556(.A1(new_n11538_), .A2(new_n7406_), .B(new_n11537_), .ZN(new_n11539_));
  NAND2_X1   g08557(.A1(new_n5625_), .A2(new_n3183_), .ZN(new_n11540_));
  OAI21_X1   g08558(.A1(new_n11539_), .A2(new_n11540_), .B(new_n10495_), .ZN(new_n11541_));
  OAI21_X1   g08559(.A1(new_n11541_), .A2(new_n11536_), .B(new_n11516_), .ZN(new_n11542_));
  NOR2_X1    g08560(.A1(new_n3290_), .A2(pi0038), .ZN(new_n11543_));
  NAND2_X1   g08561(.A1(new_n11542_), .A2(new_n11543_), .ZN(new_n11544_));
  NAND2_X1   g08562(.A1(new_n11543_), .A2(po1038), .ZN(new_n11545_));
  XOR2_X1    g08563(.A1(new_n11544_), .A2(new_n11545_), .Z(new_n11546_));
  NAND4_X1   g08564(.A1(new_n11515_), .A2(pi0039), .A3(pi0299), .A4(new_n11512_), .ZN(new_n11547_));
  NAND2_X1   g08565(.A1(new_n5526_), .A2(new_n10447_), .ZN(new_n11548_));
  NAND2_X1   g08566(.A1(new_n8248_), .A2(new_n2665_), .ZN(new_n11549_));
  NOR2_X1    g08567(.A1(new_n2788_), .A2(new_n6494_), .ZN(new_n11550_));
  NAND4_X1   g08568(.A1(new_n10495_), .A2(new_n11548_), .A3(new_n11549_), .A4(new_n11550_), .ZN(new_n11551_));
  AOI21_X1   g08569(.A1(new_n11547_), .A2(new_n2665_), .B(new_n11551_), .ZN(new_n11552_));
  NAND2_X1   g08570(.A1(new_n11546_), .A2(new_n11552_), .ZN(new_n11553_));
  AOI21_X1   g08571(.A1(new_n11553_), .A2(new_n3183_), .B(new_n11513_), .ZN(po0281));
  INV_X1     g08572(.I(new_n11315_), .ZN(new_n11555_));
  INV_X1     g08573(.I(pi0125), .ZN(new_n11556_));
  NOR2_X1    g08574(.A1(new_n11556_), .A2(new_n11305_), .ZN(new_n11557_));
  NOR2_X1    g08575(.A1(pi0125), .A2(pi0133), .ZN(new_n11558_));
  AOI21_X1   g08576(.A1(new_n11555_), .A2(new_n11558_), .B(new_n11557_), .ZN(new_n11559_));
  INV_X1     g08577(.I(new_n11559_), .ZN(new_n11560_));
  NOR2_X1    g08578(.A1(new_n11230_), .A2(new_n3827_), .ZN(new_n11561_));
  AOI21_X1   g08579(.A1(new_n11449_), .A2(new_n5158_), .B(new_n11561_), .ZN(new_n11562_));
  AOI22_X1   g08580(.A1(new_n11560_), .A2(pi0232), .B1(new_n11175_), .B2(new_n11562_), .ZN(new_n11563_));
  NOR2_X1    g08581(.A1(new_n11230_), .A2(new_n7342_), .ZN(new_n11564_));
  NOR2_X1    g08582(.A1(new_n11564_), .A2(pi0299), .ZN(new_n11565_));
  NAND2_X1   g08583(.A1(new_n11449_), .A2(pi0174), .ZN(new_n11566_));
  OAI21_X1   g08584(.A1(new_n11566_), .A2(new_n11565_), .B(new_n5551_), .ZN(new_n11567_));
  NAND3_X1   g08585(.A1(new_n11567_), .A2(pi0299), .A3(new_n11562_), .ZN(new_n11568_));
  NOR2_X1    g08586(.A1(new_n11568_), .A2(new_n3462_), .ZN(new_n11569_));
  INV_X1     g08587(.I(new_n11569_), .ZN(new_n11570_));
  NOR2_X1    g08588(.A1(new_n11182_), .A2(new_n5386_), .ZN(new_n11571_));
  NOR2_X1    g08589(.A1(new_n11244_), .A2(new_n11230_), .ZN(new_n11572_));
  XNOR2_X1   g08590(.A1(new_n11571_), .A2(new_n11572_), .ZN(new_n11573_));
  INV_X1     g08591(.I(new_n11573_), .ZN(new_n11574_));
  NAND2_X1   g08592(.A1(new_n5158_), .A2(new_n5665_), .ZN(new_n11575_));
  OAI21_X1   g08593(.A1(new_n11574_), .A2(new_n11575_), .B(new_n11561_), .ZN(new_n11576_));
  NOR2_X1    g08594(.A1(new_n11244_), .A2(new_n5373_), .ZN(new_n11577_));
  NOR2_X1    g08595(.A1(new_n11224_), .A2(new_n11577_), .ZN(new_n11578_));
  INV_X1     g08596(.I(new_n11578_), .ZN(new_n11579_));
  NOR2_X1    g08597(.A1(new_n11242_), .A2(new_n11577_), .ZN(new_n11580_));
  NAND2_X1   g08598(.A1(new_n11580_), .A2(pi0152), .ZN(new_n11581_));
  XOR2_X1    g08599(.A1(new_n11581_), .A2(new_n7779_), .Z(new_n11582_));
  NOR2_X1    g08600(.A1(new_n11582_), .A2(new_n11579_), .ZN(new_n11583_));
  NAND2_X1   g08601(.A1(new_n8174_), .A2(new_n5665_), .ZN(new_n11584_));
  NOR2_X1    g08602(.A1(new_n11196_), .A2(new_n11229_), .ZN(new_n11585_));
  OAI21_X1   g08603(.A1(new_n11239_), .A2(new_n11217_), .B(new_n11585_), .ZN(new_n11586_));
  NAND2_X1   g08604(.A1(new_n11586_), .A2(pi0172), .ZN(new_n11587_));
  XOR2_X1    g08605(.A1(new_n11587_), .A2(new_n7779_), .Z(new_n11588_));
  NOR2_X1    g08606(.A1(new_n11282_), .A2(new_n5386_), .ZN(new_n11589_));
  NOR2_X1    g08607(.A1(new_n11577_), .A2(new_n11589_), .ZN(new_n11590_));
  INV_X1     g08608(.I(new_n11590_), .ZN(new_n11591_));
  NAND4_X1   g08609(.A1(new_n11591_), .A2(pi0152), .A3(pi0172), .A4(pi0197), .ZN(new_n11592_));
  NAND4_X1   g08610(.A1(new_n11590_), .A2(pi0152), .A3(new_n3827_), .A4(pi0197), .ZN(new_n11593_));
  NAND3_X1   g08611(.A1(new_n11585_), .A2(new_n8170_), .A3(new_n11275_), .ZN(new_n11594_));
  AOI21_X1   g08612(.A1(new_n11592_), .A2(new_n11593_), .B(new_n11594_), .ZN(new_n11595_));
  NOR2_X1    g08613(.A1(new_n11595_), .A2(new_n11561_), .ZN(new_n11596_));
  NOR2_X1    g08614(.A1(pi0152), .A2(pi0197), .ZN(new_n11597_));
  NOR2_X1    g08615(.A1(new_n11485_), .A2(new_n11181_), .ZN(new_n11598_));
  AOI21_X1   g08616(.A1(new_n5386_), .A2(new_n11244_), .B(new_n11598_), .ZN(new_n11599_));
  NAND2_X1   g08617(.A1(new_n11486_), .A2(new_n5373_), .ZN(new_n11600_));
  XNOR2_X1   g08618(.A1(new_n11600_), .A2(new_n11263_), .ZN(new_n11601_));
  NAND3_X1   g08619(.A1(new_n11601_), .A2(new_n11599_), .A3(pi0051), .ZN(new_n11602_));
  NOR4_X1    g08620(.A1(new_n11588_), .A2(new_n11596_), .A3(new_n11597_), .A4(new_n11602_), .ZN(new_n11603_));
  OAI21_X1   g08621(.A1(new_n11583_), .A2(new_n11584_), .B(new_n11603_), .ZN(new_n11604_));
  NOR2_X1    g08622(.A1(new_n11192_), .A2(new_n11577_), .ZN(new_n11605_));
  NAND2_X1   g08623(.A1(new_n11605_), .A2(pi0152), .ZN(new_n11606_));
  XOR2_X1    g08624(.A1(new_n11606_), .A2(new_n7779_), .Z(new_n11607_));
  NOR2_X1    g08625(.A1(new_n11388_), .A2(new_n11196_), .ZN(new_n11608_));
  OR3_X2     g08626(.A1(new_n11607_), .A2(new_n3259_), .A3(new_n11608_), .Z(new_n11609_));
  AOI21_X1   g08627(.A1(new_n11604_), .A2(new_n11576_), .B(new_n11609_), .ZN(new_n11610_));
  NOR2_X1    g08628(.A1(new_n5641_), .A2(new_n7342_), .ZN(new_n11611_));
  NAND2_X1   g08629(.A1(new_n11608_), .A2(pi0193), .ZN(new_n11612_));
  XOR2_X1    g08630(.A1(new_n11612_), .A2(new_n11611_), .Z(new_n11613_));
  INV_X1     g08631(.I(new_n8011_), .ZN(new_n11614_));
  NOR3_X1    g08632(.A1(new_n11579_), .A2(new_n5641_), .A3(new_n7342_), .ZN(new_n11615_));
  NOR3_X1    g08633(.A1(new_n11578_), .A2(pi0145), .A3(new_n7342_), .ZN(new_n11616_));
  OAI21_X1   g08634(.A1(new_n11615_), .A2(new_n11616_), .B(new_n11599_), .ZN(new_n11617_));
  NAND3_X1   g08635(.A1(new_n11617_), .A2(new_n7378_), .A3(new_n11614_), .ZN(new_n11618_));
  NOR3_X1    g08636(.A1(new_n11574_), .A2(new_n5641_), .A3(new_n11564_), .ZN(new_n11619_));
  AOI21_X1   g08637(.A1(new_n11618_), .A2(new_n11619_), .B(pi0174), .ZN(new_n11620_));
  OAI21_X1   g08638(.A1(new_n11613_), .A2(new_n11586_), .B(new_n11620_), .ZN(new_n11621_));
  INV_X1     g08639(.I(new_n11605_), .ZN(new_n11622_));
  NAND3_X1   g08640(.A1(new_n11622_), .A2(pi0145), .A3(pi0193), .ZN(new_n11623_));
  NAND3_X1   g08641(.A1(new_n11605_), .A2(pi0145), .A3(new_n7342_), .ZN(new_n11624_));
  AOI21_X1   g08642(.A1(new_n11623_), .A2(new_n11624_), .B(new_n11580_), .ZN(new_n11625_));
  AOI21_X1   g08643(.A1(new_n11621_), .A2(new_n11625_), .B(new_n8017_), .ZN(new_n11626_));
  NAND3_X1   g08644(.A1(new_n11591_), .A2(pi0145), .A3(pi0174), .ZN(new_n11627_));
  NAND3_X1   g08645(.A1(new_n11590_), .A2(new_n5641_), .A3(pi0174), .ZN(new_n11628_));
  AOI21_X1   g08646(.A1(new_n11627_), .A2(new_n11628_), .B(new_n11244_), .ZN(new_n11629_));
  NAND2_X1   g08647(.A1(new_n11484_), .A2(pi0145), .ZN(new_n11630_));
  AOI21_X1   g08648(.A1(new_n11630_), .A2(new_n11230_), .B(new_n11161_), .ZN(new_n11631_));
  NOR2_X1    g08649(.A1(new_n11244_), .A2(new_n5386_), .ZN(new_n11632_));
  OAI21_X1   g08650(.A1(new_n11631_), .A2(pi0174), .B(new_n11632_), .ZN(new_n11633_));
  NOR3_X1    g08651(.A1(new_n11244_), .A2(new_n11275_), .A3(new_n5641_), .ZN(new_n11634_));
  NOR3_X1    g08652(.A1(new_n11196_), .A2(pi0145), .A3(new_n11275_), .ZN(new_n11635_));
  NOR2_X1    g08653(.A1(new_n7378_), .A2(new_n7342_), .ZN(new_n11636_));
  INV_X1     g08654(.I(new_n11636_), .ZN(new_n11637_));
  NOR2_X1    g08655(.A1(new_n11230_), .A2(new_n11637_), .ZN(new_n11638_));
  OAI21_X1   g08656(.A1(new_n11634_), .A2(new_n11635_), .B(new_n11638_), .ZN(new_n11639_));
  AOI21_X1   g08657(.A1(new_n11633_), .A2(new_n7342_), .B(new_n11639_), .ZN(new_n11640_));
  NOR2_X1    g08658(.A1(new_n5641_), .A2(new_n7378_), .ZN(new_n11641_));
  NAND2_X1   g08659(.A1(new_n11601_), .A2(pi0051), .ZN(new_n11642_));
  NAND2_X1   g08660(.A1(new_n11642_), .A2(pi0145), .ZN(new_n11643_));
  XOR2_X1    g08661(.A1(new_n11643_), .A2(new_n11641_), .Z(new_n11644_));
  NOR2_X1    g08662(.A1(new_n11496_), .A2(new_n11577_), .ZN(new_n11645_));
  INV_X1     g08663(.I(new_n11645_), .ZN(new_n11646_));
  NOR3_X1    g08664(.A1(new_n11644_), .A2(new_n3098_), .A3(new_n11646_), .ZN(new_n11647_));
  OAI21_X1   g08665(.A1(new_n11629_), .A2(new_n11640_), .B(new_n11647_), .ZN(new_n11648_));
  OAI21_X1   g08666(.A1(new_n11626_), .A2(new_n11648_), .B(new_n7467_), .ZN(new_n11649_));
  NOR2_X1    g08667(.A1(new_n11347_), .A2(new_n5158_), .ZN(new_n11650_));
  XOR2_X1    g08668(.A1(new_n11650_), .A2(new_n7779_), .Z(new_n11651_));
  NAND2_X1   g08669(.A1(new_n11378_), .A2(new_n11651_), .ZN(new_n11652_));
  NAND3_X1   g08670(.A1(new_n11652_), .A2(new_n3011_), .A3(new_n3362_), .ZN(new_n11653_));
  NAND2_X1   g08671(.A1(new_n11426_), .A2(new_n11351_), .ZN(new_n11654_));
  NAND2_X1   g08672(.A1(new_n11654_), .A2(new_n11230_), .ZN(new_n11655_));
  INV_X1     g08673(.I(new_n11655_), .ZN(new_n11656_));
  AOI21_X1   g08674(.A1(new_n11346_), .A2(new_n11351_), .B(new_n11205_), .ZN(new_n11657_));
  NOR2_X1    g08675(.A1(new_n11657_), .A2(new_n3827_), .ZN(new_n11658_));
  XOR2_X1    g08676(.A1(new_n11658_), .A2(new_n7779_), .Z(new_n11659_));
  NAND3_X1   g08677(.A1(new_n11659_), .A2(new_n11653_), .A3(new_n11656_), .ZN(new_n11660_));
  NOR2_X1    g08678(.A1(new_n11422_), .A2(pi0051), .ZN(new_n11661_));
  INV_X1     g08679(.I(new_n11661_), .ZN(new_n11662_));
  NOR2_X1    g08680(.A1(new_n3160_), .A2(new_n5373_), .ZN(new_n11663_));
  AOI21_X1   g08681(.A1(new_n11662_), .A2(new_n5373_), .B(new_n11663_), .ZN(new_n11664_));
  INV_X1     g08682(.I(new_n11664_), .ZN(new_n11665_));
  NOR2_X1    g08683(.A1(new_n11347_), .A2(new_n6544_), .ZN(new_n11666_));
  XOR2_X1    g08684(.A1(new_n11666_), .A2(new_n7450_), .Z(new_n11667_));
  AOI22_X1   g08685(.A1(new_n11665_), .A2(new_n11667_), .B1(new_n6544_), .B2(new_n11449_), .ZN(new_n11668_));
  NOR2_X1    g08686(.A1(new_n11668_), .A2(new_n7378_), .ZN(new_n11669_));
  XOR2_X1    g08687(.A1(new_n11669_), .A2(new_n11637_), .Z(new_n11670_));
  NOR2_X1    g08688(.A1(new_n3145_), .A2(new_n6461_), .ZN(new_n11671_));
  AOI21_X1   g08689(.A1(new_n6461_), .A2(new_n11293_), .B(new_n11665_), .ZN(new_n11672_));
  NOR2_X1    g08690(.A1(new_n11672_), .A2(new_n7378_), .ZN(new_n11673_));
  NAND2_X1   g08691(.A1(new_n11564_), .A2(pi0174), .ZN(new_n11674_));
  XNOR2_X1   g08692(.A1(new_n11673_), .A2(new_n11674_), .ZN(new_n11675_));
  NAND2_X1   g08693(.A1(new_n11675_), .A2(new_n11671_), .ZN(new_n11676_));
  AOI21_X1   g08694(.A1(new_n11676_), .A2(new_n5642_), .B(pi0299), .ZN(new_n11677_));
  NOR2_X1    g08695(.A1(new_n11429_), .A2(new_n11663_), .ZN(new_n11678_));
  AOI21_X1   g08696(.A1(new_n11656_), .A2(pi0224), .B(new_n6544_), .ZN(new_n11679_));
  AOI21_X1   g08697(.A1(new_n11679_), .A2(new_n11229_), .B(new_n6459_), .ZN(new_n11680_));
  NOR2_X1    g08698(.A1(new_n11680_), .A2(new_n11678_), .ZN(new_n11681_));
  INV_X1     g08699(.I(new_n11681_), .ZN(new_n11682_));
  NOR2_X1    g08700(.A1(new_n11423_), .A2(new_n5386_), .ZN(new_n11683_));
  NOR2_X1    g08701(.A1(new_n11683_), .A2(new_n11663_), .ZN(new_n11684_));
  INV_X1     g08702(.I(new_n11684_), .ZN(new_n11685_));
  NAND2_X1   g08703(.A1(new_n11438_), .A2(new_n7451_), .ZN(new_n11686_));
  NAND2_X1   g08704(.A1(new_n11686_), .A2(new_n11351_), .ZN(new_n11687_));
  AOI22_X1   g08705(.A1(new_n11685_), .A2(new_n6459_), .B1(new_n11293_), .B2(new_n11687_), .ZN(new_n11688_));
  NOR2_X1    g08706(.A1(new_n11688_), .A2(new_n7342_), .ZN(new_n11689_));
  XOR2_X1    g08707(.A1(new_n11689_), .A2(new_n11637_), .Z(new_n11690_));
  OAI21_X1   g08708(.A1(new_n11690_), .A2(new_n11682_), .B(new_n5642_), .ZN(new_n11691_));
  OAI21_X1   g08709(.A1(new_n6459_), .A2(new_n11353_), .B(new_n3160_), .ZN(new_n11692_));
  OAI21_X1   g08710(.A1(new_n11562_), .A2(new_n3361_), .B(new_n7811_), .ZN(new_n11693_));
  NOR2_X1    g08711(.A1(new_n11693_), .A2(new_n11692_), .ZN(new_n11694_));
  OAI21_X1   g08712(.A1(new_n11677_), .A2(new_n11691_), .B(new_n11694_), .ZN(new_n11695_));
  OAI21_X1   g08713(.A1(new_n11695_), .A2(new_n11670_), .B(new_n11660_), .ZN(new_n11696_));
  NOR2_X1    g08714(.A1(new_n11684_), .A2(pi0152), .ZN(new_n11697_));
  NOR2_X1    g08715(.A1(new_n11678_), .A2(new_n5158_), .ZN(new_n11698_));
  OAI21_X1   g08716(.A1(new_n11697_), .A2(new_n11698_), .B(pi0216), .ZN(new_n11699_));
  AOI21_X1   g08717(.A1(new_n11699_), .A2(new_n2702_), .B(new_n3827_), .ZN(new_n11700_));
  NOR4_X1    g08718(.A1(new_n11700_), .A2(pi0216), .A3(new_n3362_), .A4(new_n11562_), .ZN(new_n11701_));
  OR2_X2     g08719(.A1(new_n11701_), .A2(new_n7793_), .Z(new_n11702_));
  NOR2_X1    g08720(.A1(new_n6453_), .A2(new_n3098_), .ZN(new_n11703_));
  AOI21_X1   g08721(.A1(new_n3098_), .A2(new_n6459_), .B(new_n11703_), .ZN(new_n11704_));
  AOI21_X1   g08722(.A1(new_n3145_), .A2(new_n11361_), .B(new_n11704_), .ZN(new_n11705_));
  NAND2_X1   g08723(.A1(new_n4368_), .A2(new_n5551_), .ZN(new_n11706_));
  NAND2_X1   g08724(.A1(new_n11705_), .A2(new_n11706_), .ZN(new_n11707_));
  OAI21_X1   g08725(.A1(new_n11244_), .A2(new_n11707_), .B(new_n5551_), .ZN(new_n11708_));
  NAND4_X1   g08726(.A1(new_n11696_), .A2(new_n11700_), .A3(new_n11702_), .A4(new_n11708_), .ZN(new_n11709_));
  INV_X1     g08727(.I(new_n11568_), .ZN(new_n11710_));
  NAND2_X1   g08728(.A1(new_n11710_), .A2(pi0038), .ZN(new_n11711_));
  AOI21_X1   g08729(.A1(new_n11709_), .A2(new_n3462_), .B(new_n11711_), .ZN(new_n11712_));
  OAI21_X1   g08730(.A1(new_n11610_), .A2(new_n11649_), .B(new_n11712_), .ZN(new_n11713_));
  NAND2_X1   g08731(.A1(new_n8108_), .A2(pi0299), .ZN(new_n11714_));
  OAI21_X1   g08732(.A1(pi0140), .A2(pi0299), .B(new_n11714_), .ZN(new_n11715_));
  OAI21_X1   g08733(.A1(new_n6494_), .A2(new_n11715_), .B(pi0087), .ZN(new_n11716_));
  AOI21_X1   g08734(.A1(new_n11559_), .A2(new_n11716_), .B(new_n11408_), .ZN(new_n11717_));
  AOI21_X1   g08735(.A1(new_n11710_), .A2(new_n11717_), .B(new_n3207_), .ZN(new_n11718_));
  AOI21_X1   g08736(.A1(new_n11713_), .A2(new_n11718_), .B(new_n11570_), .ZN(new_n11719_));
  NOR2_X1    g08737(.A1(new_n11188_), .A2(new_n5386_), .ZN(new_n11720_));
  NOR2_X1    g08738(.A1(new_n11336_), .A2(new_n11217_), .ZN(new_n11721_));
  XNOR2_X1   g08739(.A1(new_n11720_), .A2(new_n11721_), .ZN(new_n11722_));
  NAND2_X1   g08740(.A1(new_n11722_), .A2(pi0172), .ZN(new_n11723_));
  XOR2_X1    g08741(.A1(new_n11723_), .A2(new_n7787_), .Z(new_n11724_));
  NOR2_X1    g08742(.A1(new_n11334_), .A2(new_n11209_), .ZN(new_n11725_));
  OAI21_X1   g08743(.A1(new_n11336_), .A2(new_n3827_), .B(new_n5386_), .ZN(new_n11726_));
  NAND4_X1   g08744(.A1(new_n11724_), .A2(pi0152), .A3(new_n11725_), .A4(new_n11726_), .ZN(new_n11727_));
  NAND2_X1   g08745(.A1(new_n11727_), .A2(new_n11342_), .ZN(new_n11728_));
  NOR2_X1    g08746(.A1(new_n11206_), .A2(new_n5373_), .ZN(new_n11729_));
  NOR2_X1    g08747(.A1(new_n11729_), .A2(new_n11205_), .ZN(new_n11730_));
  NAND2_X1   g08748(.A1(new_n11174_), .A2(new_n11730_), .ZN(new_n11731_));
  INV_X1     g08749(.I(new_n11209_), .ZN(new_n11732_));
  NAND2_X1   g08750(.A1(new_n11220_), .A2(new_n11732_), .ZN(new_n11733_));
  NAND2_X1   g08751(.A1(new_n11733_), .A2(pi0152), .ZN(new_n11734_));
  XOR2_X1    g08752(.A1(new_n11734_), .A2(new_n7779_), .Z(new_n11735_));
  OAI21_X1   g08753(.A1(new_n11735_), .A2(new_n11731_), .B(new_n5665_), .ZN(new_n11736_));
  INV_X1     g08754(.I(new_n11561_), .ZN(new_n11737_));
  NOR2_X1    g08755(.A1(new_n11245_), .A2(new_n11209_), .ZN(new_n11738_));
  INV_X1     g08756(.I(new_n11738_), .ZN(new_n11739_));
  AOI21_X1   g08757(.A1(new_n11739_), .A2(new_n5158_), .B(new_n11737_), .ZN(new_n11740_));
  NAND2_X1   g08758(.A1(new_n11736_), .A2(new_n11740_), .ZN(new_n11741_));
  INV_X1     g08759(.I(new_n11449_), .ZN(new_n11742_));
  NAND2_X1   g08760(.A1(new_n11209_), .A2(pi0172), .ZN(new_n11743_));
  AOI21_X1   g08761(.A1(new_n11743_), .A2(new_n5158_), .B(new_n11742_), .ZN(new_n11744_));
  NOR2_X1    g08762(.A1(new_n11210_), .A2(pi0172), .ZN(new_n11745_));
  NAND2_X1   g08763(.A1(new_n11449_), .A2(pi0152), .ZN(new_n11746_));
  OAI21_X1   g08764(.A1(new_n11745_), .A2(new_n11746_), .B(pi0197), .ZN(new_n11747_));
  NOR2_X1    g08765(.A1(new_n8174_), .A2(new_n3098_), .ZN(new_n11748_));
  OAI21_X1   g08766(.A1(new_n11747_), .A2(new_n11744_), .B(new_n11748_), .ZN(new_n11749_));
  AOI21_X1   g08767(.A1(new_n11215_), .A2(new_n11368_), .B(new_n11209_), .ZN(new_n11750_));
  NAND2_X1   g08768(.A1(new_n11732_), .A2(new_n11275_), .ZN(new_n11751_));
  NAND2_X1   g08769(.A1(new_n11751_), .A2(pi0172), .ZN(new_n11752_));
  XOR2_X1    g08770(.A1(new_n11752_), .A2(new_n7787_), .Z(new_n11753_));
  NAND2_X1   g08771(.A1(new_n11753_), .A2(new_n11750_), .ZN(new_n11754_));
  NAND3_X1   g08772(.A1(new_n11754_), .A2(new_n5665_), .A3(new_n11749_), .ZN(new_n11755_));
  NAND2_X1   g08773(.A1(new_n11230_), .A2(new_n5158_), .ZN(new_n11756_));
  OAI21_X1   g08774(.A1(new_n11751_), .A2(new_n11756_), .B(new_n3827_), .ZN(new_n11757_));
  NOR2_X1    g08775(.A1(new_n11209_), .A2(new_n11365_), .ZN(new_n11758_));
  INV_X1     g08776(.I(new_n11758_), .ZN(new_n11759_));
  NOR4_X1    g08777(.A1(new_n11759_), .A2(new_n5158_), .A3(new_n3098_), .A4(new_n8171_), .ZN(new_n11760_));
  NAND4_X1   g08778(.A1(new_n11741_), .A2(new_n11755_), .A3(new_n11757_), .A4(new_n11760_), .ZN(new_n11761_));
  NAND2_X1   g08779(.A1(new_n7467_), .A2(pi0152), .ZN(new_n11762_));
  AOI21_X1   g08780(.A1(new_n11761_), .A2(new_n5665_), .B(new_n11762_), .ZN(new_n11763_));
  AOI21_X1   g08781(.A1(new_n11728_), .A2(new_n11763_), .B(pi0038), .ZN(new_n11764_));
  NAND3_X1   g08782(.A1(new_n11739_), .A2(new_n5641_), .A3(new_n7378_), .ZN(new_n11765_));
  NAND2_X1   g08783(.A1(new_n11732_), .A2(new_n5641_), .ZN(new_n11766_));
  AOI21_X1   g08784(.A1(new_n11765_), .A2(pi0051), .B(new_n11766_), .ZN(new_n11767_));
  OAI21_X1   g08785(.A1(new_n11767_), .A2(new_n11342_), .B(new_n7342_), .ZN(new_n11768_));
  NAND2_X1   g08786(.A1(new_n11722_), .A2(pi0145), .ZN(new_n11769_));
  XNOR2_X1   g08787(.A1(new_n11769_), .A2(new_n11641_), .ZN(new_n11770_));
  NOR2_X1    g08788(.A1(new_n11725_), .A2(pi0174), .ZN(new_n11771_));
  AOI21_X1   g08789(.A1(new_n5641_), .A2(new_n11207_), .B(new_n11731_), .ZN(new_n11772_));
  NAND2_X1   g08790(.A1(new_n11772_), .A2(new_n10275_), .ZN(new_n11773_));
  INV_X1     g08791(.I(new_n11772_), .ZN(new_n11774_));
  NOR4_X1    g08792(.A1(new_n11774_), .A2(new_n8010_), .A3(new_n3098_), .A4(new_n11637_), .ZN(new_n11775_));
  OAI21_X1   g08793(.A1(new_n11771_), .A2(new_n11773_), .B(new_n11775_), .ZN(new_n11776_));
  AOI21_X1   g08794(.A1(new_n11770_), .A2(new_n11738_), .B(new_n11776_), .ZN(new_n11777_));
  NAND2_X1   g08795(.A1(new_n11369_), .A2(pi0145), .ZN(new_n11778_));
  NOR2_X1    g08796(.A1(new_n11566_), .A2(new_n5641_), .ZN(new_n11779_));
  XNOR2_X1   g08797(.A1(new_n11778_), .A2(new_n11779_), .ZN(new_n11780_));
  NAND2_X1   g08798(.A1(new_n11780_), .A2(pi0174), .ZN(new_n11781_));
  AOI21_X1   g08799(.A1(new_n11781_), .A2(new_n11275_), .B(new_n5641_), .ZN(new_n11782_));
  NAND2_X1   g08800(.A1(new_n11732_), .A2(pi0193), .ZN(new_n11783_));
  OAI21_X1   g08801(.A1(new_n11782_), .A2(new_n11783_), .B(new_n11614_), .ZN(new_n11784_));
  AOI21_X1   g08802(.A1(new_n11777_), .A2(new_n11768_), .B(new_n11784_), .ZN(new_n11785_));
  NAND2_X1   g08803(.A1(new_n11431_), .A2(pi0172), .ZN(new_n11786_));
  XOR2_X1    g08804(.A1(new_n11786_), .A2(new_n7779_), .Z(new_n11787_));
  OAI21_X1   g08805(.A1(new_n11787_), .A2(new_n11446_), .B(new_n7440_), .ZN(new_n11788_));
  NAND4_X1   g08806(.A1(new_n11422_), .A2(pi0152), .A3(new_n5373_), .A4(new_n11427_), .ZN(new_n11789_));
  NAND4_X1   g08807(.A1(new_n11423_), .A2(pi0152), .A3(new_n5373_), .A4(new_n11428_), .ZN(new_n11790_));
  AOI21_X1   g08808(.A1(new_n11790_), .A2(new_n11789_), .B(new_n3827_), .ZN(new_n11791_));
  AOI21_X1   g08809(.A1(new_n11788_), .A2(new_n11791_), .B(new_n3098_), .ZN(new_n11792_));
  XOR2_X1    g08810(.A1(new_n11792_), .A2(new_n7812_), .Z(new_n11793_));
  NOR2_X1    g08811(.A1(new_n7439_), .A2(pi0152), .ZN(new_n11794_));
  AOI21_X1   g08812(.A1(new_n11473_), .A2(new_n11794_), .B(new_n11737_), .ZN(new_n11795_));
  NOR3_X1    g08813(.A1(new_n11461_), .A2(pi0152), .A3(new_n11795_), .ZN(new_n11796_));
  NOR4_X1    g08814(.A1(new_n11793_), .A2(new_n7440_), .A3(new_n11737_), .A4(new_n11796_), .ZN(new_n11797_));
  OAI21_X1   g08815(.A1(new_n11797_), .A2(new_n11562_), .B(new_n11175_), .ZN(new_n11798_));
  NOR2_X1    g08816(.A1(new_n11438_), .A2(new_n7440_), .ZN(new_n11799_));
  NOR2_X1    g08817(.A1(new_n11799_), .A2(new_n3098_), .ZN(new_n11800_));
  AOI21_X1   g08818(.A1(new_n11346_), .A2(new_n7450_), .B(new_n11176_), .ZN(new_n11801_));
  INV_X1     g08819(.I(new_n11801_), .ZN(new_n11802_));
  NOR3_X1    g08820(.A1(new_n11802_), .A2(new_n3098_), .A3(new_n11176_), .ZN(new_n11803_));
  XNOR2_X1   g08821(.A1(new_n11803_), .A2(new_n11800_), .ZN(new_n11804_));
  NAND2_X1   g08822(.A1(pi0039), .A2(pi0232), .ZN(new_n11805_));
  NAND2_X1   g08823(.A1(new_n11798_), .A2(new_n11805_), .ZN(new_n11806_));
  AOI21_X1   g08824(.A1(new_n5386_), .A2(new_n11167_), .B(new_n7451_), .ZN(new_n11807_));
  NOR3_X1    g08825(.A1(new_n11430_), .A2(new_n2702_), .A3(new_n7451_), .ZN(new_n11808_));
  XNOR2_X1   g08826(.A1(new_n11808_), .A2(new_n11807_), .ZN(new_n11809_));
  INV_X1     g08827(.I(new_n11809_), .ZN(new_n11810_));
  INV_X1     g08828(.I(new_n11460_), .ZN(new_n11811_));
  NOR2_X1    g08829(.A1(new_n11811_), .A2(new_n5642_), .ZN(new_n11812_));
  OAI21_X1   g08830(.A1(new_n11810_), .A2(pi0174), .B(new_n11812_), .ZN(new_n11813_));
  NOR2_X1    g08831(.A1(pi0193), .A2(pi0299), .ZN(new_n11814_));
  NAND2_X1   g08832(.A1(new_n11802_), .A2(new_n7378_), .ZN(new_n11815_));
  NAND3_X1   g08833(.A1(new_n11815_), .A2(pi0180), .A3(new_n11472_), .ZN(new_n11816_));
  AOI21_X1   g08834(.A1(new_n11813_), .A2(new_n11814_), .B(new_n11816_), .ZN(new_n11817_));
  NAND2_X1   g08835(.A1(new_n11802_), .A2(new_n11230_), .ZN(new_n11818_));
  NOR2_X1    g08836(.A1(new_n7451_), .A2(new_n5386_), .ZN(new_n11819_));
  INV_X1     g08837(.I(new_n11819_), .ZN(new_n11820_));
  AOI21_X1   g08838(.A1(new_n11820_), .A2(new_n11167_), .B(new_n2702_), .ZN(new_n11821_));
  AOI21_X1   g08839(.A1(new_n11443_), .A2(new_n7450_), .B(new_n11821_), .ZN(new_n11822_));
  NOR2_X1    g08840(.A1(new_n11822_), .A2(new_n7378_), .ZN(new_n11823_));
  XOR2_X1    g08841(.A1(new_n11823_), .A2(new_n7886_), .Z(new_n11824_));
  OAI21_X1   g08842(.A1(new_n11824_), .A2(new_n11818_), .B(new_n7342_), .ZN(new_n11825_));
  NOR2_X1    g08843(.A1(new_n11817_), .A2(new_n11825_), .ZN(new_n11826_));
  INV_X1     g08844(.I(new_n11821_), .ZN(new_n11827_));
  NOR2_X1    g08845(.A1(new_n11422_), .A2(new_n7451_), .ZN(new_n11828_));
  XOR2_X1    g08846(.A1(new_n11828_), .A2(new_n11820_), .Z(new_n11829_));
  OAI21_X1   g08847(.A1(new_n11829_), .A2(new_n8639_), .B(new_n11827_), .ZN(new_n11830_));
  NOR2_X1    g08848(.A1(new_n11472_), .A2(pi0051), .ZN(new_n11831_));
  INV_X1     g08849(.I(new_n11831_), .ZN(new_n11832_));
  NAND2_X1   g08850(.A1(new_n11832_), .A2(new_n5373_), .ZN(new_n11833_));
  NAND2_X1   g08851(.A1(new_n11833_), .A2(new_n11802_), .ZN(new_n11834_));
  NAND2_X1   g08852(.A1(new_n11834_), .A2(pi0180), .ZN(new_n11835_));
  XOR2_X1    g08853(.A1(new_n11835_), .A2(new_n7885_), .Z(new_n11836_));
  NOR3_X1    g08854(.A1(new_n11826_), .A2(new_n11830_), .A3(new_n11836_), .ZN(new_n11837_));
  NAND2_X1   g08855(.A1(new_n11208_), .A2(new_n11706_), .ZN(new_n11838_));
  AOI21_X1   g08856(.A1(new_n11806_), .A2(new_n11837_), .B(new_n11838_), .ZN(new_n11839_));
  NOR2_X1    g08857(.A1(new_n11209_), .A2(new_n11229_), .ZN(new_n11840_));
  OAI21_X1   g08858(.A1(pi0145), .A2(new_n11166_), .B(new_n11274_), .ZN(new_n11841_));
  NAND2_X1   g08859(.A1(new_n11166_), .A2(pi0174), .ZN(new_n11842_));
  NAND4_X1   g08860(.A1(new_n11840_), .A2(pi0193), .A3(new_n11841_), .A4(new_n11842_), .ZN(new_n11843_));
  NAND2_X1   g08861(.A1(new_n11843_), .A2(new_n7378_), .ZN(new_n11844_));
  OAI21_X1   g08862(.A1(new_n11710_), .A2(new_n3133_), .B(new_n11175_), .ZN(new_n11845_));
  NOR2_X1    g08863(.A1(new_n11569_), .A2(new_n11501_), .ZN(new_n11846_));
  NAND2_X1   g08864(.A1(new_n11559_), .A2(new_n11716_), .ZN(new_n11847_));
  NAND3_X1   g08865(.A1(new_n7240_), .A2(new_n3455_), .A3(new_n8108_), .ZN(new_n11848_));
  NOR2_X1    g08866(.A1(new_n11322_), .A2(new_n6494_), .ZN(new_n11849_));
  NAND4_X1   g08867(.A1(new_n11710_), .A2(new_n11847_), .A3(new_n11848_), .A4(new_n11849_), .ZN(new_n11850_));
  NOR2_X1    g08868(.A1(new_n11850_), .A2(new_n11846_), .ZN(new_n11851_));
  NAND4_X1   g08869(.A1(new_n11844_), .A2(new_n11758_), .A3(new_n11845_), .A4(new_n11851_), .ZN(new_n11852_));
  NOR4_X1    g08870(.A1(new_n11764_), .A2(new_n11785_), .A3(new_n11839_), .A4(new_n11852_), .ZN(new_n11853_));
  OAI21_X1   g08871(.A1(new_n11719_), .A2(po1038), .B(new_n11853_), .ZN(new_n11854_));
  AOI21_X1   g08872(.A1(new_n11854_), .A2(new_n3455_), .B(new_n11563_), .ZN(po0282));
  OAI21_X1   g08873(.A1(new_n11751_), .A2(pi0189), .B(pi0178), .ZN(new_n11856_));
  OAI21_X1   g08874(.A1(new_n11856_), .A2(new_n5643_), .B(new_n8642_), .ZN(new_n11857_));
  NAND2_X1   g08875(.A1(new_n11857_), .A2(new_n11750_), .ZN(new_n11858_));
  NAND2_X1   g08876(.A1(pi0178), .A2(pi0189), .ZN(new_n11859_));
  NOR2_X1    g08877(.A1(new_n11245_), .A2(new_n8642_), .ZN(new_n11860_));
  XNOR2_X1   g08878(.A1(new_n11860_), .A2(new_n11859_), .ZN(new_n11861_));
  NOR3_X1    g08879(.A1(new_n8643_), .A2(pi0178), .A3(pi0181), .ZN(new_n11862_));
  OAI21_X1   g08880(.A1(new_n11328_), .A2(new_n11862_), .B(new_n9488_), .ZN(new_n11863_));
  AOI21_X1   g08881(.A1(new_n11861_), .A2(new_n11221_), .B(new_n11863_), .ZN(new_n11864_));
  NOR2_X1    g08882(.A1(pi0153), .A2(pi0166), .ZN(new_n11865_));
  INV_X1     g08883(.I(new_n11865_), .ZN(new_n11866_));
  NOR2_X1    g08884(.A1(new_n5373_), .A2(new_n4808_), .ZN(new_n11867_));
  NAND2_X1   g08885(.A1(pi0051), .A2(pi0166), .ZN(new_n11868_));
  OAI21_X1   g08886(.A1(new_n11731_), .A2(new_n11868_), .B(new_n11867_), .ZN(new_n11869_));
  OR3_X2     g08887(.A1(new_n11731_), .A2(new_n11867_), .A3(new_n11868_), .Z(new_n11870_));
  NAND3_X1   g08888(.A1(new_n11870_), .A2(new_n2837_), .A3(new_n11869_), .ZN(new_n11871_));
  AOI21_X1   g08889(.A1(new_n11871_), .A2(new_n10692_), .B(new_n11866_), .ZN(new_n11872_));
  NAND2_X1   g08890(.A1(new_n11209_), .A2(pi0153), .ZN(new_n11873_));
  AOI21_X1   g08891(.A1(new_n11873_), .A2(new_n4808_), .B(new_n11742_), .ZN(new_n11874_));
  NOR2_X1    g08892(.A1(new_n11449_), .A2(pi0051), .ZN(new_n11875_));
  NOR2_X1    g08893(.A1(new_n5373_), .A2(new_n2702_), .ZN(new_n11876_));
  NAND4_X1   g08894(.A1(new_n8443_), .A2(pi0051), .A3(new_n11167_), .A4(pi0153), .ZN(new_n11877_));
  XOR2_X1    g08895(.A1(new_n11877_), .A2(new_n11876_), .Z(new_n11878_));
  INV_X1     g08896(.I(new_n11878_), .ZN(new_n11879_));
  NOR2_X1    g08897(.A1(new_n11879_), .A2(new_n11875_), .ZN(new_n11880_));
  NAND2_X1   g08898(.A1(new_n2837_), .A2(new_n10692_), .ZN(new_n11881_));
  OAI21_X1   g08899(.A1(new_n11210_), .A2(new_n11881_), .B(new_n11880_), .ZN(new_n11882_));
  NOR2_X1    g08900(.A1(new_n11733_), .A2(new_n8110_), .ZN(new_n11883_));
  OAI21_X1   g08901(.A1(new_n11874_), .A2(new_n11882_), .B(new_n11883_), .ZN(new_n11884_));
  OAI21_X1   g08902(.A1(new_n11884_), .A2(new_n11872_), .B(new_n4808_), .ZN(new_n11885_));
  NAND3_X1   g08903(.A1(new_n11885_), .A2(new_n11209_), .A3(new_n11738_), .ZN(new_n11886_));
  OAI21_X1   g08904(.A1(new_n11864_), .A2(new_n11886_), .B(new_n11858_), .ZN(new_n11887_));
  INV_X1     g08905(.I(new_n11725_), .ZN(new_n11888_));
  NAND2_X1   g08906(.A1(new_n11722_), .A2(pi0189), .ZN(new_n11889_));
  XNOR2_X1   g08907(.A1(new_n11889_), .A2(new_n11859_), .ZN(new_n11890_));
  OAI21_X1   g08908(.A1(new_n11759_), .A2(new_n11868_), .B(new_n11867_), .ZN(new_n11891_));
  NOR3_X1    g08909(.A1(new_n11759_), .A2(new_n11867_), .A3(new_n11868_), .ZN(new_n11892_));
  NOR2_X1    g08910(.A1(new_n11892_), .A2(pi0153), .ZN(new_n11893_));
  AOI21_X1   g08911(.A1(new_n10692_), .A2(new_n11865_), .B(new_n8178_), .ZN(new_n11894_));
  NAND2_X1   g08912(.A1(new_n11750_), .A2(new_n11894_), .ZN(new_n11895_));
  AOI21_X1   g08913(.A1(new_n11893_), .A2(new_n11891_), .B(new_n11895_), .ZN(new_n11896_));
  NOR2_X1    g08914(.A1(new_n11896_), .A2(pi0166), .ZN(new_n11897_));
  NOR4_X1    g08915(.A1(new_n11890_), .A2(new_n11888_), .A3(new_n11751_), .A4(new_n11897_), .ZN(new_n11898_));
  AOI21_X1   g08916(.A1(new_n11898_), .A2(new_n11887_), .B(pi0157), .ZN(new_n11899_));
  NAND2_X1   g08917(.A1(pi0153), .A2(pi0166), .ZN(new_n11900_));
  NAND2_X1   g08918(.A1(new_n11722_), .A2(pi0153), .ZN(new_n11901_));
  XNOR2_X1   g08919(.A1(new_n11901_), .A2(new_n11900_), .ZN(new_n11902_));
  NOR2_X1    g08920(.A1(new_n11208_), .A2(new_n8442_), .ZN(new_n11903_));
  NOR4_X1    g08921(.A1(new_n11902_), .A2(pi0153), .A3(new_n11888_), .A4(new_n11903_), .ZN(new_n11904_));
  OAI21_X1   g08922(.A1(new_n11904_), .A2(new_n11388_), .B(pi0166), .ZN(new_n11905_));
  INV_X1     g08923(.I(new_n11840_), .ZN(new_n11906_));
  OAI21_X1   g08924(.A1(new_n11731_), .A2(new_n8642_), .B(new_n7510_), .ZN(new_n11907_));
  NAND3_X1   g08925(.A1(new_n11906_), .A2(new_n8642_), .A3(new_n11907_), .ZN(new_n11908_));
  NAND2_X1   g08926(.A1(new_n11245_), .A2(new_n11908_), .ZN(new_n11909_));
  NOR2_X1    g08927(.A1(new_n11906_), .A2(pi0189), .ZN(new_n11910_));
  NOR2_X1    g08928(.A1(new_n11910_), .A2(new_n7510_), .ZN(new_n11911_));
  NAND2_X1   g08929(.A1(new_n11210_), .A2(pi0189), .ZN(new_n11912_));
  AOI21_X1   g08930(.A1(new_n11911_), .A2(new_n11912_), .B(new_n5643_), .ZN(new_n11913_));
  AOI21_X1   g08931(.A1(new_n11913_), .A2(new_n11909_), .B(new_n9474_), .ZN(new_n11914_));
  OAI21_X1   g08932(.A1(new_n11899_), .A2(new_n11905_), .B(new_n11914_), .ZN(new_n11915_));
  NAND2_X1   g08933(.A1(new_n11198_), .A2(new_n8643_), .ZN(new_n11916_));
  NOR2_X1    g08934(.A1(new_n11336_), .A2(new_n8644_), .ZN(new_n11917_));
  XOR2_X1    g08935(.A1(new_n11916_), .A2(new_n11917_), .Z(new_n11918_));
  NOR2_X1    g08936(.A1(new_n7510_), .A2(new_n8642_), .ZN(new_n11919_));
  OAI21_X1   g08937(.A1(new_n11856_), .A2(new_n11759_), .B(new_n5643_), .ZN(new_n11920_));
  OAI21_X1   g08938(.A1(new_n11920_), .A2(new_n11919_), .B(pi0178), .ZN(new_n11921_));
  NOR2_X1    g08939(.A1(new_n11918_), .A2(new_n11921_), .ZN(new_n11922_));
  AOI21_X1   g08940(.A1(new_n11915_), .A2(new_n11922_), .B(new_n5551_), .ZN(new_n11923_));
  XOR2_X1    g08941(.A1(new_n11923_), .A2(new_n11361_), .Z(new_n11924_));
  NOR2_X1    g08942(.A1(new_n11924_), .A2(new_n11336_), .ZN(new_n11925_));
  NOR3_X1    g08943(.A1(pi0121), .A2(pi0125), .A3(pi0133), .ZN(new_n11926_));
  NOR2_X1    g08944(.A1(new_n11313_), .A2(pi0126), .ZN(new_n11927_));
  AOI21_X1   g08945(.A1(new_n11927_), .A2(new_n11926_), .B(pi0132), .ZN(new_n11928_));
  XOR2_X1    g08946(.A1(new_n11928_), .A2(new_n11313_), .Z(new_n11929_));
  NAND2_X1   g08947(.A1(new_n11929_), .A2(new_n3133_), .ZN(new_n11930_));
  NOR2_X1    g08948(.A1(new_n5644_), .A2(new_n8642_), .ZN(new_n11931_));
  NAND2_X1   g08949(.A1(new_n11834_), .A2(pi0182), .ZN(new_n11932_));
  XOR2_X1    g08950(.A1(new_n11932_), .A2(new_n11931_), .Z(new_n11933_));
  NOR2_X1    g08951(.A1(new_n11933_), .A2(new_n11830_), .ZN(new_n11934_));
  NOR2_X1    g08952(.A1(new_n11811_), .A2(new_n5644_), .ZN(new_n11935_));
  NOR2_X1    g08953(.A1(new_n11801_), .A2(pi0189), .ZN(new_n11936_));
  NAND3_X1   g08954(.A1(new_n11472_), .A2(pi0182), .A3(new_n9474_), .ZN(new_n11937_));
  OAI22_X1   g08955(.A1(new_n11937_), .A2(new_n11936_), .B1(pi0189), .B2(new_n11935_), .ZN(new_n11938_));
  AND3_X2    g08956(.A1(new_n11810_), .A2(new_n9487_), .A3(new_n11938_), .Z(new_n11939_));
  NOR2_X1    g08957(.A1(new_n11822_), .A2(new_n8642_), .ZN(new_n11940_));
  XNOR2_X1   g08958(.A1(new_n11940_), .A2(new_n11931_), .ZN(new_n11941_));
  NOR2_X1    g08959(.A1(new_n11941_), .A2(new_n11818_), .ZN(new_n11942_));
  OAI21_X1   g08960(.A1(new_n11934_), .A2(new_n11939_), .B(new_n11942_), .ZN(new_n11943_));
  NOR2_X1    g08961(.A1(new_n11230_), .A2(new_n2837_), .ZN(new_n11944_));
  NOR4_X1    g08962(.A1(new_n11462_), .A2(new_n5664_), .A3(new_n4808_), .A4(new_n11944_), .ZN(new_n11945_));
  NOR4_X1    g08963(.A1(new_n11461_), .A2(new_n5664_), .A3(pi0166), .A4(new_n11944_), .ZN(new_n11946_));
  OAI21_X1   g08964(.A1(new_n11945_), .A2(new_n11946_), .B(new_n11472_), .ZN(new_n11947_));
  AOI21_X1   g08965(.A1(new_n11879_), .A2(pi0299), .B(new_n7439_), .ZN(new_n11948_));
  NAND2_X1   g08966(.A1(new_n11947_), .A2(new_n11948_), .ZN(new_n11949_));
  NAND3_X1   g08967(.A1(new_n11422_), .A2(new_n9442_), .A3(new_n11427_), .ZN(new_n11950_));
  NAND3_X1   g08968(.A1(new_n11423_), .A2(new_n9442_), .A3(new_n11428_), .ZN(new_n11951_));
  NAND2_X1   g08969(.A1(new_n11951_), .A2(new_n11950_), .ZN(new_n11952_));
  NAND2_X1   g08970(.A1(new_n11431_), .A2(pi0153), .ZN(new_n11953_));
  XNOR2_X1   g08971(.A1(new_n11953_), .A2(new_n11900_), .ZN(new_n11954_));
  INV_X1     g08972(.I(new_n11446_), .ZN(new_n11955_));
  NAND2_X1   g08973(.A1(new_n11955_), .A2(pi0160), .ZN(new_n11956_));
  OAI21_X1   g08974(.A1(new_n11954_), .A2(new_n11956_), .B(new_n2837_), .ZN(new_n11957_));
  NAND3_X1   g08975(.A1(new_n11949_), .A2(new_n11952_), .A3(new_n11957_), .ZN(new_n11958_));
  AOI21_X1   g08976(.A1(new_n11943_), .A2(new_n11805_), .B(new_n11958_), .ZN(new_n11959_));
  OAI21_X1   g08977(.A1(new_n11925_), .A2(new_n11930_), .B(new_n11959_), .ZN(new_n11960_));
  INV_X1     g08978(.I(new_n11929_), .ZN(new_n11961_));
  NOR2_X1    g08979(.A1(new_n11672_), .A2(new_n8642_), .ZN(new_n11962_));
  XOR2_X1    g08980(.A1(new_n11962_), .A2(new_n11931_), .Z(new_n11963_));
  NAND2_X1   g08981(.A1(new_n11963_), .A2(new_n11671_), .ZN(new_n11964_));
  NOR2_X1    g08982(.A1(new_n11668_), .A2(new_n5644_), .ZN(new_n11965_));
  XNOR2_X1   g08983(.A1(new_n11965_), .A2(new_n11931_), .ZN(new_n11966_));
  OAI21_X1   g08984(.A1(new_n11966_), .A2(new_n11692_), .B(new_n11964_), .ZN(new_n11967_));
  AOI21_X1   g08985(.A1(new_n11880_), .A2(new_n3361_), .B(pi0216), .ZN(new_n11968_));
  OAI21_X1   g08986(.A1(new_n11968_), .A2(new_n5664_), .B(new_n3098_), .ZN(new_n11969_));
  AOI21_X1   g08987(.A1(new_n11967_), .A2(new_n9474_), .B(new_n11969_), .ZN(new_n11970_));
  NOR2_X1    g08988(.A1(new_n11347_), .A2(new_n4808_), .ZN(new_n11971_));
  XNOR2_X1   g08989(.A1(new_n11971_), .A2(new_n11900_), .ZN(new_n11972_));
  NAND2_X1   g08990(.A1(new_n11378_), .A2(new_n11972_), .ZN(new_n11973_));
  NOR2_X1    g08991(.A1(new_n11657_), .A2(new_n2837_), .ZN(new_n11974_));
  XNOR2_X1   g08992(.A1(new_n11974_), .A2(new_n11900_), .ZN(new_n11975_));
  NAND2_X1   g08993(.A1(new_n11975_), .A2(new_n11656_), .ZN(new_n11976_));
  NAND3_X1   g08994(.A1(new_n11976_), .A2(pi0160), .A3(new_n11973_), .ZN(new_n11977_));
  NAND2_X1   g08995(.A1(new_n11977_), .A2(new_n3361_), .ZN(new_n11978_));
  XOR2_X1    g08996(.A1(new_n11978_), .A2(new_n7440_), .Z(new_n11979_));
  INV_X1     g08997(.I(new_n11678_), .ZN(new_n11980_));
  OAI22_X1   g08998(.A1(new_n11684_), .A2(pi0166), .B1(new_n2702_), .B2(pi0153), .ZN(new_n11981_));
  AOI21_X1   g08999(.A1(pi0166), .A2(new_n11980_), .B(new_n11981_), .ZN(new_n11982_));
  NAND2_X1   g09000(.A1(new_n11979_), .A2(new_n11982_), .ZN(new_n11983_));
  NAND2_X1   g09001(.A1(new_n11705_), .A2(pi0232), .ZN(new_n11984_));
  OAI21_X1   g09002(.A1(new_n11970_), .A2(new_n11983_), .B(new_n11984_), .ZN(new_n11985_));
  NOR2_X1    g09003(.A1(new_n11688_), .A2(new_n5644_), .ZN(new_n11986_));
  XOR2_X1    g09004(.A1(new_n11986_), .A2(new_n11931_), .Z(new_n11987_));
  NAND3_X1   g09005(.A1(new_n11987_), .A2(new_n9487_), .A3(new_n11681_), .ZN(new_n11988_));
  AOI21_X1   g09006(.A1(new_n11964_), .A2(new_n11988_), .B(new_n11230_), .ZN(new_n11989_));
  AOI21_X1   g09007(.A1(new_n11985_), .A2(new_n11989_), .B(new_n11961_), .ZN(new_n11990_));
  NAND2_X1   g09008(.A1(new_n11605_), .A2(pi0178), .ZN(new_n11991_));
  XNOR2_X1   g09009(.A1(new_n11991_), .A2(new_n11859_), .ZN(new_n11992_));
  NOR2_X1    g09010(.A1(new_n11992_), .A2(new_n11573_), .ZN(new_n11993_));
  NAND2_X1   g09011(.A1(new_n11580_), .A2(pi0178), .ZN(new_n11994_));
  XOR2_X1    g09012(.A1(new_n11994_), .A2(new_n11859_), .Z(new_n11995_));
  NAND2_X1   g09013(.A1(new_n11995_), .A2(new_n11578_), .ZN(new_n11996_));
  NAND2_X1   g09014(.A1(new_n11196_), .A2(pi0189), .ZN(new_n11997_));
  OAI21_X1   g09015(.A1(new_n11229_), .A2(pi0178), .B(pi0181), .ZN(new_n11998_));
  OAI21_X1   g09016(.A1(new_n11997_), .A2(new_n11998_), .B(new_n8642_), .ZN(new_n11999_));
  AOI21_X1   g09017(.A1(new_n11645_), .A2(new_n11999_), .B(new_n9474_), .ZN(new_n12000_));
  NOR2_X1    g09018(.A1(new_n11997_), .A2(new_n5643_), .ZN(new_n12001_));
  OAI21_X1   g09019(.A1(new_n11645_), .A2(pi0178), .B(new_n12001_), .ZN(new_n12002_));
  AOI21_X1   g09020(.A1(new_n11996_), .A2(new_n12000_), .B(new_n12002_), .ZN(new_n12003_));
  NAND2_X1   g09021(.A1(new_n11590_), .A2(pi0189), .ZN(new_n12004_));
  XNOR2_X1   g09022(.A1(new_n12004_), .A2(new_n11859_), .ZN(new_n12005_));
  NOR2_X1    g09023(.A1(new_n11642_), .A2(new_n12005_), .ZN(new_n12006_));
  OAI21_X1   g09024(.A1(new_n11993_), .A2(new_n12003_), .B(new_n12006_), .ZN(new_n12007_));
  OAI21_X1   g09025(.A1(new_n11608_), .A2(new_n11910_), .B(new_n7510_), .ZN(new_n12008_));
  NAND3_X1   g09026(.A1(new_n12008_), .A2(pi0189), .A3(new_n11574_), .ZN(new_n12009_));
  NAND2_X1   g09027(.A1(new_n11642_), .A2(pi0189), .ZN(new_n12010_));
  NAND2_X1   g09028(.A1(new_n11585_), .A2(new_n11275_), .ZN(new_n12011_));
  NOR3_X1    g09029(.A1(new_n12011_), .A2(new_n8642_), .A3(new_n11230_), .ZN(new_n12012_));
  XNOR2_X1   g09030(.A1(new_n12010_), .A2(new_n12012_), .ZN(new_n12013_));
  NAND2_X1   g09031(.A1(new_n12013_), .A2(pi0178), .ZN(new_n12014_));
  AOI21_X1   g09032(.A1(new_n12009_), .A2(new_n5643_), .B(new_n12014_), .ZN(new_n12015_));
  NAND2_X1   g09033(.A1(new_n11586_), .A2(pi0178), .ZN(new_n12016_));
  XNOR2_X1   g09034(.A1(new_n12016_), .A2(new_n11859_), .ZN(new_n12017_));
  NAND3_X1   g09035(.A1(new_n11599_), .A2(new_n11645_), .A3(new_n11999_), .ZN(new_n12018_));
  NOR2_X1    g09036(.A1(new_n12017_), .A2(new_n12018_), .ZN(new_n12019_));
  OAI21_X1   g09037(.A1(new_n12015_), .A2(new_n9487_), .B(new_n12019_), .ZN(new_n12020_));
  NAND2_X1   g09038(.A1(new_n11586_), .A2(pi0153), .ZN(new_n12021_));
  XOR2_X1    g09039(.A1(new_n12021_), .A2(new_n11900_), .Z(new_n12022_));
  INV_X1     g09040(.I(new_n11944_), .ZN(new_n12023_));
  NAND4_X1   g09041(.A1(new_n11645_), .A2(new_n10692_), .A3(pi0166), .A4(new_n12023_), .ZN(new_n12024_));
  NAND4_X1   g09042(.A1(new_n11646_), .A2(new_n10692_), .A3(new_n4808_), .A4(new_n12023_), .ZN(new_n12025_));
  NAND2_X1   g09043(.A1(new_n12025_), .A2(new_n12024_), .ZN(new_n12026_));
  NOR2_X1    g09044(.A1(new_n11244_), .A2(new_n10692_), .ZN(new_n12027_));
  AOI22_X1   g09045(.A1(new_n12022_), .A2(new_n11599_), .B1(new_n12026_), .B2(new_n12027_), .ZN(new_n12028_));
  NAND2_X1   g09046(.A1(new_n11580_), .A2(pi0166), .ZN(new_n12029_));
  XOR2_X1    g09047(.A1(new_n12029_), .A2(new_n11900_), .Z(new_n12030_));
  NAND2_X1   g09048(.A1(new_n12030_), .A2(new_n11578_), .ZN(new_n12031_));
  OAI21_X1   g09049(.A1(new_n12031_), .A2(new_n12028_), .B(new_n8177_), .ZN(new_n12032_));
  NAND2_X1   g09050(.A1(new_n12020_), .A2(new_n12032_), .ZN(new_n12033_));
  NAND2_X1   g09051(.A1(new_n12033_), .A2(new_n12007_), .ZN(new_n12034_));
  NAND3_X1   g09052(.A1(new_n11622_), .A2(pi0153), .A3(pi0157), .ZN(new_n12035_));
  NAND3_X1   g09053(.A1(new_n11605_), .A2(new_n2837_), .A3(pi0157), .ZN(new_n12036_));
  AOI21_X1   g09054(.A1(new_n12035_), .A2(new_n12036_), .B(new_n11608_), .ZN(new_n12037_));
  NOR4_X1    g09055(.A1(new_n11573_), .A2(new_n10692_), .A3(pi0166), .A4(new_n11944_), .ZN(new_n12038_));
  NOR4_X1    g09056(.A1(new_n11574_), .A2(pi0157), .A3(pi0166), .A4(new_n11944_), .ZN(new_n12039_));
  NOR2_X1    g09057(.A1(new_n12039_), .A2(new_n12038_), .ZN(new_n12040_));
  NOR3_X1    g09058(.A1(new_n12040_), .A2(new_n4808_), .A3(new_n11642_), .ZN(new_n12041_));
  NOR2_X1    g09059(.A1(new_n12037_), .A2(new_n12041_), .ZN(new_n12042_));
  NOR2_X1    g09060(.A1(new_n2837_), .A2(new_n10692_), .ZN(new_n12043_));
  NAND2_X1   g09061(.A1(new_n11590_), .A2(pi0153), .ZN(new_n12044_));
  XOR2_X1    g09062(.A1(new_n12044_), .A2(new_n12043_), .Z(new_n12045_));
  NOR4_X1    g09063(.A1(new_n12042_), .A2(new_n8110_), .A3(new_n12011_), .A4(new_n12045_), .ZN(new_n12046_));
  AOI21_X1   g09064(.A1(new_n12034_), .A2(new_n12046_), .B(new_n5551_), .ZN(new_n12047_));
  XOR2_X1    g09065(.A1(new_n12047_), .A2(new_n8536_), .Z(new_n12048_));
  NAND2_X1   g09066(.A1(new_n12048_), .A2(new_n11196_), .ZN(new_n12049_));
  AOI21_X1   g09067(.A1(new_n11960_), .A2(new_n11990_), .B(new_n12049_), .ZN(new_n12050_));
  NOR2_X1    g09068(.A1(new_n3207_), .A2(new_n3132_), .ZN(new_n12051_));
  AOI21_X1   g09069(.A1(new_n11176_), .A2(new_n12051_), .B(new_n11929_), .ZN(new_n12052_));
  AOI21_X1   g09070(.A1(new_n11229_), .A2(pi0175), .B(pi0299), .ZN(new_n12053_));
  NAND2_X1   g09071(.A1(new_n11449_), .A2(pi0189), .ZN(new_n12054_));
  OAI21_X1   g09072(.A1(new_n12054_), .A2(new_n12053_), .B(new_n5551_), .ZN(new_n12055_));
  NAND3_X1   g09073(.A1(new_n11880_), .A2(pi0299), .A3(new_n12055_), .ZN(new_n12056_));
  NOR2_X1    g09074(.A1(new_n12056_), .A2(new_n3133_), .ZN(new_n12057_));
  OAI21_X1   g09075(.A1(new_n12050_), .A2(new_n12052_), .B(new_n12057_), .ZN(new_n12058_));
  NOR2_X1    g09076(.A1(new_n11875_), .A2(new_n5551_), .ZN(new_n12059_));
  OAI21_X1   g09077(.A1(new_n11929_), .A2(new_n12059_), .B(new_n11878_), .ZN(new_n12060_));
  NOR2_X1    g09078(.A1(new_n11176_), .A2(new_n5551_), .ZN(new_n12061_));
  AOI21_X1   g09079(.A1(new_n12060_), .A2(new_n12061_), .B(new_n7240_), .ZN(new_n12062_));
  NOR2_X1    g09080(.A1(new_n7240_), .A2(new_n3455_), .ZN(new_n12063_));
  XOR2_X1    g09081(.A1(new_n12062_), .A2(new_n12063_), .Z(new_n12064_));
  AOI21_X1   g09082(.A1(new_n12064_), .A2(new_n10737_), .B(po1038), .ZN(new_n12065_));
  NAND2_X1   g09083(.A1(new_n12056_), .A2(pi0087), .ZN(new_n12066_));
  NAND2_X1   g09084(.A1(new_n6493_), .A2(new_n10629_), .ZN(new_n12067_));
  XOR2_X1    g09085(.A1(new_n7492_), .A2(new_n12067_), .Z(new_n12068_));
  NOR4_X1    g09086(.A1(new_n12068_), .A2(new_n3455_), .A3(new_n10659_), .A4(new_n3288_), .ZN(new_n12069_));
  AOI22_X1   g09087(.A1(new_n12066_), .A2(new_n12069_), .B1(new_n11416_), .B2(new_n11929_), .ZN(new_n12070_));
  OAI21_X1   g09088(.A1(new_n12066_), .A2(new_n12069_), .B(new_n12070_), .ZN(new_n12071_));
  AOI21_X1   g09089(.A1(new_n12058_), .A2(new_n12065_), .B(new_n12071_), .ZN(po0283));
  INV_X1     g09090(.I(new_n2561_), .ZN(new_n12074_));
  NOR3_X1    g09091(.A1(new_n7320_), .A2(new_n3259_), .A3(new_n3183_), .ZN(new_n12105_));
  NOR2_X1    g09092(.A1(new_n12105_), .A2(pi0129), .ZN(new_n12106_));
  OAI21_X1   g09093(.A1(new_n7499_), .A2(new_n12106_), .B(new_n3184_), .ZN(new_n12107_));
  NAND2_X1   g09094(.A1(new_n3184_), .A2(pi0075), .ZN(new_n12108_));
  XOR2_X1    g09095(.A1(new_n12107_), .A2(new_n12108_), .Z(new_n12109_));
  AOI21_X1   g09096(.A1(new_n3474_), .A2(new_n7334_), .B(new_n7320_), .ZN(new_n12110_));
  AOI21_X1   g09097(.A1(new_n12109_), .A2(new_n12110_), .B(pi0092), .ZN(new_n12111_));
  INV_X1     g09098(.I(new_n6286_), .ZN(new_n12112_));
  NOR2_X1    g09099(.A1(new_n12112_), .A2(new_n7318_), .ZN(new_n12113_));
  NAND2_X1   g09100(.A1(new_n12113_), .A2(pi0075), .ZN(new_n12114_));
  OAI21_X1   g09101(.A1(new_n12111_), .A2(new_n12114_), .B(new_n10622_), .ZN(new_n12115_));
  NOR2_X1    g09102(.A1(new_n3196_), .A2(new_n3115_), .ZN(new_n12116_));
  INV_X1     g09103(.I(new_n12116_), .ZN(new_n12117_));
  NOR2_X1    g09104(.A1(new_n7320_), .A2(new_n12117_), .ZN(new_n12118_));
  NOR2_X1    g09105(.A1(new_n12113_), .A2(new_n6327_), .ZN(new_n12119_));
  NAND4_X1   g09106(.A1(new_n12113_), .A2(pi0055), .A3(new_n3287_), .A4(new_n5765_), .ZN(new_n12120_));
  OAI22_X1   g09107(.A1(new_n12120_), .A2(new_n12119_), .B1(pi0074), .B2(new_n12118_), .ZN(new_n12121_));
  NAND4_X1   g09108(.A1(new_n12115_), .A2(pi0092), .A3(pi0129), .A4(new_n12121_), .ZN(new_n12122_));
  NOR2_X1    g09109(.A1(new_n12122_), .A2(new_n3219_), .ZN(new_n12123_));
  NOR2_X1    g09110(.A1(new_n3224_), .A2(new_n7320_), .ZN(new_n12124_));
  XOR2_X1    g09111(.A1(new_n12122_), .A2(new_n3221_), .Z(new_n12125_));
  NAND2_X1   g09112(.A1(new_n12125_), .A2(new_n12124_), .ZN(new_n12126_));
  XOR2_X1    g09113(.A1(new_n12126_), .A2(new_n12123_), .Z(new_n12127_));
  NOR2_X1    g09114(.A1(new_n12127_), .A2(new_n5371_), .ZN(new_n12128_));
  XOR2_X1    g09115(.A1(new_n12127_), .A2(new_n8226_), .Z(new_n12129_));
  NAND3_X1   g09116(.A1(new_n12129_), .A2(new_n3225_), .A3(new_n12124_), .ZN(new_n12130_));
  XNOR2_X1   g09117(.A1(new_n12130_), .A2(new_n12128_), .ZN(po0284));
  NOR2_X1    g09118(.A1(new_n3461_), .A2(new_n3259_), .ZN(new_n12132_));
  XOR2_X1    g09119(.A1(new_n12132_), .A2(new_n5486_), .Z(new_n12133_));
  INV_X1     g09120(.I(new_n5507_), .ZN(new_n12134_));
  NOR2_X1    g09121(.A1(new_n12134_), .A2(new_n5537_), .ZN(new_n12135_));
  NAND2_X1   g09122(.A1(new_n8236_), .A2(new_n7337_), .ZN(new_n12136_));
  NAND4_X1   g09123(.A1(new_n7315_), .A2(new_n5530_), .A3(pi0252), .A4(new_n7337_), .ZN(new_n12137_));
  XOR2_X1    g09124(.A1(new_n12137_), .A2(new_n12136_), .Z(new_n12138_));
  NAND3_X1   g09125(.A1(new_n12138_), .A2(pi0129), .A3(new_n3160_), .ZN(new_n12139_));
  NAND2_X1   g09126(.A1(new_n12139_), .A2(new_n5499_), .ZN(new_n12140_));
  OAI22_X1   g09127(.A1(new_n12140_), .A2(new_n10619_), .B1(pi0087), .B2(new_n12135_), .ZN(new_n12141_));
  NAND2_X1   g09128(.A1(new_n12141_), .A2(new_n5492_), .ZN(new_n12142_));
  OAI21_X1   g09129(.A1(new_n5490_), .A2(new_n3258_), .B(new_n3208_), .ZN(new_n12143_));
  AOI21_X1   g09130(.A1(new_n12143_), .A2(new_n5488_), .B(new_n5767_), .ZN(new_n12144_));
  NOR4_X1    g09131(.A1(new_n5497_), .A2(new_n12144_), .A3(new_n6289_), .A4(new_n6297_), .ZN(new_n12145_));
  OAI21_X1   g09132(.A1(new_n12133_), .A2(new_n12142_), .B(new_n12145_), .ZN(new_n12146_));
  NAND2_X1   g09133(.A1(new_n5371_), .A2(new_n3229_), .ZN(new_n12147_));
  AOI21_X1   g09134(.A1(new_n12146_), .A2(new_n12147_), .B(new_n5544_), .ZN(po0286));
  INV_X1     g09135(.I(new_n11199_), .ZN(new_n12149_));
  AOI21_X1   g09136(.A1(new_n12149_), .A2(new_n5386_), .B(new_n11571_), .ZN(new_n12150_));
  INV_X1     g09137(.I(new_n12150_), .ZN(new_n12151_));
  NOR2_X1    g09138(.A1(new_n12151_), .A2(new_n5551_), .ZN(new_n12152_));
  INV_X1     g09139(.I(new_n7536_), .ZN(new_n12153_));
  NAND2_X1   g09140(.A1(new_n12153_), .A2(pi0232), .ZN(new_n12154_));
  XOR2_X1    g09141(.A1(new_n12152_), .A2(new_n12154_), .Z(new_n12155_));
  INV_X1     g09142(.I(new_n11704_), .ZN(new_n12156_));
  NAND2_X1   g09143(.A1(new_n11426_), .A2(new_n12156_), .ZN(new_n12157_));
  AOI21_X1   g09144(.A1(new_n12157_), .A2(new_n11361_), .B(new_n2702_), .ZN(new_n12158_));
  NAND2_X1   g09145(.A1(new_n11199_), .A2(new_n12158_), .ZN(new_n12159_));
  AOI21_X1   g09146(.A1(new_n12149_), .A2(new_n5551_), .B(pi0039), .ZN(new_n12160_));
  INV_X1     g09147(.I(new_n11875_), .ZN(new_n12161_));
  NOR2_X1    g09148(.A1(new_n12161_), .A2(new_n6459_), .ZN(new_n12162_));
  AOI21_X1   g09149(.A1(new_n5386_), .A2(new_n11427_), .B(new_n11683_), .ZN(new_n12163_));
  INV_X1     g09150(.I(new_n12163_), .ZN(new_n12164_));
  AOI21_X1   g09151(.A1(new_n12164_), .A2(new_n6459_), .B(new_n12162_), .ZN(new_n12165_));
  INV_X1     g09152(.I(new_n12165_), .ZN(new_n12166_));
  INV_X1     g09153(.I(pi0191), .ZN(new_n12167_));
  NOR2_X1    g09154(.A1(new_n12167_), .A2(pi0299), .ZN(new_n12168_));
  NOR2_X1    g09155(.A1(new_n12161_), .A2(new_n5700_), .ZN(new_n12169_));
  NAND2_X1   g09156(.A1(new_n12164_), .A2(new_n3100_), .ZN(new_n12170_));
  INV_X1     g09157(.I(new_n11657_), .ZN(new_n12171_));
  NOR2_X1    g09158(.A1(new_n12171_), .A2(new_n11876_), .ZN(new_n12172_));
  NAND2_X1   g09159(.A1(new_n12172_), .A2(pi0224), .ZN(new_n12173_));
  AOI21_X1   g09160(.A1(new_n12170_), .A2(new_n12173_), .B(new_n6544_), .ZN(new_n12174_));
  NOR2_X1    g09161(.A1(new_n12174_), .A2(new_n12169_), .ZN(new_n12175_));
  NAND2_X1   g09162(.A1(new_n12175_), .A2(new_n12168_), .ZN(new_n12176_));
  NAND2_X1   g09163(.A1(new_n12168_), .A2(pi0140), .ZN(new_n12177_));
  XOR2_X1    g09164(.A1(new_n12176_), .A2(new_n12177_), .Z(new_n12178_));
  NAND2_X1   g09165(.A1(new_n12178_), .A2(new_n12166_), .ZN(new_n12179_));
  AOI21_X1   g09166(.A1(new_n11426_), .A2(new_n6459_), .B(pi0051), .ZN(new_n12180_));
  NAND2_X1   g09167(.A1(new_n11679_), .A2(new_n11426_), .ZN(new_n12181_));
  NAND2_X1   g09168(.A1(new_n12181_), .A2(new_n2702_), .ZN(new_n12182_));
  NAND2_X1   g09169(.A1(new_n12182_), .A2(new_n7535_), .ZN(new_n12183_));
  NAND2_X1   g09170(.A1(new_n7535_), .A2(pi0140), .ZN(new_n12184_));
  XOR2_X1    g09171(.A1(new_n12183_), .A2(new_n12184_), .Z(new_n12185_));
  AOI21_X1   g09172(.A1(new_n12185_), .A2(new_n12180_), .B(pi0232), .ZN(new_n12186_));
  NOR2_X1    g09173(.A1(new_n5386_), .A2(new_n4474_), .ZN(new_n12187_));
  NAND3_X1   g09174(.A1(new_n11422_), .A2(new_n11427_), .A3(new_n12187_), .ZN(new_n12188_));
  NAND3_X1   g09175(.A1(new_n11423_), .A2(new_n11428_), .A3(new_n12187_), .ZN(new_n12189_));
  AOI21_X1   g09176(.A1(new_n8108_), .A2(new_n3011_), .B(new_n4474_), .ZN(new_n12190_));
  NAND2_X1   g09177(.A1(new_n12172_), .A2(new_n12190_), .ZN(new_n12191_));
  AOI21_X1   g09178(.A1(new_n12188_), .A2(new_n12189_), .B(new_n12191_), .ZN(new_n12192_));
  NAND2_X1   g09179(.A1(new_n11654_), .A2(new_n2702_), .ZN(new_n12193_));
  NOR3_X1    g09180(.A1(new_n12193_), .A2(pi0169), .A3(new_n3011_), .ZN(new_n12194_));
  AOI21_X1   g09181(.A1(new_n11449_), .A2(pi0169), .B(pi0051), .ZN(new_n12195_));
  NOR2_X1    g09182(.A1(new_n7440_), .A2(new_n8108_), .ZN(new_n12196_));
  NOR4_X1    g09183(.A1(new_n12195_), .A2(new_n3098_), .A3(new_n6451_), .A4(new_n12196_), .ZN(new_n12197_));
  OAI22_X1   g09184(.A1(new_n12192_), .A2(new_n12194_), .B1(new_n3361_), .B2(new_n12197_), .ZN(new_n12198_));
  AOI21_X1   g09185(.A1(new_n12179_), .A2(new_n12186_), .B(new_n12198_), .ZN(new_n12199_));
  AOI21_X1   g09186(.A1(new_n12199_), .A2(new_n12160_), .B(new_n3259_), .ZN(new_n12200_));
  OAI21_X1   g09187(.A1(new_n12155_), .A2(new_n12159_), .B(new_n12200_), .ZN(new_n12201_));
  XOR2_X1    g09188(.A1(new_n12201_), .A2(new_n5486_), .Z(new_n12202_));
  INV_X1     g09189(.I(new_n11926_), .ZN(new_n12203_));
  NOR2_X1    g09190(.A1(new_n12203_), .A2(pi0126), .ZN(new_n12204_));
  NAND2_X1   g09191(.A1(new_n11313_), .A2(pi0130), .ZN(new_n12205_));
  XOR2_X1    g09192(.A1(new_n12205_), .A2(new_n12204_), .Z(new_n12206_));
  NOR2_X1    g09193(.A1(new_n12206_), .A2(new_n11308_), .ZN(new_n12207_));
  INV_X1     g09194(.I(new_n12207_), .ZN(new_n12208_));
  NOR2_X1    g09195(.A1(new_n6494_), .A2(new_n12153_), .ZN(new_n12209_));
  NOR2_X1    g09196(.A1(new_n12209_), .A2(new_n11328_), .ZN(new_n12210_));
  NOR2_X1    g09197(.A1(new_n11875_), .A2(new_n12210_), .ZN(new_n12211_));
  NOR2_X1    g09198(.A1(new_n12211_), .A2(new_n3455_), .ZN(new_n12212_));
  NAND3_X1   g09199(.A1(new_n8032_), .A2(pi0087), .A3(new_n3287_), .ZN(new_n12213_));
  XOR2_X1    g09200(.A1(new_n12213_), .A2(new_n12212_), .Z(new_n12214_));
  NAND3_X1   g09201(.A1(new_n12211_), .A2(new_n3462_), .A3(new_n3207_), .ZN(new_n12215_));
  AOI21_X1   g09202(.A1(new_n12214_), .A2(new_n12208_), .B(new_n12215_), .ZN(new_n12216_));
  NAND2_X1   g09203(.A1(new_n12202_), .A2(new_n12216_), .ZN(new_n12217_));
  NOR2_X1    g09204(.A1(new_n11215_), .A2(pi0087), .ZN(new_n12218_));
  NAND2_X1   g09205(.A1(new_n6493_), .A2(pi0169), .ZN(new_n12219_));
  NOR2_X1    g09206(.A1(new_n12063_), .A2(pi0167), .ZN(new_n12220_));
  OAI22_X1   g09207(.A1(new_n12220_), .A2(new_n6494_), .B1(new_n12218_), .B2(new_n12219_), .ZN(new_n12221_));
  NOR2_X1    g09208(.A1(pi0051), .A2(pi0087), .ZN(new_n12222_));
  NOR4_X1    g09209(.A1(new_n11742_), .A2(new_n4474_), .A3(new_n7240_), .A4(new_n12222_), .ZN(new_n12223_));
  NAND3_X1   g09210(.A1(new_n12221_), .A2(new_n12207_), .A3(new_n12223_), .ZN(new_n12224_));
  NAND2_X1   g09211(.A1(new_n12211_), .A2(pi0100), .ZN(new_n12225_));
  NAND2_X1   g09212(.A1(new_n12225_), .A2(new_n3207_), .ZN(new_n12226_));
  NOR2_X1    g09213(.A1(new_n11809_), .A2(pi0051), .ZN(new_n12227_));
  AOI21_X1   g09214(.A1(new_n12227_), .A2(new_n12168_), .B(pi0140), .ZN(new_n12228_));
  NOR2_X1    g09215(.A1(new_n11801_), .A2(pi0051), .ZN(new_n12229_));
  AOI21_X1   g09216(.A1(new_n12229_), .A2(new_n7535_), .B(pi0140), .ZN(new_n12230_));
  OAI22_X1   g09217(.A1(new_n12228_), .A2(new_n11352_), .B1(new_n11833_), .B2(new_n12230_), .ZN(new_n12231_));
  AOI21_X1   g09218(.A1(new_n11804_), .A2(new_n2702_), .B(pi0232), .ZN(new_n12232_));
  NOR2_X1    g09219(.A1(new_n12232_), .A2(new_n8932_), .ZN(new_n12233_));
  INV_X1     g09220(.I(new_n12233_), .ZN(new_n12234_));
  NAND2_X1   g09221(.A1(new_n12210_), .A2(new_n8932_), .ZN(new_n12235_));
  NAND2_X1   g09222(.A1(new_n12235_), .A2(new_n3462_), .ZN(new_n12236_));
  OAI21_X1   g09223(.A1(new_n12234_), .A2(new_n12236_), .B(new_n5551_), .ZN(new_n12237_));
  NOR3_X1    g09224(.A1(new_n11441_), .A2(pi0051), .A3(new_n11351_), .ZN(new_n12238_));
  NOR3_X1    g09225(.A1(new_n12238_), .A2(new_n8108_), .A3(new_n7440_), .ZN(new_n12239_));
  NAND2_X1   g09226(.A1(new_n12196_), .A2(pi0169), .ZN(new_n12240_));
  XNOR2_X1   g09227(.A1(new_n12239_), .A2(new_n12240_), .ZN(new_n12241_));
  INV_X1     g09228(.I(new_n12187_), .ZN(new_n12242_));
  NAND4_X1   g09229(.A1(new_n11661_), .A2(new_n8108_), .A3(new_n7439_), .A4(new_n12187_), .ZN(new_n12243_));
  NAND4_X1   g09230(.A1(new_n11662_), .A2(new_n8108_), .A3(new_n7439_), .A4(new_n12242_), .ZN(new_n12244_));
  NAND2_X1   g09231(.A1(new_n12244_), .A2(new_n12243_), .ZN(new_n12245_));
  AOI21_X1   g09232(.A1(new_n12245_), .A2(new_n3160_), .B(pi0299), .ZN(new_n12246_));
  NOR2_X1    g09233(.A1(new_n11328_), .A2(new_n7439_), .ZN(new_n12247_));
  INV_X1     g09234(.I(new_n12247_), .ZN(new_n12248_));
  NOR4_X1    g09235(.A1(new_n12246_), .A2(new_n11832_), .A3(new_n12242_), .A4(new_n12248_), .ZN(new_n12249_));
  NAND4_X1   g09236(.A1(new_n12231_), .A2(new_n12237_), .A3(new_n12241_), .A4(new_n12249_), .ZN(new_n12250_));
  AOI21_X1   g09237(.A1(new_n12250_), .A2(new_n12226_), .B(new_n11499_), .ZN(new_n12251_));
  NOR2_X1    g09238(.A1(new_n12214_), .A2(new_n11417_), .ZN(new_n12252_));
  OAI21_X1   g09239(.A1(new_n12251_), .A2(new_n12207_), .B(new_n12252_), .ZN(new_n12253_));
  AOI21_X1   g09240(.A1(new_n12217_), .A2(new_n12224_), .B(new_n12253_), .ZN(po0287));
  NOR2_X1    g09241(.A1(new_n10862_), .A2(new_n3462_), .ZN(new_n12255_));
  XOR2_X1    g09242(.A1(new_n12255_), .A2(new_n3477_), .Z(new_n12256_));
  NAND3_X1   g09243(.A1(new_n12256_), .A2(new_n3235_), .A3(new_n6285_), .ZN(new_n12257_));
  NAND2_X1   g09244(.A1(new_n6286_), .A2(pi0075), .ZN(new_n12258_));
  OAI21_X1   g09245(.A1(new_n10621_), .A2(new_n7330_), .B(pi0092), .ZN(new_n12259_));
  AOI21_X1   g09246(.A1(new_n12257_), .A2(new_n12258_), .B(new_n12259_), .ZN(po0288));
  NAND3_X1   g09247(.A1(new_n11314_), .A2(new_n12204_), .A3(new_n11308_), .ZN(new_n12261_));
  OAI21_X1   g09248(.A1(new_n11308_), .A2(new_n12204_), .B(new_n12261_), .ZN(new_n12262_));
  NOR2_X1    g09249(.A1(new_n2702_), .A2(pi0151), .ZN(new_n12263_));
  AOI21_X1   g09250(.A1(new_n10681_), .A2(new_n11230_), .B(new_n12263_), .ZN(new_n12264_));
  NAND2_X1   g09251(.A1(new_n11205_), .A2(new_n12264_), .ZN(new_n12265_));
  INV_X1     g09252(.I(new_n12265_), .ZN(new_n12266_));
  AOI22_X1   g09253(.A1(new_n12266_), .A2(new_n11175_), .B1(pi0232), .B2(new_n12262_), .ZN(new_n12267_));
  NAND2_X1   g09254(.A1(new_n11229_), .A2(pi0173), .ZN(new_n12268_));
  NAND2_X1   g09255(.A1(new_n12268_), .A2(new_n3098_), .ZN(new_n12269_));
  NOR2_X1    g09256(.A1(new_n11742_), .A2(new_n10656_), .ZN(new_n12270_));
  AOI21_X1   g09257(.A1(new_n12270_), .A2(new_n12269_), .B(pi0232), .ZN(new_n12271_));
  NOR3_X1    g09258(.A1(new_n12271_), .A2(new_n3098_), .A3(new_n12265_), .ZN(new_n12272_));
  INV_X1     g09259(.I(new_n11984_), .ZN(new_n12273_));
  OAI21_X1   g09260(.A1(new_n5373_), .A2(new_n11241_), .B(new_n11247_), .ZN(new_n12274_));
  NAND2_X1   g09261(.A1(new_n12274_), .A2(pi0173), .ZN(new_n12275_));
  NOR2_X1    g09262(.A1(new_n10664_), .A2(new_n5644_), .ZN(new_n12276_));
  XOR2_X1    g09263(.A1(new_n12275_), .A2(new_n12276_), .Z(new_n12277_));
  NOR2_X1    g09264(.A1(new_n11199_), .A2(new_n3538_), .ZN(new_n12278_));
  XOR2_X1    g09265(.A1(new_n12278_), .A2(new_n10785_), .Z(new_n12279_));
  NOR2_X1    g09266(.A1(new_n11240_), .A2(new_n5373_), .ZN(new_n12280_));
  NOR2_X1    g09267(.A1(new_n12280_), .A2(pi0160), .ZN(new_n12281_));
  NOR3_X1    g09268(.A1(new_n12263_), .A2(pi0168), .A3(new_n5373_), .ZN(new_n12282_));
  NOR4_X1    g09269(.A1(new_n12281_), .A2(new_n11191_), .A3(new_n11195_), .A4(new_n12282_), .ZN(new_n12283_));
  AOI21_X1   g09270(.A1(new_n12279_), .A2(new_n12283_), .B(pi0299), .ZN(new_n12284_));
  NOR2_X1    g09271(.A1(new_n11190_), .A2(new_n5644_), .ZN(new_n12285_));
  XNOR2_X1   g09272(.A1(new_n12285_), .A2(new_n9690_), .ZN(new_n12286_));
  AOI21_X1   g09273(.A1(new_n12286_), .A2(new_n11240_), .B(pi0173), .ZN(new_n12287_));
  INV_X1     g09274(.I(new_n12274_), .ZN(new_n12288_));
  OAI21_X1   g09275(.A1(new_n5373_), .A2(new_n11240_), .B(new_n11200_), .ZN(new_n12289_));
  NAND2_X1   g09276(.A1(new_n3538_), .A2(pi0160), .ZN(new_n12290_));
  AOI21_X1   g09277(.A1(new_n11224_), .A2(pi0168), .B(new_n12290_), .ZN(new_n12291_));
  NOR2_X1    g09278(.A1(new_n11240_), .A2(new_n12291_), .ZN(new_n12292_));
  AOI21_X1   g09279(.A1(pi0051), .A2(new_n10664_), .B(new_n5386_), .ZN(new_n12293_));
  AOI21_X1   g09280(.A1(new_n11223_), .A2(new_n12293_), .B(pi0182), .ZN(new_n12294_));
  NAND3_X1   g09281(.A1(new_n8536_), .A2(pi0168), .A3(pi0182), .ZN(new_n12295_));
  NOR4_X1    g09282(.A1(new_n10681_), .A2(new_n10656_), .A3(pi0299), .A4(new_n12295_), .ZN(new_n12296_));
  OAI21_X1   g09283(.A1(new_n12294_), .A2(new_n11161_), .B(new_n12296_), .ZN(new_n12297_));
  NOR4_X1    g09284(.A1(new_n12292_), .A2(new_n11241_), .A3(new_n5386_), .A4(new_n12297_), .ZN(new_n12298_));
  OAI21_X1   g09285(.A1(new_n11485_), .A2(new_n11181_), .B(pi0168), .ZN(new_n12299_));
  OAI21_X1   g09286(.A1(new_n12280_), .A2(new_n12299_), .B(new_n3538_), .ZN(new_n12300_));
  NAND4_X1   g09287(.A1(new_n12288_), .A2(new_n12300_), .A3(new_n12289_), .A4(new_n12298_), .ZN(new_n12301_));
  NOR4_X1    g09288(.A1(new_n12277_), .A2(new_n12284_), .A3(new_n12287_), .A4(new_n12301_), .ZN(new_n12302_));
  OAI21_X1   g09289(.A1(new_n12302_), .A2(new_n11240_), .B(new_n12273_), .ZN(new_n12303_));
  NOR2_X1    g09290(.A1(new_n11668_), .A2(new_n7375_), .ZN(new_n12304_));
  NAND2_X1   g09291(.A1(pi0173), .A2(pi0183), .ZN(new_n12305_));
  XOR2_X1    g09292(.A1(new_n12304_), .A2(new_n12305_), .Z(new_n12306_));
  AOI21_X1   g09293(.A1(new_n7375_), .A2(new_n6461_), .B(new_n11293_), .ZN(new_n12308_));
  NAND2_X1   g09294(.A1(new_n11230_), .A2(new_n7375_), .ZN(new_n12309_));
  OAI21_X1   g09295(.A1(new_n11671_), .A2(new_n12309_), .B(new_n10664_), .ZN(new_n12310_));
  NOR2_X1    g09296(.A1(new_n10656_), .A2(pi0299), .ZN(new_n12311_));
  NOR2_X1    g09297(.A1(new_n7375_), .A2(new_n10656_), .ZN(new_n12312_));
  NAND4_X1   g09298(.A1(new_n6459_), .A2(pi0299), .A3(new_n12311_), .A4(new_n12312_), .ZN(new_n12313_));
  AOI21_X1   g09299(.A1(new_n11692_), .A2(new_n10664_), .B(new_n12313_), .ZN(new_n12314_));
  AND3_X2    g09300(.A1(new_n11681_), .A2(new_n12310_), .A3(new_n12314_), .Z(new_n12315_));
  OAI21_X1   g09301(.A1(new_n12315_), .A2(new_n12308_), .B(new_n11665_), .ZN(new_n12316_));
  OAI21_X1   g09302(.A1(new_n12265_), .A2(new_n3362_), .B(new_n3011_), .ZN(new_n12317_));
  AOI21_X1   g09303(.A1(new_n12317_), .A2(pi0149), .B(pi0299), .ZN(new_n12318_));
  OAI21_X1   g09304(.A1(new_n12306_), .A2(new_n12316_), .B(new_n12318_), .ZN(new_n12319_));
  NOR2_X1    g09305(.A1(new_n11347_), .A2(new_n4635_), .ZN(new_n12320_));
  XOR2_X1    g09306(.A1(new_n12320_), .A2(new_n10785_), .Z(new_n12321_));
  NAND2_X1   g09307(.A1(new_n11378_), .A2(new_n12321_), .ZN(new_n12322_));
  NOR2_X1    g09308(.A1(new_n11657_), .A2(new_n3538_), .ZN(new_n12323_));
  XOR2_X1    g09309(.A1(new_n12323_), .A2(new_n10785_), .Z(new_n12324_));
  AOI21_X1   g09310(.A1(new_n12324_), .A2(new_n11656_), .B(new_n7475_), .ZN(new_n12325_));
  AOI21_X1   g09311(.A1(new_n12325_), .A2(new_n12322_), .B(new_n3362_), .ZN(new_n12326_));
  XOR2_X1    g09312(.A1(new_n12326_), .A2(new_n7439_), .Z(new_n12327_));
  NAND2_X1   g09313(.A1(new_n11684_), .A2(pi0168), .ZN(new_n12328_));
  NAND2_X1   g09314(.A1(new_n12263_), .A2(pi0168), .ZN(new_n12329_));
  XOR2_X1    g09315(.A1(new_n12328_), .A2(new_n12329_), .Z(new_n12330_));
  NAND4_X1   g09316(.A1(new_n12319_), .A2(new_n11980_), .A3(new_n12327_), .A4(new_n12330_), .ZN(new_n12331_));
  AOI21_X1   g09317(.A1(new_n12303_), .A2(new_n5551_), .B(new_n12331_), .ZN(new_n12332_));
  NOR2_X1    g09318(.A1(new_n12332_), .A2(new_n3208_), .ZN(new_n12333_));
  NAND2_X1   g09319(.A1(new_n3207_), .A2(new_n3132_), .ZN(new_n12334_));
  XNOR2_X1   g09320(.A1(new_n12333_), .A2(new_n12334_), .ZN(new_n12335_));
  NAND2_X1   g09321(.A1(new_n12335_), .A2(new_n12272_), .ZN(new_n12336_));
  OAI21_X1   g09322(.A1(new_n7504_), .A2(new_n3455_), .B(new_n12262_), .ZN(new_n12337_));
  NAND2_X1   g09323(.A1(new_n12272_), .A2(new_n11321_), .ZN(new_n12338_));
  AOI21_X1   g09324(.A1(new_n12336_), .A2(new_n12337_), .B(new_n12338_), .ZN(new_n12339_));
  INV_X1     g09325(.I(new_n11804_), .ZN(new_n12340_));
  NAND2_X1   g09326(.A1(new_n12268_), .A2(new_n10768_), .ZN(new_n12341_));
  NAND2_X1   g09327(.A1(new_n11802_), .A2(new_n12341_), .ZN(new_n12342_));
  NOR2_X1    g09328(.A1(new_n11473_), .A2(new_n7375_), .ZN(new_n12343_));
  NOR2_X1    g09329(.A1(new_n11810_), .A2(pi0173), .ZN(new_n12344_));
  NAND2_X1   g09330(.A1(new_n11460_), .A2(pi0183), .ZN(new_n12345_));
  NOR2_X1    g09331(.A1(new_n11822_), .A2(new_n10664_), .ZN(new_n12346_));
  XOR2_X1    g09332(.A1(new_n12346_), .A2(new_n12305_), .Z(new_n12347_));
  OAI22_X1   g09333(.A1(new_n12344_), .A2(new_n12345_), .B1(new_n12347_), .B2(new_n11830_), .ZN(new_n12348_));
  AOI22_X1   g09334(.A1(new_n12348_), .A2(new_n12311_), .B1(new_n12342_), .B2(new_n12343_), .ZN(new_n12349_));
  AOI21_X1   g09335(.A1(pi0149), .A2(pi0168), .B(new_n11472_), .ZN(new_n12350_));
  NAND2_X1   g09336(.A1(new_n12264_), .A2(new_n7439_), .ZN(new_n12351_));
  OAI21_X1   g09337(.A1(new_n12350_), .A2(new_n12351_), .B(new_n4635_), .ZN(new_n12352_));
  OAI21_X1   g09338(.A1(new_n2702_), .A2(pi0151), .B(new_n11655_), .ZN(new_n12353_));
  NAND3_X1   g09339(.A1(new_n12352_), .A2(new_n11430_), .A3(new_n12353_), .ZN(new_n12354_));
  OAI21_X1   g09340(.A1(new_n11427_), .A2(new_n10681_), .B(new_n3538_), .ZN(new_n12355_));
  NOR2_X1    g09341(.A1(new_n11423_), .A2(new_n10681_), .ZN(new_n12356_));
  AOI21_X1   g09342(.A1(new_n12356_), .A2(new_n12355_), .B(pi0149), .ZN(new_n12357_));
  NAND2_X1   g09343(.A1(new_n12354_), .A2(new_n12357_), .ZN(new_n12358_));
  INV_X1     g09344(.I(new_n10785_), .ZN(new_n12359_));
  NAND2_X1   g09345(.A1(new_n11431_), .A2(pi0151), .ZN(new_n12360_));
  XOR2_X1    g09346(.A1(new_n12360_), .A2(new_n12359_), .Z(new_n12361_));
  NOR3_X1    g09347(.A1(new_n11175_), .A2(pi0299), .A3(new_n9241_), .ZN(new_n12362_));
  NOR2_X1    g09348(.A1(new_n12265_), .A2(new_n12362_), .ZN(new_n12363_));
  NAND4_X1   g09349(.A1(new_n12361_), .A2(new_n11955_), .A3(new_n12358_), .A4(new_n12363_), .ZN(new_n12364_));
  OAI21_X1   g09350(.A1(new_n12349_), .A2(new_n12364_), .B(pi0039), .ZN(new_n12365_));
  XOR2_X1    g09351(.A1(new_n12365_), .A2(new_n11361_), .Z(new_n12366_));
  NAND2_X1   g09352(.A1(new_n12366_), .A2(new_n12340_), .ZN(new_n12367_));
  INV_X1     g09353(.I(new_n12272_), .ZN(new_n12368_));
  NAND2_X1   g09354(.A1(new_n12368_), .A2(new_n12334_), .ZN(new_n12369_));
  AOI21_X1   g09355(.A1(new_n12369_), .A2(new_n11175_), .B(new_n3132_), .ZN(new_n12370_));
  NAND2_X1   g09356(.A1(new_n11369_), .A2(pi0151), .ZN(new_n12371_));
  XOR2_X1    g09357(.A1(new_n12371_), .A2(new_n12359_), .Z(new_n12372_));
  NAND2_X1   g09358(.A1(new_n11275_), .A2(new_n4635_), .ZN(new_n12373_));
  INV_X1     g09359(.I(new_n11729_), .ZN(new_n12374_));
  NAND2_X1   g09360(.A1(new_n12374_), .A2(new_n5664_), .ZN(new_n12375_));
  NOR3_X1    g09361(.A1(new_n11207_), .A2(new_n3538_), .A3(new_n11230_), .ZN(new_n12376_));
  NAND4_X1   g09362(.A1(new_n12372_), .A2(new_n12373_), .A3(new_n12375_), .A4(new_n12376_), .ZN(new_n12377_));
  OAI21_X1   g09363(.A1(new_n2702_), .A2(pi0173), .B(new_n12311_), .ZN(new_n12378_));
  OAI21_X1   g09364(.A1(new_n11729_), .A2(new_n12378_), .B(new_n11275_), .ZN(new_n12379_));
  NAND4_X1   g09365(.A1(new_n12266_), .A2(pi0168), .A3(pi0182), .A4(pi0232), .ZN(new_n12380_));
  AOI21_X1   g09366(.A1(new_n11207_), .A2(new_n12341_), .B(new_n12380_), .ZN(new_n12381_));
  OAI21_X1   g09367(.A1(new_n12374_), .A2(new_n3538_), .B(new_n11742_), .ZN(new_n12382_));
  NAND4_X1   g09368(.A1(new_n12382_), .A2(new_n11730_), .A3(new_n12379_), .A4(new_n12381_), .ZN(new_n12384_));
  AOI21_X1   g09369(.A1(new_n12377_), .A2(new_n3098_), .B(new_n12384_), .ZN(new_n12385_));
  NOR2_X1    g09370(.A1(new_n12272_), .A2(new_n11322_), .ZN(new_n12386_));
  NOR3_X1    g09371(.A1(po1038), .A2(pi0087), .A3(pi0164), .ZN(new_n12387_));
  NOR4_X1    g09372(.A1(new_n12262_), .A2(new_n5551_), .A3(new_n5386_), .A4(new_n12387_), .ZN(new_n12388_));
  OAI21_X1   g09373(.A1(new_n7504_), .A2(new_n3455_), .B(new_n12388_), .ZN(new_n12389_));
  NOR3_X1    g09374(.A1(new_n11207_), .A2(new_n12386_), .A3(new_n12389_), .ZN(new_n12390_));
  OAI21_X1   g09375(.A1(new_n12385_), .A2(pi0039), .B(new_n12390_), .ZN(new_n12391_));
  AOI21_X1   g09376(.A1(new_n12367_), .A2(new_n12370_), .B(new_n12391_), .ZN(new_n12392_));
  OAI21_X1   g09377(.A1(new_n12339_), .A2(po1038), .B(new_n12392_), .ZN(new_n12393_));
  AOI21_X1   g09378(.A1(new_n12393_), .A2(new_n3455_), .B(new_n12267_), .ZN(po0289));
  OAI21_X1   g09379(.A1(new_n5373_), .A2(new_n11282_), .B(new_n11193_), .ZN(new_n12395_));
  NOR3_X1    g09380(.A1(new_n12395_), .A2(pi0039), .A3(new_n7459_), .ZN(new_n12396_));
  NAND3_X1   g09381(.A1(new_n7520_), .A2(new_n3183_), .A3(pi0176), .ZN(new_n12397_));
  XOR2_X1    g09382(.A1(new_n12396_), .A2(new_n12397_), .Z(new_n12398_));
  OAI21_X1   g09383(.A1(new_n12340_), .A2(pi0232), .B(pi0039), .ZN(new_n12399_));
  OAI21_X1   g09384(.A1(pi0039), .A2(new_n11175_), .B(new_n7522_), .ZN(new_n12400_));
  OAI21_X1   g09385(.A1(new_n11174_), .A2(new_n12400_), .B(new_n3259_), .ZN(new_n12401_));
  NOR3_X1    g09386(.A1(new_n11473_), .A2(new_n5641_), .A3(new_n5551_), .ZN(new_n12402_));
  AOI21_X1   g09387(.A1(new_n12402_), .A2(new_n11801_), .B(pi0299), .ZN(new_n12403_));
  AOI21_X1   g09388(.A1(new_n11799_), .A2(new_n11175_), .B(pi0197), .ZN(new_n12404_));
  NOR3_X1    g09389(.A1(new_n12403_), .A2(new_n11352_), .A3(new_n12404_), .ZN(new_n12405_));
  NAND2_X1   g09390(.A1(new_n12405_), .A2(new_n12401_), .ZN(new_n12406_));
  OAI21_X1   g09391(.A1(new_n12399_), .A2(new_n12406_), .B(new_n3462_), .ZN(new_n12407_));
  NOR2_X1    g09392(.A1(new_n11176_), .A2(new_n3259_), .ZN(new_n12408_));
  AOI21_X1   g09393(.A1(new_n12407_), .A2(new_n12408_), .B(new_n11500_), .ZN(new_n12409_));
  NAND2_X1   g09394(.A1(new_n11322_), .A2(pi0087), .ZN(new_n12410_));
  NAND2_X1   g09395(.A1(new_n6493_), .A2(new_n7475_), .ZN(new_n12411_));
  XNOR2_X1   g09396(.A1(new_n7492_), .A2(new_n12411_), .ZN(new_n12412_));
  AOI21_X1   g09397(.A1(new_n11315_), .A2(new_n11556_), .B(pi0133), .ZN(new_n12413_));
  INV_X1     g09398(.I(new_n12413_), .ZN(new_n12414_));
  NOR2_X1    g09399(.A1(new_n12414_), .A2(new_n7375_), .ZN(new_n12415_));
  NAND2_X1   g09400(.A1(new_n12414_), .A2(new_n11416_), .ZN(new_n12416_));
  NOR2_X1    g09401(.A1(new_n7240_), .A2(new_n6494_), .ZN(new_n12418_));
  AOI22_X1   g09402(.A1(new_n12412_), .A2(new_n12415_), .B1(new_n12416_), .B2(new_n12418_), .ZN(new_n12419_));
  OAI21_X1   g09403(.A1(new_n12409_), .A2(new_n12410_), .B(new_n12419_), .ZN(new_n12420_));
  NOR3_X1    g09404(.A1(new_n3336_), .A2(new_n5551_), .A3(new_n3098_), .ZN(new_n12421_));
  INV_X1     g09405(.I(new_n12421_), .ZN(new_n12422_));
  NAND2_X1   g09406(.A1(new_n11031_), .A2(new_n5641_), .ZN(new_n12423_));
  NAND2_X1   g09407(.A1(new_n11351_), .A2(pi0221), .ZN(new_n12424_));
  AOI21_X1   g09408(.A1(pi0197), .A2(pi0216), .B(new_n6540_), .ZN(new_n12425_));
  AOI22_X1   g09409(.A1(new_n12425_), .A2(new_n12424_), .B1(new_n12423_), .B2(new_n11353_), .ZN(new_n12426_));
  NOR2_X1    g09410(.A1(new_n12426_), .A2(new_n3145_), .ZN(new_n12427_));
  NOR2_X1    g09411(.A1(new_n3145_), .A2(new_n5551_), .ZN(new_n12428_));
  XOR2_X1    g09412(.A1(new_n12427_), .A2(new_n12428_), .Z(new_n12429_));
  NOR2_X1    g09413(.A1(new_n3287_), .A2(new_n3132_), .ZN(new_n12430_));
  NAND2_X1   g09414(.A1(new_n3183_), .A2(new_n7459_), .ZN(new_n12431_));
  NAND2_X1   g09415(.A1(new_n12431_), .A2(pi0039), .ZN(new_n12432_));
  NOR4_X1    g09416(.A1(new_n11704_), .A2(new_n12422_), .A3(new_n12430_), .A4(new_n12432_), .ZN(new_n12433_));
  NAND2_X1   g09417(.A1(new_n12429_), .A2(new_n12433_), .ZN(new_n12434_));
  OAI21_X1   g09418(.A1(new_n11282_), .A2(new_n12434_), .B(new_n12422_), .ZN(new_n12435_));
  AOI21_X1   g09419(.A1(new_n3455_), .A2(new_n12414_), .B(new_n11282_), .ZN(new_n12436_));
  NAND4_X1   g09420(.A1(new_n12395_), .A2(new_n12420_), .A3(new_n12435_), .A4(new_n12436_), .ZN(new_n12437_));
  NOR2_X1    g09421(.A1(new_n12398_), .A2(new_n12437_), .ZN(po0290));
  NOR3_X1    g09422(.A1(new_n6494_), .A2(new_n3989_), .A3(new_n3098_), .ZN(new_n12439_));
  NOR3_X1    g09423(.A1(new_n6494_), .A2(pi0171), .A3(pi0299), .ZN(new_n12440_));
  OAI21_X1   g09424(.A1(new_n12439_), .A2(new_n12440_), .B(pi0192), .ZN(new_n12441_));
  INV_X1     g09425(.I(new_n12441_), .ZN(new_n12442_));
  NOR2_X1    g09426(.A1(new_n12442_), .A2(new_n11328_), .ZN(new_n12443_));
  NOR4_X1    g09427(.A1(new_n12203_), .A2(pi0126), .A3(pi0130), .A4(pi0132), .ZN(new_n12444_));
  INV_X1     g09428(.I(new_n12444_), .ZN(new_n12445_));
  NOR2_X1    g09429(.A1(new_n12445_), .A2(pi0136), .ZN(new_n12446_));
  NAND2_X1   g09430(.A1(new_n12446_), .A2(new_n11311_), .ZN(new_n12447_));
  NAND2_X1   g09431(.A1(new_n12447_), .A2(pi0134), .ZN(new_n12448_));
  NAND2_X1   g09432(.A1(pi0192), .A2(pi0299), .ZN(new_n12449_));
  INV_X1     g09433(.I(pi0192), .ZN(new_n12450_));
  NOR2_X1    g09434(.A1(new_n5386_), .A2(new_n3989_), .ZN(new_n12456_));
  NAND2_X1   g09435(.A1(new_n12247_), .A2(new_n12456_), .ZN(new_n12457_));
  INV_X1     g09436(.I(new_n12456_), .ZN(new_n12458_));
  NOR2_X1    g09437(.A1(new_n3160_), .A2(new_n5386_), .ZN(new_n12459_));
  AOI21_X1   g09438(.A1(new_n12459_), .A2(pi0171), .B(new_n7439_), .ZN(new_n12460_));
  OR3_X2     g09439(.A1(new_n11662_), .A2(new_n12458_), .A3(new_n12460_), .Z(new_n12461_));
  AOI21_X1   g09440(.A1(new_n12461_), .A2(new_n3098_), .B(new_n12457_), .ZN(new_n12462_));
  NAND2_X1   g09441(.A1(new_n3183_), .A2(new_n7489_), .ZN(new_n12463_));
  INV_X1     g09442(.I(new_n12232_), .ZN(new_n12464_));
  AOI21_X1   g09443(.A1(new_n12227_), .A2(new_n11352_), .B(new_n12450_), .ZN(new_n12465_));
  XOR2_X1    g09444(.A1(new_n12465_), .A2(new_n12449_), .Z(new_n12466_));
  NAND2_X1   g09445(.A1(new_n11833_), .A2(new_n12229_), .ZN(new_n12467_));
  OAI22_X1   g09446(.A1(new_n12466_), .A2(new_n12467_), .B1(new_n5551_), .B2(new_n12464_), .ZN(new_n12468_));
  AND2_X2    g09447(.A1(new_n12468_), .A2(new_n12462_), .Z(new_n12469_));
  NAND2_X1   g09448(.A1(new_n12161_), .A2(new_n12051_), .ZN(new_n12470_));
  NAND2_X1   g09449(.A1(new_n12470_), .A2(new_n12443_), .ZN(new_n12471_));
  OAI21_X1   g09450(.A1(new_n12471_), .A2(new_n11175_), .B(new_n3133_), .ZN(new_n12472_));
  AOI21_X1   g09451(.A1(new_n12469_), .A2(new_n12463_), .B(new_n12472_), .ZN(new_n12473_));
  NOR2_X1    g09452(.A1(new_n12238_), .A2(new_n7440_), .ZN(new_n12474_));
  NOR2_X1    g09453(.A1(new_n7440_), .A2(new_n3989_), .ZN(new_n12475_));
  XOR2_X1    g09454(.A1(new_n12474_), .A2(new_n12475_), .Z(new_n12476_));
  NAND2_X1   g09455(.A1(new_n12476_), .A2(new_n11831_), .ZN(new_n12477_));
  AOI21_X1   g09456(.A1(new_n12477_), .A2(new_n3098_), .B(new_n12457_), .ZN(new_n12478_));
  NAND2_X1   g09457(.A1(new_n3183_), .A2(new_n7489_), .ZN(new_n12479_));
  NAND3_X1   g09458(.A1(new_n12468_), .A2(new_n12478_), .A3(new_n12479_), .ZN(new_n12480_));
  OAI21_X1   g09459(.A1(new_n12473_), .A2(new_n12480_), .B(new_n12448_), .ZN(new_n12481_));
  NAND3_X1   g09460(.A1(new_n12481_), .A2(new_n11321_), .A3(new_n12443_), .ZN(new_n12482_));
  INV_X1     g09461(.I(new_n12448_), .ZN(new_n12483_));
  NAND3_X1   g09462(.A1(new_n11167_), .A2(pi0232), .A3(new_n12456_), .ZN(new_n12484_));
  NAND2_X1   g09463(.A1(po1038), .A2(new_n12222_), .ZN(new_n12485_));
  AOI21_X1   g09464(.A1(new_n12485_), .A2(new_n12484_), .B(new_n11167_), .ZN(new_n12486_));
  AOI21_X1   g09465(.A1(new_n12483_), .A2(new_n12486_), .B(po1038), .ZN(new_n12487_));
  NAND3_X1   g09466(.A1(pi0171), .A2(pi0232), .A3(pi0299), .ZN(new_n12488_));
  NAND3_X1   g09467(.A1(new_n3989_), .A2(new_n3098_), .A3(pi0232), .ZN(new_n12489_));
  AOI21_X1   g09468(.A1(new_n12489_), .A2(new_n12488_), .B(new_n12450_), .ZN(new_n12490_));
  NAND3_X1   g09469(.A1(new_n12151_), .A2(pi0039), .A3(new_n12490_), .ZN(new_n12491_));
  NAND3_X1   g09470(.A1(new_n12150_), .A2(new_n3183_), .A3(new_n12490_), .ZN(new_n12492_));
  AOI21_X1   g09471(.A1(new_n12491_), .A2(new_n12492_), .B(new_n12149_), .ZN(new_n12493_));
  INV_X1     g09472(.I(new_n12180_), .ZN(new_n12494_));
  NOR2_X1    g09473(.A1(pi0192), .A2(pi0299), .ZN(new_n12495_));
  NOR2_X1    g09474(.A1(new_n3183_), .A2(new_n7489_), .ZN(new_n12496_));
  OAI21_X1   g09475(.A1(new_n12494_), .A2(new_n12496_), .B(new_n12495_), .ZN(new_n12497_));
  NOR3_X1    g09476(.A1(new_n11423_), .A2(new_n11428_), .A3(new_n12458_), .ZN(new_n12498_));
  NOR3_X1    g09477(.A1(new_n11422_), .A2(new_n11427_), .A3(new_n12458_), .ZN(new_n12499_));
  NOR2_X1    g09478(.A1(pi0164), .A2(pi0216), .ZN(new_n12500_));
  NOR4_X1    g09479(.A1(new_n12171_), .A2(new_n3989_), .A3(new_n11876_), .A4(new_n12500_), .ZN(new_n12501_));
  OAI21_X1   g09480(.A1(new_n12498_), .A2(new_n12499_), .B(new_n12501_), .ZN(new_n12502_));
  NAND2_X1   g09481(.A1(new_n3989_), .A2(pi0216), .ZN(new_n12503_));
  OAI21_X1   g09482(.A1(new_n12193_), .A2(new_n12503_), .B(new_n12502_), .ZN(new_n12504_));
  NOR2_X1    g09483(.A1(new_n3011_), .A2(pi0164), .ZN(new_n12505_));
  NOR3_X1    g09484(.A1(new_n3362_), .A2(new_n2702_), .A3(new_n12505_), .ZN(new_n12506_));
  NOR2_X1    g09485(.A1(new_n11167_), .A2(new_n3098_), .ZN(new_n12507_));
  OAI21_X1   g09486(.A1(new_n12506_), .A2(new_n12456_), .B(new_n12507_), .ZN(new_n12508_));
  AOI21_X1   g09487(.A1(new_n12508_), .A2(new_n3362_), .B(new_n5551_), .ZN(new_n12509_));
  AOI22_X1   g09488(.A1(new_n12166_), .A2(new_n12497_), .B1(new_n12504_), .B2(new_n12509_), .ZN(new_n12510_));
  INV_X1     g09489(.I(new_n12175_), .ZN(new_n12511_));
  OAI21_X1   g09490(.A1(new_n12182_), .A2(new_n7489_), .B(new_n12495_), .ZN(new_n12512_));
  OAI21_X1   g09491(.A1(new_n12443_), .A2(new_n11875_), .B(new_n11321_), .ZN(new_n12513_));
  AOI21_X1   g09492(.A1(new_n12448_), .A2(new_n12513_), .B(new_n12471_), .ZN(new_n12514_));
  NAND4_X1   g09493(.A1(new_n12511_), .A2(new_n12158_), .A3(new_n12512_), .A4(new_n12514_), .ZN(new_n12515_));
  NOR2_X1    g09494(.A1(new_n12515_), .A2(new_n12510_), .ZN(new_n12516_));
  OAI21_X1   g09495(.A1(new_n12493_), .A2(new_n3132_), .B(new_n12516_), .ZN(new_n12517_));
  AOI21_X1   g09496(.A1(new_n12482_), .A2(new_n12487_), .B(new_n12517_), .ZN(po0291));
  NOR2_X1    g09497(.A1(new_n5386_), .A2(new_n4150_), .ZN(new_n12519_));
  INV_X1     g09498(.I(new_n12519_), .ZN(new_n12520_));
  AOI21_X1   g09499(.A1(new_n11328_), .A2(new_n8648_), .B(new_n12520_), .ZN(new_n12521_));
  INV_X1     g09500(.I(pi0194), .ZN(new_n12522_));
  NAND2_X1   g09501(.A1(new_n6494_), .A2(new_n12522_), .ZN(new_n12523_));
  OAI21_X1   g09502(.A1(new_n12521_), .A2(new_n12523_), .B(pi0299), .ZN(new_n12524_));
  NOR3_X1    g09503(.A1(new_n12149_), .A2(new_n4150_), .A3(new_n8648_), .ZN(new_n12525_));
  AOI21_X1   g09504(.A1(new_n12525_), .A2(new_n12160_), .B(pi0170), .ZN(new_n12526_));
  NAND2_X1   g09505(.A1(new_n12150_), .A2(new_n5551_), .ZN(new_n12527_));
  NOR2_X1    g09506(.A1(new_n3259_), .A2(new_n12522_), .ZN(new_n12528_));
  NOR2_X1    g09507(.A1(new_n11875_), .A2(new_n12528_), .ZN(new_n12529_));
  OAI21_X1   g09508(.A1(new_n11328_), .A2(new_n6494_), .B(new_n3098_), .ZN(new_n12530_));
  NAND2_X1   g09509(.A1(new_n12530_), .A2(pi0170), .ZN(new_n12531_));
  NOR3_X1    g09510(.A1(new_n12529_), .A2(new_n3259_), .A3(new_n12531_), .ZN(new_n12532_));
  AOI21_X1   g09511(.A1(new_n12527_), .A2(pi0299), .B(new_n12532_), .ZN(new_n12533_));
  NAND2_X1   g09512(.A1(pi0185), .A2(pi0299), .ZN(new_n12534_));
  NAND2_X1   g09513(.A1(new_n12175_), .A2(pi0185), .ZN(new_n12535_));
  XOR2_X1    g09514(.A1(new_n12535_), .A2(new_n12534_), .Z(new_n12536_));
  NOR2_X1    g09515(.A1(new_n12172_), .A2(new_n3011_), .ZN(new_n12537_));
  NOR2_X1    g09516(.A1(new_n4150_), .A2(new_n3011_), .ZN(new_n12538_));
  XOR2_X1    g09517(.A1(new_n12537_), .A2(new_n12538_), .Z(new_n12539_));
  NAND2_X1   g09518(.A1(new_n11428_), .A2(new_n12520_), .ZN(new_n12540_));
  NAND3_X1   g09519(.A1(new_n6453_), .A2(new_n4150_), .A3(new_n5386_), .ZN(new_n12541_));
  NAND3_X1   g09520(.A1(new_n11422_), .A2(new_n12540_), .A3(new_n12541_), .ZN(new_n12542_));
  NAND2_X1   g09521(.A1(new_n12542_), .A2(new_n7440_), .ZN(new_n12543_));
  OAI21_X1   g09522(.A1(new_n12520_), .A2(new_n11166_), .B(new_n2702_), .ZN(new_n12544_));
  NAND4_X1   g09523(.A1(new_n3361_), .A2(pi0150), .A3(pi0216), .A4(pi0299), .ZN(new_n12545_));
  OR3_X2     g09524(.A1(new_n12542_), .A2(new_n12544_), .A3(new_n12545_), .Z(new_n12546_));
  AOI21_X1   g09525(.A1(new_n12546_), .A2(new_n12543_), .B(new_n12193_), .ZN(new_n12547_));
  AND2_X2    g09526(.A1(new_n12158_), .A2(pi0232), .Z(new_n12548_));
  AOI21_X1   g09527(.A1(new_n12539_), .A2(new_n12547_), .B(new_n12548_), .ZN(new_n12549_));
  INV_X1     g09528(.I(new_n12521_), .ZN(new_n12550_));
  NOR4_X1    g09529(.A1(new_n12549_), .A2(new_n12165_), .A3(new_n12529_), .A4(new_n12550_), .ZN(new_n12551_));
  NAND2_X1   g09530(.A1(new_n12536_), .A2(new_n12551_), .ZN(new_n12552_));
  OAI21_X1   g09531(.A1(new_n12533_), .A2(new_n12552_), .B(new_n3259_), .ZN(new_n12553_));
  INV_X1     g09532(.I(new_n12526_), .ZN(new_n12554_));
  NAND2_X1   g09533(.A1(new_n12182_), .A2(pi0185), .ZN(new_n12555_));
  XOR2_X1    g09534(.A1(new_n12555_), .A2(new_n12534_), .Z(new_n12556_));
  NOR2_X1    g09535(.A1(new_n12549_), .A2(new_n12494_), .ZN(new_n12557_));
  NAND4_X1   g09536(.A1(new_n12554_), .A2(new_n12151_), .A3(new_n12556_), .A4(new_n12557_), .ZN(new_n12558_));
  NOR2_X1    g09537(.A1(new_n12446_), .A2(new_n11311_), .ZN(new_n12559_));
  NOR2_X1    g09538(.A1(new_n12447_), .A2(new_n11310_), .ZN(new_n12560_));
  NOR2_X1    g09539(.A1(new_n3207_), .A2(pi0100), .ZN(new_n12562_));
  OAI21_X1   g09540(.A1(new_n12161_), .A2(new_n12524_), .B(new_n3462_), .ZN(new_n12563_));
  NAND2_X1   g09541(.A1(new_n11199_), .A2(new_n12563_), .ZN(new_n12564_));
  AOI21_X1   g09542(.A1(new_n12558_), .A2(new_n3098_), .B(new_n12564_), .ZN(new_n12565_));
  NOR2_X1    g09543(.A1(new_n12560_), .A2(new_n12559_), .ZN(new_n12566_));
  NOR2_X1    g09544(.A1(new_n12566_), .A2(new_n12485_), .ZN(new_n12567_));
  NOR2_X1    g09545(.A1(new_n12485_), .A2(new_n11167_), .ZN(new_n12568_));
  XNOR2_X1   g09546(.A1(new_n12567_), .A2(new_n12568_), .ZN(new_n12569_));
  NAND2_X1   g09547(.A1(new_n6493_), .A2(pi0170), .ZN(new_n12570_));
  OAI21_X1   g09548(.A1(new_n12569_), .A2(new_n12570_), .B(new_n7240_), .ZN(new_n12571_));
  AOI21_X1   g09549(.A1(new_n12565_), .A2(new_n12553_), .B(new_n12571_), .ZN(new_n12572_));
  AOI21_X1   g09550(.A1(new_n12161_), .A2(new_n12562_), .B(new_n12524_), .ZN(new_n12573_));
  OAI21_X1   g09551(.A1(new_n12550_), .A2(new_n8931_), .B(new_n12522_), .ZN(new_n12574_));
  OAI21_X1   g09552(.A1(new_n12531_), .A2(new_n8931_), .B(pi0194), .ZN(new_n12575_));
  NAND2_X1   g09553(.A1(new_n12575_), .A2(new_n12574_), .ZN(new_n12576_));
  NAND2_X1   g09554(.A1(pi0150), .A2(pi0299), .ZN(new_n12577_));
  NAND2_X1   g09555(.A1(new_n7439_), .A2(pi0170), .ZN(new_n12578_));
  XOR2_X1    g09556(.A1(new_n12474_), .A2(new_n12578_), .Z(new_n12579_));
  OAI21_X1   g09557(.A1(new_n12579_), .A2(new_n11832_), .B(pi0299), .ZN(new_n12580_));
  XOR2_X1    g09558(.A1(new_n12580_), .A2(new_n12577_), .Z(new_n12581_));
  NAND2_X1   g09559(.A1(new_n12459_), .A2(pi0170), .ZN(new_n12582_));
  NAND2_X1   g09560(.A1(new_n12582_), .A2(new_n7440_), .ZN(new_n12583_));
  NAND4_X1   g09561(.A1(new_n12581_), .A2(new_n11661_), .A3(new_n12519_), .A4(new_n12583_), .ZN(new_n12584_));
  NAND2_X1   g09562(.A1(new_n12247_), .A2(new_n12519_), .ZN(new_n12585_));
  AOI21_X1   g09563(.A1(new_n12584_), .A2(new_n12576_), .B(new_n12585_), .ZN(new_n12586_));
  INV_X1     g09564(.I(new_n12227_), .ZN(new_n12587_));
  OAI21_X1   g09565(.A1(new_n12587_), .A2(new_n12575_), .B(new_n10659_), .ZN(new_n12588_));
  NAND3_X1   g09566(.A1(new_n12588_), .A2(pi0299), .A3(new_n11351_), .ZN(new_n12589_));
  OAI21_X1   g09567(.A1(new_n11833_), .A2(new_n10659_), .B(new_n12229_), .ZN(new_n12590_));
  AOI21_X1   g09568(.A1(new_n12589_), .A2(new_n12574_), .B(new_n12590_), .ZN(new_n12591_));
  OAI21_X1   g09569(.A1(new_n12586_), .A2(new_n12591_), .B(pi0232), .ZN(new_n12592_));
  NAND2_X1   g09570(.A1(new_n12234_), .A2(new_n12576_), .ZN(new_n12593_));
  NAND2_X1   g09571(.A1(new_n12592_), .A2(new_n12593_), .ZN(new_n12594_));
  NAND2_X1   g09572(.A1(new_n12594_), .A2(new_n12573_), .ZN(new_n12595_));
  NAND2_X1   g09573(.A1(new_n12573_), .A2(pi0100), .ZN(new_n12596_));
  XOR2_X1    g09574(.A1(new_n12595_), .A2(new_n12596_), .Z(new_n12597_));
  AOI21_X1   g09575(.A1(new_n12597_), .A2(new_n11175_), .B(new_n12566_), .ZN(new_n12598_));
  NOR4_X1    g09576(.A1(new_n12598_), .A2(new_n11408_), .A3(new_n12524_), .A4(new_n12572_), .ZN(po0292));
  NAND2_X1   g09577(.A1(new_n11310_), .A2(new_n11312_), .ZN(new_n12600_));
  OAI21_X1   g09578(.A1(new_n12445_), .A2(new_n12600_), .B(new_n11311_), .ZN(new_n12601_));
  XOR2_X1    g09579(.A1(new_n12601_), .A2(new_n11310_), .Z(new_n12602_));
  INV_X1     g09580(.I(new_n12602_), .ZN(new_n12603_));
  NOR2_X1    g09581(.A1(new_n8068_), .A2(new_n5551_), .ZN(new_n12604_));
  XOR2_X1    g09582(.A1(new_n12152_), .A2(new_n12604_), .Z(new_n12605_));
  NAND2_X1   g09583(.A1(new_n12182_), .A2(new_n8067_), .ZN(new_n12606_));
  NAND2_X1   g09584(.A1(new_n8067_), .A2(pi0184), .ZN(new_n12607_));
  XNOR2_X1   g09585(.A1(new_n12606_), .A2(new_n12607_), .ZN(new_n12608_));
  NOR2_X1    g09586(.A1(new_n7439_), .A2(new_n11412_), .ZN(new_n12609_));
  OAI21_X1   g09587(.A1(pi0051), .A2(pi0148), .B(pi0287), .ZN(new_n12610_));
  NOR2_X1    g09588(.A1(new_n12609_), .A2(new_n12610_), .ZN(new_n12611_));
  AOI21_X1   g09589(.A1(new_n11426_), .A2(new_n12611_), .B(pi0299), .ZN(new_n12612_));
  OAI21_X1   g09590(.A1(new_n12608_), .A2(new_n12494_), .B(new_n12612_), .ZN(new_n12613_));
  NAND3_X1   g09591(.A1(new_n6453_), .A2(new_n9456_), .A3(new_n3362_), .ZN(new_n12614_));
  AOI21_X1   g09592(.A1(new_n12172_), .A2(new_n12614_), .B(pi0148), .ZN(new_n12615_));
  NOR3_X1    g09593(.A1(new_n12163_), .A2(new_n12615_), .A3(new_n6453_), .ZN(new_n12616_));
  AOI21_X1   g09594(.A1(new_n12613_), .A2(new_n12616_), .B(new_n12548_), .ZN(new_n12617_));
  INV_X1     g09595(.I(pi0141), .ZN(new_n12618_));
  NOR2_X1    g09596(.A1(new_n12618_), .A2(pi0299), .ZN(new_n12619_));
  INV_X1     g09597(.I(new_n12619_), .ZN(new_n12620_));
  NOR3_X1    g09598(.A1(new_n12175_), .A2(new_n9471_), .A3(new_n12620_), .ZN(new_n12621_));
  NOR3_X1    g09599(.A1(new_n12511_), .A2(pi0184), .A3(new_n12620_), .ZN(new_n12622_));
  OAI21_X1   g09600(.A1(new_n12622_), .A2(new_n12621_), .B(new_n12166_), .ZN(new_n12623_));
  OAI21_X1   g09601(.A1(new_n12623_), .A2(new_n12617_), .B(new_n3133_), .ZN(new_n12624_));
  NAND4_X1   g09602(.A1(new_n12605_), .A2(new_n11199_), .A3(new_n12160_), .A4(new_n12624_), .ZN(new_n12625_));
  AOI21_X1   g09603(.A1(new_n8069_), .A2(new_n11167_), .B(pi0051), .ZN(new_n12626_));
  NAND2_X1   g09604(.A1(new_n12626_), .A2(new_n3132_), .ZN(new_n12627_));
  AOI21_X1   g09605(.A1(new_n12625_), .A2(new_n3208_), .B(new_n12627_), .ZN(new_n12628_));
  INV_X1     g09606(.I(new_n12626_), .ZN(new_n12629_));
  NOR2_X1    g09607(.A1(new_n12629_), .A2(new_n11408_), .ZN(new_n12630_));
  OAI21_X1   g09608(.A1(new_n12628_), .A2(new_n12603_), .B(new_n12630_), .ZN(new_n12631_));
  OAI21_X1   g09609(.A1(new_n6494_), .A2(new_n4329_), .B(new_n11167_), .ZN(new_n12632_));
  OAI21_X1   g09610(.A1(new_n12485_), .A2(new_n12632_), .B(new_n12602_), .ZN(new_n12633_));
  AOI21_X1   g09611(.A1(new_n12633_), .A2(new_n11215_), .B(po1038), .ZN(new_n12634_));
  AOI21_X1   g09612(.A1(new_n12229_), .A2(new_n8067_), .B(pi0184), .ZN(new_n12635_));
  NOR2_X1    g09613(.A1(new_n11833_), .A2(new_n12635_), .ZN(new_n12636_));
  OAI21_X1   g09614(.A1(new_n12587_), .A2(new_n12620_), .B(new_n9471_), .ZN(new_n12637_));
  AOI21_X1   g09615(.A1(new_n12637_), .A2(new_n11351_), .B(new_n12636_), .ZN(new_n12638_));
  NAND2_X1   g09616(.A1(new_n11799_), .A2(new_n2702_), .ZN(new_n12639_));
  NAND2_X1   g09617(.A1(new_n12639_), .A2(new_n4329_), .ZN(new_n12640_));
  OAI21_X1   g09618(.A1(new_n12248_), .A2(new_n5373_), .B(pi0148), .ZN(new_n12641_));
  NOR2_X1    g09619(.A1(new_n7439_), .A2(pi0051), .ZN(new_n12642_));
  AOI22_X1   g09620(.A1(new_n12641_), .A2(new_n12642_), .B1(new_n5401_), .B2(new_n11412_), .ZN(new_n12643_));
  NAND3_X1   g09621(.A1(new_n11441_), .A2(new_n12640_), .A3(new_n12643_), .ZN(new_n12644_));
  NAND3_X1   g09622(.A1(pi0148), .A2(pi0232), .A3(pi0299), .ZN(new_n12645_));
  AOI21_X1   g09623(.A1(new_n12644_), .A2(new_n11328_), .B(new_n12645_), .ZN(new_n12646_));
  OAI21_X1   g09624(.A1(new_n12233_), .A2(pi0100), .B(new_n12646_), .ZN(new_n12647_));
  NOR3_X1    g09625(.A1(new_n12603_), .A2(new_n11321_), .A3(new_n12626_), .ZN(new_n12648_));
  NAND2_X1   g09626(.A1(new_n3207_), .A2(new_n11166_), .ZN(new_n12649_));
  OAI22_X1   g09627(.A1(new_n12638_), .A2(new_n12647_), .B1(new_n12648_), .B2(new_n12649_), .ZN(new_n12650_));
  NAND2_X1   g09628(.A1(new_n12629_), .A2(new_n11167_), .ZN(new_n12651_));
  NAND4_X1   g09629(.A1(new_n12650_), .A2(pi0100), .A3(new_n8931_), .A4(new_n12651_), .ZN(new_n12652_));
  AOI21_X1   g09630(.A1(new_n12631_), .A2(new_n12634_), .B(new_n12652_), .ZN(po0293));
  NOR2_X1    g09631(.A1(po1038), .A2(pi0299), .ZN(new_n12654_));
  INV_X1     g09632(.I(new_n12654_), .ZN(new_n12655_));
  NAND3_X1   g09633(.A1(new_n9365_), .A2(new_n2777_), .A3(pi0299), .ZN(new_n12656_));
  NAND3_X1   g09634(.A1(new_n12655_), .A2(new_n12656_), .A3(new_n9423_), .ZN(new_n12657_));
  NAND2_X1   g09635(.A1(po1038), .A2(pi0198), .ZN(new_n12658_));
  NOR3_X1    g09636(.A1(new_n9366_), .A2(pi0210), .A3(new_n12658_), .ZN(new_n12659_));
  AOI21_X1   g09637(.A1(new_n12657_), .A2(new_n12659_), .B(new_n11543_), .ZN(new_n12660_));
  OAI21_X1   g09638(.A1(new_n12660_), .A2(new_n8639_), .B(pi0039), .ZN(new_n12661_));
  NAND2_X1   g09639(.A1(new_n8536_), .A2(pi0137), .ZN(new_n12662_));
  XOR2_X1    g09640(.A1(new_n12661_), .A2(new_n12662_), .Z(po0294));
  NAND2_X1   g09641(.A1(new_n9221_), .A2(new_n5385_), .ZN(new_n12664_));
  OAI21_X1   g09642(.A1(new_n12664_), .A2(new_n7451_), .B(new_n12619_), .ZN(new_n12665_));
  NOR2_X1    g09643(.A1(new_n4329_), .A2(new_n3098_), .ZN(new_n12666_));
  AOI21_X1   g09644(.A1(new_n6448_), .A2(new_n12666_), .B(new_n5551_), .ZN(new_n12667_));
  NAND2_X1   g09645(.A1(new_n12665_), .A2(new_n12667_), .ZN(new_n12668_));
  NAND4_X1   g09646(.A1(new_n9283_), .A2(new_n12668_), .A3(pi0232), .A4(new_n12620_), .ZN(new_n12669_));
  NAND2_X1   g09647(.A1(new_n12669_), .A2(new_n8346_), .ZN(new_n12670_));
  XNOR2_X1   g09648(.A1(new_n12670_), .A2(new_n9285_), .ZN(new_n12671_));
  NOR2_X1    g09649(.A1(new_n7424_), .A2(new_n3138_), .ZN(new_n12672_));
  INV_X1     g09650(.I(new_n12672_), .ZN(new_n12673_));
  NOR3_X1    g09651(.A1(new_n12671_), .A2(new_n8069_), .A3(new_n12673_), .ZN(new_n12674_));
  NAND3_X1   g09652(.A1(new_n7675_), .A2(pi0299), .A3(new_n5373_), .ZN(new_n12675_));
  NAND3_X1   g09653(.A1(new_n7676_), .A2(new_n3098_), .A3(new_n5373_), .ZN(new_n12676_));
  NAND2_X1   g09654(.A1(new_n12676_), .A2(new_n12675_), .ZN(new_n12677_));
  NAND2_X1   g09655(.A1(new_n12677_), .A2(new_n8131_), .ZN(new_n12678_));
  NOR2_X1    g09656(.A1(new_n7775_), .A2(new_n5386_), .ZN(new_n12679_));
  INV_X1     g09657(.I(new_n8131_), .ZN(new_n12683_));
  NOR2_X1    g09658(.A1(new_n7854_), .A2(new_n3098_), .ZN(new_n12684_));
  XOR2_X1    g09659(.A1(new_n12684_), .A2(new_n6216_), .Z(new_n12685_));
  OAI21_X1   g09660(.A1(new_n12685_), .A2(new_n12683_), .B(new_n3183_), .ZN(new_n12686_));
  INV_X1     g09661(.I(new_n12686_), .ZN(new_n12687_));
  NOR2_X1    g09662(.A1(new_n8131_), .A2(pi0299), .ZN(new_n12688_));
  NOR2_X1    g09663(.A1(new_n12678_), .A2(new_n12618_), .ZN(new_n12689_));
  INV_X1     g09664(.I(new_n10805_), .ZN(new_n12690_));
  NOR2_X1    g09665(.A1(new_n7613_), .A2(new_n9746_), .ZN(new_n12691_));
  NAND4_X1   g09666(.A1(new_n12691_), .A2(new_n7450_), .A3(new_n7634_), .A4(new_n7576_), .ZN(new_n12692_));
  INV_X1     g09667(.I(new_n12692_), .ZN(new_n12693_));
  NOR2_X1    g09668(.A1(new_n12693_), .A2(new_n12690_), .ZN(new_n12694_));
  INV_X1     g09669(.I(new_n12694_), .ZN(new_n12695_));
  AOI21_X1   g09670(.A1(new_n7613_), .A2(new_n7439_), .B(new_n5454_), .ZN(new_n12696_));
  INV_X1     g09671(.I(new_n12696_), .ZN(new_n12697_));
  AOI21_X1   g09672(.A1(new_n12697_), .A2(new_n9746_), .B(new_n7604_), .ZN(new_n12698_));
  INV_X1     g09673(.I(new_n12698_), .ZN(new_n12699_));
  AOI21_X1   g09674(.A1(new_n12695_), .A2(new_n12699_), .B(pi0232), .ZN(new_n12700_));
  AOI21_X1   g09675(.A1(new_n12700_), .A2(pi0039), .B(pi0232), .ZN(new_n12701_));
  NOR3_X1    g09676(.A1(new_n12692_), .A2(new_n7624_), .A3(new_n10805_), .ZN(new_n12702_));
  NOR2_X1    g09677(.A1(new_n12694_), .A2(new_n12618_), .ZN(new_n12703_));
  NOR2_X1    g09678(.A1(new_n7618_), .A2(new_n12691_), .ZN(new_n12704_));
  INV_X1     g09679(.I(new_n12704_), .ZN(new_n12705_));
  NAND3_X1   g09680(.A1(new_n12705_), .A2(pi0148), .A3(new_n7603_), .ZN(new_n12706_));
  NAND4_X1   g09681(.A1(new_n12706_), .A2(new_n12699_), .A3(pi0148), .A4(new_n12619_), .ZN(new_n12707_));
  XNOR2_X1   g09682(.A1(new_n12707_), .A2(new_n12703_), .ZN(new_n12708_));
  NAND2_X1   g09683(.A1(new_n12708_), .A2(new_n12702_), .ZN(new_n12709_));
  OAI21_X1   g09684(.A1(new_n6313_), .A2(new_n7943_), .B(new_n7933_), .ZN(new_n12710_));
  NOR2_X1    g09685(.A1(new_n8103_), .A2(new_n3258_), .ZN(new_n12711_));
  OAI21_X1   g09686(.A1(new_n7933_), .A2(new_n12711_), .B(pi0092), .ZN(new_n12712_));
  OAI21_X1   g09687(.A1(new_n3258_), .A2(new_n12712_), .B(new_n12710_), .ZN(new_n12713_));
  OAI21_X1   g09688(.A1(new_n7576_), .A2(new_n3694_), .B(new_n3132_), .ZN(new_n12714_));
  OAI21_X1   g09689(.A1(new_n12714_), .A2(new_n3303_), .B(new_n3455_), .ZN(new_n12715_));
  AND3_X2    g09690(.A1(new_n12713_), .A2(new_n3132_), .A3(new_n12715_), .Z(new_n12716_));
  OAI21_X1   g09691(.A1(new_n12709_), .A2(new_n12701_), .B(new_n12716_), .ZN(new_n12717_));
  OAI21_X1   g09692(.A1(new_n12689_), .A2(new_n12717_), .B(new_n3225_), .ZN(new_n12718_));
  NAND2_X1   g09693(.A1(new_n12718_), .A2(new_n8104_), .ZN(new_n12719_));
  NAND2_X1   g09694(.A1(new_n12719_), .A2(pi0138), .ZN(new_n12720_));
  NOR2_X1    g09695(.A1(new_n9783_), .A2(pi0118), .ZN(new_n12721_));
  NAND2_X1   g09696(.A1(new_n12721_), .A2(new_n7955_), .ZN(new_n12722_));
  INV_X1     g09697(.I(new_n12722_), .ZN(new_n12723_));
  NAND2_X1   g09698(.A1(new_n12723_), .A2(pi0138), .ZN(new_n12724_));
  XOR2_X1    g09699(.A1(new_n12720_), .A2(new_n12724_), .Z(new_n12725_));
  NAND2_X1   g09700(.A1(new_n12719_), .A2(new_n12723_), .ZN(new_n12726_));
  OAI21_X1   g09701(.A1(pi0195), .A2(pi0196), .B(new_n7954_), .ZN(new_n12727_));
  NOR2_X1    g09702(.A1(new_n12722_), .A2(new_n12727_), .ZN(new_n12728_));
  XNOR2_X1   g09703(.A1(new_n12726_), .A2(new_n12728_), .ZN(new_n12729_));
  OAI21_X1   g09704(.A1(new_n12729_), .A2(new_n12725_), .B(new_n12674_), .ZN(po0295));
  NOR2_X1    g09705(.A1(pi0169), .A2(pi0299), .ZN(new_n12731_));
  OAI21_X1   g09706(.A1(new_n6448_), .A2(new_n12731_), .B(pi0232), .ZN(new_n12732_));
  INV_X1     g09707(.I(new_n12732_), .ZN(new_n12733_));
  NAND2_X1   g09708(.A1(new_n9281_), .A2(pi0191), .ZN(new_n12734_));
  NAND2_X1   g09709(.A1(pi0191), .A2(pi0299), .ZN(new_n12735_));
  XOR2_X1    g09710(.A1(new_n12734_), .A2(new_n12735_), .Z(new_n12736_));
  NOR4_X1    g09711(.A1(new_n9283_), .A2(new_n5551_), .A3(new_n7451_), .A4(new_n12664_), .ZN(new_n12737_));
  NAND2_X1   g09712(.A1(new_n12737_), .A2(new_n12736_), .ZN(new_n12738_));
  NAND2_X1   g09713(.A1(new_n12738_), .A2(new_n12733_), .ZN(new_n12739_));
  NAND3_X1   g09714(.A1(new_n12737_), .A2(new_n12736_), .A3(new_n12732_), .ZN(new_n12740_));
  NAND3_X1   g09715(.A1(new_n12739_), .A2(new_n8346_), .A3(new_n12740_), .ZN(new_n12741_));
  XNOR2_X1   g09716(.A1(new_n12741_), .A2(new_n9285_), .ZN(new_n12742_));
  NOR3_X1    g09717(.A1(new_n12742_), .A2(new_n12209_), .A3(new_n12673_), .ZN(new_n12743_));
  INV_X1     g09718(.I(new_n12712_), .ZN(new_n12744_));
  INV_X1     g09719(.I(new_n12679_), .ZN(new_n12745_));
  NOR2_X1    g09720(.A1(new_n12187_), .A2(new_n3098_), .ZN(new_n12746_));
  AOI21_X1   g09721(.A1(new_n7855_), .A2(new_n12746_), .B(pi0169), .ZN(new_n12747_));
  OAI21_X1   g09722(.A1(new_n12745_), .A2(new_n12747_), .B(new_n5551_), .ZN(new_n12748_));
  INV_X1     g09723(.I(new_n12688_), .ZN(new_n12749_));
  NOR3_X1    g09724(.A1(new_n12686_), .A2(new_n12167_), .A3(new_n12749_), .ZN(new_n12750_));
  AOI21_X1   g09725(.A1(new_n12750_), .A2(new_n12748_), .B(pi0191), .ZN(new_n12751_));
  INV_X1     g09726(.I(new_n12700_), .ZN(new_n12752_));
  INV_X1     g09727(.I(new_n12702_), .ZN(new_n12753_));
  NAND2_X1   g09728(.A1(new_n12753_), .A2(pi0191), .ZN(new_n12754_));
  NAND2_X1   g09729(.A1(new_n12695_), .A2(new_n12167_), .ZN(new_n12755_));
  AOI21_X1   g09730(.A1(new_n12755_), .A2(new_n12754_), .B(new_n5551_), .ZN(new_n12756_));
  AOI21_X1   g09731(.A1(new_n12704_), .A2(new_n7439_), .B(new_n7613_), .ZN(new_n12757_));
  NOR2_X1    g09732(.A1(new_n12757_), .A2(new_n4474_), .ZN(new_n12758_));
  OAI21_X1   g09733(.A1(new_n12756_), .A2(new_n7605_), .B(new_n12758_), .ZN(new_n12759_));
  AOI21_X1   g09734(.A1(new_n12759_), .A2(new_n3417_), .B(new_n12752_), .ZN(new_n12760_));
  NOR2_X1    g09735(.A1(new_n12714_), .A2(new_n3455_), .ZN(new_n12761_));
  OAI21_X1   g09736(.A1(new_n12710_), .A2(new_n3258_), .B(new_n3303_), .ZN(new_n12762_));
  OAI21_X1   g09737(.A1(new_n12760_), .A2(new_n12761_), .B(new_n12762_), .ZN(new_n12763_));
  OR2_X2     g09738(.A1(new_n12678_), .A2(new_n12763_), .Z(new_n12764_));
  OAI22_X1   g09739(.A1(new_n12764_), .A2(new_n12751_), .B1(new_n3226_), .B2(new_n10754_), .ZN(new_n12765_));
  NAND2_X1   g09740(.A1(new_n12765_), .A2(new_n12744_), .ZN(new_n12766_));
  NAND2_X1   g09741(.A1(new_n12766_), .A2(pi0139), .ZN(new_n12767_));
  NAND2_X1   g09742(.A1(new_n12721_), .A2(pi0139), .ZN(new_n12768_));
  XOR2_X1    g09743(.A1(new_n12767_), .A2(new_n12768_), .Z(new_n12769_));
  NAND2_X1   g09744(.A1(new_n12766_), .A2(new_n12721_), .ZN(new_n12770_));
  NAND3_X1   g09745(.A1(new_n7955_), .A2(new_n7956_), .A3(new_n7957_), .ZN(new_n12771_));
  NAND3_X1   g09746(.A1(new_n12721_), .A2(pi0138), .A3(new_n12771_), .ZN(new_n12772_));
  XOR2_X1    g09747(.A1(new_n12770_), .A2(new_n12772_), .Z(new_n12773_));
  OAI21_X1   g09748(.A1(new_n12769_), .A2(new_n12773_), .B(new_n12743_), .ZN(po0296));
  INV_X1     g09749(.I(pi0790), .ZN(new_n12775_));
  INV_X1     g09750(.I(pi0787), .ZN(new_n12776_));
  INV_X1     g09751(.I(pi0792), .ZN(new_n12777_));
  NOR2_X1    g09752(.A1(new_n5407_), .A2(pi0287), .ZN(new_n12778_));
  INV_X1     g09753(.I(new_n12778_), .ZN(new_n12779_));
  NOR2_X1    g09754(.A1(new_n3145_), .A2(new_n12779_), .ZN(new_n12780_));
  NAND3_X1   g09755(.A1(new_n12780_), .A2(pi0120), .A3(new_n9992_), .ZN(new_n12781_));
  NAND2_X1   g09756(.A1(new_n3160_), .A2(new_n12778_), .ZN(new_n12782_));
  NAND3_X1   g09757(.A1(new_n12782_), .A2(new_n10925_), .A3(new_n9992_), .ZN(new_n12783_));
  AOI21_X1   g09758(.A1(new_n12783_), .A2(new_n12781_), .B(new_n3145_), .ZN(new_n12784_));
  NOR2_X1    g09759(.A1(new_n10925_), .A2(new_n2726_), .ZN(new_n12785_));
  OAI21_X1   g09760(.A1(new_n3160_), .A2(new_n12785_), .B(new_n9992_), .ZN(new_n12786_));
  OAI21_X1   g09761(.A1(new_n12786_), .A2(new_n10925_), .B(new_n2984_), .ZN(new_n12787_));
  NOR3_X1    g09762(.A1(new_n8325_), .A2(new_n5401_), .A3(new_n3143_), .ZN(new_n12788_));
  NAND3_X1   g09763(.A1(new_n2711_), .A2(pi1092), .A3(new_n12788_), .ZN(new_n12789_));
  AOI21_X1   g09764(.A1(new_n12789_), .A2(new_n2722_), .B(new_n5683_), .ZN(new_n12790_));
  NOR2_X1    g09765(.A1(pi0287), .A2(pi0824), .ZN(new_n12791_));
  AOI21_X1   g09766(.A1(new_n3145_), .A2(new_n12791_), .B(new_n5408_), .ZN(new_n12792_));
  NOR2_X1    g09767(.A1(new_n12790_), .A2(new_n12792_), .ZN(new_n12793_));
  NOR2_X1    g09768(.A1(new_n3145_), .A2(new_n2723_), .ZN(new_n12794_));
  NOR2_X1    g09769(.A1(new_n12794_), .A2(new_n10925_), .ZN(new_n12795_));
  INV_X1     g09770(.I(new_n12795_), .ZN(new_n12796_));
  INV_X1     g09771(.I(new_n12785_), .ZN(new_n12797_));
  NOR2_X1    g09772(.A1(new_n2983_), .A2(new_n2723_), .ZN(new_n12798_));
  INV_X1     g09773(.I(new_n12798_), .ZN(new_n12799_));
  OAI21_X1   g09774(.A1(new_n12782_), .A2(new_n12799_), .B(new_n12797_), .ZN(new_n12800_));
  NAND3_X1   g09775(.A1(new_n2495_), .A2(new_n12788_), .A3(new_n2709_), .ZN(new_n12801_));
  NOR3_X1    g09776(.A1(new_n3160_), .A2(pi0287), .A3(pi0824), .ZN(new_n12802_));
  OAI21_X1   g09777(.A1(new_n6431_), .A2(pi1092), .B(pi0829), .ZN(new_n12803_));
  OAI22_X1   g09778(.A1(new_n12802_), .A2(new_n5408_), .B1(new_n12801_), .B2(new_n12803_), .ZN(new_n12804_));
  NAND3_X1   g09779(.A1(new_n12790_), .A2(new_n12800_), .A3(new_n12804_), .ZN(new_n12805_));
  AOI22_X1   g09780(.A1(new_n12805_), .A2(new_n12796_), .B1(new_n12793_), .B2(new_n12787_), .ZN(new_n12806_));
  NOR3_X1    g09781(.A1(new_n12782_), .A2(new_n10925_), .A3(new_n2723_), .ZN(new_n12807_));
  NOR3_X1    g09782(.A1(new_n12780_), .A2(pi0120), .A3(new_n2723_), .ZN(new_n12808_));
  OAI21_X1   g09783(.A1(new_n12807_), .A2(new_n12808_), .B(new_n3160_), .ZN(new_n12809_));
  OAI21_X1   g09784(.A1(new_n12801_), .A2(new_n2979_), .B(new_n2722_), .ZN(new_n12810_));
  NAND2_X1   g09785(.A1(new_n12810_), .A2(pi0824), .ZN(new_n12811_));
  INV_X1     g09786(.I(new_n12792_), .ZN(new_n12812_));
  NAND3_X1   g09787(.A1(new_n12811_), .A2(new_n12787_), .A3(new_n12812_), .ZN(new_n12813_));
  AOI21_X1   g09788(.A1(new_n12780_), .A2(new_n12798_), .B(new_n12785_), .ZN(new_n12814_));
  NOR2_X1    g09789(.A1(new_n12801_), .A2(new_n12803_), .ZN(new_n12815_));
  NOR2_X1    g09790(.A1(new_n12815_), .A2(new_n12792_), .ZN(new_n12816_));
  NOR3_X1    g09791(.A1(new_n12811_), .A2(new_n12816_), .A3(new_n12814_), .ZN(new_n12817_));
  OAI21_X1   g09792(.A1(new_n12795_), .A2(new_n12817_), .B(new_n12813_), .ZN(new_n12818_));
  NOR4_X1    g09793(.A1(new_n12818_), .A2(new_n5386_), .A3(new_n5796_), .A4(new_n12809_), .ZN(new_n12819_));
  NOR4_X1    g09794(.A1(new_n12806_), .A2(new_n5386_), .A3(new_n5796_), .A4(new_n12784_), .ZN(new_n12820_));
  NOR2_X1    g09795(.A1(new_n12820_), .A2(new_n12819_), .ZN(new_n12821_));
  NAND2_X1   g09796(.A1(new_n5635_), .A2(pi0681), .ZN(new_n12822_));
  AOI21_X1   g09797(.A1(new_n12821_), .A2(new_n5635_), .B(new_n12822_), .ZN(new_n12823_));
  NAND4_X1   g09798(.A1(new_n12806_), .A2(new_n5373_), .A3(new_n5383_), .A4(new_n12784_), .ZN(new_n12824_));
  NAND4_X1   g09799(.A1(new_n12818_), .A2(new_n5373_), .A3(new_n5383_), .A4(new_n12809_), .ZN(new_n12825_));
  NAND2_X1   g09800(.A1(new_n12824_), .A2(new_n12825_), .ZN(new_n12826_));
  NOR3_X1    g09801(.A1(new_n12826_), .A2(pi0681), .A3(new_n5377_), .ZN(new_n12827_));
  OAI21_X1   g09802(.A1(new_n12823_), .A2(new_n12827_), .B(new_n12806_), .ZN(new_n12828_));
  NOR2_X1    g09803(.A1(new_n12826_), .A2(new_n5632_), .ZN(new_n12829_));
  INV_X1     g09804(.I(new_n12829_), .ZN(new_n12830_));
  NAND3_X1   g09805(.A1(new_n12828_), .A2(new_n5453_), .A3(new_n12830_), .ZN(new_n12831_));
  NOR2_X1    g09806(.A1(new_n3313_), .A2(new_n3111_), .ZN(new_n12832_));
  INV_X1     g09807(.I(new_n12832_), .ZN(new_n12833_));
  AOI21_X1   g09808(.A1(new_n12831_), .A2(new_n3312_), .B(new_n12833_), .ZN(new_n12834_));
  NAND3_X1   g09809(.A1(new_n12826_), .A2(pi0681), .A3(new_n5635_), .ZN(new_n12835_));
  NAND3_X1   g09810(.A1(new_n12821_), .A2(new_n5632_), .A3(new_n5635_), .ZN(new_n12836_));
  AOI21_X1   g09811(.A1(new_n12836_), .A2(new_n12835_), .B(new_n12818_), .ZN(new_n12837_));
  NOR3_X1    g09812(.A1(new_n12837_), .A2(new_n5452_), .A3(new_n12829_), .ZN(new_n12838_));
  NOR3_X1    g09813(.A1(new_n12838_), .A2(pi0215), .A3(new_n3313_), .ZN(new_n12839_));
  OAI21_X1   g09814(.A1(new_n12839_), .A2(new_n12834_), .B(new_n12784_), .ZN(new_n12840_));
  INV_X1     g09815(.I(pi0616), .ZN(new_n12841_));
  NOR2_X1    g09816(.A1(pi0661), .A2(pi0681), .ZN(new_n12842_));
  INV_X1     g09817(.I(new_n12842_), .ZN(new_n12843_));
  NOR2_X1    g09818(.A1(new_n12843_), .A2(pi0662), .ZN(new_n12844_));
  INV_X1     g09819(.I(new_n12844_), .ZN(new_n12845_));
  NAND2_X1   g09820(.A1(new_n12784_), .A2(new_n12845_), .ZN(new_n12846_));
  NOR2_X1    g09821(.A1(new_n12846_), .A2(new_n12841_), .ZN(new_n12847_));
  NAND2_X1   g09822(.A1(new_n12784_), .A2(pi0680), .ZN(new_n12848_));
  NOR2_X1    g09823(.A1(new_n12844_), .A2(pi0616), .ZN(new_n12849_));
  NOR2_X1    g09824(.A1(new_n12848_), .A2(new_n12849_), .ZN(new_n12850_));
  NOR2_X1    g09825(.A1(new_n12809_), .A2(new_n5386_), .ZN(new_n12851_));
  INV_X1     g09826(.I(new_n12851_), .ZN(new_n12852_));
  NOR3_X1    g09827(.A1(new_n3145_), .A2(new_n10925_), .A3(new_n2723_), .ZN(new_n12853_));
  OAI21_X1   g09828(.A1(new_n12853_), .A2(new_n11073_), .B(new_n5409_), .ZN(new_n12854_));
  INV_X1     g09829(.I(new_n12854_), .ZN(new_n12855_));
  OAI21_X1   g09830(.A1(new_n12782_), .A2(new_n2723_), .B(new_n10925_), .ZN(new_n12856_));
  AOI21_X1   g09831(.A1(new_n3145_), .A2(new_n12797_), .B(new_n2723_), .ZN(new_n12857_));
  NOR2_X1    g09832(.A1(pi0120), .A2(pi0824), .ZN(new_n12858_));
  INV_X1     g09833(.I(new_n12858_), .ZN(new_n12859_));
  OAI21_X1   g09834(.A1(new_n12857_), .A2(new_n12859_), .B(new_n5409_), .ZN(new_n12860_));
  OAI21_X1   g09835(.A1(new_n12860_), .A2(new_n12856_), .B(new_n2726_), .ZN(new_n12861_));
  NAND2_X1   g09836(.A1(new_n12861_), .A2(new_n12855_), .ZN(new_n12862_));
  NAND2_X1   g09837(.A1(new_n12862_), .A2(new_n5386_), .ZN(new_n12863_));
  NAND3_X1   g09838(.A1(new_n12863_), .A2(new_n12852_), .A3(pi0680), .ZN(new_n12864_));
  AOI21_X1   g09839(.A1(new_n12864_), .A2(new_n12850_), .B(new_n12847_), .ZN(new_n12865_));
  NOR2_X1    g09840(.A1(new_n12865_), .A2(new_n5632_), .ZN(new_n12866_));
  INV_X1     g09841(.I(new_n12866_), .ZN(new_n12867_));
  INV_X1     g09842(.I(pi0614), .ZN(new_n12868_));
  NOR2_X1    g09843(.A1(new_n12868_), .A2(new_n12841_), .ZN(new_n12869_));
  INV_X1     g09844(.I(new_n12869_), .ZN(new_n12870_));
  AOI21_X1   g09845(.A1(new_n12780_), .A2(new_n9992_), .B(pi0120), .ZN(new_n12871_));
  AOI21_X1   g09846(.A1(new_n12786_), .A2(new_n12858_), .B(new_n5410_), .ZN(new_n12872_));
  AOI21_X1   g09847(.A1(new_n12872_), .A2(new_n12871_), .B(pi1091), .ZN(new_n12873_));
  NOR2_X1    g09848(.A1(new_n5386_), .A2(new_n5380_), .ZN(new_n12874_));
  INV_X1     g09849(.I(new_n12874_), .ZN(new_n12875_));
  NOR4_X1    g09850(.A1(new_n12873_), .A2(new_n12809_), .A3(new_n12854_), .A4(new_n12875_), .ZN(new_n12876_));
  NAND2_X1   g09851(.A1(new_n12872_), .A2(new_n12871_), .ZN(new_n12877_));
  AOI21_X1   g09852(.A1(new_n12877_), .A2(new_n2726_), .B(new_n12854_), .ZN(new_n12878_));
  NOR3_X1    g09853(.A1(new_n12878_), .A2(new_n12784_), .A3(new_n12875_), .ZN(new_n12879_));
  NOR2_X1    g09854(.A1(new_n12879_), .A2(new_n12876_), .ZN(new_n12880_));
  AOI21_X1   g09855(.A1(new_n12880_), .A2(pi0614), .B(new_n12870_), .ZN(new_n12881_));
  NAND4_X1   g09856(.A1(new_n12861_), .A2(new_n12784_), .A3(new_n12855_), .A4(new_n12874_), .ZN(new_n12882_));
  NAND3_X1   g09857(.A1(new_n12862_), .A2(new_n12809_), .A3(new_n12874_), .ZN(new_n12883_));
  NAND2_X1   g09858(.A1(new_n12883_), .A2(new_n12882_), .ZN(new_n12884_));
  NOR3_X1    g09859(.A1(new_n12884_), .A2(new_n12868_), .A3(pi0616), .ZN(new_n12885_));
  OAI21_X1   g09860(.A1(new_n12881_), .A2(new_n12885_), .B(new_n12784_), .ZN(new_n12886_));
  INV_X1     g09861(.I(new_n12849_), .ZN(new_n12887_));
  NOR3_X1    g09862(.A1(new_n12880_), .A2(new_n12868_), .A3(new_n12887_), .ZN(new_n12888_));
  NOR3_X1    g09863(.A1(new_n12884_), .A2(pi0614), .A3(new_n12887_), .ZN(new_n12889_));
  AOI21_X1   g09864(.A1(new_n5386_), .A2(new_n12862_), .B(new_n12851_), .ZN(new_n12890_));
  NOR3_X1    g09865(.A1(new_n12809_), .A2(pi0616), .A3(new_n12845_), .ZN(new_n12891_));
  INV_X1     g09866(.I(new_n12891_), .ZN(new_n12892_));
  AOI21_X1   g09867(.A1(new_n12890_), .A2(pi0680), .B(new_n12892_), .ZN(new_n12893_));
  OAI21_X1   g09868(.A1(new_n12888_), .A2(new_n12889_), .B(new_n12893_), .ZN(new_n12894_));
  AOI21_X1   g09869(.A1(new_n12894_), .A2(new_n12886_), .B(new_n5375_), .ZN(new_n12895_));
  NOR4_X1    g09870(.A1(new_n12862_), .A2(new_n12809_), .A3(new_n12870_), .A4(new_n12875_), .ZN(new_n12896_));
  NOR4_X1    g09871(.A1(new_n12879_), .A2(new_n12784_), .A3(new_n12870_), .A4(new_n12876_), .ZN(new_n12897_));
  NOR2_X1    g09872(.A1(new_n12897_), .A2(new_n12896_), .ZN(new_n12898_));
  NOR2_X1    g09873(.A1(new_n12898_), .A2(new_n5632_), .ZN(new_n12899_));
  NAND3_X1   g09874(.A1(new_n12895_), .A2(new_n12867_), .A3(new_n12899_), .ZN(new_n12900_));
  NAND3_X1   g09875(.A1(new_n12884_), .A2(pi0614), .A3(pi0616), .ZN(new_n12901_));
  NAND3_X1   g09876(.A1(new_n12880_), .A2(pi0614), .A3(new_n12841_), .ZN(new_n12902_));
  AOI21_X1   g09877(.A1(new_n12902_), .A2(new_n12901_), .B(new_n12809_), .ZN(new_n12903_));
  NAND3_X1   g09878(.A1(new_n12884_), .A2(pi0614), .A3(new_n12849_), .ZN(new_n12904_));
  NAND3_X1   g09879(.A1(new_n12880_), .A2(new_n12868_), .A3(new_n12849_), .ZN(new_n12905_));
  NAND2_X1   g09880(.A1(new_n12864_), .A2(new_n12891_), .ZN(new_n12906_));
  AOI21_X1   g09881(.A1(new_n12905_), .A2(new_n12904_), .B(new_n12906_), .ZN(new_n12907_));
  OAI21_X1   g09882(.A1(new_n12903_), .A2(new_n12907_), .B(pi0680), .ZN(new_n12908_));
  INV_X1     g09883(.I(new_n12899_), .ZN(new_n12909_));
  OAI21_X1   g09884(.A1(new_n12908_), .A2(new_n12909_), .B(new_n12866_), .ZN(new_n12910_));
  NAND2_X1   g09885(.A1(new_n12900_), .A2(new_n12910_), .ZN(new_n12911_));
  NOR2_X1    g09886(.A1(new_n5386_), .A2(new_n5634_), .ZN(new_n12912_));
  NAND2_X1   g09887(.A1(new_n12878_), .A2(new_n12912_), .ZN(new_n12913_));
  AOI21_X1   g09888(.A1(new_n12898_), .A2(new_n12912_), .B(new_n12913_), .ZN(new_n12914_));
  INV_X1     g09889(.I(new_n12896_), .ZN(new_n12915_));
  NAND4_X1   g09890(.A1(new_n12883_), .A2(new_n12809_), .A3(new_n12869_), .A4(new_n12882_), .ZN(new_n12916_));
  NAND4_X1   g09891(.A1(new_n12916_), .A2(new_n12862_), .A3(new_n12915_), .A4(new_n12912_), .ZN(new_n12917_));
  INV_X1     g09892(.I(new_n12917_), .ZN(new_n12918_));
  NOR2_X1    g09893(.A1(new_n12914_), .A2(new_n12918_), .ZN(new_n12919_));
  NOR2_X1    g09894(.A1(new_n5374_), .A2(new_n5632_), .ZN(new_n12920_));
  NAND2_X1   g09895(.A1(new_n12809_), .A2(new_n5386_), .ZN(new_n12921_));
  OAI21_X1   g09896(.A1(new_n5386_), .A2(new_n12862_), .B(new_n12921_), .ZN(new_n12922_));
  NOR2_X1    g09897(.A1(new_n12884_), .A2(pi0614), .ZN(new_n12923_));
  AOI21_X1   g09898(.A1(new_n12923_), .A2(new_n12841_), .B(new_n12922_), .ZN(new_n12924_));
  NAND2_X1   g09899(.A1(new_n12924_), .A2(new_n12920_), .ZN(new_n12925_));
  AOI21_X1   g09900(.A1(new_n12919_), .A2(new_n12920_), .B(new_n12925_), .ZN(new_n12926_));
  NAND2_X1   g09901(.A1(new_n12916_), .A2(new_n12915_), .ZN(new_n12927_));
  NAND3_X1   g09902(.A1(new_n12927_), .A2(new_n12878_), .A3(new_n12912_), .ZN(new_n12928_));
  NOR2_X1    g09903(.A1(new_n12784_), .A2(new_n5373_), .ZN(new_n12929_));
  AOI21_X1   g09904(.A1(new_n5373_), .A2(new_n12878_), .B(new_n12929_), .ZN(new_n12930_));
  NAND3_X1   g09905(.A1(new_n12880_), .A2(new_n12868_), .A3(new_n12841_), .ZN(new_n12931_));
  NAND2_X1   g09906(.A1(new_n12931_), .A2(new_n12930_), .ZN(new_n12932_));
  NAND4_X1   g09907(.A1(new_n12928_), .A2(new_n12932_), .A3(new_n12917_), .A4(new_n12920_), .ZN(new_n12933_));
  INV_X1     g09908(.I(new_n12933_), .ZN(new_n12934_));
  NOR2_X1    g09909(.A1(new_n12926_), .A2(new_n12934_), .ZN(new_n12935_));
  AOI21_X1   g09910(.A1(new_n12935_), .A2(new_n5452_), .B(new_n5455_), .ZN(new_n12936_));
  NAND2_X1   g09911(.A1(new_n12928_), .A2(new_n12917_), .ZN(new_n12937_));
  NAND3_X1   g09912(.A1(new_n12937_), .A2(new_n12920_), .A3(new_n12924_), .ZN(new_n12938_));
  NAND4_X1   g09913(.A1(new_n12938_), .A2(new_n5452_), .A3(new_n5455_), .A4(new_n12933_), .ZN(new_n12939_));
  INV_X1     g09914(.I(new_n12939_), .ZN(new_n12940_));
  OAI21_X1   g09915(.A1(new_n12936_), .A2(new_n12940_), .B(new_n12911_), .ZN(new_n12941_));
  NOR2_X1    g09916(.A1(new_n12935_), .A2(new_n5452_), .ZN(new_n12942_));
  NOR2_X1    g09917(.A1(new_n12942_), .A2(new_n3855_), .ZN(new_n12943_));
  NAND2_X1   g09918(.A1(new_n12941_), .A2(new_n12943_), .ZN(new_n12944_));
  AOI21_X1   g09919(.A1(new_n12818_), .A2(new_n5386_), .B(new_n12851_), .ZN(new_n12945_));
  NOR2_X1    g09920(.A1(new_n5794_), .A2(new_n5379_), .ZN(new_n12946_));
  INV_X1     g09921(.I(new_n12946_), .ZN(new_n12947_));
  NOR3_X1    g09922(.A1(new_n12945_), .A2(new_n12809_), .A3(new_n12947_), .ZN(new_n12948_));
  OAI21_X1   g09923(.A1(new_n12806_), .A2(new_n5373_), .B(new_n12852_), .ZN(new_n12949_));
  NOR3_X1    g09924(.A1(new_n12949_), .A2(new_n12784_), .A3(new_n12947_), .ZN(new_n12950_));
  NOR2_X1    g09925(.A1(new_n12950_), .A2(new_n12948_), .ZN(new_n12951_));
  NOR4_X1    g09926(.A1(new_n12809_), .A2(pi0614), .A3(new_n12841_), .A4(new_n5636_), .ZN(new_n12952_));
  AOI21_X1   g09927(.A1(new_n12949_), .A2(new_n12952_), .B(pi0616), .ZN(new_n12953_));
  OAI21_X1   g09928(.A1(new_n12951_), .A2(new_n12953_), .B(pi0681), .ZN(new_n12954_));
  NOR4_X1    g09929(.A1(new_n12945_), .A2(new_n12809_), .A3(new_n12870_), .A4(new_n12947_), .ZN(new_n12955_));
  INV_X1     g09930(.I(new_n12955_), .ZN(new_n12956_));
  NAND3_X1   g09931(.A1(new_n12949_), .A2(new_n12784_), .A3(new_n12946_), .ZN(new_n12957_));
  NAND3_X1   g09932(.A1(new_n12945_), .A2(new_n12809_), .A3(new_n12946_), .ZN(new_n12958_));
  NAND4_X1   g09933(.A1(new_n12957_), .A2(new_n12958_), .A3(new_n12809_), .A4(new_n12869_), .ZN(new_n12959_));
  NAND2_X1   g09934(.A1(new_n12959_), .A2(new_n12956_), .ZN(new_n12960_));
  NAND3_X1   g09935(.A1(new_n12784_), .A2(pi0614), .A3(new_n12845_), .ZN(new_n12961_));
  NAND2_X1   g09936(.A1(new_n12845_), .A2(new_n12868_), .ZN(new_n12962_));
  NAND4_X1   g09937(.A1(new_n12949_), .A2(pi0680), .A3(new_n12784_), .A4(new_n12962_), .ZN(new_n12963_));
  NAND3_X1   g09938(.A1(new_n12963_), .A2(pi0681), .A3(new_n12961_), .ZN(new_n12964_));
  INV_X1     g09939(.I(new_n12964_), .ZN(new_n12965_));
  NAND3_X1   g09940(.A1(new_n12960_), .A2(new_n12954_), .A3(new_n12965_), .ZN(new_n12966_));
  NAND2_X1   g09941(.A1(new_n12957_), .A2(new_n12958_), .ZN(new_n12967_));
  INV_X1     g09942(.I(new_n12953_), .ZN(new_n12968_));
  AOI21_X1   g09943(.A1(new_n12967_), .A2(new_n12968_), .B(new_n5632_), .ZN(new_n12969_));
  NOR4_X1    g09944(.A1(new_n12950_), .A2(new_n12948_), .A3(new_n12784_), .A4(new_n12870_), .ZN(new_n12970_));
  NOR2_X1    g09945(.A1(new_n12970_), .A2(new_n12955_), .ZN(new_n12971_));
  OAI21_X1   g09946(.A1(new_n12971_), .A2(new_n12964_), .B(new_n12969_), .ZN(new_n12972_));
  NAND2_X1   g09947(.A1(new_n12972_), .A2(new_n12966_), .ZN(new_n12973_));
  NOR2_X1    g09948(.A1(new_n12837_), .A2(new_n12829_), .ZN(new_n12974_));
  AOI21_X1   g09949(.A1(new_n3313_), .A2(new_n5453_), .B(new_n5451_), .ZN(new_n12975_));
  NAND2_X1   g09950(.A1(new_n12973_), .A2(new_n12975_), .ZN(new_n12976_));
  AOI21_X1   g09951(.A1(new_n12944_), .A2(new_n12840_), .B(new_n12976_), .ZN(new_n12977_));
  NOR3_X1    g09952(.A1(new_n12971_), .A2(new_n12969_), .A3(new_n12964_), .ZN(new_n12978_));
  AOI21_X1   g09953(.A1(new_n12960_), .A2(new_n12965_), .B(new_n12954_), .ZN(new_n12979_));
  NOR2_X1    g09954(.A1(new_n12979_), .A2(new_n12978_), .ZN(new_n12980_));
  NOR2_X1    g09955(.A1(new_n5397_), .A2(new_n3092_), .ZN(new_n12981_));
  INV_X1     g09956(.I(new_n12981_), .ZN(new_n12982_));
  AOI21_X1   g09957(.A1(new_n12980_), .A2(new_n5398_), .B(new_n12982_), .ZN(new_n12983_));
  NAND4_X1   g09958(.A1(new_n12972_), .A2(new_n12966_), .A3(new_n3092_), .A4(new_n5398_), .ZN(new_n12984_));
  INV_X1     g09959(.I(new_n12984_), .ZN(new_n12985_));
  OAI21_X1   g09960(.A1(new_n12983_), .A2(new_n12985_), .B(new_n12974_), .ZN(new_n12986_));
  NOR2_X1    g09961(.A1(new_n12809_), .A2(new_n3092_), .ZN(new_n12987_));
  NOR2_X1    g09962(.A1(new_n12987_), .A2(pi0223), .ZN(new_n12988_));
  AOI21_X1   g09963(.A1(new_n12938_), .A2(new_n12933_), .B(new_n5398_), .ZN(new_n12989_));
  AOI21_X1   g09964(.A1(new_n12900_), .A2(new_n12910_), .B(new_n5397_), .ZN(new_n12990_));
  NOR3_X1    g09965(.A1(new_n12990_), .A2(new_n3090_), .A3(new_n12989_), .ZN(new_n12991_));
  AOI21_X1   g09966(.A1(new_n12991_), .A2(pi0299), .B(new_n12988_), .ZN(new_n12992_));
  NOR2_X1    g09967(.A1(new_n8352_), .A2(new_n9231_), .ZN(new_n12993_));
  NOR2_X1    g09968(.A1(new_n12993_), .A2(pi0047), .ZN(new_n12994_));
  NOR2_X1    g09969(.A1(new_n2676_), .A2(new_n2798_), .ZN(new_n12995_));
  INV_X1     g09970(.I(new_n12995_), .ZN(new_n12996_));
  NOR2_X1    g09971(.A1(new_n12996_), .A2(new_n2692_), .ZN(new_n12997_));
  NOR2_X1    g09972(.A1(new_n8952_), .A2(new_n2672_), .ZN(new_n12998_));
  NOR2_X1    g09973(.A1(new_n9153_), .A2(pi0102), .ZN(new_n12999_));
  NAND2_X1   g09974(.A1(pi0098), .A2(pi0102), .ZN(new_n13000_));
  AOI21_X1   g09975(.A1(new_n2453_), .A2(new_n13000_), .B(new_n2492_), .ZN(new_n13001_));
  INV_X1     g09976(.I(new_n13001_), .ZN(new_n13002_));
  NOR2_X1    g09977(.A1(new_n12999_), .A2(new_n13002_), .ZN(new_n13003_));
  NAND2_X1   g09978(.A1(new_n13003_), .A2(pi0088), .ZN(new_n13004_));
  NOR2_X1    g09979(.A1(new_n13004_), .A2(new_n12998_), .ZN(new_n13005_));
  OAI21_X1   g09980(.A1(new_n12997_), .A2(new_n12994_), .B(new_n13005_), .ZN(new_n13006_));
  AOI21_X1   g09981(.A1(new_n3721_), .A2(new_n2499_), .B(new_n8367_), .ZN(new_n13007_));
  OAI21_X1   g09982(.A1(new_n13003_), .A2(pi0088), .B(new_n8952_), .ZN(new_n13008_));
  NOR3_X1    g09983(.A1(new_n2750_), .A2(new_n2486_), .A3(new_n3721_), .ZN(new_n13010_));
  NOR2_X1    g09984(.A1(new_n13007_), .A2(new_n13010_), .ZN(new_n13011_));
  AOI21_X1   g09985(.A1(new_n2981_), .A2(new_n2436_), .B(new_n2794_), .ZN(new_n13012_));
  NAND2_X1   g09986(.A1(new_n5557_), .A2(new_n13012_), .ZN(new_n13013_));
  AOI21_X1   g09987(.A1(new_n13013_), .A2(new_n5683_), .B(new_n2794_), .ZN(new_n13014_));
  INV_X1     g09988(.I(new_n13014_), .ZN(new_n13015_));
  NOR3_X1    g09989(.A1(new_n13015_), .A2(new_n13006_), .A3(new_n13011_), .ZN(new_n13016_));
  NOR3_X1    g09990(.A1(new_n2460_), .A2(new_n7277_), .A3(pi0088), .ZN(new_n13017_));
  NAND2_X1   g09991(.A1(new_n13003_), .A2(new_n13017_), .ZN(new_n13018_));
  NOR2_X1    g09992(.A1(new_n7668_), .A2(pi0040), .ZN(new_n13019_));
  AOI21_X1   g09993(.A1(new_n13018_), .A2(new_n13019_), .B(new_n7270_), .ZN(new_n13020_));
  NOR2_X1    g09994(.A1(new_n3142_), .A2(new_n3721_), .ZN(new_n13021_));
  INV_X1     g09995(.I(new_n13021_), .ZN(new_n13022_));
  NOR2_X1    g09996(.A1(new_n2502_), .A2(new_n3721_), .ZN(new_n13023_));
  NOR2_X1    g09997(.A1(new_n5556_), .A2(new_n2692_), .ZN(new_n13024_));
  AOI21_X1   g09998(.A1(new_n2499_), .A2(new_n2486_), .B(new_n2692_), .ZN(new_n13025_));
  AOI21_X1   g09999(.A1(new_n13024_), .A2(new_n13025_), .B(new_n12995_), .ZN(new_n13026_));
  NAND4_X1   g10000(.A1(new_n12999_), .A2(new_n2900_), .A3(new_n7267_), .A4(new_n13017_), .ZN(new_n13027_));
  OAI21_X1   g10001(.A1(new_n13027_), .A2(new_n13002_), .B(new_n2673_), .ZN(new_n13028_));
  NAND2_X1   g10002(.A1(new_n13028_), .A2(new_n12993_), .ZN(new_n13029_));
  NOR2_X1    g10003(.A1(new_n13029_), .A2(new_n13026_), .ZN(new_n13030_));
  AOI21_X1   g10004(.A1(pi0824), .A2(pi0950), .B(new_n2979_), .ZN(new_n13031_));
  NAND4_X1   g10005(.A1(new_n13030_), .A2(new_n13022_), .A3(new_n13023_), .A4(new_n13031_), .ZN(new_n13032_));
  OAI21_X1   g10006(.A1(new_n13020_), .A2(new_n8380_), .B(new_n3721_), .ZN(new_n13033_));
  OAI21_X1   g10007(.A1(new_n13029_), .A2(new_n13026_), .B(new_n13023_), .ZN(new_n13034_));
  NAND2_X1   g10008(.A1(new_n5683_), .A2(pi0829), .ZN(new_n13035_));
  AOI21_X1   g10009(.A1(new_n13013_), .A2(new_n13035_), .B(new_n2794_), .ZN(new_n13036_));
  NAND3_X1   g10010(.A1(new_n13034_), .A2(new_n13033_), .A3(new_n13036_), .ZN(new_n13037_));
  NAND3_X1   g10011(.A1(new_n13037_), .A2(new_n13032_), .A3(new_n2984_), .ZN(new_n13038_));
  NAND2_X1   g10012(.A1(new_n13038_), .A2(new_n13016_), .ZN(new_n13039_));
  INV_X1     g10013(.I(new_n13039_), .ZN(new_n13040_));
  NAND3_X1   g10014(.A1(new_n13030_), .A2(new_n13022_), .A3(new_n13023_), .ZN(new_n13041_));
  NOR2_X1    g10015(.A1(new_n10461_), .A2(new_n2979_), .ZN(po1106));
  INV_X1     g10016(.I(po1106), .ZN(new_n13043_));
  OAI21_X1   g10017(.A1(new_n13041_), .A2(new_n13043_), .B(new_n2730_), .ZN(new_n13044_));
  NAND2_X1   g10018(.A1(new_n13024_), .A2(new_n13025_), .ZN(new_n13045_));
  NAND2_X1   g10019(.A1(new_n13045_), .A2(new_n12996_), .ZN(new_n13046_));
  NAND4_X1   g10020(.A1(new_n13046_), .A2(new_n12993_), .A3(new_n13023_), .A4(new_n13028_), .ZN(new_n13047_));
  INV_X1     g10021(.I(new_n13031_), .ZN(new_n13048_));
  NOR3_X1    g10022(.A1(new_n13047_), .A2(new_n13021_), .A3(new_n13048_), .ZN(new_n13049_));
  OAI21_X1   g10023(.A1(new_n13049_), .A2(new_n13016_), .B(new_n6940_), .ZN(new_n13050_));
  OAI21_X1   g10024(.A1(new_n13050_), .A2(new_n13044_), .B(new_n2983_), .ZN(new_n13051_));
  AOI21_X1   g10025(.A1(new_n13040_), .A2(new_n13051_), .B(new_n3072_), .ZN(new_n13052_));
  NOR2_X1    g10026(.A1(new_n13047_), .A2(new_n13021_), .ZN(new_n13053_));
  AOI21_X1   g10027(.A1(new_n13053_), .A2(po1106), .B(new_n2729_), .ZN(new_n13054_));
  NOR2_X1    g10028(.A1(new_n7679_), .A2(pi0040), .ZN(new_n13055_));
  AOI21_X1   g10029(.A1(new_n13008_), .A2(new_n13055_), .B(new_n3721_), .ZN(new_n13056_));
  NOR2_X1    g10030(.A1(new_n8380_), .A2(new_n6403_), .ZN(new_n13057_));
  AOI21_X1   g10031(.A1(new_n13056_), .A2(new_n13057_), .B(new_n13007_), .ZN(new_n13058_));
  NOR3_X1    g10032(.A1(new_n13058_), .A2(new_n13006_), .A3(new_n2984_), .ZN(new_n13059_));
  OAI21_X1   g10033(.A1(new_n13059_), .A2(new_n13031_), .B(new_n13053_), .ZN(new_n13060_));
  AOI21_X1   g10034(.A1(new_n13060_), .A2(new_n2983_), .B(new_n13054_), .ZN(new_n13061_));
  NOR2_X1    g10035(.A1(new_n13060_), .A2(pi1091), .ZN(new_n13062_));
  NOR2_X1    g10036(.A1(new_n13061_), .A2(new_n13062_), .ZN(new_n13063_));
  NOR2_X1    g10037(.A1(new_n13063_), .A2(pi0198), .ZN(new_n13064_));
  NOR2_X1    g10038(.A1(new_n13064_), .A2(new_n13052_), .ZN(new_n13065_));
  NOR2_X1    g10039(.A1(new_n13065_), .A2(pi0299), .ZN(new_n13066_));
  AOI21_X1   g10040(.A1(new_n13040_), .A2(new_n13051_), .B(new_n2777_), .ZN(new_n13067_));
  NOR2_X1    g10041(.A1(new_n13063_), .A2(pi0210), .ZN(new_n13068_));
  OAI21_X1   g10042(.A1(new_n13068_), .A2(new_n13067_), .B(pi0299), .ZN(new_n13069_));
  INV_X1     g10043(.I(new_n13069_), .ZN(new_n13070_));
  OAI21_X1   g10044(.A1(new_n13066_), .A2(new_n13070_), .B(pi0039), .ZN(new_n13071_));
  NOR3_X1    g10045(.A1(new_n12992_), .A2(new_n12986_), .A3(new_n13071_), .ZN(new_n13072_));
  OAI21_X1   g10046(.A1(new_n12977_), .A2(new_n3183_), .B(new_n13072_), .ZN(new_n13073_));
  NOR3_X1    g10047(.A1(new_n12908_), .A2(new_n12866_), .A3(new_n12909_), .ZN(new_n13074_));
  AOI21_X1   g10048(.A1(new_n12895_), .A2(new_n12899_), .B(new_n12867_), .ZN(new_n13075_));
  NOR2_X1    g10049(.A1(new_n13075_), .A2(new_n13074_), .ZN(new_n13076_));
  INV_X1     g10050(.I(new_n5451_), .ZN(new_n13077_));
  NAND2_X1   g10051(.A1(new_n12938_), .A2(new_n12933_), .ZN(new_n13078_));
  NAND3_X1   g10052(.A1(new_n13078_), .A2(new_n13077_), .A3(new_n5452_), .ZN(new_n13079_));
  AOI21_X1   g10053(.A1(new_n13079_), .A2(new_n12939_), .B(new_n13076_), .ZN(new_n13080_));
  NAND2_X1   g10054(.A1(new_n13078_), .A2(new_n5453_), .ZN(new_n13081_));
  NAND2_X1   g10055(.A1(new_n13081_), .A2(new_n3695_), .ZN(new_n13082_));
  OAI21_X1   g10056(.A1(new_n13080_), .A2(new_n13082_), .B(new_n12840_), .ZN(new_n13083_));
  INV_X1     g10057(.I(new_n12976_), .ZN(new_n13084_));
  NAND2_X1   g10058(.A1(new_n13083_), .A2(new_n13084_), .ZN(new_n13085_));
  INV_X1     g10059(.I(new_n12974_), .ZN(new_n13086_));
  NAND3_X1   g10060(.A1(new_n12973_), .A2(new_n3091_), .A3(new_n5398_), .ZN(new_n13087_));
  AOI21_X1   g10061(.A1(new_n13087_), .A2(new_n12984_), .B(new_n13086_), .ZN(new_n13088_));
  INV_X1     g10062(.I(new_n12988_), .ZN(new_n13089_));
  OAI21_X1   g10063(.A1(new_n12926_), .A2(new_n12934_), .B(new_n5397_), .ZN(new_n13090_));
  OAI21_X1   g10064(.A1(new_n13075_), .A2(new_n13074_), .B(new_n5398_), .ZN(new_n13091_));
  NAND4_X1   g10065(.A1(new_n13091_), .A2(pi0223), .A3(new_n13090_), .A4(pi0299), .ZN(new_n13092_));
  NAND2_X1   g10066(.A1(new_n13092_), .A2(new_n13089_), .ZN(new_n13093_));
  INV_X1     g10067(.I(new_n13071_), .ZN(new_n13094_));
  NAND3_X1   g10068(.A1(new_n13093_), .A2(new_n13088_), .A3(new_n13094_), .ZN(new_n13095_));
  NAND3_X1   g10069(.A1(new_n13085_), .A2(new_n13095_), .A3(pi0039), .ZN(new_n13096_));
  NAND2_X1   g10070(.A1(new_n13073_), .A2(new_n13096_), .ZN(new_n13097_));
  NAND2_X1   g10071(.A1(new_n13097_), .A2(pi0761), .ZN(new_n13098_));
  INV_X1     g10072(.I(pi0761), .ZN(new_n13099_));
  NOR2_X1    g10073(.A1(new_n7971_), .A2(new_n13099_), .ZN(new_n13100_));
  INV_X1     g10074(.I(new_n13100_), .ZN(new_n13101_));
  NAND2_X1   g10075(.A1(pi0621), .A2(pi1091), .ZN(new_n13102_));
  NAND2_X1   g10076(.A1(new_n13102_), .A2(pi0603), .ZN(new_n13103_));
  NOR2_X1    g10077(.A1(new_n13103_), .A2(new_n2723_), .ZN(new_n13104_));
  INV_X1     g10078(.I(new_n13104_), .ZN(new_n13105_));
  NOR2_X1    g10079(.A1(new_n5504_), .A2(new_n13105_), .ZN(new_n13106_));
  INV_X1     g10080(.I(new_n13106_), .ZN(new_n13107_));
  NOR2_X1    g10081(.A1(new_n5504_), .A2(new_n2723_), .ZN(new_n13108_));
  INV_X1     g10082(.I(new_n13108_), .ZN(new_n13109_));
  OAI21_X1   g10083(.A1(new_n13107_), .A2(new_n13109_), .B(new_n13101_), .ZN(new_n13110_));
  AOI21_X1   g10084(.A1(new_n13110_), .A2(pi0038), .B(new_n3290_), .ZN(new_n13111_));
  OAI21_X1   g10085(.A1(new_n13098_), .A2(pi0038), .B(new_n13111_), .ZN(new_n13112_));
  NAND2_X1   g10086(.A1(new_n3290_), .A2(new_n7971_), .ZN(new_n13113_));
  NAND2_X1   g10087(.A1(new_n13112_), .A2(new_n13113_), .ZN(new_n13114_));
  INV_X1     g10088(.I(new_n13114_), .ZN(new_n13115_));
  NOR2_X1    g10089(.A1(new_n5794_), .A2(pi0665), .ZN(new_n13116_));
  INV_X1     g10090(.I(new_n13116_), .ZN(new_n13117_));
  AOI21_X1   g10091(.A1(new_n13038_), .A2(new_n13016_), .B(new_n2728_), .ZN(new_n13118_));
  NOR2_X1    g10092(.A1(new_n13118_), .A2(new_n13054_), .ZN(new_n13119_));
  INV_X1     g10093(.I(new_n13119_), .ZN(new_n13120_));
  AOI21_X1   g10094(.A1(new_n13061_), .A2(pi0621), .B(pi0198), .ZN(new_n13121_));
  AOI21_X1   g10095(.A1(new_n13121_), .A2(pi0198), .B(pi0621), .ZN(new_n13122_));
  NOR2_X1    g10096(.A1(new_n13122_), .A2(new_n13120_), .ZN(new_n13123_));
  INV_X1     g10097(.I(pi0665), .ZN(new_n13124_));
  AOI21_X1   g10098(.A1(new_n13061_), .A2(new_n13124_), .B(new_n13062_), .ZN(new_n13125_));
  OR2_X2     g10099(.A1(new_n13125_), .A2(pi0198), .Z(new_n13126_));
  AOI21_X1   g10100(.A1(pi0035), .A2(new_n12995_), .B(new_n12994_), .ZN(new_n13127_));
  NOR3_X1    g10101(.A1(new_n13127_), .A2(new_n12998_), .A3(new_n13004_), .ZN(new_n13128_));
  INV_X1     g10102(.I(new_n13011_), .ZN(new_n13129_));
  NAND3_X1   g10103(.A1(new_n13128_), .A2(new_n13129_), .A3(new_n13014_), .ZN(new_n13130_));
  AOI21_X1   g10104(.A1(new_n13130_), .A2(new_n13032_), .B(new_n6941_), .ZN(new_n13131_));
  AOI21_X1   g10105(.A1(new_n13119_), .A2(new_n13124_), .B(new_n13131_), .ZN(new_n13132_));
  OR2_X2     g10106(.A1(new_n13132_), .A2(new_n3072_), .Z(new_n13133_));
  NAND2_X1   g10107(.A1(new_n13133_), .A2(new_n13126_), .ZN(new_n13134_));
  NAND3_X1   g10108(.A1(new_n13134_), .A2(pi0603), .A3(new_n13123_), .ZN(new_n13135_));
  XOR2_X1    g10109(.A1(new_n13135_), .A2(new_n13117_), .Z(new_n13136_));
  NAND2_X1   g10110(.A1(new_n13136_), .A2(pi0680), .ZN(new_n13137_));
  INV_X1     g10111(.I(new_n13137_), .ZN(new_n13138_));
  NOR2_X1    g10112(.A1(new_n13125_), .A2(pi0210), .ZN(new_n13139_));
  NOR2_X1    g10113(.A1(new_n13132_), .A2(new_n2777_), .ZN(new_n13140_));
  NOR2_X1    g10114(.A1(new_n13140_), .A2(new_n13139_), .ZN(new_n13141_));
  INV_X1     g10115(.I(pi0621), .ZN(new_n13142_));
  NOR4_X1    g10116(.A1(new_n13118_), .A2(new_n2777_), .A3(new_n13142_), .A4(new_n13054_), .ZN(new_n13143_));
  NOR3_X1    g10117(.A1(new_n13119_), .A2(pi0210), .A3(new_n13142_), .ZN(new_n13144_));
  OAI21_X1   g10118(.A1(new_n13144_), .A2(new_n13143_), .B(new_n13061_), .ZN(new_n13145_));
  NOR3_X1    g10119(.A1(new_n13141_), .A2(new_n5794_), .A3(new_n13145_), .ZN(new_n13146_));
  NAND2_X1   g10120(.A1(new_n13146_), .A2(new_n13117_), .ZN(new_n13147_));
  INV_X1     g10121(.I(new_n13147_), .ZN(new_n13148_));
  NOR2_X1    g10122(.A1(new_n13146_), .A2(new_n13117_), .ZN(new_n13149_));
  NOR2_X1    g10123(.A1(new_n13148_), .A2(new_n13149_), .ZN(new_n13150_));
  NOR3_X1    g10124(.A1(new_n13150_), .A2(new_n3098_), .A3(new_n5375_), .ZN(new_n13151_));
  AOI21_X1   g10125(.A1(new_n13138_), .A2(new_n3098_), .B(new_n13151_), .ZN(new_n13152_));
  NOR3_X1    g10126(.A1(new_n13120_), .A2(new_n2777_), .A3(new_n13124_), .ZN(new_n13153_));
  NOR3_X1    g10127(.A1(new_n13119_), .A2(pi0210), .A3(new_n13124_), .ZN(new_n13154_));
  OAI21_X1   g10128(.A1(new_n13153_), .A2(new_n13154_), .B(new_n13061_), .ZN(new_n13155_));
  AOI21_X1   g10129(.A1(new_n5375_), .A2(new_n13069_), .B(new_n13155_), .ZN(new_n13156_));
  NOR3_X1    g10130(.A1(new_n13120_), .A2(new_n3072_), .A3(new_n13124_), .ZN(new_n13157_));
  NOR3_X1    g10131(.A1(new_n13119_), .A2(pi0198), .A3(new_n13124_), .ZN(new_n13158_));
  OAI21_X1   g10132(.A1(new_n13157_), .A2(new_n13158_), .B(new_n13061_), .ZN(new_n13159_));
  AOI21_X1   g10133(.A1(new_n13131_), .A2(new_n13054_), .B(new_n2728_), .ZN(new_n13160_));
  OAI21_X1   g10134(.A1(new_n13160_), .A2(new_n13039_), .B(pi0198), .ZN(new_n13161_));
  OAI21_X1   g10135(.A1(pi0198), .A2(new_n13063_), .B(new_n13161_), .ZN(new_n13162_));
  NAND2_X1   g10136(.A1(new_n13162_), .A2(pi0299), .ZN(new_n13163_));
  AOI21_X1   g10137(.A1(new_n13163_), .A2(new_n5375_), .B(new_n13159_), .ZN(new_n13164_));
  NOR2_X1    g10138(.A1(new_n13164_), .A2(new_n13156_), .ZN(new_n13165_));
  AOI21_X1   g10139(.A1(new_n13061_), .A2(new_n13142_), .B(new_n13062_), .ZN(new_n13166_));
  INV_X1     g10140(.I(new_n13166_), .ZN(new_n13167_));
  NOR2_X1    g10141(.A1(new_n13131_), .A2(new_n13142_), .ZN(new_n13168_));
  NAND2_X1   g10142(.A1(new_n13168_), .A2(pi0198), .ZN(new_n13169_));
  INV_X1     g10143(.I(new_n13169_), .ZN(new_n13170_));
  NAND3_X1   g10144(.A1(new_n13167_), .A2(new_n13161_), .A3(new_n13170_), .ZN(new_n13171_));
  OAI21_X1   g10145(.A1(new_n13166_), .A2(new_n13169_), .B(new_n13052_), .ZN(new_n13172_));
  NAND3_X1   g10146(.A1(new_n13171_), .A2(new_n13172_), .A3(pi0603), .ZN(new_n13173_));
  INV_X1     g10147(.I(new_n13173_), .ZN(new_n13174_));
  NOR2_X1    g10148(.A1(new_n13166_), .A2(pi0210), .ZN(new_n13175_));
  NOR2_X1    g10149(.A1(new_n13160_), .A2(new_n13039_), .ZN(new_n13176_));
  NOR3_X1    g10150(.A1(new_n13176_), .A2(new_n2777_), .A3(new_n13168_), .ZN(new_n13177_));
  OAI21_X1   g10151(.A1(new_n13177_), .A2(new_n13175_), .B(pi0603), .ZN(new_n13178_));
  NOR2_X1    g10152(.A1(new_n13178_), .A2(new_n3098_), .ZN(new_n13179_));
  AOI21_X1   g10153(.A1(new_n13174_), .A2(new_n3098_), .B(new_n13179_), .ZN(new_n13180_));
  NOR2_X1    g10154(.A1(new_n13180_), .A2(new_n5375_), .ZN(new_n13181_));
  OAI21_X1   g10155(.A1(new_n13181_), .A2(new_n13165_), .B(pi0761), .ZN(new_n13182_));
  XOR2_X1    g10156(.A1(new_n13182_), .A2(new_n13100_), .Z(new_n13183_));
  OAI21_X1   g10157(.A1(new_n13152_), .A2(new_n13183_), .B(new_n3211_), .ZN(new_n13184_));
  OAI21_X1   g10158(.A1(new_n13122_), .A2(new_n13120_), .B(new_n3098_), .ZN(new_n13185_));
  AOI21_X1   g10159(.A1(new_n13171_), .A2(new_n13172_), .B(new_n5794_), .ZN(new_n13186_));
  NAND2_X1   g10160(.A1(new_n13186_), .A2(new_n13185_), .ZN(new_n13187_));
  AOI21_X1   g10161(.A1(new_n5794_), .A2(new_n13069_), .B(new_n13145_), .ZN(new_n13188_));
  NAND3_X1   g10162(.A1(new_n13164_), .A2(new_n13156_), .A3(new_n13188_), .ZN(new_n13189_));
  NOR2_X1    g10163(.A1(new_n13189_), .A2(new_n13187_), .ZN(new_n13190_));
  INV_X1     g10164(.I(new_n13190_), .ZN(new_n13191_));
  INV_X1     g10165(.I(new_n13178_), .ZN(new_n13192_));
  NAND2_X1   g10166(.A1(new_n13192_), .A2(pi0299), .ZN(new_n13193_));
  OAI21_X1   g10167(.A1(pi0299), .A2(new_n13173_), .B(new_n13193_), .ZN(new_n13194_));
  NAND3_X1   g10168(.A1(new_n13134_), .A2(pi0299), .A3(pi0680), .ZN(new_n13195_));
  NAND4_X1   g10169(.A1(new_n13133_), .A2(new_n13126_), .A3(new_n3098_), .A4(pi0680), .ZN(new_n13196_));
  AOI21_X1   g10170(.A1(new_n13195_), .A2(new_n13196_), .B(new_n13141_), .ZN(new_n13197_));
  NOR2_X1    g10171(.A1(new_n13197_), .A2(new_n13194_), .ZN(new_n13198_));
  NAND3_X1   g10172(.A1(new_n13198_), .A2(pi0140), .A3(pi0761), .ZN(new_n13199_));
  INV_X1     g10173(.I(new_n13198_), .ZN(new_n13200_));
  NAND3_X1   g10174(.A1(new_n13200_), .A2(pi0140), .A3(new_n13099_), .ZN(new_n13201_));
  AOI21_X1   g10175(.A1(new_n13201_), .A2(new_n13199_), .B(new_n13191_), .ZN(new_n13202_));
  INV_X1     g10176(.I(new_n13103_), .ZN(new_n13203_));
  NAND2_X1   g10177(.A1(pi0665), .A2(pi1091), .ZN(new_n13204_));
  NAND2_X1   g10178(.A1(new_n13204_), .A2(pi0680), .ZN(new_n13205_));
  INV_X1     g10179(.I(new_n13205_), .ZN(new_n13206_));
  NOR2_X1    g10180(.A1(new_n13203_), .A2(new_n13206_), .ZN(new_n13207_));
  NAND2_X1   g10181(.A1(new_n12794_), .A2(new_n13207_), .ZN(new_n13208_));
  INV_X1     g10182(.I(new_n13208_), .ZN(new_n13209_));
  INV_X1     g10183(.I(new_n13204_), .ZN(new_n13210_));
  NOR2_X1    g10184(.A1(new_n13203_), .A2(new_n13210_), .ZN(new_n13211_));
  INV_X1     g10185(.I(new_n13211_), .ZN(new_n13212_));
  NOR2_X1    g10186(.A1(new_n13212_), .A2(new_n5375_), .ZN(new_n13213_));
  NOR2_X1    g10187(.A1(new_n13205_), .A2(new_n2723_), .ZN(new_n13218_));
  INV_X1     g10188(.I(new_n13218_), .ZN(new_n13219_));
  NOR2_X1    g10189(.A1(new_n13219_), .A2(new_n13203_), .ZN(new_n13220_));
  NOR2_X1    g10190(.A1(new_n13220_), .A2(new_n13104_), .ZN(new_n13221_));
  NAND2_X1   g10191(.A1(new_n13209_), .A2(pi0140), .ZN(new_n13222_));
  NAND2_X1   g10192(.A1(new_n13222_), .A2(pi0038), .ZN(new_n13223_));
  XOR2_X1    g10193(.A1(new_n13223_), .A2(new_n3262_), .Z(new_n13224_));
  INV_X1     g10194(.I(new_n13224_), .ZN(new_n13225_));
  INV_X1     g10195(.I(pi0738), .ZN(new_n13226_));
  NOR2_X1    g10196(.A1(new_n7971_), .A2(new_n13226_), .ZN(new_n13227_));
  AOI22_X1   g10197(.A1(new_n13184_), .A2(new_n13202_), .B1(new_n13225_), .B2(new_n13227_), .ZN(new_n13228_));
  NOR2_X1    g10198(.A1(new_n12817_), .A2(new_n12795_), .ZN(new_n13229_));
  INV_X1     g10199(.I(new_n13102_), .ZN(new_n13230_));
  NAND2_X1   g10200(.A1(new_n13229_), .A2(new_n13230_), .ZN(new_n13231_));
  NOR2_X1    g10201(.A1(new_n13231_), .A2(pi0665), .ZN(new_n13232_));
  INV_X1     g10202(.I(new_n13232_), .ZN(new_n13233_));
  NOR2_X1    g10203(.A1(new_n12844_), .A2(new_n5375_), .ZN(new_n13234_));
  NOR2_X1    g10204(.A1(new_n12795_), .A2(pi0665), .ZN(new_n13235_));
  NAND2_X1   g10205(.A1(new_n12813_), .A2(new_n13235_), .ZN(new_n13236_));
  NAND2_X1   g10206(.A1(new_n13236_), .A2(new_n12817_), .ZN(new_n13237_));
  NOR2_X1    g10207(.A1(new_n13237_), .A2(new_n5636_), .ZN(new_n13238_));
  NAND2_X1   g10208(.A1(new_n13238_), .A2(new_n13234_), .ZN(new_n13239_));
  AOI21_X1   g10209(.A1(new_n13239_), .A2(new_n5794_), .B(new_n13233_), .ZN(new_n13240_));
  INV_X1     g10210(.I(new_n13240_), .ZN(new_n13241_));
  AOI21_X1   g10211(.A1(new_n12813_), .A2(new_n13235_), .B(new_n12805_), .ZN(new_n13242_));
  NOR2_X1    g10212(.A1(new_n12809_), .A2(new_n5373_), .ZN(new_n13243_));
  OAI21_X1   g10213(.A1(new_n12813_), .A2(new_n5386_), .B(new_n12796_), .ZN(new_n13244_));
  AND2_X2    g10214(.A1(new_n13244_), .A2(new_n12817_), .Z(new_n13245_));
  NOR2_X1    g10215(.A1(new_n12809_), .A2(new_n13210_), .ZN(new_n13246_));
  AOI22_X1   g10216(.A1(new_n13245_), .A2(new_n13246_), .B1(new_n13242_), .B2(new_n13243_), .ZN(new_n13247_));
  NAND2_X1   g10217(.A1(new_n13232_), .A2(pi0603), .ZN(new_n13248_));
  OAI21_X1   g10218(.A1(new_n13247_), .A2(pi0603), .B(new_n13248_), .ZN(new_n13249_));
  NOR2_X1    g10219(.A1(pi0614), .A2(pi0642), .ZN(new_n13250_));
  INV_X1     g10220(.I(new_n13250_), .ZN(new_n13251_));
  NOR2_X1    g10221(.A1(new_n13251_), .A2(new_n12841_), .ZN(new_n13252_));
  NAND2_X1   g10222(.A1(new_n12805_), .A2(new_n12796_), .ZN(new_n13253_));
  NOR2_X1    g10223(.A1(new_n13253_), .A2(new_n13102_), .ZN(new_n13254_));
  NAND2_X1   g10224(.A1(new_n12784_), .A2(new_n5386_), .ZN(new_n13255_));
  OAI21_X1   g10225(.A1(new_n13255_), .A2(new_n13102_), .B(new_n5794_), .ZN(new_n13256_));
  NAND3_X1   g10226(.A1(new_n13254_), .A2(new_n5373_), .A3(new_n13256_), .ZN(new_n13257_));
  INV_X1     g10227(.I(new_n13246_), .ZN(new_n13258_));
  NAND2_X1   g10228(.A1(new_n13237_), .A2(new_n13258_), .ZN(new_n13259_));
  NAND2_X1   g10229(.A1(new_n13257_), .A2(new_n13259_), .ZN(new_n13260_));
  NAND2_X1   g10230(.A1(new_n13244_), .A2(new_n12817_), .ZN(new_n13261_));
  NAND2_X1   g10231(.A1(new_n13261_), .A2(new_n13255_), .ZN(new_n13262_));
  INV_X1     g10232(.I(new_n13262_), .ZN(new_n13263_));
  NAND3_X1   g10233(.A1(new_n13260_), .A2(new_n13263_), .A3(pi0603), .ZN(new_n13264_));
  INV_X1     g10234(.I(new_n13264_), .ZN(new_n13265_));
  NAND3_X1   g10235(.A1(new_n13265_), .A2(new_n13249_), .A3(new_n13252_), .ZN(new_n13266_));
  INV_X1     g10236(.I(new_n13249_), .ZN(new_n13267_));
  NAND3_X1   g10237(.A1(new_n13267_), .A2(new_n13252_), .A3(new_n13264_), .ZN(new_n13268_));
  NAND3_X1   g10238(.A1(new_n13268_), .A2(new_n13266_), .A3(new_n12845_), .ZN(new_n13269_));
  NAND2_X1   g10239(.A1(new_n12784_), .A2(new_n13230_), .ZN(new_n13270_));
  NAND3_X1   g10240(.A1(new_n13254_), .A2(pi0603), .A3(new_n5373_), .ZN(new_n13271_));
  NAND3_X1   g10241(.A1(new_n13231_), .A2(pi0603), .A3(new_n5386_), .ZN(new_n13272_));
  AOI21_X1   g10242(.A1(new_n13272_), .A2(new_n13271_), .B(new_n13270_), .ZN(new_n13273_));
  INV_X1     g10243(.I(new_n13273_), .ZN(new_n13274_));
  NOR2_X1    g10244(.A1(new_n12809_), .A2(new_n13203_), .ZN(new_n13275_));
  INV_X1     g10245(.I(new_n13275_), .ZN(new_n13276_));
  NOR2_X1    g10246(.A1(new_n13276_), .A2(new_n13210_), .ZN(new_n13277_));
  AOI21_X1   g10247(.A1(new_n13277_), .A2(new_n13251_), .B(pi0616), .ZN(new_n13278_));
  OAI21_X1   g10248(.A1(new_n13258_), .A2(pi0603), .B(new_n13117_), .ZN(new_n13279_));
  NOR3_X1    g10249(.A1(new_n13278_), .A2(new_n13250_), .A3(new_n13279_), .ZN(new_n13280_));
  NOR2_X1    g10250(.A1(new_n13274_), .A2(new_n13280_), .ZN(new_n13281_));
  NOR2_X1    g10251(.A1(new_n5386_), .A2(new_n5794_), .ZN(new_n13282_));
  INV_X1     g10252(.I(new_n13282_), .ZN(new_n13283_));
  NAND2_X1   g10253(.A1(new_n12818_), .A2(pi0603), .ZN(new_n13284_));
  XOR2_X1    g10254(.A1(new_n13284_), .A2(new_n13283_), .Z(new_n13285_));
  NAND2_X1   g10255(.A1(new_n13285_), .A2(new_n12784_), .ZN(new_n13286_));
  NOR2_X1    g10256(.A1(new_n13117_), .A2(new_n13102_), .ZN(new_n13287_));
  NOR2_X1    g10257(.A1(new_n5378_), .A2(new_n13287_), .ZN(new_n13288_));
  NOR2_X1    g10258(.A1(new_n12809_), .A2(new_n13204_), .ZN(new_n13289_));
  NAND2_X1   g10259(.A1(new_n13229_), .A2(new_n13210_), .ZN(new_n13290_));
  AOI21_X1   g10260(.A1(new_n13290_), .A2(new_n5373_), .B(new_n13283_), .ZN(new_n13291_));
  INV_X1     g10261(.I(new_n13290_), .ZN(new_n13292_));
  NOR3_X1    g10262(.A1(new_n13292_), .A2(pi0603), .A3(new_n5386_), .ZN(new_n13293_));
  OAI21_X1   g10263(.A1(new_n13293_), .A2(new_n13291_), .B(new_n13289_), .ZN(new_n13294_));
  AOI21_X1   g10264(.A1(new_n13286_), .A2(new_n13288_), .B(new_n13294_), .ZN(new_n13295_));
  INV_X1     g10265(.I(new_n13234_), .ZN(new_n13296_));
  INV_X1     g10266(.I(new_n13277_), .ZN(new_n13297_));
  AOI21_X1   g10267(.A1(new_n13297_), .A2(pi0616), .B(new_n13296_), .ZN(new_n13298_));
  AOI22_X1   g10268(.A1(new_n13295_), .A2(new_n13298_), .B1(new_n12949_), .B2(new_n13281_), .ZN(new_n13299_));
  NAND2_X1   g10269(.A1(new_n13299_), .A2(new_n5398_), .ZN(new_n13300_));
  INV_X1     g10270(.I(new_n13221_), .ZN(new_n13301_));
  AOI21_X1   g10271(.A1(new_n12987_), .A2(new_n13203_), .B(pi0223), .ZN(new_n13302_));
  NOR3_X1    g10272(.A1(new_n12809_), .A2(new_n3091_), .A3(new_n13301_), .ZN(new_n13303_));
  AOI22_X1   g10273(.A1(new_n13300_), .A2(new_n13303_), .B1(new_n13241_), .B2(new_n13269_), .ZN(new_n13304_));
  OAI21_X1   g10274(.A1(new_n13304_), .A2(new_n5397_), .B(pi0299), .ZN(new_n13305_));
  INV_X1     g10275(.I(new_n13299_), .ZN(new_n13306_));
  AOI21_X1   g10276(.A1(new_n13306_), .A2(new_n5454_), .B(new_n3312_), .ZN(new_n13307_));
  INV_X1     g10277(.I(new_n13307_), .ZN(new_n13308_));
  INV_X1     g10278(.I(new_n5456_), .ZN(new_n13309_));
  NOR2_X1    g10279(.A1(new_n13203_), .A2(new_n2723_), .ZN(new_n13310_));
  NAND3_X1   g10280(.A1(new_n13279_), .A2(new_n12930_), .A3(new_n13310_), .ZN(new_n13311_));
  INV_X1     g10281(.I(new_n13311_), .ZN(new_n13312_));
  NOR2_X1    g10282(.A1(new_n13312_), .A2(new_n12841_), .ZN(new_n13313_));
  NAND3_X1   g10283(.A1(new_n12855_), .A2(new_n12871_), .A3(new_n13230_), .ZN(new_n13314_));
  INV_X1     g10284(.I(new_n13314_), .ZN(new_n13315_));
  INV_X1     g10285(.I(new_n13270_), .ZN(new_n13316_));
  NAND3_X1   g10286(.A1(new_n13316_), .A2(pi0603), .A3(new_n5373_), .ZN(new_n13317_));
  NAND3_X1   g10287(.A1(new_n13270_), .A2(pi0603), .A3(new_n5386_), .ZN(new_n13318_));
  NAND2_X1   g10288(.A1(new_n13317_), .A2(new_n13318_), .ZN(new_n13319_));
  NAND2_X1   g10289(.A1(new_n13319_), .A2(new_n13315_), .ZN(new_n13320_));
  AOI21_X1   g10290(.A1(new_n13320_), .A2(new_n13279_), .B(pi0642), .ZN(new_n13321_));
  NOR2_X1    g10291(.A1(new_n13311_), .A2(new_n12841_), .ZN(new_n13322_));
  OAI21_X1   g10292(.A1(new_n13321_), .A2(new_n13322_), .B(pi0614), .ZN(new_n13323_));
  INV_X1     g10293(.I(new_n13213_), .ZN(new_n13324_));
  NOR2_X1    g10294(.A1(new_n13234_), .A2(new_n12845_), .ZN(new_n13325_));
  OAI21_X1   g10295(.A1(new_n12878_), .A2(new_n13324_), .B(new_n13325_), .ZN(new_n13326_));
  NAND2_X1   g10296(.A1(new_n13323_), .A2(new_n13326_), .ZN(new_n13327_));
  NAND2_X1   g10297(.A1(new_n13327_), .A2(new_n13313_), .ZN(new_n13328_));
  AOI21_X1   g10298(.A1(new_n13328_), .A2(pi0215), .B(new_n13309_), .ZN(new_n13329_));
  NAND2_X1   g10299(.A1(new_n13328_), .A2(pi0215), .ZN(new_n13330_));
  NOR2_X1    g10300(.A1(new_n13330_), .A2(new_n5456_), .ZN(new_n13331_));
  INV_X1     g10301(.I(new_n13279_), .ZN(new_n13332_));
  INV_X1     g10302(.I(new_n13298_), .ZN(new_n13333_));
  INV_X1     g10303(.I(new_n12890_), .ZN(new_n13334_));
  NAND3_X1   g10304(.A1(new_n13320_), .A2(new_n5378_), .A3(new_n13334_), .ZN(new_n13335_));
  NOR2_X1    g10305(.A1(new_n13251_), .A2(pi0616), .ZN(new_n13336_));
  NOR2_X1    g10306(.A1(new_n13276_), .A2(new_n13336_), .ZN(new_n13337_));
  OAI21_X1   g10307(.A1(new_n12784_), .A2(pi0603), .B(new_n13336_), .ZN(new_n13338_));
  AOI21_X1   g10308(.A1(new_n13319_), .A2(new_n13315_), .B(new_n13338_), .ZN(new_n13339_));
  NOR2_X1    g10309(.A1(new_n13339_), .A2(new_n13337_), .ZN(new_n13340_));
  OAI21_X1   g10310(.A1(new_n13340_), .A2(new_n13210_), .B(new_n12841_), .ZN(new_n13341_));
  OAI22_X1   g10311(.A1(new_n13341_), .A2(new_n13332_), .B1(new_n13333_), .B2(new_n13335_), .ZN(new_n13342_));
  NOR2_X1    g10312(.A1(new_n12809_), .A2(new_n3313_), .ZN(new_n13343_));
  NAND2_X1   g10313(.A1(new_n13343_), .A2(new_n13213_), .ZN(new_n13344_));
  AND3_X2    g10314(.A1(new_n13342_), .A2(new_n3111_), .A3(new_n13344_), .Z(new_n13345_));
  OAI21_X1   g10315(.A1(new_n13331_), .A2(new_n13329_), .B(new_n13345_), .ZN(new_n13346_));
  NAND2_X1   g10316(.A1(new_n13346_), .A2(new_n13308_), .ZN(new_n13347_));
  INV_X1     g10317(.I(new_n13328_), .ZN(new_n13348_));
  NAND3_X1   g10318(.A1(new_n13348_), .A2(pi0223), .A3(new_n5398_), .ZN(new_n13349_));
  NAND3_X1   g10319(.A1(new_n13328_), .A2(pi0223), .A3(new_n5397_), .ZN(new_n13350_));
  NAND2_X1   g10320(.A1(new_n13268_), .A2(new_n13266_), .ZN(new_n13351_));
  NAND2_X1   g10321(.A1(new_n13240_), .A2(new_n5454_), .ZN(new_n13352_));
  AOI21_X1   g10322(.A1(new_n13352_), .A2(new_n12845_), .B(new_n3098_), .ZN(new_n13353_));
  NAND3_X1   g10323(.A1(new_n13351_), .A2(new_n13342_), .A3(new_n13353_), .ZN(new_n13354_));
  AOI21_X1   g10324(.A1(new_n13349_), .A2(new_n13350_), .B(new_n13354_), .ZN(new_n13355_));
  NAND3_X1   g10325(.A1(new_n13347_), .A2(new_n13305_), .A3(new_n13355_), .ZN(new_n13356_));
  AOI21_X1   g10326(.A1(new_n13347_), .A2(new_n13355_), .B(new_n13305_), .ZN(new_n13357_));
  INV_X1     g10327(.I(new_n13357_), .ZN(new_n13358_));
  NAND2_X1   g10328(.A1(new_n13358_), .A2(new_n13356_), .ZN(new_n13359_));
  AOI21_X1   g10329(.A1(new_n13359_), .A2(pi0140), .B(new_n13099_), .ZN(new_n13360_));
  NOR2_X1    g10330(.A1(new_n13242_), .A2(new_n13246_), .ZN(new_n13361_));
  AOI21_X1   g10331(.A1(new_n12949_), .A2(new_n5378_), .B(new_n13361_), .ZN(new_n13362_));
  NOR2_X1    g10332(.A1(new_n12809_), .A2(new_n13103_), .ZN(new_n13363_));
  INV_X1     g10333(.I(new_n13363_), .ZN(new_n13364_));
  INV_X1     g10334(.I(new_n13336_), .ZN(new_n13365_));
  NOR3_X1    g10335(.A1(new_n12818_), .A2(new_n5386_), .A3(new_n13103_), .ZN(new_n13366_));
  NOR3_X1    g10336(.A1(new_n12806_), .A2(new_n5373_), .A3(new_n13103_), .ZN(new_n13367_));
  OAI21_X1   g10337(.A1(new_n13367_), .A2(new_n13366_), .B(new_n12784_), .ZN(new_n13368_));
  NOR3_X1    g10338(.A1(new_n13368_), .A2(new_n5375_), .A3(new_n13365_), .ZN(new_n13369_));
  NAND3_X1   g10339(.A1(new_n12806_), .A2(new_n5373_), .A3(new_n13203_), .ZN(new_n13370_));
  NAND3_X1   g10340(.A1(new_n12818_), .A2(new_n5386_), .A3(new_n13203_), .ZN(new_n13371_));
  AOI21_X1   g10341(.A1(new_n13370_), .A2(new_n13371_), .B(new_n12809_), .ZN(new_n13372_));
  NOR3_X1    g10342(.A1(new_n13372_), .A2(pi0680), .A3(new_n13365_), .ZN(new_n13373_));
  NOR2_X1    g10343(.A1(new_n13369_), .A2(new_n13373_), .ZN(new_n13374_));
  OAI22_X1   g10344(.A1(new_n13374_), .A2(new_n13364_), .B1(new_n13103_), .B2(new_n13362_), .ZN(new_n13375_));
  AOI21_X1   g10345(.A1(new_n13372_), .A2(new_n13336_), .B(new_n13279_), .ZN(new_n13376_));
  NAND2_X1   g10346(.A1(new_n13142_), .A2(pi0603), .ZN(new_n13377_));
  NAND2_X1   g10347(.A1(new_n13210_), .A2(new_n13377_), .ZN(new_n13378_));
  INV_X1     g10348(.I(new_n13378_), .ZN(new_n13379_));
  NOR2_X1    g10349(.A1(new_n12809_), .A2(new_n13379_), .ZN(new_n13380_));
  INV_X1     g10350(.I(new_n13380_), .ZN(new_n13381_));
  NOR2_X1    g10351(.A1(new_n13381_), .A2(new_n13336_), .ZN(new_n13382_));
  NOR4_X1    g10352(.A1(new_n13274_), .A2(new_n13376_), .A3(new_n13296_), .A4(new_n13382_), .ZN(new_n13383_));
  NAND2_X1   g10353(.A1(new_n13375_), .A2(new_n13383_), .ZN(new_n13384_));
  OAI21_X1   g10354(.A1(new_n13384_), .A2(new_n5397_), .B(new_n3092_), .ZN(new_n13385_));
  NAND2_X1   g10355(.A1(new_n12878_), .A2(new_n5386_), .ZN(new_n13386_));
  NOR2_X1    g10356(.A1(new_n13386_), .A2(new_n13365_), .ZN(new_n13387_));
  INV_X1     g10357(.I(new_n13387_), .ZN(new_n13388_));
  NAND2_X1   g10358(.A1(new_n13363_), .A2(new_n12862_), .ZN(new_n13389_));
  NAND2_X1   g10359(.A1(new_n12930_), .A2(new_n13363_), .ZN(new_n13390_));
  AND3_X2    g10360(.A1(new_n13390_), .A2(new_n5636_), .A3(new_n13389_), .Z(new_n13391_));
  NOR2_X1    g10361(.A1(new_n13391_), .A2(new_n13388_), .ZN(new_n13392_));
  NOR3_X1    g10362(.A1(new_n13392_), .A2(pi0223), .A3(new_n5398_), .ZN(new_n13393_));
  AOI21_X1   g10363(.A1(new_n13386_), .A2(new_n13246_), .B(new_n12845_), .ZN(new_n13394_));
  INV_X1     g10364(.I(new_n13394_), .ZN(new_n13395_));
  NOR2_X1    g10365(.A1(new_n12862_), .A2(new_n5373_), .ZN(new_n13396_));
  AOI21_X1   g10366(.A1(new_n13396_), .A2(new_n5383_), .B(new_n13258_), .ZN(new_n13397_));
  NOR2_X1    g10367(.A1(new_n12922_), .A2(new_n13258_), .ZN(new_n13398_));
  INV_X1     g10368(.I(new_n13398_), .ZN(new_n13399_));
  NOR4_X1    g10369(.A1(new_n13399_), .A2(new_n13395_), .A3(new_n5375_), .A4(new_n13397_), .ZN(new_n13400_));
  NAND2_X1   g10370(.A1(new_n13400_), .A2(pi0299), .ZN(new_n13401_));
  OAI21_X1   g10371(.A1(new_n13393_), .A2(new_n13401_), .B(new_n5397_), .ZN(new_n13402_));
  NAND2_X1   g10372(.A1(new_n13386_), .A2(new_n13363_), .ZN(new_n13403_));
  NAND3_X1   g10373(.A1(new_n13390_), .A2(new_n5636_), .A3(new_n13403_), .ZN(new_n13404_));
  NAND2_X1   g10374(.A1(new_n13404_), .A2(new_n13387_), .ZN(new_n13405_));
  INV_X1     g10375(.I(new_n13397_), .ZN(new_n13406_));
  INV_X1     g10376(.I(new_n13403_), .ZN(new_n13407_));
  NOR2_X1    g10377(.A1(new_n13296_), .A2(new_n13365_), .ZN(new_n13408_));
  OAI21_X1   g10378(.A1(new_n13406_), .A2(new_n13408_), .B(new_n13407_), .ZN(new_n13409_));
  NOR2_X1    g10379(.A1(new_n13405_), .A2(new_n13409_), .ZN(new_n13410_));
  OAI21_X1   g10380(.A1(new_n13410_), .A2(pi0680), .B(new_n13394_), .ZN(new_n13411_));
  NOR2_X1    g10381(.A1(new_n3092_), .A2(new_n3090_), .ZN(new_n13412_));
  NOR2_X1    g10382(.A1(new_n12784_), .A2(new_n13412_), .ZN(new_n13413_));
  NOR3_X1    g10383(.A1(new_n13411_), .A2(new_n13301_), .A3(new_n13413_), .ZN(new_n13414_));
  NAND2_X1   g10384(.A1(new_n13402_), .A2(new_n13414_), .ZN(new_n13415_));
  NOR2_X1    g10385(.A1(new_n12806_), .A2(new_n5636_), .ZN(new_n13416_));
  AOI21_X1   g10386(.A1(new_n12826_), .A2(new_n5636_), .B(new_n13416_), .ZN(new_n13417_));
  NOR2_X1    g10387(.A1(new_n13417_), .A2(new_n13103_), .ZN(new_n13418_));
  OAI21_X1   g10388(.A1(new_n13234_), .A2(new_n13238_), .B(new_n13418_), .ZN(new_n13419_));
  AOI21_X1   g10389(.A1(new_n13103_), .A2(new_n13361_), .B(new_n13263_), .ZN(new_n13420_));
  INV_X1     g10390(.I(new_n13420_), .ZN(new_n13421_));
  NOR2_X1    g10391(.A1(new_n13232_), .A2(new_n5794_), .ZN(new_n13422_));
  OAI21_X1   g10392(.A1(new_n13253_), .A2(pi0621), .B(new_n12813_), .ZN(new_n13423_));
  NAND2_X1   g10393(.A1(new_n13423_), .A2(pi0603), .ZN(new_n13424_));
  OAI21_X1   g10394(.A1(new_n13247_), .A2(new_n13424_), .B(new_n13422_), .ZN(new_n13425_));
  NOR3_X1    g10395(.A1(new_n13247_), .A2(new_n13422_), .A3(new_n13424_), .ZN(new_n13426_));
  NOR2_X1    g10396(.A1(new_n13426_), .A2(new_n13296_), .ZN(new_n13427_));
  NOR2_X1    g10397(.A1(new_n13296_), .A2(new_n13365_), .ZN(new_n13428_));
  INV_X1     g10398(.I(new_n13428_), .ZN(new_n13429_));
  AOI21_X1   g10399(.A1(new_n13427_), .A2(new_n13425_), .B(new_n13429_), .ZN(new_n13430_));
  AND3_X2    g10400(.A1(new_n13427_), .A2(new_n13425_), .A3(new_n13429_), .Z(new_n13431_));
  OAI21_X1   g10401(.A1(new_n13431_), .A2(new_n13430_), .B(new_n13421_), .ZN(new_n13432_));
  NAND3_X1   g10402(.A1(new_n13432_), .A2(new_n5397_), .A3(new_n13419_), .ZN(new_n13433_));
  AOI21_X1   g10403(.A1(new_n13385_), .A2(new_n13415_), .B(new_n13433_), .ZN(new_n13434_));
  INV_X1     g10404(.I(new_n13384_), .ZN(new_n13435_));
  INV_X1     g10405(.I(new_n13419_), .ZN(new_n13436_));
  NOR2_X1    g10406(.A1(new_n13436_), .A2(new_n5455_), .ZN(new_n13437_));
  INV_X1     g10407(.I(new_n13437_), .ZN(new_n13438_));
  NOR2_X1    g10408(.A1(new_n13432_), .A2(new_n5455_), .ZN(new_n13439_));
  NAND3_X1   g10409(.A1(new_n13439_), .A2(new_n13435_), .A3(new_n13438_), .ZN(new_n13440_));
  INV_X1     g10410(.I(new_n13440_), .ZN(new_n13441_));
  AOI21_X1   g10411(.A1(new_n13439_), .A2(new_n13435_), .B(new_n13438_), .ZN(new_n13442_));
  NAND2_X1   g10412(.A1(new_n13411_), .A2(pi0215), .ZN(new_n13443_));
  XOR2_X1    g10413(.A1(new_n13443_), .A2(new_n13309_), .Z(new_n13444_));
  INV_X1     g10414(.I(new_n13392_), .ZN(new_n13445_));
  NOR2_X1    g10415(.A1(new_n3312_), .A2(pi0215), .ZN(new_n13446_));
  INV_X1     g10416(.I(new_n13446_), .ZN(new_n13447_));
  NOR2_X1    g10417(.A1(new_n12784_), .A2(new_n13447_), .ZN(new_n13448_));
  NOR4_X1    g10418(.A1(new_n13445_), .A2(new_n13301_), .A3(new_n13400_), .A4(new_n13448_), .ZN(new_n13449_));
  NAND2_X1   g10419(.A1(new_n13444_), .A2(new_n13449_), .ZN(new_n13450_));
  INV_X1     g10420(.I(new_n13450_), .ZN(new_n13451_));
  OAI22_X1   g10421(.A1(new_n13441_), .A2(new_n13442_), .B1(new_n13451_), .B2(new_n3312_), .ZN(new_n13452_));
  AOI21_X1   g10422(.A1(new_n13452_), .A2(pi0299), .B(new_n13434_), .ZN(new_n13453_));
  NAND3_X1   g10423(.A1(new_n13453_), .A2(pi0140), .A3(pi0761), .ZN(new_n13454_));
  NAND2_X1   g10424(.A1(new_n13385_), .A2(new_n13415_), .ZN(new_n13455_));
  INV_X1     g10425(.I(new_n13432_), .ZN(new_n13456_));
  NOR2_X1    g10426(.A1(new_n13456_), .A2(new_n13436_), .ZN(new_n13457_));
  NAND3_X1   g10427(.A1(new_n13457_), .A2(new_n13455_), .A3(new_n5397_), .ZN(new_n13458_));
  INV_X1     g10428(.I(new_n13442_), .ZN(new_n13459_));
  AOI22_X1   g10429(.A1(new_n13459_), .A2(new_n13440_), .B1(new_n3313_), .B2(new_n13450_), .ZN(new_n13460_));
  OAI21_X1   g10430(.A1(new_n13460_), .A2(new_n3098_), .B(new_n13458_), .ZN(new_n13461_));
  NAND3_X1   g10431(.A1(new_n13461_), .A2(pi0140), .A3(new_n13099_), .ZN(new_n13462_));
  NOR2_X1    g10432(.A1(new_n12780_), .A2(pi0120), .ZN(new_n13463_));
  NOR2_X1    g10433(.A1(new_n3091_), .A2(pi0223), .ZN(new_n13464_));
  NAND2_X1   g10434(.A1(new_n13208_), .A2(new_n13464_), .ZN(new_n13465_));
  INV_X1     g10435(.I(new_n5481_), .ZN(new_n13466_));
  NOR3_X1    g10436(.A1(new_n12855_), .A2(new_n2726_), .A3(new_n12871_), .ZN(new_n13467_));
  NAND2_X1   g10437(.A1(new_n13467_), .A2(pi0665), .ZN(new_n13468_));
  NAND2_X1   g10438(.A1(new_n13289_), .A2(new_n5373_), .ZN(new_n13469_));
  OAI21_X1   g10439(.A1(new_n5373_), .A2(new_n13468_), .B(new_n13469_), .ZN(new_n13470_));
  NOR2_X1    g10440(.A1(new_n13470_), .A2(new_n5378_), .ZN(new_n13471_));
  NAND2_X1   g10441(.A1(pi0603), .A2(pi0621), .ZN(new_n13472_));
  NOR2_X1    g10442(.A1(new_n5378_), .A2(new_n13206_), .ZN(new_n13473_));
  OAI21_X1   g10443(.A1(new_n13471_), .A2(new_n13472_), .B(new_n13473_), .ZN(new_n13474_));
  NAND2_X1   g10444(.A1(new_n13340_), .A2(new_n13474_), .ZN(new_n13475_));
  NAND2_X1   g10445(.A1(new_n13475_), .A2(pi0223), .ZN(new_n13476_));
  XOR2_X1    g10446(.A1(new_n13476_), .A2(new_n13466_), .Z(new_n13477_));
  INV_X1     g10447(.I(new_n13340_), .ZN(new_n13478_));
  NAND2_X1   g10448(.A1(new_n13243_), .A2(new_n13210_), .ZN(new_n13479_));
  NAND2_X1   g10449(.A1(new_n13479_), .A2(new_n13468_), .ZN(new_n13480_));
  AOI21_X1   g10450(.A1(new_n13478_), .A2(new_n13480_), .B(new_n13296_), .ZN(new_n13481_));
  INV_X1     g10451(.I(new_n13467_), .ZN(new_n13482_));
  NAND3_X1   g10452(.A1(new_n12930_), .A2(pi0680), .A3(new_n13310_), .ZN(new_n13483_));
  AOI21_X1   g10453(.A1(new_n13483_), .A2(new_n5796_), .B(new_n13482_), .ZN(new_n13484_));
  INV_X1     g10454(.I(new_n13468_), .ZN(new_n13485_));
  AOI22_X1   g10455(.A1(new_n13485_), .A2(pi0603), .B1(pi0621), .B2(pi0680), .ZN(new_n13486_));
  NOR2_X1    g10456(.A1(new_n13486_), .A2(new_n5636_), .ZN(new_n13487_));
  OAI21_X1   g10457(.A1(new_n13481_), .A2(new_n13484_), .B(new_n13487_), .ZN(new_n13488_));
  NOR2_X1    g10458(.A1(new_n13488_), .A2(new_n3098_), .ZN(new_n13489_));
  AOI22_X1   g10459(.A1(new_n13477_), .A2(new_n13489_), .B1(new_n13463_), .B2(new_n13465_), .ZN(new_n13490_));
  NOR2_X1    g10460(.A1(new_n13274_), .A2(new_n13338_), .ZN(new_n13491_));
  INV_X1     g10461(.I(new_n13337_), .ZN(new_n13492_));
  NAND2_X1   g10462(.A1(new_n13492_), .A2(new_n5375_), .ZN(new_n13493_));
  NAND2_X1   g10463(.A1(new_n13289_), .A2(new_n13377_), .ZN(new_n13494_));
  OAI21_X1   g10464(.A1(new_n13494_), .A2(new_n13336_), .B(new_n13234_), .ZN(new_n13495_));
  NAND3_X1   g10465(.A1(new_n13495_), .A2(new_n13204_), .A3(new_n13338_), .ZN(new_n13496_));
  AOI22_X1   g10466(.A1(new_n13491_), .A2(new_n13493_), .B1(new_n13273_), .B2(new_n13496_), .ZN(new_n13497_));
  OAI21_X1   g10467(.A1(new_n13290_), .A2(new_n5373_), .B(new_n13469_), .ZN(new_n13498_));
  INV_X1     g10468(.I(new_n13498_), .ZN(new_n13499_));
  NOR4_X1    g10469(.A1(new_n13497_), .A2(new_n5636_), .A3(new_n13378_), .A4(new_n13499_), .ZN(new_n13500_));
  OAI21_X1   g10470(.A1(new_n13290_), .A2(new_n5636_), .B(new_n5794_), .ZN(new_n13501_));
  NAND3_X1   g10471(.A1(new_n13501_), .A2(pi0621), .A3(new_n13234_), .ZN(new_n13502_));
  NAND2_X1   g10472(.A1(new_n13502_), .A2(new_n13378_), .ZN(new_n13503_));
  NAND4_X1   g10473(.A1(new_n13290_), .A2(new_n5386_), .A3(new_n5383_), .A4(new_n13479_), .ZN(new_n13504_));
  NOR2_X1    g10474(.A1(new_n13504_), .A2(new_n5375_), .ZN(new_n13505_));
  NAND2_X1   g10475(.A1(new_n13503_), .A2(new_n13505_), .ZN(new_n13506_));
  AOI21_X1   g10476(.A1(new_n13506_), .A2(new_n12821_), .B(new_n13103_), .ZN(new_n13507_));
  NOR2_X1    g10477(.A1(new_n13507_), .A2(new_n5397_), .ZN(new_n13508_));
  XOR2_X1    g10478(.A1(new_n13508_), .A2(new_n12981_), .Z(new_n13509_));
  NAND2_X1   g10479(.A1(new_n13509_), .A2(new_n13500_), .ZN(new_n13510_));
  NOR2_X1    g10480(.A1(new_n13510_), .A2(new_n13490_), .ZN(new_n13511_));
  NAND2_X1   g10481(.A1(new_n13208_), .A2(new_n13446_), .ZN(new_n13512_));
  NAND2_X1   g10482(.A1(new_n13475_), .A2(pi0215), .ZN(new_n13513_));
  XOR2_X1    g10483(.A1(new_n13513_), .A2(new_n13309_), .Z(new_n13514_));
  AOI22_X1   g10484(.A1(new_n13514_), .A2(new_n13489_), .B1(new_n13463_), .B2(new_n13512_), .ZN(new_n13515_));
  NOR2_X1    g10485(.A1(new_n5455_), .A2(new_n3313_), .ZN(new_n13516_));
  NOR2_X1    g10486(.A1(new_n13507_), .A2(new_n5455_), .ZN(new_n13517_));
  XOR2_X1    g10487(.A1(new_n13517_), .A2(new_n13516_), .Z(new_n13518_));
  NAND2_X1   g10488(.A1(new_n13518_), .A2(new_n13500_), .ZN(new_n13519_));
  NOR2_X1    g10489(.A1(new_n13519_), .A2(new_n13515_), .ZN(new_n13520_));
  NOR2_X1    g10490(.A1(new_n13511_), .A2(new_n13520_), .ZN(new_n13521_));
  NAND2_X1   g10491(.A1(new_n13521_), .A2(pi0039), .ZN(new_n13522_));
  AOI21_X1   g10492(.A1(new_n13454_), .A2(new_n13462_), .B(new_n13522_), .ZN(new_n13523_));
  NAND2_X1   g10493(.A1(new_n12784_), .A2(new_n13212_), .ZN(new_n13524_));
  INV_X1     g10494(.I(new_n13524_), .ZN(new_n13525_));
  NOR2_X1    g10495(.A1(new_n13525_), .A2(new_n12841_), .ZN(new_n13526_));
  INV_X1     g10496(.I(new_n13526_), .ZN(new_n13527_));
  NAND3_X1   g10497(.A1(new_n12806_), .A2(new_n12784_), .A3(new_n13282_), .ZN(new_n13528_));
  NAND3_X1   g10498(.A1(new_n12818_), .A2(new_n12809_), .A3(new_n13282_), .ZN(new_n13529_));
  NAND2_X1   g10499(.A1(new_n13528_), .A2(new_n13529_), .ZN(new_n13530_));
  NAND3_X1   g10500(.A1(new_n13530_), .A2(pi0642), .A3(new_n13211_), .ZN(new_n13531_));
  NAND4_X1   g10501(.A1(new_n13528_), .A2(new_n13529_), .A3(pi0642), .A4(new_n13212_), .ZN(new_n13532_));
  AOI21_X1   g10502(.A1(new_n13531_), .A2(new_n13532_), .B(new_n12809_), .ZN(new_n13533_));
  NOR2_X1    g10503(.A1(new_n13533_), .A2(new_n12868_), .ZN(new_n13534_));
  XOR2_X1    g10504(.A1(new_n13534_), .A2(new_n12870_), .Z(new_n13535_));
  OAI21_X1   g10505(.A1(new_n13535_), .A2(new_n13524_), .B(new_n13527_), .ZN(new_n13536_));
  NAND2_X1   g10506(.A1(new_n13536_), .A2(new_n13234_), .ZN(new_n13537_));
  NOR2_X1    g10507(.A1(new_n12960_), .A2(pi0680), .ZN(new_n13538_));
  NOR2_X1    g10508(.A1(new_n13538_), .A2(new_n13295_), .ZN(new_n13539_));
  NAND2_X1   g10509(.A1(new_n13501_), .A2(pi0621), .ZN(new_n13540_));
  NOR3_X1    g10510(.A1(new_n12813_), .A2(new_n5794_), .A3(new_n13142_), .ZN(new_n13541_));
  INV_X1     g10511(.I(new_n13541_), .ZN(new_n13542_));
  OAI22_X1   g10512(.A1(new_n13540_), .A2(new_n12821_), .B1(new_n5375_), .B2(new_n13542_), .ZN(new_n13543_));
  NAND2_X1   g10513(.A1(new_n13543_), .A2(new_n13234_), .ZN(new_n13544_));
  AOI21_X1   g10514(.A1(new_n13544_), .A2(new_n12821_), .B(new_n13212_), .ZN(new_n13545_));
  NAND3_X1   g10515(.A1(new_n13539_), .A2(new_n13545_), .A3(new_n5454_), .ZN(new_n13546_));
  AOI21_X1   g10516(.A1(new_n13537_), .A2(new_n5454_), .B(new_n13546_), .ZN(new_n13547_));
  INV_X1     g10517(.I(new_n13547_), .ZN(new_n13548_));
  NAND3_X1   g10518(.A1(new_n13537_), .A2(new_n5454_), .A3(new_n13546_), .ZN(new_n13549_));
  NAND2_X1   g10519(.A1(new_n13548_), .A2(new_n13549_), .ZN(new_n13550_));
  NAND2_X1   g10520(.A1(new_n13403_), .A2(new_n5379_), .ZN(new_n13551_));
  NAND2_X1   g10521(.A1(new_n13389_), .A2(new_n13468_), .ZN(new_n13552_));
  NOR2_X1    g10522(.A1(new_n13479_), .A2(new_n5794_), .ZN(new_n13553_));
  NAND2_X1   g10523(.A1(new_n13552_), .A2(new_n13553_), .ZN(new_n13554_));
  NAND2_X1   g10524(.A1(new_n13524_), .A2(pi0642), .ZN(new_n13555_));
  NAND3_X1   g10525(.A1(new_n13554_), .A2(new_n13551_), .A3(new_n13555_), .ZN(new_n13556_));
  NAND4_X1   g10526(.A1(new_n13556_), .A2(pi0614), .A3(pi0616), .A4(new_n13470_), .ZN(new_n13557_));
  NAND2_X1   g10527(.A1(new_n13556_), .A2(new_n13470_), .ZN(new_n13558_));
  NAND3_X1   g10528(.A1(new_n13558_), .A2(pi0614), .A3(new_n12870_), .ZN(new_n13559_));
  AOI21_X1   g10529(.A1(new_n13559_), .A2(new_n13557_), .B(new_n13524_), .ZN(new_n13560_));
  NOR2_X1    g10530(.A1(new_n12927_), .A2(pi0680), .ZN(new_n13561_));
  NOR3_X1    g10531(.A1(new_n13470_), .A2(new_n5636_), .A3(new_n13407_), .ZN(new_n13562_));
  NOR3_X1    g10532(.A1(new_n13561_), .A2(new_n13562_), .A3(new_n13296_), .ZN(new_n13563_));
  OAI21_X1   g10533(.A1(new_n13560_), .A2(new_n13563_), .B(new_n13526_), .ZN(new_n13564_));
  AOI21_X1   g10534(.A1(new_n13564_), .A2(pi0215), .B(new_n13309_), .ZN(new_n13565_));
  INV_X1     g10535(.I(new_n13564_), .ZN(new_n13566_));
  NOR3_X1    g10536(.A1(new_n13566_), .A2(new_n3111_), .A3(new_n5454_), .ZN(new_n13567_));
  NAND2_X1   g10537(.A1(new_n13390_), .A2(new_n13336_), .ZN(new_n13568_));
  NOR3_X1    g10538(.A1(new_n13554_), .A2(new_n13365_), .A3(new_n13480_), .ZN(new_n13569_));
  XOR2_X1    g10539(.A1(new_n13569_), .A2(new_n13568_), .Z(new_n13570_));
  OAI22_X1   g10540(.A1(new_n13570_), .A2(new_n13552_), .B1(new_n5636_), .B2(new_n13296_), .ZN(new_n13571_));
  OAI21_X1   g10541(.A1(pi0680), .A2(new_n12924_), .B(new_n13571_), .ZN(new_n13572_));
  NOR2_X1    g10542(.A1(new_n12784_), .A2(new_n12832_), .ZN(new_n13573_));
  NOR3_X1    g10543(.A1(new_n13572_), .A2(new_n13324_), .A3(new_n13573_), .ZN(new_n13574_));
  OAI21_X1   g10544(.A1(new_n13565_), .A2(new_n13567_), .B(new_n13574_), .ZN(new_n13575_));
  NAND2_X1   g10545(.A1(new_n13575_), .A2(new_n3313_), .ZN(new_n13576_));
  NAND2_X1   g10546(.A1(new_n13550_), .A2(new_n13576_), .ZN(new_n13577_));
  NAND3_X1   g10547(.A1(new_n13566_), .A2(pi0223), .A3(new_n5398_), .ZN(new_n13578_));
  NAND3_X1   g10548(.A1(new_n13564_), .A2(pi0223), .A3(new_n5397_), .ZN(new_n13579_));
  AOI21_X1   g10549(.A1(new_n13578_), .A2(new_n13579_), .B(new_n13572_), .ZN(new_n13580_));
  NAND2_X1   g10550(.A1(new_n12784_), .A2(new_n13324_), .ZN(new_n13581_));
  AOI21_X1   g10551(.A1(new_n13581_), .A2(new_n3091_), .B(pi0223), .ZN(new_n13582_));
  INV_X1     g10552(.I(new_n13582_), .ZN(new_n13583_));
  NOR2_X1    g10553(.A1(new_n13580_), .A2(new_n13583_), .ZN(new_n13584_));
  AOI21_X1   g10554(.A1(new_n13545_), .A2(new_n5397_), .B(new_n3091_), .ZN(new_n13585_));
  NOR3_X1    g10555(.A1(new_n13585_), .A2(new_n5398_), .A3(new_n13539_), .ZN(new_n13586_));
  NOR3_X1    g10556(.A1(new_n13584_), .A2(new_n13537_), .A3(new_n13586_), .ZN(new_n13587_));
  NAND3_X1   g10557(.A1(new_n13587_), .A2(pi0140), .A3(pi0299), .ZN(new_n13588_));
  NOR3_X1    g10558(.A1(new_n13587_), .A2(pi0140), .A3(new_n3098_), .ZN(new_n13589_));
  INV_X1     g10559(.I(new_n13589_), .ZN(new_n13590_));
  AOI21_X1   g10560(.A1(new_n13590_), .A2(new_n13588_), .B(new_n13577_), .ZN(new_n13591_));
  OAI21_X1   g10561(.A1(new_n13523_), .A2(new_n13360_), .B(new_n13591_), .ZN(new_n13592_));
  OAI21_X1   g10562(.A1(new_n13592_), .A2(new_n13228_), .B(new_n3289_), .ZN(new_n13593_));
  NAND2_X1   g10563(.A1(new_n13098_), .A2(pi0738), .ZN(new_n13594_));
  NAND2_X1   g10564(.A1(pi0038), .A2(pi0738), .ZN(new_n13595_));
  XOR2_X1    g10565(.A1(new_n13594_), .A2(new_n13595_), .Z(new_n13596_));
  AND3_X2    g10566(.A1(new_n13110_), .A2(pi0140), .A3(new_n3289_), .Z(new_n13597_));
  NAND3_X1   g10567(.A1(new_n13593_), .A2(new_n13596_), .A3(new_n13597_), .ZN(new_n13598_));
  INV_X1     g10568(.I(new_n13228_), .ZN(new_n13599_));
  INV_X1     g10569(.I(new_n13360_), .ZN(new_n13600_));
  AOI21_X1   g10570(.A1(new_n13461_), .A2(pi0140), .B(new_n13101_), .ZN(new_n13601_));
  INV_X1     g10571(.I(new_n13462_), .ZN(new_n13602_));
  INV_X1     g10572(.I(new_n13522_), .ZN(new_n13603_));
  OAI21_X1   g10573(.A1(new_n13602_), .A2(new_n13601_), .B(new_n13603_), .ZN(new_n13604_));
  AOI22_X1   g10574(.A1(new_n13548_), .A2(new_n13549_), .B1(new_n13575_), .B2(new_n3313_), .ZN(new_n13605_));
  INV_X1     g10575(.I(new_n13588_), .ZN(new_n13606_));
  OAI21_X1   g10576(.A1(new_n13606_), .A2(new_n13589_), .B(new_n13605_), .ZN(new_n13607_));
  AOI21_X1   g10577(.A1(new_n13604_), .A2(new_n13600_), .B(new_n13607_), .ZN(new_n13608_));
  AOI21_X1   g10578(.A1(new_n13599_), .A2(new_n13608_), .B(new_n3290_), .ZN(new_n13609_));
  NAND2_X1   g10579(.A1(new_n13596_), .A2(new_n13597_), .ZN(new_n13610_));
  NAND2_X1   g10580(.A1(new_n13609_), .A2(new_n13610_), .ZN(new_n13611_));
  NAND3_X1   g10581(.A1(new_n13611_), .A2(new_n13598_), .A3(pi1153), .ZN(new_n13612_));
  INV_X1     g10582(.I(pi0625), .ZN(new_n13613_));
  INV_X1     g10583(.I(pi1153), .ZN(new_n13614_));
  NOR2_X1    g10584(.A1(new_n13613_), .A2(new_n13614_), .ZN(new_n13615_));
  NAND2_X1   g10585(.A1(new_n13612_), .A2(new_n13615_), .ZN(new_n13616_));
  NOR2_X1    g10586(.A1(new_n13609_), .A2(new_n13610_), .ZN(new_n13617_));
  AOI21_X1   g10587(.A1(new_n13596_), .A2(new_n13597_), .B(new_n13593_), .ZN(new_n13618_));
  NOR3_X1    g10588(.A1(new_n13617_), .A2(new_n13618_), .A3(new_n13614_), .ZN(new_n13619_));
  INV_X1     g10589(.I(new_n13615_), .ZN(new_n13620_));
  NAND2_X1   g10590(.A1(new_n13619_), .A2(new_n13620_), .ZN(new_n13621_));
  AOI21_X1   g10591(.A1(new_n13621_), .A2(new_n13616_), .B(new_n13115_), .ZN(new_n13622_));
  AOI21_X1   g10592(.A1(new_n13073_), .A2(new_n13096_), .B(pi0038), .ZN(new_n13623_));
  NOR2_X1    g10593(.A1(new_n7499_), .A2(new_n2723_), .ZN(new_n13624_));
  INV_X1     g10594(.I(new_n13624_), .ZN(new_n13625_));
  NOR2_X1    g10595(.A1(new_n13625_), .A2(new_n3259_), .ZN(new_n13626_));
  OAI21_X1   g10596(.A1(new_n13623_), .A2(new_n13626_), .B(new_n3289_), .ZN(new_n13627_));
  NAND2_X1   g10597(.A1(new_n13627_), .A2(new_n7971_), .ZN(new_n13628_));
  INV_X1     g10598(.I(new_n13628_), .ZN(new_n13629_));
  AOI21_X1   g10599(.A1(new_n13085_), .A2(pi0039), .B(new_n13095_), .ZN(new_n13630_));
  NOR3_X1    g10600(.A1(new_n12977_), .A2(new_n13072_), .A3(new_n3183_), .ZN(new_n13631_));
  NOR2_X1    g10601(.A1(new_n13631_), .A2(new_n13630_), .ZN(new_n13632_));
  INV_X1     g10602(.I(new_n13626_), .ZN(new_n13633_));
  OAI21_X1   g10603(.A1(new_n13632_), .A2(pi0038), .B(new_n13633_), .ZN(new_n13634_));
  NAND2_X1   g10604(.A1(new_n7971_), .A2(pi0738), .ZN(new_n13635_));
  OAI21_X1   g10605(.A1(new_n13634_), .A2(new_n13635_), .B(new_n3289_), .ZN(new_n13636_));
  NAND3_X1   g10606(.A1(new_n12960_), .A2(pi0680), .A3(new_n12844_), .ZN(new_n13637_));
  NAND2_X1   g10607(.A1(new_n12844_), .A2(pi0680), .ZN(new_n13638_));
  NAND3_X1   g10608(.A1(new_n12971_), .A2(new_n12844_), .A3(new_n13638_), .ZN(new_n13639_));
  AOI21_X1   g10609(.A1(new_n13639_), .A2(new_n13637_), .B(new_n13499_), .ZN(new_n13640_));
  AOI21_X1   g10610(.A1(new_n13289_), .A2(new_n5796_), .B(new_n5375_), .ZN(new_n13641_));
  INV_X1     g10611(.I(new_n13641_), .ZN(new_n13642_));
  AOI21_X1   g10612(.A1(new_n13498_), .A2(new_n5383_), .B(new_n13642_), .ZN(new_n13643_));
  OAI21_X1   g10613(.A1(new_n13643_), .A2(new_n12844_), .B(pi0680), .ZN(new_n13644_));
  NOR2_X1    g10614(.A1(new_n12971_), .A2(new_n13644_), .ZN(new_n13645_));
  NAND2_X1   g10615(.A1(new_n13504_), .A2(pi0680), .ZN(new_n13646_));
  XNOR2_X1   g10616(.A1(new_n13646_), .A2(new_n13638_), .ZN(new_n13647_));
  OAI22_X1   g10617(.A1(new_n13647_), .A2(new_n13290_), .B1(pi0680), .B2(new_n12826_), .ZN(new_n13648_));
  OAI21_X1   g10618(.A1(new_n13648_), .A2(new_n3091_), .B(new_n5397_), .ZN(new_n13649_));
  OAI21_X1   g10619(.A1(new_n13649_), .A2(new_n13645_), .B(new_n13640_), .ZN(new_n13650_));
  AOI21_X1   g10620(.A1(new_n12987_), .A2(new_n13205_), .B(pi0223), .ZN(new_n13651_));
  NOR2_X1    g10621(.A1(new_n13641_), .A2(new_n5378_), .ZN(new_n13652_));
  NOR2_X1    g10622(.A1(new_n13470_), .A2(new_n13652_), .ZN(new_n13653_));
  NOR2_X1    g10623(.A1(new_n13561_), .A2(new_n13653_), .ZN(new_n13654_));
  INV_X1     g10624(.I(new_n13654_), .ZN(new_n13655_));
  OAI21_X1   g10625(.A1(new_n13479_), .A2(new_n5383_), .B(pi0680), .ZN(new_n13656_));
  NOR3_X1    g10626(.A1(new_n12932_), .A2(new_n5375_), .A3(new_n13468_), .ZN(new_n13657_));
  NAND2_X1   g10627(.A1(new_n13657_), .A2(new_n13656_), .ZN(new_n13658_));
  INV_X1     g10628(.I(new_n13656_), .ZN(new_n13659_));
  NAND3_X1   g10629(.A1(new_n12924_), .A2(pi0680), .A3(new_n13485_), .ZN(new_n13660_));
  NAND2_X1   g10630(.A1(new_n13660_), .A2(new_n13659_), .ZN(new_n13661_));
  AOI21_X1   g10631(.A1(new_n13658_), .A2(new_n13661_), .B(new_n13653_), .ZN(new_n13662_));
  NAND3_X1   g10632(.A1(new_n13662_), .A2(pi0223), .A3(new_n5398_), .ZN(new_n13663_));
  NOR2_X1    g10633(.A1(new_n13660_), .A2(new_n13659_), .ZN(new_n13664_));
  NOR2_X1    g10634(.A1(new_n13657_), .A2(new_n13656_), .ZN(new_n13665_));
  OAI22_X1   g10635(.A1(new_n13665_), .A2(new_n13664_), .B1(new_n13470_), .B2(new_n13652_), .ZN(new_n13666_));
  NAND3_X1   g10636(.A1(new_n13666_), .A2(pi0223), .A3(new_n13466_), .ZN(new_n13667_));
  AOI21_X1   g10637(.A1(new_n13667_), .A2(new_n13663_), .B(new_n13655_), .ZN(new_n13668_));
  AOI21_X1   g10638(.A1(new_n13668_), .A2(pi0299), .B(new_n13651_), .ZN(new_n13669_));
  XOR2_X1    g10639(.A1(new_n13646_), .A2(new_n13638_), .Z(new_n13670_));
  NOR2_X1    g10640(.A1(new_n12826_), .A2(pi0680), .ZN(new_n13671_));
  AOI21_X1   g10641(.A1(new_n13670_), .A2(new_n13292_), .B(new_n13671_), .ZN(new_n13672_));
  OAI21_X1   g10642(.A1(new_n13672_), .A2(new_n5454_), .B(new_n3313_), .ZN(new_n13673_));
  NOR2_X1    g10643(.A1(new_n13645_), .A2(new_n5454_), .ZN(new_n13674_));
  NAND2_X1   g10644(.A1(new_n13673_), .A2(new_n13674_), .ZN(new_n13675_));
  OAI21_X1   g10645(.A1(pi0120), .A2(new_n12778_), .B(new_n3160_), .ZN(new_n13676_));
  INV_X1     g10646(.I(new_n13676_), .ZN(new_n13677_));
  NOR2_X1    g10647(.A1(new_n13677_), .A2(new_n13447_), .ZN(new_n13678_));
  NOR2_X1    g10648(.A1(new_n13206_), .A2(new_n2723_), .ZN(new_n13679_));
  INV_X1     g10649(.I(new_n13679_), .ZN(new_n13680_));
  AOI21_X1   g10650(.A1(new_n13666_), .A2(pi0215), .B(new_n13309_), .ZN(new_n13681_));
  NOR3_X1    g10651(.A1(new_n13662_), .A2(new_n3111_), .A3(new_n5454_), .ZN(new_n13682_));
  OAI21_X1   g10652(.A1(new_n13681_), .A2(new_n13682_), .B(new_n13654_), .ZN(new_n13683_));
  OAI22_X1   g10653(.A1(new_n13683_), .A2(new_n3098_), .B1(new_n13678_), .B2(new_n13680_), .ZN(new_n13684_));
  NAND3_X1   g10654(.A1(new_n13684_), .A2(new_n13640_), .A3(new_n13675_), .ZN(new_n13685_));
  OAI21_X1   g10655(.A1(new_n13650_), .A2(new_n13669_), .B(new_n13685_), .ZN(new_n13686_));
  NOR2_X1    g10656(.A1(new_n3183_), .A2(new_n7971_), .ZN(new_n13687_));
  NAND2_X1   g10657(.A1(new_n13259_), .A2(new_n12949_), .ZN(new_n13688_));
  AOI21_X1   g10658(.A1(new_n13688_), .A2(new_n12844_), .B(new_n5375_), .ZN(new_n13689_));
  NOR2_X1    g10659(.A1(new_n13246_), .A2(new_n5383_), .ZN(new_n13690_));
  AOI21_X1   g10660(.A1(new_n13688_), .A2(new_n5383_), .B(new_n13690_), .ZN(new_n13691_));
  OAI21_X1   g10661(.A1(new_n13691_), .A2(new_n12844_), .B(new_n13689_), .ZN(new_n13692_));
  NOR2_X1    g10662(.A1(new_n13238_), .A2(new_n13206_), .ZN(new_n13693_));
  AOI21_X1   g10663(.A1(new_n12821_), .A2(new_n13693_), .B(new_n12845_), .ZN(new_n13694_));
  NOR3_X1    g10664(.A1(new_n12809_), .A2(new_n3092_), .A3(new_n13205_), .ZN(new_n13695_));
  NAND2_X1   g10665(.A1(new_n13695_), .A2(new_n3092_), .ZN(new_n13696_));
  AOI21_X1   g10666(.A1(new_n13694_), .A2(new_n5397_), .B(new_n13696_), .ZN(new_n13697_));
  NOR2_X1    g10667(.A1(new_n13697_), .A2(new_n5398_), .ZN(new_n13698_));
  OR2_X2     g10668(.A1(new_n13698_), .A2(new_n13692_), .Z(new_n13699_));
  NOR2_X1    g10669(.A1(new_n12930_), .A2(new_n5398_), .ZN(new_n13700_));
  INV_X1     g10670(.I(new_n13700_), .ZN(new_n13701_));
  NAND3_X1   g10671(.A1(new_n13701_), .A2(pi0680), .A3(new_n13397_), .ZN(new_n13702_));
  NOR3_X1    g10672(.A1(new_n13702_), .A2(new_n3090_), .A3(new_n13394_), .ZN(new_n13703_));
  AOI21_X1   g10673(.A1(new_n13703_), .A2(pi0299), .B(pi0223), .ZN(new_n13704_));
  AOI21_X1   g10674(.A1(new_n13694_), .A2(new_n5455_), .B(new_n3313_), .ZN(new_n13705_));
  NAND2_X1   g10675(.A1(new_n13689_), .A2(new_n5454_), .ZN(new_n13706_));
  NOR2_X1    g10676(.A1(new_n12809_), .A2(new_n13205_), .ZN(new_n13707_));
  NAND3_X1   g10677(.A1(new_n13707_), .A2(new_n3312_), .A3(new_n12844_), .ZN(new_n13708_));
  AOI21_X1   g10678(.A1(new_n13706_), .A2(new_n13691_), .B(new_n13708_), .ZN(new_n13709_));
  XOR2_X1    g10679(.A1(new_n13709_), .A2(new_n13705_), .Z(new_n13710_));
  NAND2_X1   g10680(.A1(new_n12922_), .A2(new_n5454_), .ZN(new_n13711_));
  AOI21_X1   g10681(.A1(new_n5375_), .A2(new_n13397_), .B(new_n13711_), .ZN(new_n13712_));
  NAND3_X1   g10682(.A1(new_n13712_), .A2(pi0215), .A3(new_n13395_), .ZN(new_n13713_));
  OAI21_X1   g10683(.A1(new_n13713_), .A2(new_n3098_), .B(new_n3111_), .ZN(new_n13714_));
  NAND2_X1   g10684(.A1(new_n13710_), .A2(new_n13714_), .ZN(new_n13715_));
  OAI21_X1   g10685(.A1(new_n13699_), .A2(new_n13704_), .B(new_n13715_), .ZN(new_n13716_));
  NAND2_X1   g10686(.A1(new_n13716_), .A2(pi0039), .ZN(new_n13717_));
  XOR2_X1    g10687(.A1(new_n13717_), .A2(new_n13687_), .Z(new_n13718_));
  NOR2_X1    g10688(.A1(new_n5504_), .A2(new_n13219_), .ZN(new_n13719_));
  NOR2_X1    g10689(.A1(new_n13719_), .A2(new_n3259_), .ZN(new_n13720_));
  INV_X1     g10690(.I(new_n13720_), .ZN(new_n13721_));
  OAI21_X1   g10691(.A1(new_n13721_), .A2(new_n13226_), .B(new_n7971_), .ZN(new_n13722_));
  NOR2_X1    g10692(.A1(new_n13109_), .A2(new_n3259_), .ZN(new_n13723_));
  NAND2_X1   g10693(.A1(new_n13722_), .A2(new_n13723_), .ZN(new_n13724_));
  OAI21_X1   g10694(.A1(new_n13718_), .A2(new_n13686_), .B(new_n13724_), .ZN(new_n13725_));
  NOR2_X1    g10695(.A1(new_n13165_), .A2(new_n7971_), .ZN(new_n13726_));
  XNOR2_X1   g10696(.A1(new_n13726_), .A2(new_n13687_), .ZN(new_n13727_));
  NAND3_X1   g10697(.A1(new_n13197_), .A2(pi0140), .A3(new_n3289_), .ZN(new_n13728_));
  NOR2_X1    g10698(.A1(new_n13727_), .A2(new_n13728_), .ZN(new_n13729_));
  NAND2_X1   g10699(.A1(new_n13725_), .A2(new_n13729_), .ZN(new_n13730_));
  XNOR2_X1   g10700(.A1(new_n13730_), .A2(new_n13636_), .ZN(new_n13731_));
  AOI21_X1   g10701(.A1(new_n13731_), .A2(pi0625), .B(new_n13620_), .ZN(new_n13732_));
  XOR2_X1    g10702(.A1(new_n13730_), .A2(new_n13636_), .Z(new_n13733_));
  NOR3_X1    g10703(.A1(new_n13733_), .A2(new_n13613_), .A3(new_n13615_), .ZN(new_n13734_));
  OAI21_X1   g10704(.A1(new_n13732_), .A2(new_n13734_), .B(new_n13629_), .ZN(new_n13735_));
  NAND2_X1   g10705(.A1(new_n13735_), .A2(pi0608), .ZN(new_n13736_));
  OAI21_X1   g10706(.A1(new_n13622_), .A2(new_n13736_), .B(pi0778), .ZN(new_n13737_));
  NAND3_X1   g10707(.A1(new_n13611_), .A2(new_n13598_), .A3(pi0625), .ZN(new_n13738_));
  NAND2_X1   g10708(.A1(new_n13738_), .A2(new_n13615_), .ZN(new_n13739_));
  NOR3_X1    g10709(.A1(new_n13617_), .A2(new_n13618_), .A3(new_n13613_), .ZN(new_n13740_));
  NAND2_X1   g10710(.A1(new_n13740_), .A2(new_n13620_), .ZN(new_n13741_));
  NAND2_X1   g10711(.A1(new_n13741_), .A2(new_n13739_), .ZN(new_n13742_));
  NOR2_X1    g10712(.A1(new_n13733_), .A2(new_n13614_), .ZN(new_n13743_));
  NOR2_X1    g10713(.A1(new_n13743_), .A2(new_n13620_), .ZN(new_n13744_));
  NAND2_X1   g10714(.A1(new_n13731_), .A2(pi1153), .ZN(new_n13745_));
  NOR2_X1    g10715(.A1(new_n13745_), .A2(new_n13615_), .ZN(new_n13746_));
  OAI21_X1   g10716(.A1(new_n13746_), .A2(new_n13744_), .B(new_n13629_), .ZN(new_n13747_));
  INV_X1     g10717(.I(pi0778), .ZN(new_n13748_));
  NOR2_X1    g10718(.A1(new_n13748_), .A2(pi0608), .ZN(new_n13749_));
  INV_X1     g10719(.I(new_n13749_), .ZN(new_n13750_));
  AOI21_X1   g10720(.A1(new_n13611_), .A2(new_n13598_), .B(new_n13750_), .ZN(new_n13751_));
  NAND2_X1   g10721(.A1(new_n13747_), .A2(new_n13751_), .ZN(new_n13752_));
  AOI21_X1   g10722(.A1(new_n13742_), .A2(new_n13114_), .B(new_n13752_), .ZN(new_n13753_));
  NAND2_X1   g10723(.A1(new_n13737_), .A2(new_n13753_), .ZN(new_n13754_));
  NOR2_X1    g10724(.A1(new_n13619_), .A2(new_n13620_), .ZN(new_n13755_));
  NOR2_X1    g10725(.A1(new_n13612_), .A2(new_n13615_), .ZN(new_n13756_));
  OAI21_X1   g10726(.A1(new_n13755_), .A2(new_n13756_), .B(new_n13114_), .ZN(new_n13757_));
  INV_X1     g10727(.I(new_n13736_), .ZN(new_n13758_));
  AOI21_X1   g10728(.A1(new_n13757_), .A2(new_n13758_), .B(new_n13748_), .ZN(new_n13759_));
  NOR2_X1    g10729(.A1(new_n13740_), .A2(new_n13620_), .ZN(new_n13760_));
  NOR2_X1    g10730(.A1(new_n13738_), .A2(new_n13615_), .ZN(new_n13761_));
  OAI21_X1   g10731(.A1(new_n13760_), .A2(new_n13761_), .B(new_n13114_), .ZN(new_n13762_));
  NAND3_X1   g10732(.A1(new_n13762_), .A2(new_n13747_), .A3(new_n13751_), .ZN(new_n13763_));
  NAND2_X1   g10733(.A1(new_n13759_), .A2(new_n13763_), .ZN(new_n13764_));
  NAND2_X1   g10734(.A1(new_n13764_), .A2(new_n13754_), .ZN(new_n13765_));
  INV_X1     g10735(.I(pi0609), .ZN(new_n13766_));
  NAND2_X1   g10736(.A1(new_n13735_), .A2(pi0778), .ZN(new_n13767_));
  NOR3_X1    g10737(.A1(new_n13747_), .A2(new_n13748_), .A3(new_n13731_), .ZN(new_n13768_));
  NAND2_X1   g10738(.A1(new_n13768_), .A2(new_n13767_), .ZN(new_n13769_));
  AND2_X2    g10739(.A1(new_n13735_), .A2(pi0778), .Z(new_n13770_));
  NAND2_X1   g10740(.A1(new_n13733_), .A2(pi0778), .ZN(new_n13771_));
  OAI21_X1   g10741(.A1(new_n13747_), .A2(new_n13771_), .B(new_n13770_), .ZN(new_n13772_));
  NAND2_X1   g10742(.A1(new_n13772_), .A2(new_n13769_), .ZN(new_n13773_));
  XNOR2_X1   g10743(.A1(pi0608), .A2(pi1153), .ZN(new_n13774_));
  NOR2_X1    g10744(.A1(new_n13774_), .A2(new_n13748_), .ZN(new_n13775_));
  INV_X1     g10745(.I(new_n13775_), .ZN(new_n13776_));
  NAND3_X1   g10746(.A1(new_n13112_), .A2(new_n13113_), .A3(new_n13776_), .ZN(new_n13777_));
  INV_X1     g10747(.I(pi1155), .ZN(new_n13778_));
  NOR2_X1    g10748(.A1(new_n13775_), .A2(pi0609), .ZN(new_n13779_));
  NOR2_X1    g10749(.A1(new_n13779_), .A2(new_n13778_), .ZN(new_n13780_));
  NAND2_X1   g10750(.A1(new_n13628_), .A2(new_n13780_), .ZN(new_n13781_));
  AOI21_X1   g10751(.A1(new_n13781_), .A2(new_n13777_), .B(new_n13766_), .ZN(new_n13782_));
  INV_X1     g10752(.I(pi0660), .ZN(new_n13783_));
  NOR2_X1    g10753(.A1(new_n13783_), .A2(new_n13778_), .ZN(new_n13784_));
  INV_X1     g10754(.I(new_n13784_), .ZN(new_n13785_));
  NOR2_X1    g10755(.A1(new_n13782_), .A2(new_n13785_), .ZN(new_n13786_));
  INV_X1     g10756(.I(new_n13786_), .ZN(new_n13787_));
  OAI21_X1   g10757(.A1(new_n13773_), .A2(new_n13787_), .B(new_n13766_), .ZN(new_n13788_));
  AOI21_X1   g10758(.A1(new_n13772_), .A2(new_n13769_), .B(new_n13766_), .ZN(new_n13789_));
  INV_X1     g10759(.I(new_n13777_), .ZN(new_n13790_));
  OAI21_X1   g10760(.A1(new_n13629_), .A2(new_n13778_), .B(new_n13766_), .ZN(new_n13791_));
  NAND2_X1   g10761(.A1(new_n13791_), .A2(new_n13790_), .ZN(new_n13792_));
  NOR2_X1    g10762(.A1(pi0660), .A2(pi1155), .ZN(new_n13793_));
  NAND2_X1   g10763(.A1(new_n13792_), .A2(new_n13793_), .ZN(new_n13794_));
  OAI21_X1   g10764(.A1(new_n13789_), .A2(new_n13794_), .B(new_n13766_), .ZN(new_n13795_));
  NAND4_X1   g10765(.A1(new_n13765_), .A2(new_n13795_), .A3(new_n13788_), .A4(pi0785), .ZN(new_n13796_));
  NAND2_X1   g10766(.A1(new_n13765_), .A2(new_n13788_), .ZN(new_n13797_));
  NAND3_X1   g10767(.A1(new_n13765_), .A2(new_n13795_), .A3(pi0785), .ZN(new_n13798_));
  NAND3_X1   g10768(.A1(new_n13798_), .A2(new_n13797_), .A3(pi0785), .ZN(new_n13799_));
  NAND2_X1   g10769(.A1(new_n13799_), .A2(new_n13796_), .ZN(new_n13800_));
  INV_X1     g10770(.I(pi0785), .ZN(new_n13801_));
  XNOR2_X1   g10771(.A1(pi0660), .A2(pi1155), .ZN(new_n13802_));
  NOR2_X1    g10772(.A1(new_n13802_), .A2(new_n13801_), .ZN(new_n13803_));
  AOI21_X1   g10773(.A1(new_n13772_), .A2(new_n13769_), .B(new_n13803_), .ZN(new_n13804_));
  INV_X1     g10774(.I(new_n13803_), .ZN(new_n13805_));
  NOR2_X1    g10775(.A1(new_n13628_), .A2(new_n13805_), .ZN(new_n13806_));
  NOR2_X1    g10776(.A1(new_n13804_), .A2(new_n13806_), .ZN(new_n13807_));
  NOR2_X1    g10777(.A1(new_n13782_), .A2(new_n13801_), .ZN(new_n13808_));
  NOR2_X1    g10778(.A1(new_n13628_), .A2(new_n13776_), .ZN(new_n13809_));
  AOI21_X1   g10779(.A1(new_n13114_), .A2(new_n13776_), .B(new_n13809_), .ZN(new_n13810_));
  NOR4_X1    g10780(.A1(new_n13808_), .A2(new_n13801_), .A3(new_n13792_), .A4(new_n13810_), .ZN(new_n13811_));
  INV_X1     g10781(.I(new_n13808_), .ZN(new_n13812_));
  NOR3_X1    g10782(.A1(new_n13792_), .A2(new_n13801_), .A3(new_n13810_), .ZN(new_n13813_));
  NOR2_X1    g10783(.A1(new_n13813_), .A2(new_n13812_), .ZN(new_n13814_));
  NOR2_X1    g10784(.A1(new_n13814_), .A2(new_n13811_), .ZN(new_n13815_));
  INV_X1     g10785(.I(pi0618), .ZN(new_n13816_));
  INV_X1     g10786(.I(pi1154), .ZN(new_n13817_));
  NOR2_X1    g10787(.A1(new_n13816_), .A2(new_n13817_), .ZN(new_n13818_));
  INV_X1     g10788(.I(new_n13818_), .ZN(new_n13819_));
  AOI21_X1   g10789(.A1(new_n13815_), .A2(pi0618), .B(new_n13819_), .ZN(new_n13820_));
  NOR4_X1    g10790(.A1(new_n13814_), .A2(new_n13816_), .A3(pi1154), .A4(new_n13811_), .ZN(new_n13821_));
  OAI21_X1   g10791(.A1(new_n13820_), .A2(new_n13821_), .B(new_n13629_), .ZN(new_n13822_));
  INV_X1     g10792(.I(pi0627), .ZN(new_n13823_));
  NOR2_X1    g10793(.A1(new_n13823_), .A2(new_n13817_), .ZN(new_n13824_));
  NAND2_X1   g10794(.A1(new_n13822_), .A2(new_n13824_), .ZN(new_n13825_));
  INV_X1     g10795(.I(new_n13825_), .ZN(new_n13826_));
  AOI21_X1   g10796(.A1(new_n13807_), .A2(new_n13826_), .B(pi0618), .ZN(new_n13827_));
  INV_X1     g10797(.I(new_n13827_), .ZN(new_n13828_));
  NAND2_X1   g10798(.A1(new_n13813_), .A2(new_n13812_), .ZN(new_n13829_));
  OR2_X2     g10799(.A1(new_n13810_), .A2(new_n13801_), .Z(new_n13830_));
  OAI21_X1   g10800(.A1(new_n13830_), .A2(new_n13792_), .B(new_n13808_), .ZN(new_n13831_));
  NAND2_X1   g10801(.A1(new_n13831_), .A2(new_n13829_), .ZN(new_n13832_));
  NAND3_X1   g10802(.A1(new_n13832_), .A2(pi0618), .A3(pi1154), .ZN(new_n13833_));
  NAND3_X1   g10803(.A1(new_n13815_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n13834_));
  AOI21_X1   g10804(.A1(new_n13833_), .A2(new_n13834_), .B(new_n13628_), .ZN(new_n13835_));
  NOR2_X1    g10805(.A1(pi0627), .A2(pi1154), .ZN(new_n13836_));
  INV_X1     g10806(.I(new_n13836_), .ZN(new_n13837_));
  NOR2_X1    g10807(.A1(new_n13835_), .A2(new_n13837_), .ZN(new_n13838_));
  OAI21_X1   g10808(.A1(new_n13807_), .A2(new_n13816_), .B(new_n13838_), .ZN(new_n13839_));
  NAND2_X1   g10809(.A1(new_n13839_), .A2(new_n13816_), .ZN(new_n13840_));
  NAND4_X1   g10810(.A1(new_n13800_), .A2(pi0781), .A3(new_n13828_), .A4(new_n13840_), .ZN(new_n13841_));
  INV_X1     g10811(.I(new_n13796_), .ZN(new_n13842_));
  XOR2_X1    g10812(.A1(new_n13737_), .A2(new_n13753_), .Z(new_n13843_));
  INV_X1     g10813(.I(new_n13769_), .ZN(new_n13844_));
  NOR2_X1    g10814(.A1(new_n13768_), .A2(new_n13767_), .ZN(new_n13845_));
  NOR2_X1    g10815(.A1(new_n13844_), .A2(new_n13845_), .ZN(new_n13846_));
  AOI21_X1   g10816(.A1(new_n13846_), .A2(new_n13786_), .B(pi0609), .ZN(new_n13847_));
  OAI21_X1   g10817(.A1(new_n13843_), .A2(new_n13847_), .B(pi0785), .ZN(new_n13848_));
  OAI21_X1   g10818(.A1(new_n13844_), .A2(new_n13845_), .B(pi0609), .ZN(new_n13849_));
  INV_X1     g10819(.I(new_n13794_), .ZN(new_n13850_));
  AOI21_X1   g10820(.A1(new_n13849_), .A2(new_n13850_), .B(pi0609), .ZN(new_n13851_));
  NOR3_X1    g10821(.A1(new_n13843_), .A2(new_n13851_), .A3(new_n13801_), .ZN(new_n13852_));
  NOR2_X1    g10822(.A1(new_n13852_), .A2(new_n13848_), .ZN(new_n13853_));
  OAI21_X1   g10823(.A1(new_n13853_), .A2(new_n13842_), .B(new_n13828_), .ZN(new_n13854_));
  INV_X1     g10824(.I(pi0781), .ZN(new_n13855_));
  AOI21_X1   g10825(.A1(new_n13839_), .A2(new_n13816_), .B(new_n13855_), .ZN(new_n13856_));
  OAI21_X1   g10826(.A1(new_n13853_), .A2(new_n13842_), .B(new_n13856_), .ZN(new_n13857_));
  NAND3_X1   g10827(.A1(new_n13854_), .A2(new_n13857_), .A3(pi0781), .ZN(new_n13858_));
  NAND2_X1   g10828(.A1(new_n13858_), .A2(new_n13841_), .ZN(new_n13859_));
  INV_X1     g10829(.I(pi0619), .ZN(new_n13860_));
  NAND2_X1   g10830(.A1(new_n13822_), .A2(pi0781), .ZN(new_n13861_));
  NOR2_X1    g10831(.A1(new_n13815_), .A2(new_n13855_), .ZN(new_n13862_));
  NAND3_X1   g10832(.A1(new_n13861_), .A2(new_n13835_), .A3(new_n13862_), .ZN(new_n13863_));
  NAND2_X1   g10833(.A1(new_n13835_), .A2(new_n13862_), .ZN(new_n13864_));
  NAND3_X1   g10834(.A1(new_n13864_), .A2(pi0781), .A3(new_n13822_), .ZN(new_n13865_));
  NAND2_X1   g10835(.A1(new_n13865_), .A2(new_n13863_), .ZN(new_n13866_));
  NAND3_X1   g10836(.A1(new_n13866_), .A2(pi0619), .A3(pi1159), .ZN(new_n13867_));
  INV_X1     g10837(.I(pi1159), .ZN(new_n13868_));
  NAND2_X1   g10838(.A1(new_n13833_), .A2(new_n13834_), .ZN(new_n13869_));
  NAND2_X1   g10839(.A1(new_n13869_), .A2(new_n13629_), .ZN(new_n13870_));
  NOR4_X1    g10840(.A1(new_n13870_), .A2(new_n13822_), .A3(new_n13855_), .A4(new_n13815_), .ZN(new_n13871_));
  AOI21_X1   g10841(.A1(new_n13835_), .A2(new_n13862_), .B(new_n13861_), .ZN(new_n13872_));
  NOR2_X1    g10842(.A1(new_n13872_), .A2(new_n13871_), .ZN(new_n13873_));
  NAND3_X1   g10843(.A1(new_n13873_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n13874_));
  AOI21_X1   g10844(.A1(new_n13874_), .A2(new_n13867_), .B(new_n13628_), .ZN(new_n13875_));
  NOR2_X1    g10845(.A1(new_n13817_), .A2(pi0627), .ZN(new_n13876_));
  NOR2_X1    g10846(.A1(new_n13823_), .A2(pi1154), .ZN(new_n13877_));
  NOR2_X1    g10847(.A1(new_n13876_), .A2(new_n13877_), .ZN(new_n13878_));
  NOR2_X1    g10848(.A1(new_n13878_), .A2(new_n13855_), .ZN(new_n13879_));
  INV_X1     g10849(.I(new_n13879_), .ZN(new_n13880_));
  NOR2_X1    g10850(.A1(new_n13629_), .A2(new_n13880_), .ZN(new_n13881_));
  AOI21_X1   g10851(.A1(new_n13807_), .A2(new_n13880_), .B(new_n13881_), .ZN(new_n13882_));
  NAND2_X1   g10852(.A1(new_n13882_), .A2(new_n13860_), .ZN(new_n13883_));
  INV_X1     g10853(.I(pi0648), .ZN(new_n13884_));
  NOR2_X1    g10854(.A1(new_n13884_), .A2(new_n13868_), .ZN(new_n13885_));
  NAND2_X1   g10855(.A1(new_n13883_), .A2(new_n13885_), .ZN(new_n13886_));
  OAI21_X1   g10856(.A1(new_n13875_), .A2(new_n13886_), .B(new_n13860_), .ZN(new_n13887_));
  NAND3_X1   g10857(.A1(new_n13866_), .A2(pi0619), .A3(pi1159), .ZN(new_n13888_));
  NAND4_X1   g10858(.A1(new_n13865_), .A2(new_n13863_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n13889_));
  AOI21_X1   g10859(.A1(new_n13888_), .A2(new_n13889_), .B(new_n13628_), .ZN(new_n13890_));
  NAND2_X1   g10860(.A1(new_n13882_), .A2(pi0619), .ZN(new_n13891_));
  NOR2_X1    g10861(.A1(pi0648), .A2(pi1159), .ZN(new_n13892_));
  NAND2_X1   g10862(.A1(new_n13891_), .A2(new_n13892_), .ZN(new_n13893_));
  OAI21_X1   g10863(.A1(new_n13890_), .A2(new_n13893_), .B(new_n13860_), .ZN(new_n13894_));
  NAND4_X1   g10864(.A1(new_n13859_), .A2(pi0789), .A3(new_n13887_), .A4(new_n13894_), .ZN(new_n13895_));
  INV_X1     g10865(.I(pi0789), .ZN(new_n13896_));
  AOI21_X1   g10866(.A1(new_n13859_), .A2(new_n13887_), .B(new_n13896_), .ZN(new_n13897_));
  NAND3_X1   g10867(.A1(new_n13859_), .A2(pi0789), .A3(new_n13894_), .ZN(new_n13898_));
  NAND2_X1   g10868(.A1(new_n13897_), .A2(new_n13898_), .ZN(new_n13899_));
  NAND2_X1   g10869(.A1(new_n13899_), .A2(new_n13895_), .ZN(new_n13900_));
  INV_X1     g10870(.I(pi0626), .ZN(new_n13901_));
  NAND4_X1   g10871(.A1(new_n13875_), .A2(new_n13890_), .A3(pi0789), .A4(new_n13866_), .ZN(new_n13902_));
  NOR2_X1    g10872(.A1(new_n13860_), .A2(new_n13868_), .ZN(new_n13903_));
  INV_X1     g10873(.I(new_n13903_), .ZN(new_n13904_));
  AOI21_X1   g10874(.A1(new_n13873_), .A2(pi0619), .B(new_n13904_), .ZN(new_n13905_));
  NOR3_X1    g10875(.A1(new_n13866_), .A2(new_n13860_), .A3(new_n13903_), .ZN(new_n13906_));
  OAI21_X1   g10876(.A1(new_n13905_), .A2(new_n13906_), .B(new_n13629_), .ZN(new_n13907_));
  NOR2_X1    g10877(.A1(new_n13873_), .A2(new_n13896_), .ZN(new_n13908_));
  NAND2_X1   g10878(.A1(new_n13890_), .A2(new_n13908_), .ZN(new_n13909_));
  NAND3_X1   g10879(.A1(new_n13909_), .A2(pi0789), .A3(new_n13907_), .ZN(new_n13910_));
  NAND2_X1   g10880(.A1(new_n13910_), .A2(new_n13902_), .ZN(new_n13911_));
  NAND3_X1   g10881(.A1(new_n13911_), .A2(pi0626), .A3(pi1158), .ZN(new_n13912_));
  NAND4_X1   g10882(.A1(new_n13910_), .A2(new_n13901_), .A3(pi1158), .A4(new_n13902_), .ZN(new_n13913_));
  AOI21_X1   g10883(.A1(new_n13912_), .A2(new_n13913_), .B(new_n13628_), .ZN(new_n13914_));
  NOR2_X1    g10884(.A1(new_n13868_), .A2(pi0648), .ZN(new_n13915_));
  NOR2_X1    g10885(.A1(new_n13884_), .A2(pi1159), .ZN(new_n13916_));
  NOR2_X1    g10886(.A1(new_n13915_), .A2(new_n13916_), .ZN(new_n13917_));
  NOR2_X1    g10887(.A1(new_n13917_), .A2(new_n13896_), .ZN(new_n13918_));
  INV_X1     g10888(.I(new_n13918_), .ZN(new_n13919_));
  NOR2_X1    g10889(.A1(new_n13628_), .A2(new_n13919_), .ZN(new_n13920_));
  AOI21_X1   g10890(.A1(new_n13882_), .A2(new_n13919_), .B(new_n13920_), .ZN(new_n13921_));
  INV_X1     g10891(.I(pi0641), .ZN(new_n13922_));
  NOR2_X1    g10892(.A1(new_n13922_), .A2(pi1158), .ZN(new_n13923_));
  INV_X1     g10893(.I(new_n13923_), .ZN(new_n13924_));
  AOI21_X1   g10894(.A1(new_n13921_), .A2(new_n13901_), .B(new_n13924_), .ZN(new_n13925_));
  INV_X1     g10895(.I(new_n13925_), .ZN(new_n13926_));
  OAI21_X1   g10896(.A1(new_n13914_), .A2(new_n13926_), .B(new_n13901_), .ZN(new_n13927_));
  NAND3_X1   g10897(.A1(new_n13911_), .A2(pi0626), .A3(pi1158), .ZN(new_n13928_));
  INV_X1     g10898(.I(pi1158), .ZN(new_n13929_));
  NAND4_X1   g10899(.A1(new_n13910_), .A2(pi0626), .A3(new_n13929_), .A4(new_n13902_), .ZN(new_n13930_));
  AOI21_X1   g10900(.A1(new_n13928_), .A2(new_n13930_), .B(new_n13628_), .ZN(new_n13931_));
  AND2_X2    g10901(.A1(new_n13882_), .A2(new_n13919_), .Z(new_n13932_));
  NAND4_X1   g10902(.A1(new_n13927_), .A2(new_n13900_), .A3(pi0626), .A4(pi0788), .ZN(new_n13936_));
  INV_X1     g10903(.I(pi0788), .ZN(new_n13937_));
  AOI21_X1   g10904(.A1(new_n13927_), .A2(new_n13900_), .B(new_n13937_), .ZN(new_n13938_));
  NAND3_X1   g10905(.A1(new_n13900_), .A2(pi0626), .A3(pi0788), .ZN(new_n13939_));
  NAND2_X1   g10906(.A1(new_n13938_), .A2(new_n13939_), .ZN(new_n13940_));
  NAND2_X1   g10907(.A1(new_n13940_), .A2(new_n13936_), .ZN(new_n13941_));
  INV_X1     g10908(.I(pi0628), .ZN(new_n13942_));
  NAND4_X1   g10909(.A1(new_n13914_), .A2(new_n13931_), .A3(pi0788), .A4(new_n13911_), .ZN(new_n13943_));
  AOI21_X1   g10910(.A1(new_n13873_), .A2(pi1159), .B(new_n13904_), .ZN(new_n13944_));
  INV_X1     g10911(.I(new_n13889_), .ZN(new_n13945_));
  OAI21_X1   g10912(.A1(new_n13944_), .A2(new_n13945_), .B(new_n13629_), .ZN(new_n13946_));
  NOR4_X1    g10913(.A1(new_n13946_), .A2(new_n13907_), .A3(new_n13896_), .A4(new_n13873_), .ZN(new_n13947_));
  NAND2_X1   g10914(.A1(new_n13907_), .A2(pi0789), .ZN(new_n13948_));
  INV_X1     g10915(.I(new_n13908_), .ZN(new_n13949_));
  NOR2_X1    g10916(.A1(new_n13946_), .A2(new_n13949_), .ZN(new_n13950_));
  NOR2_X1    g10917(.A1(new_n13950_), .A2(new_n13948_), .ZN(new_n13951_));
  NOR2_X1    g10918(.A1(new_n13951_), .A2(new_n13947_), .ZN(new_n13952_));
  NOR2_X1    g10919(.A1(new_n13901_), .A2(new_n13929_), .ZN(new_n13953_));
  INV_X1     g10920(.I(new_n13953_), .ZN(new_n13954_));
  AOI21_X1   g10921(.A1(new_n13952_), .A2(pi1158), .B(new_n13954_), .ZN(new_n13955_));
  INV_X1     g10922(.I(new_n13913_), .ZN(new_n13956_));
  OAI21_X1   g10923(.A1(new_n13955_), .A2(new_n13956_), .B(new_n13629_), .ZN(new_n13957_));
  NOR2_X1    g10924(.A1(new_n13952_), .A2(new_n13937_), .ZN(new_n13958_));
  NAND2_X1   g10925(.A1(new_n13931_), .A2(new_n13958_), .ZN(new_n13959_));
  NAND3_X1   g10926(.A1(new_n13959_), .A2(pi0788), .A3(new_n13957_), .ZN(new_n13960_));
  NAND2_X1   g10927(.A1(new_n13960_), .A2(new_n13943_), .ZN(new_n13961_));
  NOR2_X1    g10928(.A1(new_n13929_), .A2(pi0641), .ZN(new_n13962_));
  NOR2_X1    g10929(.A1(new_n13922_), .A2(pi1158), .ZN(new_n13963_));
  NOR2_X1    g10930(.A1(new_n13962_), .A2(new_n13963_), .ZN(new_n13964_));
  NOR2_X1    g10931(.A1(new_n13964_), .A2(new_n13937_), .ZN(new_n13965_));
  INV_X1     g10932(.I(new_n13965_), .ZN(new_n13966_));
  NOR2_X1    g10933(.A1(new_n13629_), .A2(new_n13966_), .ZN(new_n13967_));
  AOI21_X1   g10934(.A1(new_n13921_), .A2(new_n13966_), .B(new_n13967_), .ZN(new_n13968_));
  INV_X1     g10935(.I(pi1156), .ZN(new_n13969_));
  NOR2_X1    g10936(.A1(new_n13942_), .A2(new_n13969_), .ZN(new_n13970_));
  INV_X1     g10937(.I(new_n13970_), .ZN(new_n13971_));
  AOI21_X1   g10938(.A1(new_n13968_), .A2(pi0628), .B(new_n13971_), .ZN(new_n13972_));
  NOR3_X1    g10939(.A1(new_n13932_), .A2(new_n13920_), .A3(new_n13965_), .ZN(new_n13973_));
  NOR4_X1    g10940(.A1(new_n13973_), .A2(new_n13942_), .A3(pi1156), .A4(new_n13967_), .ZN(new_n13974_));
  OAI21_X1   g10941(.A1(new_n13974_), .A2(new_n13972_), .B(new_n13629_), .ZN(new_n13975_));
  INV_X1     g10942(.I(pi0629), .ZN(new_n13976_));
  NOR2_X1    g10943(.A1(new_n13976_), .A2(new_n13969_), .ZN(new_n13977_));
  AND2_X2    g10944(.A1(new_n13975_), .A2(new_n13977_), .Z(new_n13978_));
  INV_X1     g10945(.I(new_n13978_), .ZN(new_n13979_));
  OAI21_X1   g10946(.A1(new_n13961_), .A2(new_n13979_), .B(new_n13942_), .ZN(new_n13980_));
  AOI21_X1   g10947(.A1(new_n13941_), .A2(new_n13980_), .B(new_n12777_), .ZN(new_n13981_));
  AOI21_X1   g10948(.A1(new_n13968_), .A2(pi1156), .B(new_n13971_), .ZN(new_n13982_));
  NOR4_X1    g10949(.A1(new_n13973_), .A2(pi0628), .A3(new_n13969_), .A4(new_n13967_), .ZN(new_n13983_));
  OAI21_X1   g10950(.A1(new_n13983_), .A2(new_n13982_), .B(new_n13629_), .ZN(new_n13984_));
  NOR2_X1    g10951(.A1(pi0629), .A2(pi1156), .ZN(new_n13985_));
  NAND3_X1   g10952(.A1(new_n13941_), .A2(pi0628), .A3(pi0792), .ZN(new_n13988_));
  XOR2_X1    g10953(.A1(new_n13981_), .A2(new_n13988_), .Z(new_n13989_));
  NOR2_X1    g10954(.A1(new_n13969_), .A2(pi0629), .ZN(new_n13990_));
  NOR2_X1    g10955(.A1(new_n13976_), .A2(pi1156), .ZN(new_n13991_));
  NOR2_X1    g10956(.A1(new_n13990_), .A2(new_n13991_), .ZN(new_n13992_));
  NOR2_X1    g10957(.A1(new_n13992_), .A2(new_n12777_), .ZN(new_n13993_));
  INV_X1     g10958(.I(new_n13993_), .ZN(new_n13994_));
  NOR2_X1    g10959(.A1(new_n13629_), .A2(new_n13994_), .ZN(new_n13995_));
  INV_X1     g10960(.I(new_n13995_), .ZN(new_n13996_));
  NAND3_X1   g10961(.A1(new_n13960_), .A2(new_n13943_), .A3(new_n13994_), .ZN(new_n13997_));
  NAND2_X1   g10962(.A1(new_n13997_), .A2(new_n13996_), .ZN(new_n13998_));
  NOR4_X1    g10963(.A1(new_n13975_), .A2(new_n13984_), .A3(new_n12777_), .A4(new_n13968_), .ZN(new_n13999_));
  NAND2_X1   g10964(.A1(new_n13975_), .A2(pi0792), .ZN(new_n14000_));
  NOR3_X1    g10965(.A1(new_n13984_), .A2(new_n12777_), .A3(new_n13968_), .ZN(new_n14001_));
  NOR2_X1    g10966(.A1(new_n14001_), .A2(new_n14000_), .ZN(new_n14002_));
  NOR2_X1    g10967(.A1(new_n14002_), .A2(new_n13999_), .ZN(new_n14003_));
  NAND2_X1   g10968(.A1(new_n14003_), .A2(pi0647), .ZN(new_n14004_));
  INV_X1     g10969(.I(pi0647), .ZN(new_n14005_));
  INV_X1     g10970(.I(pi1157), .ZN(new_n14006_));
  NOR2_X1    g10971(.A1(new_n14005_), .A2(new_n14006_), .ZN(new_n14007_));
  INV_X1     g10972(.I(new_n14007_), .ZN(new_n14008_));
  XOR2_X1    g10973(.A1(new_n14004_), .A2(new_n14008_), .Z(new_n14009_));
  INV_X1     g10974(.I(pi0630), .ZN(new_n14010_));
  NOR2_X1    g10975(.A1(new_n14010_), .A2(new_n14006_), .ZN(new_n14011_));
  INV_X1     g10976(.I(new_n14011_), .ZN(new_n14012_));
  AOI21_X1   g10977(.A1(new_n14009_), .A2(new_n13629_), .B(new_n14012_), .ZN(new_n14013_));
  AOI21_X1   g10978(.A1(new_n14013_), .A2(new_n13998_), .B(pi0647), .ZN(new_n14014_));
  INV_X1     g10979(.I(new_n13943_), .ZN(new_n14015_));
  NAND2_X1   g10980(.A1(new_n13957_), .A2(pi0788), .ZN(new_n14016_));
  AOI21_X1   g10981(.A1(new_n13952_), .A2(pi0626), .B(new_n13954_), .ZN(new_n14017_));
  INV_X1     g10982(.I(new_n13930_), .ZN(new_n14018_));
  OAI21_X1   g10983(.A1(new_n14017_), .A2(new_n14018_), .B(new_n13629_), .ZN(new_n14019_));
  NOR3_X1    g10984(.A1(new_n14019_), .A2(new_n13937_), .A3(new_n13952_), .ZN(new_n14020_));
  NOR2_X1    g10985(.A1(new_n14020_), .A2(new_n14016_), .ZN(new_n14021_));
  NOR3_X1    g10986(.A1(new_n14021_), .A2(new_n14015_), .A3(new_n13993_), .ZN(new_n14022_));
  NOR3_X1    g10987(.A1(new_n14022_), .A2(new_n14005_), .A3(new_n13995_), .ZN(new_n14023_));
  AOI21_X1   g10988(.A1(new_n14003_), .A2(pi1157), .B(new_n14008_), .ZN(new_n14024_));
  NOR4_X1    g10989(.A1(new_n14002_), .A2(pi0647), .A3(new_n14006_), .A4(new_n13999_), .ZN(new_n14025_));
  OAI21_X1   g10990(.A1(new_n14024_), .A2(new_n14025_), .B(new_n13629_), .ZN(new_n14026_));
  NOR2_X1    g10991(.A1(pi0630), .A2(pi1157), .ZN(new_n14027_));
  NAND2_X1   g10992(.A1(new_n14026_), .A2(new_n14027_), .ZN(new_n14028_));
  OAI21_X1   g10993(.A1(new_n14023_), .A2(new_n14028_), .B(new_n14005_), .ZN(new_n14029_));
  INV_X1     g10994(.I(new_n14029_), .ZN(new_n14030_));
  NOR4_X1    g10995(.A1(new_n13989_), .A2(new_n12776_), .A3(new_n14014_), .A4(new_n14030_), .ZN(new_n14031_));
  NAND4_X1   g10996(.A1(new_n13941_), .A2(new_n13980_), .A3(pi0628), .A4(pi0792), .ZN(new_n14032_));
  NAND2_X1   g10997(.A1(new_n13981_), .A2(new_n13988_), .ZN(new_n14033_));
  AOI21_X1   g10998(.A1(new_n14033_), .A2(new_n14032_), .B(new_n14014_), .ZN(new_n14034_));
  NAND2_X1   g10999(.A1(new_n14029_), .A2(pi0787), .ZN(new_n14035_));
  AOI21_X1   g11000(.A1(new_n14032_), .A2(new_n14033_), .B(new_n14035_), .ZN(new_n14036_));
  NOR3_X1    g11001(.A1(new_n14036_), .A2(new_n14034_), .A3(new_n12776_), .ZN(new_n14037_));
  OAI21_X1   g11002(.A1(new_n14037_), .A2(new_n14031_), .B(new_n12775_), .ZN(new_n14038_));
  NOR2_X1    g11003(.A1(new_n9992_), .A2(pi0140), .ZN(new_n14039_));
  AOI21_X1   g11004(.A1(new_n13218_), .A2(new_n13226_), .B(new_n14039_), .ZN(new_n14040_));
  INV_X1     g11005(.I(new_n14040_), .ZN(new_n14041_));
  NOR3_X1    g11006(.A1(new_n13219_), .A2(pi0625), .A3(pi0738), .ZN(new_n14042_));
  NAND3_X1   g11007(.A1(new_n14041_), .A2(new_n14042_), .A3(new_n14039_), .ZN(new_n14043_));
  NOR3_X1    g11008(.A1(new_n14042_), .A2(new_n13614_), .A3(new_n14040_), .ZN(new_n14044_));
  XOR2_X1    g11009(.A1(new_n14043_), .A2(new_n14044_), .Z(new_n14045_));
  NAND2_X1   g11010(.A1(new_n14041_), .A2(new_n13748_), .ZN(new_n14046_));
  OAI21_X1   g11011(.A1(new_n14045_), .A2(new_n13748_), .B(new_n14046_), .ZN(new_n14047_));
  NOR2_X1    g11012(.A1(new_n13805_), .A2(new_n2723_), .ZN(new_n14048_));
  INV_X1     g11013(.I(new_n14048_), .ZN(new_n14049_));
  NAND2_X1   g11014(.A1(new_n14047_), .A2(new_n14049_), .ZN(new_n14050_));
  NOR2_X1    g11015(.A1(new_n13880_), .A2(new_n2723_), .ZN(new_n14051_));
  NOR2_X1    g11016(.A1(new_n14050_), .A2(new_n14051_), .ZN(new_n14052_));
  NAND2_X1   g11017(.A1(new_n14052_), .A2(new_n9992_), .ZN(new_n14053_));
  AOI21_X1   g11018(.A1(new_n14053_), .A2(new_n13966_), .B(new_n13919_), .ZN(new_n14054_));
  NOR2_X1    g11019(.A1(new_n13969_), .A2(pi0628), .ZN(new_n14055_));
  NOR2_X1    g11020(.A1(new_n13942_), .A2(pi1156), .ZN(new_n14056_));
  NOR2_X1    g11021(.A1(new_n14055_), .A2(new_n14056_), .ZN(new_n14057_));
  NOR2_X1    g11022(.A1(new_n14057_), .A2(new_n12777_), .ZN(new_n14058_));
  INV_X1     g11023(.I(new_n14058_), .ZN(new_n14059_));
  NOR2_X1    g11024(.A1(new_n14059_), .A2(new_n2723_), .ZN(new_n14060_));
  INV_X1     g11025(.I(new_n14060_), .ZN(new_n14061_));
  NAND2_X1   g11026(.A1(new_n14054_), .A2(new_n14061_), .ZN(new_n14062_));
  NAND2_X1   g11027(.A1(new_n14062_), .A2(pi0647), .ZN(new_n14063_));
  XOR2_X1    g11028(.A1(new_n14063_), .A2(new_n14008_), .Z(new_n14064_));
  NAND2_X1   g11029(.A1(new_n14064_), .A2(new_n14039_), .ZN(new_n14065_));
  NAND2_X1   g11030(.A1(new_n14065_), .A2(pi0787), .ZN(new_n14066_));
  NAND2_X1   g11031(.A1(new_n14062_), .A2(pi1157), .ZN(new_n14067_));
  XOR2_X1    g11032(.A1(new_n14067_), .A2(new_n14008_), .Z(new_n14068_));
  NAND2_X1   g11033(.A1(new_n14068_), .A2(new_n14039_), .ZN(new_n14069_));
  NOR3_X1    g11034(.A1(new_n14069_), .A2(new_n12776_), .A3(new_n14062_), .ZN(new_n14070_));
  XOR2_X1    g11035(.A1(new_n14070_), .A2(new_n14066_), .Z(new_n14071_));
  INV_X1     g11036(.I(new_n14052_), .ZN(new_n14072_));
  NOR3_X1    g11037(.A1(new_n14040_), .A2(new_n13613_), .A3(new_n13203_), .ZN(new_n14073_));
  INV_X1     g11038(.I(new_n14039_), .ZN(new_n14074_));
  NAND2_X1   g11039(.A1(new_n14074_), .A2(new_n13614_), .ZN(new_n14075_));
  OAI21_X1   g11040(.A1(new_n14042_), .A2(new_n14075_), .B(pi0608), .ZN(new_n14076_));
  OAI21_X1   g11041(.A1(new_n13105_), .A2(pi0761), .B(new_n14074_), .ZN(new_n14077_));
  NAND3_X1   g11042(.A1(new_n14076_), .A2(new_n13614_), .A3(new_n14077_), .ZN(new_n14078_));
  AOI21_X1   g11043(.A1(new_n14078_), .A2(new_n14073_), .B(new_n13748_), .ZN(new_n14079_));
  NOR2_X1    g11044(.A1(new_n14040_), .A2(new_n13203_), .ZN(new_n14080_));
  INV_X1     g11045(.I(pi0608), .ZN(new_n14081_));
  NOR2_X1    g11046(.A1(new_n14081_), .A2(new_n13614_), .ZN(new_n14082_));
  INV_X1     g11047(.I(new_n14082_), .ZN(new_n14083_));
  NAND2_X1   g11048(.A1(new_n14041_), .A2(new_n14083_), .ZN(new_n14084_));
  NOR4_X1    g11049(.A1(new_n14075_), .A2(pi0625), .A3(pi0738), .A4(new_n13219_), .ZN(new_n14085_));
  AOI21_X1   g11050(.A1(new_n14084_), .A2(new_n14085_), .B(new_n14073_), .ZN(new_n14086_));
  NOR4_X1    g11051(.A1(new_n14086_), .A2(new_n13748_), .A3(new_n14080_), .A4(new_n14077_), .ZN(new_n14087_));
  XOR2_X1    g11052(.A1(new_n14087_), .A2(new_n14079_), .Z(new_n14088_));
  NAND2_X1   g11053(.A1(new_n14088_), .A2(new_n13801_), .ZN(new_n14089_));
  NOR2_X1    g11054(.A1(new_n13766_), .A2(new_n13778_), .ZN(new_n14090_));
  NOR2_X1    g11055(.A1(new_n14088_), .A2(new_n13778_), .ZN(new_n14091_));
  XOR2_X1    g11056(.A1(new_n14091_), .A2(new_n14090_), .Z(new_n14092_));
  NAND2_X1   g11057(.A1(new_n14092_), .A2(new_n14047_), .ZN(new_n14093_));
  NAND2_X1   g11058(.A1(new_n9992_), .A2(pi0609), .ZN(new_n14094_));
  INV_X1     g11059(.I(new_n14077_), .ZN(new_n14095_));
  NOR2_X1    g11060(.A1(new_n13776_), .A2(new_n2723_), .ZN(new_n14096_));
  NOR2_X1    g11061(.A1(new_n14095_), .A2(new_n14096_), .ZN(new_n14097_));
  AOI21_X1   g11062(.A1(new_n14097_), .A2(new_n14094_), .B(pi1155), .ZN(new_n14098_));
  NOR2_X1    g11063(.A1(new_n14098_), .A2(new_n13783_), .ZN(new_n14099_));
  NAND2_X1   g11064(.A1(new_n14093_), .A2(new_n14099_), .ZN(new_n14100_));
  NOR2_X1    g11065(.A1(new_n13775_), .A2(new_n13766_), .ZN(new_n14101_));
  INV_X1     g11066(.I(new_n14101_), .ZN(new_n14102_));
  NAND2_X1   g11067(.A1(new_n14095_), .A2(pi1155), .ZN(new_n14103_));
  AOI21_X1   g11068(.A1(new_n14103_), .A2(new_n2723_), .B(new_n14102_), .ZN(new_n14104_));
  NOR2_X1    g11069(.A1(new_n14104_), .A2(pi0660), .ZN(new_n14105_));
  NAND2_X1   g11070(.A1(new_n14100_), .A2(new_n14105_), .ZN(new_n14106_));
  NOR2_X1    g11071(.A1(new_n14088_), .A2(new_n13766_), .ZN(new_n14107_));
  XOR2_X1    g11072(.A1(new_n14107_), .A2(new_n14090_), .Z(new_n14108_));
  NAND4_X1   g11073(.A1(new_n14106_), .A2(pi0785), .A3(new_n14047_), .A4(new_n14108_), .ZN(new_n14109_));
  NAND2_X1   g11074(.A1(new_n14109_), .A2(new_n14089_), .ZN(new_n14110_));
  NAND2_X1   g11075(.A1(new_n14110_), .A2(new_n13855_), .ZN(new_n14111_));
  NOR2_X1    g11076(.A1(new_n14110_), .A2(new_n13816_), .ZN(new_n14112_));
  XOR2_X1    g11077(.A1(new_n14112_), .A2(new_n13818_), .Z(new_n14113_));
  NAND3_X1   g11078(.A1(new_n14113_), .A2(new_n14047_), .A3(new_n14049_), .ZN(new_n14114_));
  NOR2_X1    g11079(.A1(new_n14098_), .A2(new_n13801_), .ZN(new_n14115_));
  NAND3_X1   g11080(.A1(new_n14104_), .A2(pi0785), .A3(new_n14097_), .ZN(new_n14116_));
  XOR2_X1    g11081(.A1(new_n14116_), .A2(new_n14115_), .Z(new_n14117_));
  NOR2_X1    g11082(.A1(new_n14117_), .A2(new_n13817_), .ZN(new_n14118_));
  OAI21_X1   g11083(.A1(new_n14118_), .A2(new_n9992_), .B(pi0618), .ZN(new_n14119_));
  NAND3_X1   g11084(.A1(new_n14114_), .A2(new_n13823_), .A3(new_n14119_), .ZN(new_n14120_));
  OAI21_X1   g11085(.A1(new_n14118_), .A2(pi0618), .B(new_n9992_), .ZN(new_n14121_));
  NAND3_X1   g11086(.A1(new_n14120_), .A2(new_n13823_), .A3(new_n14121_), .ZN(new_n14122_));
  NOR2_X1    g11087(.A1(new_n14110_), .A2(new_n13817_), .ZN(new_n14123_));
  XOR2_X1    g11088(.A1(new_n14123_), .A2(new_n13819_), .Z(new_n14124_));
  NOR3_X1    g11089(.A1(new_n14124_), .A2(new_n13855_), .A3(new_n14050_), .ZN(new_n14125_));
  NAND2_X1   g11090(.A1(new_n14122_), .A2(new_n14125_), .ZN(new_n14126_));
  NAND2_X1   g11091(.A1(new_n14126_), .A2(new_n14111_), .ZN(new_n14127_));
  NOR2_X1    g11092(.A1(new_n14127_), .A2(new_n13860_), .ZN(new_n14128_));
  XOR2_X1    g11093(.A1(new_n14128_), .A2(new_n13904_), .Z(new_n14129_));
  NOR2_X1    g11094(.A1(new_n14129_), .A2(new_n14072_), .ZN(new_n14130_));
  NAND2_X1   g11095(.A1(new_n14121_), .A2(pi0781), .ZN(new_n14131_));
  NOR3_X1    g11096(.A1(new_n14119_), .A2(new_n13855_), .A3(new_n14117_), .ZN(new_n14132_));
  XOR2_X1    g11097(.A1(new_n14132_), .A2(new_n14131_), .Z(new_n14133_));
  NAND2_X1   g11098(.A1(new_n14133_), .A2(pi1159), .ZN(new_n14134_));
  XOR2_X1    g11099(.A1(new_n14134_), .A2(new_n13904_), .Z(new_n14135_));
  NAND2_X1   g11100(.A1(new_n14135_), .A2(new_n14039_), .ZN(new_n14136_));
  NAND2_X1   g11101(.A1(new_n14136_), .A2(new_n13884_), .ZN(new_n14137_));
  INV_X1     g11102(.I(new_n14127_), .ZN(new_n14138_));
  NOR2_X1    g11103(.A1(new_n13929_), .A2(pi0626), .ZN(new_n14139_));
  NOR2_X1    g11104(.A1(new_n13901_), .A2(pi1158), .ZN(new_n14140_));
  NOR2_X1    g11105(.A1(new_n14139_), .A2(new_n14140_), .ZN(new_n14141_));
  NOR2_X1    g11106(.A1(new_n14141_), .A2(new_n13937_), .ZN(new_n14142_));
  NOR2_X1    g11107(.A1(new_n13965_), .A2(new_n14142_), .ZN(new_n14143_));
  AOI21_X1   g11108(.A1(new_n14138_), .A2(new_n14143_), .B(pi0789), .ZN(new_n14144_));
  OAI21_X1   g11109(.A1(new_n14130_), .A2(new_n14137_), .B(new_n14144_), .ZN(new_n14145_));
  NOR2_X1    g11110(.A1(new_n14127_), .A2(new_n13868_), .ZN(new_n14146_));
  XOR2_X1    g11111(.A1(new_n14146_), .A2(new_n13903_), .Z(new_n14147_));
  NAND2_X1   g11112(.A1(new_n14147_), .A2(new_n14052_), .ZN(new_n14148_));
  NAND2_X1   g11113(.A1(new_n14133_), .A2(pi0619), .ZN(new_n14149_));
  XOR2_X1    g11114(.A1(new_n14149_), .A2(new_n13904_), .Z(new_n14150_));
  NAND2_X1   g11115(.A1(new_n14150_), .A2(new_n14039_), .ZN(new_n14151_));
  NAND4_X1   g11116(.A1(new_n14145_), .A2(pi0648), .A3(new_n14148_), .A4(new_n14151_), .ZN(new_n14152_));
  INV_X1     g11117(.I(new_n14141_), .ZN(new_n14153_));
  NAND2_X1   g11118(.A1(new_n14151_), .A2(pi0789), .ZN(new_n14154_));
  NOR3_X1    g11119(.A1(new_n14136_), .A2(new_n13896_), .A3(new_n14133_), .ZN(new_n14155_));
  XOR2_X1    g11120(.A1(new_n14155_), .A2(new_n14154_), .Z(new_n14156_));
  NAND2_X1   g11121(.A1(new_n14156_), .A2(new_n14153_), .ZN(new_n14157_));
  NAND2_X1   g11122(.A1(new_n14153_), .A2(new_n14039_), .ZN(new_n14158_));
  XOR2_X1    g11123(.A1(new_n14157_), .A2(new_n14158_), .Z(new_n14159_));
  NOR2_X1    g11124(.A1(pi0641), .A2(pi1158), .ZN(new_n14160_));
  NOR3_X1    g11125(.A1(new_n13922_), .A2(new_n13929_), .A3(pi0626), .ZN(new_n14161_));
  AOI21_X1   g11126(.A1(pi0626), .A2(new_n14160_), .B(new_n14161_), .ZN(new_n14162_));
  NOR2_X1    g11127(.A1(new_n13919_), .A2(new_n2723_), .ZN(new_n14163_));
  INV_X1     g11128(.I(new_n14163_), .ZN(new_n14164_));
  AOI21_X1   g11129(.A1(new_n14072_), .A2(new_n14162_), .B(new_n14164_), .ZN(new_n14165_));
  AOI21_X1   g11130(.A1(new_n14165_), .A2(new_n13929_), .B(pi0641), .ZN(new_n14166_));
  OAI21_X1   g11131(.A1(new_n13929_), .A2(new_n14165_), .B(new_n14166_), .ZN(new_n14167_));
  NAND2_X1   g11132(.A1(new_n14159_), .A2(new_n14167_), .ZN(new_n14168_));
  NAND2_X1   g11133(.A1(new_n14168_), .A2(pi0788), .ZN(new_n14169_));
  NAND2_X1   g11134(.A1(new_n14152_), .A2(new_n14169_), .ZN(new_n14170_));
  NOR2_X1    g11135(.A1(new_n14170_), .A2(pi0792), .ZN(new_n14171_));
  NAND2_X1   g11136(.A1(new_n14170_), .A2(pi1156), .ZN(new_n14172_));
  XOR2_X1    g11137(.A1(new_n14172_), .A2(new_n13971_), .Z(new_n14173_));
  NAND2_X1   g11138(.A1(new_n14159_), .A2(pi0788), .ZN(new_n14174_));
  OAI21_X1   g11139(.A1(pi0788), .A2(new_n14156_), .B(new_n14174_), .ZN(new_n14175_));
  NOR2_X1    g11140(.A1(new_n2723_), .A2(pi0628), .ZN(new_n14176_));
  OR2_X2     g11141(.A1(new_n14054_), .A2(new_n13977_), .Z(new_n14177_));
  NAND4_X1   g11142(.A1(new_n14173_), .A2(new_n14175_), .A3(new_n14176_), .A4(new_n14177_), .ZN(new_n14178_));
  NAND2_X1   g11143(.A1(new_n14170_), .A2(pi0628), .ZN(new_n14179_));
  XOR2_X1    g11144(.A1(new_n14179_), .A2(new_n13971_), .Z(new_n14180_));
  NOR2_X1    g11145(.A1(new_n2723_), .A2(new_n13942_), .ZN(new_n14181_));
  NAND4_X1   g11146(.A1(new_n14180_), .A2(new_n14175_), .A3(new_n14177_), .A4(new_n14181_), .ZN(new_n14182_));
  AOI21_X1   g11147(.A1(new_n14178_), .A2(new_n14182_), .B(new_n12777_), .ZN(new_n14183_));
  OAI21_X1   g11148(.A1(new_n14183_), .A2(new_n14171_), .B(new_n12776_), .ZN(new_n14184_));
  NOR2_X1    g11149(.A1(new_n14175_), .A2(new_n13993_), .ZN(new_n14185_));
  AOI21_X1   g11150(.A1(new_n13993_), .A2(new_n14074_), .B(new_n14185_), .ZN(new_n14186_));
  NOR2_X1    g11151(.A1(new_n14183_), .A2(new_n14171_), .ZN(new_n14187_));
  NAND2_X1   g11152(.A1(new_n14187_), .A2(pi1157), .ZN(new_n14188_));
  XOR2_X1    g11153(.A1(new_n14188_), .A2(new_n14007_), .Z(new_n14189_));
  NOR2_X1    g11154(.A1(new_n14189_), .A2(new_n14186_), .ZN(new_n14190_));
  NAND2_X1   g11155(.A1(new_n14065_), .A2(pi0630), .ZN(new_n14191_));
  NOR2_X1    g11156(.A1(new_n14190_), .A2(new_n14191_), .ZN(new_n14192_));
  NAND2_X1   g11157(.A1(new_n14069_), .A2(new_n14010_), .ZN(new_n14193_));
  NAND2_X1   g11158(.A1(new_n14187_), .A2(pi0647), .ZN(new_n14194_));
  XOR2_X1    g11159(.A1(new_n14194_), .A2(new_n14007_), .Z(new_n14195_));
  NOR3_X1    g11160(.A1(new_n14195_), .A2(new_n12776_), .A3(new_n14186_), .ZN(new_n14196_));
  OAI21_X1   g11161(.A1(new_n14192_), .A2(new_n14193_), .B(new_n14196_), .ZN(new_n14197_));
  NAND2_X1   g11162(.A1(new_n14197_), .A2(new_n14184_), .ZN(new_n14198_));
  NAND3_X1   g11163(.A1(new_n14198_), .A2(pi0644), .A3(pi0715), .ZN(new_n14199_));
  INV_X1     g11164(.I(pi0715), .ZN(new_n14200_));
  NAND4_X1   g11165(.A1(new_n14197_), .A2(pi0644), .A3(new_n14200_), .A4(new_n14184_), .ZN(new_n14201_));
  AOI21_X1   g11166(.A1(new_n14199_), .A2(new_n14201_), .B(new_n14071_), .ZN(new_n14202_));
  INV_X1     g11167(.I(pi1160), .ZN(new_n14203_));
  INV_X1     g11168(.I(pi0644), .ZN(new_n14204_));
  NOR2_X1    g11169(.A1(new_n14204_), .A2(new_n14200_), .ZN(new_n14205_));
  NOR2_X1    g11170(.A1(new_n14006_), .A2(pi0630), .ZN(new_n14206_));
  INV_X1     g11171(.I(new_n14206_), .ZN(new_n14207_));
  NOR2_X1    g11172(.A1(new_n14010_), .A2(pi1157), .ZN(new_n14208_));
  INV_X1     g11173(.I(new_n14208_), .ZN(new_n14209_));
  AOI21_X1   g11174(.A1(new_n14207_), .A2(new_n14209_), .B(new_n12776_), .ZN(new_n14210_));
  INV_X1     g11175(.I(new_n14210_), .ZN(new_n14211_));
  NOR2_X1    g11176(.A1(new_n14211_), .A2(new_n14074_), .ZN(new_n14212_));
  AOI21_X1   g11177(.A1(new_n14186_), .A2(new_n14211_), .B(new_n14212_), .ZN(new_n14213_));
  NAND2_X1   g11178(.A1(new_n14213_), .A2(pi0715), .ZN(new_n14214_));
  XOR2_X1    g11179(.A1(new_n14214_), .A2(new_n14205_), .Z(new_n14215_));
  OAI21_X1   g11180(.A1(new_n14215_), .A2(new_n14074_), .B(new_n14203_), .ZN(new_n14216_));
  INV_X1     g11181(.I(new_n14205_), .ZN(new_n14217_));
  NAND2_X1   g11182(.A1(new_n14213_), .A2(pi0644), .ZN(new_n14218_));
  XOR2_X1    g11183(.A1(new_n14218_), .A2(new_n14217_), .Z(new_n14219_));
  AOI21_X1   g11184(.A1(new_n14219_), .A2(new_n14039_), .B(pi1160), .ZN(new_n14220_));
  OAI21_X1   g11185(.A1(new_n14202_), .A2(new_n14216_), .B(new_n14220_), .ZN(new_n14221_));
  NAND3_X1   g11186(.A1(new_n14198_), .A2(pi0644), .A3(pi0715), .ZN(new_n14222_));
  NAND4_X1   g11187(.A1(new_n14197_), .A2(new_n14204_), .A3(pi0715), .A4(new_n14184_), .ZN(new_n14223_));
  AOI21_X1   g11188(.A1(new_n14222_), .A2(new_n14223_), .B(new_n14071_), .ZN(new_n14224_));
  NAND4_X1   g11189(.A1(new_n14221_), .A2(pi0790), .A3(new_n14224_), .A4(pi0832), .ZN(new_n14225_));
  NAND2_X1   g11190(.A1(new_n14221_), .A2(new_n14224_), .ZN(new_n14226_));
  NAND3_X1   g11191(.A1(new_n14226_), .A2(new_n12775_), .A3(pi0832), .ZN(new_n14227_));
  AOI21_X1   g11192(.A1(po1038), .A2(new_n7971_), .B(pi0832), .ZN(new_n14228_));
  NAND2_X1   g11193(.A1(new_n14198_), .A2(new_n14228_), .ZN(new_n14229_));
  AOI21_X1   g11194(.A1(new_n14227_), .A2(new_n14225_), .B(new_n14229_), .ZN(new_n14230_));
  AOI21_X1   g11195(.A1(new_n14038_), .A2(new_n7240_), .B(new_n14230_), .ZN(new_n14231_));
  NOR2_X1    g11196(.A1(new_n14037_), .A2(new_n14031_), .ZN(new_n14232_));
  AOI21_X1   g11197(.A1(new_n14232_), .A2(pi0715), .B(new_n14217_), .ZN(new_n14233_));
  NOR4_X1    g11198(.A1(new_n14037_), .A2(new_n14031_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n14234_));
  NOR2_X1    g11199(.A1(new_n14233_), .A2(new_n14234_), .ZN(new_n14235_));
  OAI21_X1   g11200(.A1(new_n12776_), .A2(new_n14034_), .B(new_n14036_), .ZN(new_n14236_));
  NOR2_X1    g11201(.A1(new_n14034_), .A2(new_n12776_), .ZN(new_n14237_));
  NAND2_X1   g11202(.A1(new_n14033_), .A2(new_n14032_), .ZN(new_n14238_));
  NAND3_X1   g11203(.A1(new_n14238_), .A2(pi0787), .A3(new_n14029_), .ZN(new_n14239_));
  NAND2_X1   g11204(.A1(new_n14237_), .A2(new_n14239_), .ZN(new_n14240_));
  NOR2_X1    g11205(.A1(new_n13998_), .A2(new_n14210_), .ZN(new_n14241_));
  AOI21_X1   g11206(.A1(new_n13629_), .A2(new_n14210_), .B(new_n14241_), .ZN(new_n14242_));
  NOR2_X1    g11207(.A1(new_n14200_), .A2(new_n14203_), .ZN(new_n14243_));
  OAI21_X1   g11208(.A1(new_n13628_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n14244_));
  NAND2_X1   g11209(.A1(new_n14242_), .A2(new_n14244_), .ZN(new_n14245_));
  NAND2_X1   g11210(.A1(new_n14009_), .A2(new_n13629_), .ZN(new_n14246_));
  NOR4_X1    g11211(.A1(new_n14246_), .A2(new_n12776_), .A3(new_n14003_), .A4(new_n14026_), .ZN(new_n14247_));
  NAND2_X1   g11212(.A1(new_n14246_), .A2(pi0787), .ZN(new_n14248_));
  NOR3_X1    g11213(.A1(new_n14026_), .A2(new_n12776_), .A3(new_n14003_), .ZN(new_n14249_));
  NOR2_X1    g11214(.A1(new_n14248_), .A2(new_n14249_), .ZN(new_n14250_));
  NOR4_X1    g11215(.A1(new_n14250_), .A2(new_n14204_), .A3(pi0715), .A4(new_n14247_), .ZN(new_n14251_));
  AOI21_X1   g11216(.A1(new_n14251_), .A2(new_n14245_), .B(pi0644), .ZN(new_n14252_));
  AOI21_X1   g11217(.A1(new_n14240_), .A2(new_n14236_), .B(new_n14252_), .ZN(new_n14253_));
  NOR2_X1    g11218(.A1(new_n14203_), .A2(pi0715), .ZN(new_n14254_));
  INV_X1     g11219(.I(new_n14254_), .ZN(new_n14255_));
  OAI21_X1   g11220(.A1(new_n13629_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n14256_));
  OAI21_X1   g11221(.A1(new_n14250_), .A2(new_n14247_), .B(new_n14256_), .ZN(new_n14257_));
  NOR2_X1    g11222(.A1(new_n14257_), .A2(new_n14242_), .ZN(new_n14258_));
  OAI21_X1   g11223(.A1(new_n14253_), .A2(pi0790), .B(new_n14258_), .ZN(new_n14259_));
  NOR3_X1    g11224(.A1(new_n14235_), .A2(new_n14231_), .A3(new_n14259_), .ZN(po0297));
  INV_X1     g11225(.I(pi0706), .ZN(new_n14261_));
  INV_X1     g11226(.I(new_n13521_), .ZN(new_n14262_));
  INV_X1     g11227(.I(pi0749), .ZN(new_n14263_));
  NOR3_X1    g11228(.A1(new_n13461_), .A2(new_n12618_), .A3(new_n14263_), .ZN(new_n14264_));
  NOR3_X1    g11229(.A1(new_n13453_), .A2(pi0141), .A3(new_n14263_), .ZN(new_n14265_));
  NOR2_X1    g11230(.A1(new_n14265_), .A2(new_n14264_), .ZN(new_n14266_));
  NOR2_X1    g11231(.A1(new_n14266_), .A2(new_n14262_), .ZN(new_n14267_));
  INV_X1     g11232(.I(new_n13151_), .ZN(new_n14268_));
  OAI21_X1   g11233(.A1(pi0299), .A2(new_n13137_), .B(new_n14268_), .ZN(new_n14269_));
  NOR2_X1    g11234(.A1(new_n13181_), .A2(new_n13165_), .ZN(new_n14270_));
  NAND3_X1   g11235(.A1(new_n14270_), .A2(pi0141), .A3(pi0749), .ZN(new_n14271_));
  INV_X1     g11236(.I(new_n14270_), .ZN(new_n14272_));
  NAND3_X1   g11237(.A1(new_n14272_), .A2(pi0141), .A3(new_n14263_), .ZN(new_n14273_));
  NAND2_X1   g11238(.A1(new_n14273_), .A2(new_n14271_), .ZN(new_n14274_));
  NAND2_X1   g11239(.A1(new_n14269_), .A2(new_n14274_), .ZN(new_n14275_));
  NAND3_X1   g11240(.A1(new_n13198_), .A2(pi0141), .A3(pi0749), .ZN(new_n14276_));
  NAND3_X1   g11241(.A1(new_n13200_), .A2(new_n12618_), .A3(pi0749), .ZN(new_n14277_));
  NAND2_X1   g11242(.A1(new_n14277_), .A2(new_n14276_), .ZN(new_n14278_));
  NAND2_X1   g11243(.A1(new_n14278_), .A2(new_n13190_), .ZN(new_n14279_));
  AOI21_X1   g11244(.A1(new_n14275_), .A2(new_n3211_), .B(new_n14279_), .ZN(new_n14280_));
  NOR3_X1    g11245(.A1(new_n14267_), .A2(new_n14280_), .A3(pi0039), .ZN(new_n14281_));
  NAND2_X1   g11246(.A1(new_n13587_), .A2(new_n3098_), .ZN(new_n14282_));
  NAND2_X1   g11247(.A1(new_n13605_), .A2(pi0299), .ZN(new_n14283_));
  NAND2_X1   g11248(.A1(new_n14283_), .A2(new_n14282_), .ZN(new_n14284_));
  INV_X1     g11249(.I(new_n14284_), .ZN(new_n14285_));
  NOR3_X1    g11250(.A1(new_n14285_), .A2(new_n12618_), .A3(new_n14263_), .ZN(new_n14286_));
  NOR3_X1    g11251(.A1(new_n14284_), .A2(new_n12618_), .A3(pi0749), .ZN(new_n14287_));
  OAI21_X1   g11252(.A1(new_n14286_), .A2(new_n14287_), .B(new_n13359_), .ZN(new_n14288_));
  AOI22_X1   g11253(.A1(pi0141), .A2(new_n13106_), .B1(new_n13108_), .B2(pi0749), .ZN(new_n14289_));
  INV_X1     g11254(.I(new_n14289_), .ZN(new_n14290_));
  INV_X1     g11255(.I(new_n12794_), .ZN(new_n14291_));
  NOR2_X1    g11256(.A1(new_n13213_), .A2(pi0038), .ZN(new_n14292_));
  AOI21_X1   g11257(.A1(new_n14291_), .A2(new_n14292_), .B(new_n3183_), .ZN(new_n14293_));
  AOI21_X1   g11258(.A1(new_n14290_), .A2(new_n14293_), .B(new_n14261_), .ZN(new_n14294_));
  OAI21_X1   g11259(.A1(new_n14288_), .A2(new_n14281_), .B(new_n14294_), .ZN(new_n14295_));
  NOR2_X1    g11260(.A1(new_n3289_), .A2(new_n12618_), .ZN(new_n14296_));
  NAND3_X1   g11261(.A1(new_n14295_), .A2(new_n3289_), .A3(new_n14296_), .ZN(new_n14297_));
  NOR2_X1    g11262(.A1(new_n13066_), .A2(new_n13070_), .ZN(new_n14298_));
  NOR2_X1    g11263(.A1(new_n14298_), .A2(pi0039), .ZN(new_n14299_));
  INV_X1     g11264(.I(new_n14299_), .ZN(new_n14300_));
  NOR2_X1    g11265(.A1(new_n13194_), .A2(pi0039), .ZN(new_n14301_));
  NAND2_X1   g11266(.A1(new_n12930_), .A2(new_n13310_), .ZN(new_n14302_));
  OAI21_X1   g11267(.A1(new_n13467_), .A2(new_n5796_), .B(new_n5636_), .ZN(new_n14303_));
  INV_X1     g11268(.I(new_n13310_), .ZN(new_n14304_));
  NOR3_X1    g11269(.A1(new_n12878_), .A2(new_n5636_), .A3(new_n14304_), .ZN(new_n14305_));
  INV_X1     g11270(.I(new_n14305_), .ZN(new_n14306_));
  OAI21_X1   g11271(.A1(new_n14302_), .A2(new_n14303_), .B(new_n14306_), .ZN(new_n14307_));
  NOR2_X1    g11272(.A1(new_n14307_), .A2(new_n3090_), .ZN(new_n14308_));
  NOR2_X1    g11273(.A1(new_n14308_), .A2(new_n13466_), .ZN(new_n14309_));
  NOR3_X1    g11274(.A1(new_n14307_), .A2(new_n3090_), .A3(new_n5481_), .ZN(new_n14310_));
  NOR2_X1    g11275(.A1(new_n14309_), .A2(new_n14310_), .ZN(new_n14311_));
  NAND2_X1   g11276(.A1(new_n13478_), .A2(new_n5636_), .ZN(new_n14312_));
  NAND3_X1   g11277(.A1(new_n14312_), .A2(pi0299), .A3(new_n13335_), .ZN(new_n14313_));
  OAI21_X1   g11278(.A1(new_n14313_), .A2(new_n14311_), .B(new_n3090_), .ZN(new_n14314_));
  INV_X1     g11279(.I(new_n13416_), .ZN(new_n14315_));
  OAI21_X1   g11280(.A1(new_n12821_), .A2(new_n5378_), .B(new_n14315_), .ZN(new_n14316_));
  OAI21_X1   g11281(.A1(pi0603), .A2(new_n13262_), .B(new_n13257_), .ZN(new_n14317_));
  AOI21_X1   g11282(.A1(new_n13423_), .A2(new_n5794_), .B(new_n13254_), .ZN(new_n14318_));
  NAND2_X1   g11283(.A1(new_n14317_), .A2(new_n14318_), .ZN(new_n14319_));
  NAND2_X1   g11284(.A1(new_n14319_), .A2(new_n14316_), .ZN(new_n14320_));
  OAI21_X1   g11285(.A1(new_n13273_), .A2(new_n12945_), .B(new_n5378_), .ZN(new_n14321_));
  INV_X1     g11286(.I(new_n14321_), .ZN(new_n14322_));
  INV_X1     g11287(.I(new_n13338_), .ZN(new_n14323_));
  NAND2_X1   g11288(.A1(new_n13492_), .A2(new_n5636_), .ZN(new_n14324_));
  NAND3_X1   g11289(.A1(new_n13273_), .A2(new_n14323_), .A3(new_n14324_), .ZN(new_n14325_));
  NAND2_X1   g11290(.A1(new_n13275_), .A2(new_n3091_), .ZN(new_n14326_));
  NOR2_X1    g11291(.A1(new_n14325_), .A2(new_n14326_), .ZN(new_n14327_));
  OAI21_X1   g11292(.A1(new_n12981_), .A2(new_n14322_), .B(new_n14327_), .ZN(new_n14328_));
  AOI21_X1   g11293(.A1(new_n14328_), .A2(new_n5397_), .B(new_n14320_), .ZN(new_n14329_));
  AOI21_X1   g11294(.A1(new_n14314_), .A2(new_n14329_), .B(new_n3183_), .ZN(new_n14330_));
  INV_X1     g11295(.I(new_n13185_), .ZN(new_n14331_));
  NOR3_X1    g11296(.A1(new_n13052_), .A2(new_n13166_), .A3(new_n13169_), .ZN(new_n14332_));
  AOI21_X1   g11297(.A1(new_n13167_), .A2(new_n13170_), .B(new_n13161_), .ZN(new_n14333_));
  OAI21_X1   g11298(.A1(new_n14333_), .A2(new_n14332_), .B(pi0603), .ZN(new_n14334_));
  OAI21_X1   g11299(.A1(new_n13061_), .A2(new_n13062_), .B(new_n2777_), .ZN(new_n14335_));
  OAI21_X1   g11300(.A1(new_n2777_), .A2(new_n13176_), .B(new_n14335_), .ZN(new_n14336_));
  AOI21_X1   g11301(.A1(new_n14336_), .A2(pi0299), .B(pi0603), .ZN(new_n14337_));
  OAI22_X1   g11302(.A1(new_n14334_), .A2(new_n14331_), .B1(new_n13145_), .B2(new_n14337_), .ZN(new_n14338_));
  INV_X1     g11303(.I(new_n14320_), .ZN(new_n14339_));
  NOR2_X1    g11304(.A1(new_n14307_), .A2(new_n3111_), .ZN(new_n14340_));
  NOR2_X1    g11305(.A1(new_n14340_), .A2(new_n13309_), .ZN(new_n14341_));
  NOR3_X1    g11306(.A1(new_n14307_), .A2(new_n3111_), .A3(new_n5456_), .ZN(new_n14342_));
  NOR2_X1    g11307(.A1(new_n14341_), .A2(new_n14342_), .ZN(new_n14343_));
  OAI21_X1   g11308(.A1(new_n14313_), .A2(new_n14343_), .B(new_n3111_), .ZN(new_n14344_));
  NOR2_X1    g11309(.A1(new_n14322_), .A2(new_n13516_), .ZN(new_n14345_));
  NAND4_X1   g11310(.A1(new_n13491_), .A2(new_n3312_), .A3(new_n13275_), .A4(new_n14324_), .ZN(new_n14346_));
  OAI21_X1   g11311(.A1(new_n14346_), .A2(new_n14345_), .B(new_n5455_), .ZN(new_n14347_));
  NAND4_X1   g11312(.A1(new_n14344_), .A2(pi0039), .A3(new_n14339_), .A4(new_n14347_), .ZN(new_n14348_));
  NOR3_X1    g11313(.A1(new_n14348_), .A2(new_n14338_), .A3(new_n14330_), .ZN(new_n14349_));
  INV_X1     g11314(.I(new_n14311_), .ZN(new_n14350_));
  OAI21_X1   g11315(.A1(new_n5378_), .A2(new_n13340_), .B(new_n13335_), .ZN(new_n14351_));
  NOR2_X1    g11316(.A1(new_n14351_), .A2(new_n3098_), .ZN(new_n14352_));
  AOI21_X1   g11317(.A1(new_n14352_), .A2(new_n14350_), .B(pi0223), .ZN(new_n14353_));
  INV_X1     g11318(.I(new_n14329_), .ZN(new_n14354_));
  OAI21_X1   g11319(.A1(new_n14354_), .A2(new_n14353_), .B(pi0039), .ZN(new_n14355_));
  AOI21_X1   g11320(.A1(new_n13185_), .A2(new_n13186_), .B(new_n13188_), .ZN(new_n14356_));
  INV_X1     g11321(.I(new_n14343_), .ZN(new_n14357_));
  AOI21_X1   g11322(.A1(new_n14352_), .A2(new_n14357_), .B(pi0215), .ZN(new_n14358_));
  NAND2_X1   g11323(.A1(new_n14347_), .A2(new_n14339_), .ZN(new_n14359_));
  NOR3_X1    g11324(.A1(new_n14359_), .A2(new_n3183_), .A3(new_n14358_), .ZN(new_n14360_));
  AOI21_X1   g11325(.A1(new_n14356_), .A2(new_n14360_), .B(new_n14355_), .ZN(new_n14361_));
  NOR2_X1    g11326(.A1(new_n14361_), .A2(new_n14349_), .ZN(new_n14362_));
  AOI21_X1   g11327(.A1(new_n12618_), .A2(new_n14263_), .B(new_n14300_), .ZN(new_n14363_));
  NOR2_X1    g11328(.A1(new_n14363_), .A2(pi0038), .ZN(new_n14364_));
  NOR2_X1    g11329(.A1(new_n12992_), .A2(new_n12986_), .ZN(new_n14365_));
  NOR2_X1    g11330(.A1(new_n12977_), .A2(new_n14365_), .ZN(new_n14366_));
  OAI21_X1   g11331(.A1(new_n13405_), .A2(new_n3111_), .B(new_n12930_), .ZN(new_n14367_));
  AOI21_X1   g11332(.A1(new_n14367_), .A2(new_n5454_), .B(pi0299), .ZN(new_n14368_));
  NAND3_X1   g11333(.A1(new_n13418_), .A2(new_n3312_), .A3(new_n5454_), .ZN(new_n14369_));
  NAND2_X1   g11334(.A1(new_n14316_), .A2(new_n13203_), .ZN(new_n14370_));
  INV_X1     g11335(.I(new_n13516_), .ZN(new_n14371_));
  NAND3_X1   g11336(.A1(new_n14370_), .A2(new_n5454_), .A3(new_n14371_), .ZN(new_n14372_));
  NAND2_X1   g11337(.A1(new_n14372_), .A2(new_n14369_), .ZN(new_n14373_));
  NOR2_X1    g11338(.A1(new_n13365_), .A2(new_n5636_), .ZN(new_n14374_));
  NAND2_X1   g11339(.A1(new_n13364_), .A2(new_n14374_), .ZN(new_n14375_));
  NAND2_X1   g11340(.A1(new_n13372_), .A2(new_n14374_), .ZN(new_n14376_));
  XOR2_X1    g11341(.A1(new_n14376_), .A2(new_n14375_), .Z(new_n14377_));
  NOR2_X1    g11342(.A1(new_n13678_), .A2(new_n13105_), .ZN(new_n14378_));
  NAND3_X1   g11343(.A1(new_n14373_), .A2(new_n14377_), .A3(new_n14378_), .ZN(new_n14379_));
  NOR2_X1    g11344(.A1(new_n14379_), .A2(new_n14368_), .ZN(new_n14380_));
  INV_X1     g11345(.I(new_n13302_), .ZN(new_n14381_));
  XNOR2_X1   g11346(.A1(new_n14376_), .A2(new_n14375_), .ZN(new_n14382_));
  NAND3_X1   g11347(.A1(new_n13418_), .A2(new_n3091_), .A3(new_n5398_), .ZN(new_n14383_));
  NAND3_X1   g11348(.A1(new_n14370_), .A2(new_n3092_), .A3(new_n5398_), .ZN(new_n14384_));
  AOI21_X1   g11349(.A1(new_n14383_), .A2(new_n14384_), .B(new_n14382_), .ZN(new_n14385_));
  AOI21_X1   g11350(.A1(new_n13405_), .A2(new_n3565_), .B(new_n13701_), .ZN(new_n14386_));
  OAI21_X1   g11351(.A1(new_n14385_), .A2(new_n14381_), .B(new_n14386_), .ZN(new_n14387_));
  INV_X1     g11352(.I(new_n14387_), .ZN(new_n14388_));
  NOR2_X1    g11353(.A1(new_n14388_), .A2(new_n14380_), .ZN(new_n14389_));
  AOI22_X1   g11354(.A1(new_n14366_), .A2(pi0141), .B1(pi0749), .B2(new_n14389_), .ZN(new_n14390_));
  NOR3_X1    g11355(.A1(new_n14390_), .A2(new_n3183_), .A3(new_n14364_), .ZN(new_n14391_));
  NOR2_X1    g11356(.A1(new_n14290_), .A2(new_n3259_), .ZN(new_n14392_));
  NOR2_X1    g11357(.A1(new_n14391_), .A2(new_n14392_), .ZN(new_n14393_));
  INV_X1     g11358(.I(new_n14393_), .ZN(new_n14394_));
  AOI21_X1   g11359(.A1(new_n14297_), .A2(new_n14261_), .B(new_n14394_), .ZN(new_n14395_));
  AOI21_X1   g11360(.A1(new_n13097_), .A2(new_n3259_), .B(new_n13626_), .ZN(new_n14396_));
  AOI21_X1   g11361(.A1(new_n13720_), .A2(pi0706), .B(pi0141), .ZN(new_n14397_));
  NAND2_X1   g11362(.A1(new_n12618_), .A2(new_n14261_), .ZN(new_n14398_));
  NAND3_X1   g11363(.A1(new_n3290_), .A2(pi0141), .A3(new_n14398_), .ZN(new_n14399_));
  OAI22_X1   g11364(.A1(new_n14396_), .A2(new_n14399_), .B1(new_n13109_), .B2(new_n14397_), .ZN(new_n14400_));
  NAND2_X1   g11365(.A1(new_n13715_), .A2(pi0039), .ZN(new_n14401_));
  NOR3_X1    g11366(.A1(new_n13699_), .A2(new_n3183_), .A3(new_n13704_), .ZN(new_n14402_));
  NAND2_X1   g11367(.A1(new_n13197_), .A2(new_n14402_), .ZN(new_n14403_));
  XNOR2_X1   g11368(.A1(new_n14403_), .A2(new_n14401_), .ZN(new_n14404_));
  NOR2_X1    g11369(.A1(new_n13669_), .A2(new_n13650_), .ZN(new_n14405_));
  NAND2_X1   g11370(.A1(new_n13675_), .A2(new_n13640_), .ZN(new_n14406_));
  NOR2_X1    g11371(.A1(new_n13678_), .A2(new_n13680_), .ZN(new_n14407_));
  NAND3_X1   g11372(.A1(new_n13662_), .A2(pi0215), .A3(new_n5454_), .ZN(new_n14408_));
  NAND3_X1   g11373(.A1(new_n13666_), .A2(pi0215), .A3(new_n5455_), .ZN(new_n14409_));
  AOI21_X1   g11374(.A1(new_n14409_), .A2(new_n14408_), .B(new_n13655_), .ZN(new_n14410_));
  AOI21_X1   g11375(.A1(new_n14410_), .A2(pi0299), .B(new_n14407_), .ZN(new_n14411_));
  OAI21_X1   g11376(.A1(new_n14411_), .A2(new_n14406_), .B(pi0039), .ZN(new_n14412_));
  NAND4_X1   g11377(.A1(new_n14412_), .A2(new_n14405_), .A3(pi0039), .A4(new_n13165_), .ZN(new_n14413_));
  INV_X1     g11378(.I(new_n13650_), .ZN(new_n14414_));
  INV_X1     g11379(.I(new_n13651_), .ZN(new_n14415_));
  AOI21_X1   g11380(.A1(new_n13666_), .A2(pi0223), .B(new_n13466_), .ZN(new_n14416_));
  NOR3_X1    g11381(.A1(new_n13662_), .A2(new_n3090_), .A3(new_n5398_), .ZN(new_n14417_));
  OAI21_X1   g11382(.A1(new_n14416_), .A2(new_n14417_), .B(new_n13654_), .ZN(new_n14418_));
  OAI21_X1   g11383(.A1(new_n14418_), .A2(new_n3098_), .B(new_n14415_), .ZN(new_n14419_));
  NAND4_X1   g11384(.A1(new_n14419_), .A2(new_n14414_), .A3(pi0039), .A4(new_n13165_), .ZN(new_n14420_));
  NAND3_X1   g11385(.A1(new_n13685_), .A2(new_n14420_), .A3(pi0039), .ZN(new_n14421_));
  NAND2_X1   g11386(.A1(new_n14421_), .A2(new_n14413_), .ZN(new_n14422_));
  NAND3_X1   g11387(.A1(new_n14422_), .A2(pi0038), .A3(pi0141), .ZN(new_n14423_));
  XNOR2_X1   g11388(.A1(new_n14420_), .A2(new_n14412_), .ZN(new_n14424_));
  NAND3_X1   g11389(.A1(new_n14424_), .A2(new_n3259_), .A3(pi0141), .ZN(new_n14425_));
  AOI21_X1   g11390(.A1(new_n14425_), .A2(new_n14423_), .B(new_n14404_), .ZN(new_n14426_));
  NAND2_X1   g11391(.A1(new_n14426_), .A2(new_n14400_), .ZN(new_n14427_));
  INV_X1     g11392(.I(new_n13627_), .ZN(new_n14428_));
  NOR2_X1    g11393(.A1(pi0625), .A2(pi1153), .ZN(new_n14429_));
  INV_X1     g11394(.I(new_n14429_), .ZN(new_n14430_));
  NOR2_X1    g11395(.A1(new_n14428_), .A2(new_n14430_), .ZN(new_n14431_));
  OR3_X2     g11396(.A1(new_n14431_), .A2(new_n12618_), .A3(new_n14081_), .Z(new_n14432_));
  NOR2_X1    g11397(.A1(new_n14392_), .A2(new_n3290_), .ZN(new_n14433_));
  INV_X1     g11398(.I(new_n14433_), .ZN(new_n14434_));
  NOR2_X1    g11399(.A1(new_n3290_), .A2(new_n12618_), .ZN(new_n14435_));
  NAND3_X1   g11400(.A1(new_n14391_), .A2(new_n14434_), .A3(new_n14435_), .ZN(new_n14436_));
  NAND2_X1   g11401(.A1(new_n14391_), .A2(new_n14435_), .ZN(new_n14437_));
  NAND2_X1   g11402(.A1(new_n14437_), .A2(new_n14433_), .ZN(new_n14438_));
  NAND2_X1   g11403(.A1(new_n14438_), .A2(new_n14436_), .ZN(new_n14439_));
  NAND2_X1   g11404(.A1(pi0625), .A2(pi1153), .ZN(new_n14441_));
  AOI21_X1   g11405(.A1(new_n14432_), .A2(new_n14427_), .B(new_n14441_), .ZN(new_n14442_));
  NAND3_X1   g11406(.A1(new_n14395_), .A2(pi0625), .A3(pi0778), .ZN(new_n14446_));
  OAI21_X1   g11407(.A1(pi0625), .A2(new_n14442_), .B(new_n14395_), .ZN(new_n14447_));
  NAND3_X1   g11408(.A1(new_n14395_), .A2(pi0625), .A3(pi0778), .ZN(new_n14448_));
  NAND3_X1   g11409(.A1(new_n14447_), .A2(pi0778), .A3(new_n14448_), .ZN(new_n14449_));
  NAND2_X1   g11410(.A1(new_n14449_), .A2(new_n14446_), .ZN(new_n14450_));
  NAND3_X1   g11411(.A1(new_n14426_), .A2(new_n13748_), .A3(new_n14400_), .ZN(new_n14451_));
  XNOR2_X1   g11412(.A1(pi0625), .A2(pi1153), .ZN(new_n14452_));
  AOI21_X1   g11413(.A1(new_n14426_), .A2(new_n14400_), .B(new_n14452_), .ZN(new_n14453_));
  NAND2_X1   g11414(.A1(new_n13627_), .A2(new_n12618_), .ZN(new_n14454_));
  NOR2_X1    g11415(.A1(new_n14454_), .A2(new_n14452_), .ZN(new_n14455_));
  XNOR2_X1   g11416(.A1(new_n14453_), .A2(new_n14455_), .ZN(new_n14456_));
  OAI21_X1   g11417(.A1(new_n14456_), .A2(new_n13748_), .B(new_n14451_), .ZN(new_n14457_));
  INV_X1     g11418(.I(new_n14436_), .ZN(new_n14458_));
  AOI21_X1   g11419(.A1(new_n14391_), .A2(new_n14435_), .B(new_n14434_), .ZN(new_n14459_));
  NOR3_X1    g11420(.A1(new_n14458_), .A2(new_n13775_), .A3(new_n14459_), .ZN(new_n14460_));
  NAND2_X1   g11421(.A1(new_n14454_), .A2(new_n13780_), .ZN(new_n14461_));
  INV_X1     g11422(.I(new_n14461_), .ZN(new_n14462_));
  OAI21_X1   g11423(.A1(new_n14457_), .A2(new_n13785_), .B(new_n13766_), .ZN(new_n14463_));
  NAND2_X1   g11424(.A1(new_n14457_), .A2(pi0609), .ZN(new_n14464_));
  INV_X1     g11425(.I(new_n13793_), .ZN(new_n14465_));
  NAND3_X1   g11426(.A1(new_n14438_), .A2(new_n13776_), .A3(new_n14436_), .ZN(new_n14466_));
  NOR2_X1    g11427(.A1(new_n14101_), .A2(new_n13778_), .ZN(new_n14467_));
  AOI21_X1   g11428(.A1(new_n14454_), .A2(new_n14467_), .B(pi0609), .ZN(new_n14468_));
  NOR2_X1    g11429(.A1(new_n14466_), .A2(new_n14468_), .ZN(new_n14469_));
  NOR2_X1    g11430(.A1(new_n14469_), .A2(new_n14465_), .ZN(new_n14470_));
  AOI21_X1   g11431(.A1(new_n14464_), .A2(new_n14470_), .B(pi0609), .ZN(new_n14471_));
  INV_X1     g11432(.I(new_n14471_), .ZN(new_n14472_));
  NAND4_X1   g11433(.A1(new_n14450_), .A2(pi0785), .A3(new_n14463_), .A4(new_n14472_), .ZN(new_n14473_));
  NAND2_X1   g11434(.A1(new_n14450_), .A2(new_n14463_), .ZN(new_n14474_));
  NAND3_X1   g11435(.A1(new_n14450_), .A2(pi0785), .A3(new_n14472_), .ZN(new_n14475_));
  NAND3_X1   g11436(.A1(new_n14475_), .A2(new_n14474_), .A3(pi0785), .ZN(new_n14476_));
  NAND2_X1   g11437(.A1(new_n14476_), .A2(new_n14473_), .ZN(new_n14477_));
  INV_X1     g11438(.I(new_n14454_), .ZN(new_n14478_));
  OAI21_X1   g11439(.A1(new_n14460_), .A2(new_n14462_), .B(pi0609), .ZN(new_n14479_));
  INV_X1     g11440(.I(new_n14468_), .ZN(new_n14480_));
  NAND2_X1   g11441(.A1(new_n14460_), .A2(new_n14480_), .ZN(new_n14481_));
  NOR2_X1    g11442(.A1(new_n14454_), .A2(new_n13776_), .ZN(new_n14482_));
  AOI21_X1   g11443(.A1(new_n14439_), .A2(new_n13776_), .B(new_n14482_), .ZN(new_n14483_));
  NOR4_X1    g11444(.A1(new_n14479_), .A2(new_n14481_), .A3(new_n14483_), .A4(new_n13801_), .ZN(new_n14484_));
  NAND2_X1   g11445(.A1(new_n14479_), .A2(pi0785), .ZN(new_n14485_));
  NOR3_X1    g11446(.A1(new_n14481_), .A2(new_n14483_), .A3(new_n13801_), .ZN(new_n14486_));
  NOR2_X1    g11447(.A1(new_n14486_), .A2(new_n14485_), .ZN(new_n14487_));
  NOR2_X1    g11448(.A1(new_n14487_), .A2(new_n14484_), .ZN(new_n14488_));
  AOI21_X1   g11449(.A1(new_n14488_), .A2(pi0618), .B(new_n13819_), .ZN(new_n14489_));
  AOI21_X1   g11450(.A1(new_n14466_), .A2(new_n14461_), .B(new_n13766_), .ZN(new_n14490_));
  OAI21_X1   g11451(.A1(new_n14458_), .A2(new_n14459_), .B(new_n13776_), .ZN(new_n14491_));
  INV_X1     g11452(.I(new_n14482_), .ZN(new_n14492_));
  NAND2_X1   g11453(.A1(new_n14491_), .A2(new_n14492_), .ZN(new_n14493_));
  NAND4_X1   g11454(.A1(new_n14490_), .A2(new_n14493_), .A3(new_n14469_), .A4(pi0785), .ZN(new_n14494_));
  NOR2_X1    g11455(.A1(new_n14490_), .A2(new_n13801_), .ZN(new_n14495_));
  NAND3_X1   g11456(.A1(new_n14493_), .A2(new_n14469_), .A3(pi0785), .ZN(new_n14496_));
  NAND2_X1   g11457(.A1(new_n14496_), .A2(new_n14495_), .ZN(new_n14497_));
  NAND2_X1   g11458(.A1(new_n14497_), .A2(new_n14494_), .ZN(new_n14498_));
  NOR3_X1    g11459(.A1(new_n14498_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n14499_));
  OAI21_X1   g11460(.A1(new_n14489_), .A2(new_n14499_), .B(new_n14478_), .ZN(new_n14500_));
  INV_X1     g11461(.I(new_n13824_), .ZN(new_n14501_));
  NOR2_X1    g11462(.A1(new_n14454_), .A2(new_n13805_), .ZN(new_n14502_));
  AOI21_X1   g11463(.A1(new_n14457_), .A2(new_n13805_), .B(new_n14502_), .ZN(new_n14503_));
  NOR2_X1    g11464(.A1(new_n14503_), .A2(pi0618), .ZN(new_n14504_));
  NOR2_X1    g11465(.A1(new_n14504_), .A2(new_n14501_), .ZN(new_n14505_));
  AOI21_X1   g11466(.A1(new_n14500_), .A2(new_n14505_), .B(pi0618), .ZN(new_n14506_));
  INV_X1     g11467(.I(new_n14506_), .ZN(new_n14507_));
  NAND3_X1   g11468(.A1(new_n14498_), .A2(pi0618), .A3(pi1154), .ZN(new_n14508_));
  NAND4_X1   g11469(.A1(new_n14497_), .A2(new_n13816_), .A3(pi1154), .A4(new_n14494_), .ZN(new_n14509_));
  AOI21_X1   g11470(.A1(new_n14508_), .A2(new_n14509_), .B(new_n14454_), .ZN(new_n14510_));
  OAI21_X1   g11471(.A1(new_n14503_), .A2(new_n13816_), .B(new_n13836_), .ZN(new_n14511_));
  OAI21_X1   g11472(.A1(new_n14510_), .A2(new_n14511_), .B(new_n13816_), .ZN(new_n14512_));
  NAND4_X1   g11473(.A1(new_n14477_), .A2(pi0781), .A3(new_n14507_), .A4(new_n14512_), .ZN(new_n14513_));
  NAND2_X1   g11474(.A1(new_n14477_), .A2(new_n14507_), .ZN(new_n14514_));
  NAND3_X1   g11475(.A1(new_n14477_), .A2(pi0781), .A3(new_n14512_), .ZN(new_n14515_));
  NAND3_X1   g11476(.A1(new_n14515_), .A2(new_n14514_), .A3(pi0781), .ZN(new_n14516_));
  NAND2_X1   g11477(.A1(new_n14516_), .A2(new_n14513_), .ZN(new_n14517_));
  NAND3_X1   g11478(.A1(new_n14498_), .A2(pi0618), .A3(pi1154), .ZN(new_n14518_));
  NAND3_X1   g11479(.A1(new_n14488_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n14519_));
  AOI21_X1   g11480(.A1(new_n14519_), .A2(new_n14518_), .B(new_n14454_), .ZN(new_n14520_));
  NOR2_X1    g11481(.A1(new_n14520_), .A2(new_n13855_), .ZN(new_n14521_));
  NOR2_X1    g11482(.A1(new_n14488_), .A2(new_n13855_), .ZN(new_n14522_));
  NAND2_X1   g11483(.A1(new_n14510_), .A2(new_n14522_), .ZN(new_n14523_));
  NOR2_X1    g11484(.A1(new_n14521_), .A2(new_n14523_), .ZN(new_n14524_));
  NAND2_X1   g11485(.A1(new_n14500_), .A2(pi0781), .ZN(new_n14525_));
  AOI21_X1   g11486(.A1(new_n14488_), .A2(pi1154), .B(new_n13819_), .ZN(new_n14526_));
  INV_X1     g11487(.I(new_n14509_), .ZN(new_n14527_));
  NOR2_X1    g11488(.A1(new_n14526_), .A2(new_n14527_), .ZN(new_n14528_));
  NOR4_X1    g11489(.A1(new_n14528_), .A2(new_n13855_), .A3(new_n14454_), .A4(new_n14488_), .ZN(new_n14529_));
  NOR2_X1    g11490(.A1(new_n14529_), .A2(new_n14525_), .ZN(new_n14530_));
  NOR2_X1    g11491(.A1(new_n14530_), .A2(new_n14524_), .ZN(new_n14531_));
  AOI21_X1   g11492(.A1(new_n14531_), .A2(pi0619), .B(new_n13904_), .ZN(new_n14532_));
  NAND4_X1   g11493(.A1(new_n14520_), .A2(new_n14510_), .A3(pi0781), .A4(new_n14498_), .ZN(new_n14533_));
  NAND2_X1   g11494(.A1(new_n14521_), .A2(new_n14523_), .ZN(new_n14534_));
  NAND2_X1   g11495(.A1(new_n14534_), .A2(new_n14533_), .ZN(new_n14535_));
  NOR3_X1    g11496(.A1(new_n14535_), .A2(new_n13860_), .A3(pi1159), .ZN(new_n14536_));
  OAI21_X1   g11497(.A1(new_n14532_), .A2(new_n14536_), .B(new_n14478_), .ZN(new_n14537_));
  INV_X1     g11498(.I(new_n13885_), .ZN(new_n14538_));
  NOR2_X1    g11499(.A1(new_n14478_), .A2(new_n13880_), .ZN(new_n14539_));
  AOI21_X1   g11500(.A1(new_n14503_), .A2(new_n13880_), .B(new_n14539_), .ZN(new_n14540_));
  AOI21_X1   g11501(.A1(new_n14540_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n14541_));
  NAND2_X1   g11502(.A1(new_n14537_), .A2(new_n14541_), .ZN(new_n14542_));
  NAND2_X1   g11503(.A1(new_n14542_), .A2(new_n13860_), .ZN(new_n14543_));
  AOI21_X1   g11504(.A1(new_n14543_), .A2(new_n14517_), .B(new_n13896_), .ZN(new_n14544_));
  NAND3_X1   g11505(.A1(new_n14535_), .A2(pi0619), .A3(pi1159), .ZN(new_n14545_));
  NAND4_X1   g11506(.A1(new_n14534_), .A2(new_n13860_), .A3(pi1159), .A4(new_n14533_), .ZN(new_n14546_));
  AOI21_X1   g11507(.A1(new_n14545_), .A2(new_n14546_), .B(new_n14454_), .ZN(new_n14547_));
  NAND2_X1   g11508(.A1(new_n14540_), .A2(pi0619), .ZN(new_n14548_));
  NAND2_X1   g11509(.A1(new_n14548_), .A2(new_n13892_), .ZN(new_n14549_));
  OAI21_X1   g11510(.A1(new_n14547_), .A2(new_n14549_), .B(new_n13860_), .ZN(new_n14550_));
  NAND3_X1   g11511(.A1(new_n14517_), .A2(pi0789), .A3(new_n14550_), .ZN(new_n14551_));
  XNOR2_X1   g11512(.A1(new_n14544_), .A2(new_n14551_), .ZN(new_n14552_));
  NAND3_X1   g11513(.A1(new_n14535_), .A2(pi0619), .A3(pi1159), .ZN(new_n14553_));
  NAND3_X1   g11514(.A1(new_n14531_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n14554_));
  AOI21_X1   g11515(.A1(new_n14554_), .A2(new_n14553_), .B(new_n14454_), .ZN(new_n14555_));
  NAND4_X1   g11516(.A1(new_n14555_), .A2(new_n14547_), .A3(pi0789), .A4(new_n14535_), .ZN(new_n14556_));
  NOR2_X1    g11517(.A1(new_n14531_), .A2(new_n13896_), .ZN(new_n14557_));
  NAND2_X1   g11518(.A1(new_n14547_), .A2(new_n14557_), .ZN(new_n14558_));
  NAND3_X1   g11519(.A1(new_n14558_), .A2(pi0789), .A3(new_n14537_), .ZN(new_n14559_));
  NAND2_X1   g11520(.A1(new_n14559_), .A2(new_n14556_), .ZN(new_n14560_));
  NAND3_X1   g11521(.A1(new_n14560_), .A2(pi0626), .A3(pi1158), .ZN(new_n14561_));
  NAND4_X1   g11522(.A1(new_n14559_), .A2(new_n13901_), .A3(pi1158), .A4(new_n14556_), .ZN(new_n14562_));
  AOI21_X1   g11523(.A1(new_n14561_), .A2(new_n14562_), .B(new_n14454_), .ZN(new_n14563_));
  NOR2_X1    g11524(.A1(new_n14454_), .A2(new_n13919_), .ZN(new_n14564_));
  AOI21_X1   g11525(.A1(new_n14540_), .A2(new_n13919_), .B(new_n14564_), .ZN(new_n14565_));
  AOI21_X1   g11526(.A1(new_n14565_), .A2(new_n13901_), .B(new_n13924_), .ZN(new_n14566_));
  INV_X1     g11527(.I(new_n14566_), .ZN(new_n14567_));
  OAI21_X1   g11528(.A1(new_n14563_), .A2(new_n14567_), .B(new_n13901_), .ZN(new_n14568_));
  NAND3_X1   g11529(.A1(new_n14560_), .A2(pi0626), .A3(pi1158), .ZN(new_n14569_));
  NAND4_X1   g11530(.A1(new_n14559_), .A2(pi0626), .A3(new_n13929_), .A4(new_n14556_), .ZN(new_n14570_));
  AOI21_X1   g11531(.A1(new_n14569_), .A2(new_n14570_), .B(new_n14454_), .ZN(new_n14571_));
  NAND4_X1   g11532(.A1(new_n14568_), .A2(pi0626), .A3(new_n14552_), .A4(pi0788), .ZN(new_n14575_));
  NAND2_X1   g11533(.A1(new_n14568_), .A2(new_n14552_), .ZN(new_n14576_));
  NOR2_X1    g11534(.A1(new_n13901_), .A2(new_n13937_), .ZN(new_n14577_));
  NAND2_X1   g11535(.A1(new_n14552_), .A2(new_n14577_), .ZN(new_n14578_));
  NAND3_X1   g11536(.A1(new_n14576_), .A2(pi0788), .A3(new_n14578_), .ZN(new_n14579_));
  NAND2_X1   g11537(.A1(new_n14579_), .A2(new_n14575_), .ZN(new_n14580_));
  NAND4_X1   g11538(.A1(new_n14563_), .A2(new_n14571_), .A3(pi0788), .A4(new_n14560_), .ZN(new_n14581_));
  AOI21_X1   g11539(.A1(new_n14531_), .A2(pi1159), .B(new_n13904_), .ZN(new_n14582_));
  INV_X1     g11540(.I(new_n14546_), .ZN(new_n14583_));
  OAI21_X1   g11541(.A1(new_n14582_), .A2(new_n14583_), .B(new_n14478_), .ZN(new_n14584_));
  NOR4_X1    g11542(.A1(new_n14537_), .A2(new_n14584_), .A3(new_n13896_), .A4(new_n14531_), .ZN(new_n14585_));
  NAND2_X1   g11543(.A1(new_n14537_), .A2(pi0789), .ZN(new_n14586_));
  INV_X1     g11544(.I(new_n14557_), .ZN(new_n14587_));
  NOR2_X1    g11545(.A1(new_n14584_), .A2(new_n14587_), .ZN(new_n14588_));
  NOR2_X1    g11546(.A1(new_n14588_), .A2(new_n14586_), .ZN(new_n14589_));
  NOR2_X1    g11547(.A1(new_n14589_), .A2(new_n14585_), .ZN(new_n14590_));
  AOI21_X1   g11548(.A1(new_n14590_), .A2(pi1158), .B(new_n13954_), .ZN(new_n14591_));
  INV_X1     g11549(.I(new_n14562_), .ZN(new_n14592_));
  OAI21_X1   g11550(.A1(new_n14591_), .A2(new_n14592_), .B(new_n14478_), .ZN(new_n14593_));
  NOR2_X1    g11551(.A1(new_n14590_), .A2(new_n13937_), .ZN(new_n14594_));
  NAND2_X1   g11552(.A1(new_n14571_), .A2(new_n14594_), .ZN(new_n14595_));
  NAND3_X1   g11553(.A1(new_n14595_), .A2(pi0788), .A3(new_n14593_), .ZN(new_n14596_));
  NAND2_X1   g11554(.A1(new_n14596_), .A2(new_n14581_), .ZN(new_n14597_));
  NOR2_X1    g11555(.A1(new_n14478_), .A2(new_n13966_), .ZN(new_n14598_));
  AOI21_X1   g11556(.A1(new_n14565_), .A2(new_n13966_), .B(new_n14598_), .ZN(new_n14599_));
  NAND2_X1   g11557(.A1(new_n14599_), .A2(pi0628), .ZN(new_n14600_));
  XOR2_X1    g11558(.A1(new_n14600_), .A2(new_n13971_), .Z(new_n14601_));
  NAND2_X1   g11559(.A1(new_n14601_), .A2(new_n14478_), .ZN(new_n14602_));
  NAND2_X1   g11560(.A1(new_n14602_), .A2(new_n13977_), .ZN(new_n14603_));
  OAI21_X1   g11561(.A1(new_n14597_), .A2(new_n14603_), .B(new_n13942_), .ZN(new_n14604_));
  AOI21_X1   g11562(.A1(new_n14580_), .A2(new_n14604_), .B(new_n12777_), .ZN(new_n14605_));
  NOR2_X1    g11563(.A1(new_n13942_), .A2(new_n12777_), .ZN(new_n14606_));
  INV_X1     g11564(.I(new_n14599_), .ZN(new_n14607_));
  NOR2_X1    g11565(.A1(new_n14607_), .A2(new_n13969_), .ZN(new_n14608_));
  XOR2_X1    g11566(.A1(new_n14608_), .A2(new_n13970_), .Z(new_n14609_));
  NAND2_X1   g11567(.A1(new_n14580_), .A2(new_n14606_), .ZN(new_n14613_));
  XOR2_X1    g11568(.A1(new_n14605_), .A2(new_n14613_), .Z(new_n14614_));
  NOR2_X1    g11569(.A1(new_n14478_), .A2(new_n13994_), .ZN(new_n14615_));
  INV_X1     g11570(.I(new_n14615_), .ZN(new_n14616_));
  NAND3_X1   g11571(.A1(new_n14596_), .A2(new_n13994_), .A3(new_n14581_), .ZN(new_n14617_));
  NAND2_X1   g11572(.A1(new_n14617_), .A2(new_n14616_), .ZN(new_n14618_));
  NAND4_X1   g11573(.A1(new_n14609_), .A2(pi0792), .A3(new_n14478_), .A4(new_n14607_), .ZN(new_n14619_));
  AOI21_X1   g11574(.A1(pi0792), .A2(new_n14602_), .B(new_n14619_), .ZN(new_n14620_));
  AND3_X2    g11575(.A1(new_n14619_), .A2(pi0792), .A3(new_n14602_), .Z(new_n14621_));
  NOR2_X1    g11576(.A1(new_n14621_), .A2(new_n14620_), .ZN(new_n14622_));
  NAND2_X1   g11577(.A1(new_n14622_), .A2(pi0647), .ZN(new_n14623_));
  XOR2_X1    g11578(.A1(new_n14623_), .A2(new_n14008_), .Z(new_n14624_));
  AOI21_X1   g11579(.A1(new_n14624_), .A2(new_n14478_), .B(new_n14012_), .ZN(new_n14625_));
  AOI21_X1   g11580(.A1(new_n14618_), .A2(new_n14625_), .B(pi0647), .ZN(new_n14626_));
  INV_X1     g11581(.I(new_n14581_), .ZN(new_n14627_));
  NAND2_X1   g11582(.A1(new_n14593_), .A2(pi0788), .ZN(new_n14628_));
  AOI21_X1   g11583(.A1(new_n14590_), .A2(pi0626), .B(new_n13954_), .ZN(new_n14629_));
  INV_X1     g11584(.I(new_n14570_), .ZN(new_n14630_));
  OAI21_X1   g11585(.A1(new_n14629_), .A2(new_n14630_), .B(new_n14478_), .ZN(new_n14631_));
  INV_X1     g11586(.I(new_n14594_), .ZN(new_n14632_));
  NOR2_X1    g11587(.A1(new_n14631_), .A2(new_n14632_), .ZN(new_n14633_));
  NOR2_X1    g11588(.A1(new_n14633_), .A2(new_n14628_), .ZN(new_n14634_));
  NOR3_X1    g11589(.A1(new_n14634_), .A2(new_n13993_), .A3(new_n14627_), .ZN(new_n14635_));
  NOR3_X1    g11590(.A1(new_n14635_), .A2(new_n14005_), .A3(new_n14615_), .ZN(new_n14636_));
  AOI21_X1   g11591(.A1(new_n14622_), .A2(pi1157), .B(new_n14008_), .ZN(new_n14637_));
  NOR4_X1    g11592(.A1(new_n14621_), .A2(pi0647), .A3(new_n14006_), .A4(new_n14620_), .ZN(new_n14638_));
  OAI21_X1   g11593(.A1(new_n14637_), .A2(new_n14638_), .B(new_n14478_), .ZN(new_n14639_));
  NAND2_X1   g11594(.A1(new_n14639_), .A2(new_n14027_), .ZN(new_n14640_));
  OAI21_X1   g11595(.A1(new_n14636_), .A2(new_n14640_), .B(new_n14005_), .ZN(new_n14641_));
  INV_X1     g11596(.I(new_n14641_), .ZN(new_n14642_));
  NOR4_X1    g11597(.A1(new_n14614_), .A2(new_n12776_), .A3(new_n14626_), .A4(new_n14642_), .ZN(new_n14643_));
  NAND4_X1   g11598(.A1(new_n14580_), .A2(new_n14604_), .A3(pi0628), .A4(pi0792), .ZN(new_n14644_));
  NAND2_X1   g11599(.A1(new_n14605_), .A2(new_n14613_), .ZN(new_n14645_));
  AOI21_X1   g11600(.A1(new_n14645_), .A2(new_n14644_), .B(new_n14626_), .ZN(new_n14646_));
  NAND2_X1   g11601(.A1(new_n14641_), .A2(pi0787), .ZN(new_n14647_));
  AOI21_X1   g11602(.A1(new_n14644_), .A2(new_n14645_), .B(new_n14647_), .ZN(new_n14648_));
  NOR3_X1    g11603(.A1(new_n14648_), .A2(new_n12776_), .A3(new_n14646_), .ZN(new_n14649_));
  OAI21_X1   g11604(.A1(new_n14649_), .A2(new_n14643_), .B(new_n12775_), .ZN(new_n14650_));
  NOR2_X1    g11605(.A1(new_n9992_), .A2(pi0141), .ZN(new_n14651_));
  NAND2_X1   g11606(.A1(new_n13218_), .A2(new_n13613_), .ZN(new_n14652_));
  NOR2_X1    g11607(.A1(new_n14652_), .A2(new_n14261_), .ZN(new_n14653_));
  INV_X1     g11608(.I(new_n14651_), .ZN(new_n14654_));
  OAI21_X1   g11609(.A1(new_n13219_), .A2(new_n14261_), .B(new_n14654_), .ZN(new_n14655_));
  NAND3_X1   g11610(.A1(new_n14655_), .A2(new_n14653_), .A3(new_n14651_), .ZN(new_n14656_));
  AOI21_X1   g11611(.A1(new_n13218_), .A2(pi0706), .B(new_n14651_), .ZN(new_n14657_));
  NOR3_X1    g11612(.A1(new_n14653_), .A2(new_n13614_), .A3(new_n14657_), .ZN(new_n14658_));
  XNOR2_X1   g11613(.A1(new_n14656_), .A2(new_n14658_), .ZN(new_n14659_));
  NAND2_X1   g11614(.A1(new_n14659_), .A2(pi0778), .ZN(new_n14660_));
  NAND2_X1   g11615(.A1(new_n14655_), .A2(new_n13748_), .ZN(new_n14661_));
  NAND2_X1   g11616(.A1(new_n14660_), .A2(new_n14661_), .ZN(new_n14662_));
  INV_X1     g11617(.I(new_n14662_), .ZN(new_n14663_));
  NOR2_X1    g11618(.A1(new_n14663_), .A2(new_n14048_), .ZN(new_n14664_));
  INV_X1     g11619(.I(new_n14664_), .ZN(new_n14665_));
  NOR2_X1    g11620(.A1(new_n14665_), .A2(new_n14051_), .ZN(new_n14666_));
  NAND2_X1   g11621(.A1(new_n14666_), .A2(new_n9992_), .ZN(new_n14667_));
  AOI21_X1   g11622(.A1(new_n14667_), .A2(new_n13966_), .B(new_n13919_), .ZN(new_n14668_));
  NAND2_X1   g11623(.A1(new_n14668_), .A2(new_n14061_), .ZN(new_n14669_));
  NAND2_X1   g11624(.A1(new_n14669_), .A2(pi0647), .ZN(new_n14670_));
  XOR2_X1    g11625(.A1(new_n14670_), .A2(new_n14008_), .Z(new_n14671_));
  NAND2_X1   g11626(.A1(new_n14671_), .A2(new_n14651_), .ZN(new_n14672_));
  NAND2_X1   g11627(.A1(new_n14672_), .A2(pi0787), .ZN(new_n14673_));
  NAND2_X1   g11628(.A1(new_n14669_), .A2(pi1157), .ZN(new_n14674_));
  XOR2_X1    g11629(.A1(new_n14674_), .A2(new_n14008_), .Z(new_n14675_));
  NAND2_X1   g11630(.A1(new_n14675_), .A2(new_n14651_), .ZN(new_n14676_));
  NOR3_X1    g11631(.A1(new_n14676_), .A2(new_n12776_), .A3(new_n14669_), .ZN(new_n14677_));
  XOR2_X1    g11632(.A1(new_n14677_), .A2(new_n14673_), .Z(new_n14678_));
  INV_X1     g11633(.I(new_n14666_), .ZN(new_n14679_));
  NAND2_X1   g11634(.A1(new_n14655_), .A2(new_n13103_), .ZN(new_n14680_));
  NOR2_X1    g11635(.A1(new_n14680_), .A2(new_n13613_), .ZN(new_n14681_));
  NAND2_X1   g11636(.A1(new_n14654_), .A2(new_n13614_), .ZN(new_n14682_));
  OAI21_X1   g11637(.A1(new_n14653_), .A2(new_n14682_), .B(pi0608), .ZN(new_n14683_));
  AOI21_X1   g11638(.A1(new_n13104_), .A2(pi0749), .B(new_n14651_), .ZN(new_n14684_));
  NOR2_X1    g11639(.A1(new_n14684_), .A2(pi1153), .ZN(new_n14685_));
  NAND2_X1   g11640(.A1(new_n14683_), .A2(new_n14685_), .ZN(new_n14686_));
  AOI21_X1   g11641(.A1(new_n14686_), .A2(new_n14681_), .B(new_n13748_), .ZN(new_n14687_));
  NOR2_X1    g11642(.A1(new_n14657_), .A2(new_n14082_), .ZN(new_n14688_));
  NAND3_X1   g11643(.A1(new_n14653_), .A2(new_n13614_), .A3(new_n14654_), .ZN(new_n14689_));
  OAI22_X1   g11644(.A1(new_n14689_), .A2(new_n14688_), .B1(new_n14680_), .B2(new_n13613_), .ZN(new_n14690_));
  NAND4_X1   g11645(.A1(new_n14690_), .A2(pi0778), .A3(new_n14680_), .A4(new_n14684_), .ZN(new_n14691_));
  XNOR2_X1   g11646(.A1(new_n14691_), .A2(new_n14687_), .ZN(new_n14692_));
  NAND2_X1   g11647(.A1(new_n14692_), .A2(new_n13801_), .ZN(new_n14693_));
  INV_X1     g11648(.I(new_n14090_), .ZN(new_n14694_));
  NOR2_X1    g11649(.A1(new_n14692_), .A2(new_n13778_), .ZN(new_n14695_));
  XOR2_X1    g11650(.A1(new_n14695_), .A2(new_n14694_), .Z(new_n14696_));
  NOR2_X1    g11651(.A1(new_n14096_), .A2(new_n14684_), .ZN(new_n14697_));
  AOI21_X1   g11652(.A1(new_n14697_), .A2(new_n14094_), .B(pi1155), .ZN(new_n14698_));
  NOR2_X1    g11653(.A1(new_n14698_), .A2(new_n13783_), .ZN(new_n14699_));
  OAI21_X1   g11654(.A1(new_n14696_), .A2(new_n14663_), .B(new_n14699_), .ZN(new_n14700_));
  AOI21_X1   g11655(.A1(new_n14684_), .A2(pi1155), .B(new_n9992_), .ZN(new_n14701_));
  NOR2_X1    g11656(.A1(new_n14701_), .A2(new_n14102_), .ZN(new_n14702_));
  NOR2_X1    g11657(.A1(new_n14702_), .A2(pi0660), .ZN(new_n14703_));
  NAND2_X1   g11658(.A1(new_n14700_), .A2(new_n14703_), .ZN(new_n14704_));
  NOR2_X1    g11659(.A1(new_n14692_), .A2(new_n13766_), .ZN(new_n14705_));
  XOR2_X1    g11660(.A1(new_n14705_), .A2(new_n14090_), .Z(new_n14706_));
  NAND4_X1   g11661(.A1(new_n14704_), .A2(pi0785), .A3(new_n14662_), .A4(new_n14706_), .ZN(new_n14707_));
  NAND2_X1   g11662(.A1(new_n14707_), .A2(new_n14693_), .ZN(new_n14708_));
  NAND2_X1   g11663(.A1(new_n14708_), .A2(new_n13855_), .ZN(new_n14709_));
  NOR2_X1    g11664(.A1(new_n14708_), .A2(new_n13816_), .ZN(new_n14710_));
  XOR2_X1    g11665(.A1(new_n14710_), .A2(new_n13818_), .Z(new_n14711_));
  NOR2_X1    g11666(.A1(new_n14698_), .A2(new_n13801_), .ZN(new_n14712_));
  NAND3_X1   g11667(.A1(new_n14702_), .A2(new_n14697_), .A3(pi0785), .ZN(new_n14713_));
  XOR2_X1    g11668(.A1(new_n14712_), .A2(new_n14713_), .Z(new_n14714_));
  NOR2_X1    g11669(.A1(new_n14714_), .A2(new_n13817_), .ZN(new_n14715_));
  OAI21_X1   g11670(.A1(new_n14715_), .A2(new_n9992_), .B(pi0618), .ZN(new_n14716_));
  NAND2_X1   g11671(.A1(new_n14716_), .A2(new_n13823_), .ZN(new_n14717_));
  AOI21_X1   g11672(.A1(new_n14711_), .A2(new_n14664_), .B(new_n14717_), .ZN(new_n14718_));
  OAI21_X1   g11673(.A1(new_n14715_), .A2(pi0618), .B(new_n9992_), .ZN(new_n14719_));
  NAND2_X1   g11674(.A1(new_n14719_), .A2(new_n13823_), .ZN(new_n14720_));
  NOR2_X1    g11675(.A1(new_n14708_), .A2(new_n13817_), .ZN(new_n14721_));
  XOR2_X1    g11676(.A1(new_n14721_), .A2(new_n13819_), .Z(new_n14722_));
  NOR3_X1    g11677(.A1(new_n14722_), .A2(new_n13855_), .A3(new_n14665_), .ZN(new_n14723_));
  OAI21_X1   g11678(.A1(new_n14718_), .A2(new_n14720_), .B(new_n14723_), .ZN(new_n14724_));
  NAND2_X1   g11679(.A1(new_n14724_), .A2(new_n14709_), .ZN(new_n14725_));
  NOR2_X1    g11680(.A1(new_n14725_), .A2(new_n13860_), .ZN(new_n14726_));
  XOR2_X1    g11681(.A1(new_n14726_), .A2(new_n13904_), .Z(new_n14727_));
  NOR2_X1    g11682(.A1(new_n14727_), .A2(new_n14679_), .ZN(new_n14728_));
  NAND2_X1   g11683(.A1(new_n14719_), .A2(pi0781), .ZN(new_n14729_));
  NOR3_X1    g11684(.A1(new_n14716_), .A2(new_n13855_), .A3(new_n14714_), .ZN(new_n14730_));
  XOR2_X1    g11685(.A1(new_n14730_), .A2(new_n14729_), .Z(new_n14731_));
  NAND2_X1   g11686(.A1(new_n14731_), .A2(pi1159), .ZN(new_n14732_));
  XOR2_X1    g11687(.A1(new_n14732_), .A2(new_n13904_), .Z(new_n14733_));
  NAND2_X1   g11688(.A1(new_n14733_), .A2(new_n14651_), .ZN(new_n14734_));
  NAND2_X1   g11689(.A1(new_n14734_), .A2(new_n13884_), .ZN(new_n14735_));
  INV_X1     g11690(.I(new_n14725_), .ZN(new_n14736_));
  AOI21_X1   g11691(.A1(new_n14736_), .A2(new_n14143_), .B(pi0789), .ZN(new_n14737_));
  OAI21_X1   g11692(.A1(new_n14728_), .A2(new_n14735_), .B(new_n14737_), .ZN(new_n14738_));
  NOR2_X1    g11693(.A1(new_n14725_), .A2(new_n13868_), .ZN(new_n14739_));
  XOR2_X1    g11694(.A1(new_n14739_), .A2(new_n13903_), .Z(new_n14740_));
  NAND2_X1   g11695(.A1(new_n14740_), .A2(new_n14666_), .ZN(new_n14741_));
  NAND2_X1   g11696(.A1(new_n14731_), .A2(pi0619), .ZN(new_n14742_));
  XOR2_X1    g11697(.A1(new_n14742_), .A2(new_n13904_), .Z(new_n14743_));
  NAND2_X1   g11698(.A1(new_n14743_), .A2(new_n14651_), .ZN(new_n14744_));
  NAND4_X1   g11699(.A1(new_n14738_), .A2(pi0648), .A3(new_n14741_), .A4(new_n14744_), .ZN(new_n14745_));
  NAND2_X1   g11700(.A1(new_n14744_), .A2(pi0789), .ZN(new_n14746_));
  NOR3_X1    g11701(.A1(new_n14734_), .A2(new_n13896_), .A3(new_n14731_), .ZN(new_n14747_));
  XOR2_X1    g11702(.A1(new_n14747_), .A2(new_n14746_), .Z(new_n14748_));
  NAND2_X1   g11703(.A1(new_n14748_), .A2(new_n14153_), .ZN(new_n14749_));
  NAND2_X1   g11704(.A1(new_n14153_), .A2(new_n14651_), .ZN(new_n14750_));
  XOR2_X1    g11705(.A1(new_n14749_), .A2(new_n14750_), .Z(new_n14751_));
  AOI21_X1   g11706(.A1(new_n14679_), .A2(new_n14162_), .B(new_n14164_), .ZN(new_n14752_));
  AOI21_X1   g11707(.A1(new_n14752_), .A2(new_n13929_), .B(pi0641), .ZN(new_n14753_));
  OAI21_X1   g11708(.A1(new_n13929_), .A2(new_n14752_), .B(new_n14753_), .ZN(new_n14754_));
  NAND2_X1   g11709(.A1(new_n14751_), .A2(new_n14754_), .ZN(new_n14755_));
  NAND2_X1   g11710(.A1(new_n14755_), .A2(pi0788), .ZN(new_n14756_));
  NAND2_X1   g11711(.A1(new_n14745_), .A2(new_n14756_), .ZN(new_n14757_));
  NOR2_X1    g11712(.A1(new_n14757_), .A2(pi0792), .ZN(new_n14758_));
  NAND2_X1   g11713(.A1(new_n14757_), .A2(pi1156), .ZN(new_n14759_));
  XOR2_X1    g11714(.A1(new_n14759_), .A2(new_n13971_), .Z(new_n14760_));
  NAND2_X1   g11715(.A1(new_n14751_), .A2(pi0788), .ZN(new_n14761_));
  OAI21_X1   g11716(.A1(pi0788), .A2(new_n14748_), .B(new_n14761_), .ZN(new_n14762_));
  OR2_X2     g11717(.A1(new_n14668_), .A2(new_n13977_), .Z(new_n14763_));
  NAND4_X1   g11718(.A1(new_n14760_), .A2(new_n14176_), .A3(new_n14762_), .A4(new_n14763_), .ZN(new_n14764_));
  NAND2_X1   g11719(.A1(new_n14757_), .A2(pi0628), .ZN(new_n14765_));
  XOR2_X1    g11720(.A1(new_n14765_), .A2(new_n13971_), .Z(new_n14766_));
  NAND4_X1   g11721(.A1(new_n14766_), .A2(new_n14181_), .A3(new_n14762_), .A4(new_n14763_), .ZN(new_n14767_));
  AOI21_X1   g11722(.A1(new_n14764_), .A2(new_n14767_), .B(new_n12777_), .ZN(new_n14768_));
  NOR2_X1    g11723(.A1(new_n14768_), .A2(new_n14758_), .ZN(new_n14769_));
  NOR2_X1    g11724(.A1(new_n14762_), .A2(new_n13993_), .ZN(new_n14770_));
  AOI21_X1   g11725(.A1(new_n13993_), .A2(new_n14654_), .B(new_n14770_), .ZN(new_n14771_));
  INV_X1     g11726(.I(new_n14771_), .ZN(new_n14772_));
  NAND2_X1   g11727(.A1(new_n14769_), .A2(pi1157), .ZN(new_n14773_));
  XOR2_X1    g11728(.A1(new_n14773_), .A2(new_n14008_), .Z(new_n14774_));
  NAND2_X1   g11729(.A1(new_n14672_), .A2(pi0630), .ZN(new_n14775_));
  AOI21_X1   g11730(.A1(new_n14774_), .A2(new_n14772_), .B(new_n14775_), .ZN(new_n14776_));
  NAND2_X1   g11731(.A1(new_n14676_), .A2(new_n14010_), .ZN(new_n14777_));
  NOR2_X1    g11732(.A1(new_n14776_), .A2(new_n14777_), .ZN(new_n14778_));
  NAND2_X1   g11733(.A1(new_n14769_), .A2(pi0647), .ZN(new_n14779_));
  XOR2_X1    g11734(.A1(new_n14779_), .A2(new_n14008_), .Z(new_n14780_));
  NAND3_X1   g11735(.A1(new_n14780_), .A2(pi0787), .A3(new_n14772_), .ZN(new_n14781_));
  OAI22_X1   g11736(.A1(new_n14778_), .A2(new_n14781_), .B1(pi0787), .B2(new_n14769_), .ZN(new_n14782_));
  NAND3_X1   g11737(.A1(new_n14782_), .A2(pi0644), .A3(pi0715), .ZN(new_n14783_));
  OR3_X2     g11738(.A1(new_n14782_), .A2(new_n14204_), .A3(new_n14205_), .Z(new_n14784_));
  AOI21_X1   g11739(.A1(new_n14784_), .A2(new_n14783_), .B(new_n14678_), .ZN(new_n14785_));
  NOR2_X1    g11740(.A1(new_n14211_), .A2(new_n14654_), .ZN(new_n14786_));
  AOI21_X1   g11741(.A1(new_n14771_), .A2(new_n14211_), .B(new_n14786_), .ZN(new_n14787_));
  NAND2_X1   g11742(.A1(new_n14787_), .A2(pi0715), .ZN(new_n14788_));
  XOR2_X1    g11743(.A1(new_n14788_), .A2(new_n14205_), .Z(new_n14789_));
  OAI21_X1   g11744(.A1(new_n14789_), .A2(new_n14654_), .B(new_n14203_), .ZN(new_n14790_));
  NAND2_X1   g11745(.A1(new_n14787_), .A2(pi0644), .ZN(new_n14791_));
  XOR2_X1    g11746(.A1(new_n14791_), .A2(new_n14217_), .Z(new_n14792_));
  AOI21_X1   g11747(.A1(new_n14792_), .A2(new_n14651_), .B(pi1160), .ZN(new_n14793_));
  OAI21_X1   g11748(.A1(new_n14785_), .A2(new_n14790_), .B(new_n14793_), .ZN(new_n14794_));
  NAND3_X1   g11749(.A1(new_n14782_), .A2(pi0644), .A3(pi0715), .ZN(new_n14795_));
  OR3_X2     g11750(.A1(new_n14782_), .A2(new_n14200_), .A3(new_n14205_), .Z(new_n14796_));
  AOI21_X1   g11751(.A1(new_n14796_), .A2(new_n14795_), .B(new_n14678_), .ZN(new_n14797_));
  NAND4_X1   g11752(.A1(new_n14794_), .A2(new_n14797_), .A3(pi0790), .A4(pi0832), .ZN(new_n14798_));
  INV_X1     g11753(.I(pi0832), .ZN(new_n14799_));
  NOR2_X1    g11754(.A1(new_n12775_), .A2(new_n14799_), .ZN(new_n14800_));
  INV_X1     g11755(.I(new_n14800_), .ZN(new_n14801_));
  NAND2_X1   g11756(.A1(new_n14794_), .A2(new_n14797_), .ZN(new_n14802_));
  NAND3_X1   g11757(.A1(new_n14802_), .A2(pi0832), .A3(new_n14801_), .ZN(new_n14803_));
  AOI21_X1   g11758(.A1(po1038), .A2(new_n12618_), .B(pi0832), .ZN(new_n14804_));
  NAND2_X1   g11759(.A1(new_n14782_), .A2(new_n14804_), .ZN(new_n14805_));
  AOI21_X1   g11760(.A1(new_n14803_), .A2(new_n14798_), .B(new_n14805_), .ZN(new_n14806_));
  AOI21_X1   g11761(.A1(new_n14650_), .A2(new_n7240_), .B(new_n14806_), .ZN(new_n14807_));
  NOR2_X1    g11762(.A1(new_n14649_), .A2(new_n14643_), .ZN(new_n14808_));
  AOI21_X1   g11763(.A1(new_n14808_), .A2(pi0715), .B(new_n14217_), .ZN(new_n14809_));
  NOR4_X1    g11764(.A1(new_n14649_), .A2(new_n14643_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n14810_));
  NOR2_X1    g11765(.A1(new_n14809_), .A2(new_n14810_), .ZN(new_n14811_));
  OAI21_X1   g11766(.A1(new_n12776_), .A2(new_n14646_), .B(new_n14648_), .ZN(new_n14812_));
  NOR2_X1    g11767(.A1(new_n14646_), .A2(new_n12776_), .ZN(new_n14813_));
  OAI21_X1   g11768(.A1(new_n14614_), .A2(new_n14647_), .B(new_n14813_), .ZN(new_n14814_));
  NOR2_X1    g11769(.A1(new_n14204_), .A2(pi0715), .ZN(new_n14815_));
  NOR2_X1    g11770(.A1(new_n14618_), .A2(new_n14210_), .ZN(new_n14816_));
  AOI21_X1   g11771(.A1(new_n14210_), .A2(new_n14478_), .B(new_n14816_), .ZN(new_n14817_));
  OAI21_X1   g11772(.A1(new_n14454_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n14818_));
  NAND2_X1   g11773(.A1(new_n14817_), .A2(new_n14818_), .ZN(new_n14819_));
  NAND2_X1   g11774(.A1(new_n14624_), .A2(new_n14478_), .ZN(new_n14820_));
  NOR4_X1    g11775(.A1(new_n14820_), .A2(new_n12776_), .A3(new_n14622_), .A4(new_n14639_), .ZN(new_n14821_));
  NAND2_X1   g11776(.A1(new_n14820_), .A2(pi0787), .ZN(new_n14822_));
  NOR3_X1    g11777(.A1(new_n14639_), .A2(new_n12776_), .A3(new_n14622_), .ZN(new_n14823_));
  NOR2_X1    g11778(.A1(new_n14822_), .A2(new_n14823_), .ZN(new_n14824_));
  AOI21_X1   g11779(.A1(new_n14819_), .A2(new_n14815_), .B(pi0644), .ZN(new_n14825_));
  AOI21_X1   g11780(.A1(new_n14814_), .A2(new_n14812_), .B(new_n14825_), .ZN(new_n14826_));
  OAI21_X1   g11781(.A1(new_n14478_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n14827_));
  OAI21_X1   g11782(.A1(new_n14824_), .A2(new_n14821_), .B(new_n14827_), .ZN(new_n14828_));
  NOR2_X1    g11783(.A1(new_n14828_), .A2(new_n14817_), .ZN(new_n14829_));
  OAI21_X1   g11784(.A1(new_n14826_), .A2(pi0790), .B(new_n14829_), .ZN(new_n14830_));
  NOR3_X1    g11785(.A1(new_n14811_), .A2(new_n14807_), .A3(new_n14830_), .ZN(po0298));
  NAND2_X1   g11786(.A1(new_n13086_), .A2(pi0735), .ZN(new_n14832_));
  INV_X1     g11787(.I(pi0735), .ZN(new_n14833_));
  NOR3_X1    g11788(.A1(new_n13672_), .A2(new_n3089_), .A3(new_n14833_), .ZN(new_n14834_));
  XOR2_X1    g11789(.A1(new_n14832_), .A2(new_n14834_), .Z(new_n14835_));
  NOR2_X1    g11790(.A1(new_n3089_), .A2(new_n14833_), .ZN(new_n14836_));
  NOR2_X1    g11791(.A1(new_n12973_), .A2(new_n14833_), .ZN(new_n14837_));
  INV_X1     g11792(.I(new_n14837_), .ZN(new_n14838_));
  NOR2_X1    g11793(.A1(new_n13645_), .A2(new_n3089_), .ZN(new_n14839_));
  INV_X1     g11794(.I(new_n13640_), .ZN(new_n14840_));
  NOR3_X1    g11795(.A1(new_n14840_), .A2(new_n3089_), .A3(new_n13692_), .ZN(new_n14841_));
  XOR2_X1    g11796(.A1(new_n14841_), .A2(new_n14839_), .Z(new_n14842_));
  NAND3_X1   g11797(.A1(new_n14842_), .A2(new_n14836_), .A3(new_n14838_), .ZN(new_n14843_));
  AOI21_X1   g11798(.A1(new_n14842_), .A2(new_n14836_), .B(new_n14838_), .ZN(new_n14844_));
  INV_X1     g11799(.I(new_n14844_), .ZN(new_n14845_));
  NAND2_X1   g11800(.A1(new_n14845_), .A2(new_n14843_), .ZN(new_n14846_));
  NOR2_X1    g11801(.A1(new_n14846_), .A2(new_n5397_), .ZN(new_n14847_));
  NOR2_X1    g11802(.A1(new_n14847_), .A2(new_n12982_), .ZN(new_n14848_));
  INV_X1     g11803(.I(new_n14848_), .ZN(new_n14849_));
  NAND2_X1   g11804(.A1(new_n14847_), .A2(new_n12982_), .ZN(new_n14850_));
  AOI21_X1   g11805(.A1(new_n14849_), .A2(new_n14850_), .B(new_n14835_), .ZN(new_n14851_));
  NOR2_X1    g11806(.A1(new_n12784_), .A2(new_n3089_), .ZN(new_n14852_));
  NAND2_X1   g11807(.A1(new_n13218_), .A2(pi0735), .ZN(new_n14853_));
  INV_X1     g11808(.I(new_n14853_), .ZN(new_n14854_));
  AOI21_X1   g11809(.A1(new_n13677_), .A2(new_n14854_), .B(new_n14852_), .ZN(new_n14855_));
  INV_X1     g11810(.I(new_n14855_), .ZN(new_n14856_));
  NOR2_X1    g11811(.A1(new_n14856_), .A2(new_n3092_), .ZN(new_n14857_));
  OAI21_X1   g11812(.A1(new_n14851_), .A2(pi0223), .B(new_n14857_), .ZN(new_n14858_));
  OAI21_X1   g11813(.A1(new_n13654_), .A2(new_n3089_), .B(pi0735), .ZN(new_n14859_));
  NAND2_X1   g11814(.A1(new_n13076_), .A2(pi0142), .ZN(new_n14860_));
  NAND4_X1   g11815(.A1(new_n13406_), .A2(pi0142), .A3(pi0680), .A4(new_n13394_), .ZN(new_n14861_));
  NOR3_X1    g11816(.A1(new_n14860_), .A2(new_n14833_), .A3(new_n14861_), .ZN(new_n14862_));
  XOR2_X1    g11817(.A1(new_n14862_), .A2(new_n14859_), .Z(new_n14863_));
  AOI21_X1   g11818(.A1(new_n13666_), .A2(pi0142), .B(new_n14833_), .ZN(new_n14864_));
  NOR2_X1    g11819(.A1(new_n13078_), .A2(new_n3089_), .ZN(new_n14865_));
  NOR3_X1    g11820(.A1(new_n14861_), .A2(new_n14833_), .A3(new_n13399_), .ZN(new_n14866_));
  NAND2_X1   g11821(.A1(new_n14865_), .A2(new_n14866_), .ZN(new_n14867_));
  XOR2_X1    g11822(.A1(new_n14867_), .A2(new_n14864_), .Z(new_n14868_));
  NAND2_X1   g11823(.A1(new_n14868_), .A2(pi0223), .ZN(new_n14869_));
  XOR2_X1    g11824(.A1(new_n14869_), .A2(new_n5481_), .Z(new_n14870_));
  NOR2_X1    g11825(.A1(new_n14870_), .A2(new_n14863_), .ZN(new_n14871_));
  INV_X1     g11826(.I(new_n14871_), .ZN(new_n14872_));
  AOI21_X1   g11827(.A1(new_n14858_), .A2(new_n3097_), .B(new_n14872_), .ZN(new_n14873_));
  INV_X1     g11828(.I(new_n14298_), .ZN(new_n14874_));
  NAND2_X1   g11829(.A1(new_n3089_), .A2(new_n14833_), .ZN(new_n14875_));
  AOI21_X1   g11830(.A1(new_n14874_), .A2(new_n14875_), .B(pi0039), .ZN(new_n14876_));
  NOR2_X1    g11831(.A1(new_n3183_), .A2(new_n3089_), .ZN(new_n14877_));
  NOR3_X1    g11832(.A1(new_n9992_), .A2(pi0038), .A3(new_n3183_), .ZN(new_n14878_));
  NAND4_X1   g11833(.A1(new_n3160_), .A2(new_n3089_), .A3(new_n14853_), .A4(new_n14878_), .ZN(new_n14879_));
  NOR2_X1    g11834(.A1(new_n14876_), .A2(new_n14879_), .ZN(new_n14880_));
  NAND3_X1   g11835(.A1(new_n14846_), .A2(new_n3312_), .A3(new_n5454_), .ZN(new_n14881_));
  NAND4_X1   g11836(.A1(new_n14845_), .A2(new_n3313_), .A3(new_n5454_), .A4(new_n14843_), .ZN(new_n14882_));
  NAND2_X1   g11837(.A1(new_n14868_), .A2(pi0215), .ZN(new_n14883_));
  XOR2_X1    g11838(.A1(new_n14883_), .A2(new_n5456_), .Z(new_n14884_));
  NOR2_X1    g11839(.A1(new_n14884_), .A2(new_n14863_), .ZN(new_n14885_));
  INV_X1     g11840(.I(new_n14835_), .ZN(new_n14886_));
  AOI21_X1   g11841(.A1(new_n14855_), .A2(new_n3312_), .B(pi0215), .ZN(new_n14887_));
  NAND2_X1   g11842(.A1(new_n14886_), .A2(new_n14887_), .ZN(new_n14888_));
  INV_X1     g11843(.I(new_n14888_), .ZN(new_n14889_));
  OAI21_X1   g11844(.A1(new_n14885_), .A2(pi0299), .B(new_n14889_), .ZN(new_n14890_));
  AOI21_X1   g11845(.A1(new_n14882_), .A2(new_n14881_), .B(new_n14890_), .ZN(new_n14891_));
  OAI21_X1   g11846(.A1(new_n14873_), .A2(new_n14880_), .B(new_n14891_), .ZN(new_n14892_));
  INV_X1     g11847(.I(new_n11543_), .ZN(new_n14893_));
  NAND3_X1   g11848(.A1(new_n12973_), .A2(pi0142), .A3(new_n5454_), .ZN(new_n14894_));
  NAND3_X1   g11849(.A1(new_n12980_), .A2(pi0142), .A3(new_n5455_), .ZN(new_n14895_));
  NAND2_X1   g11850(.A1(new_n14895_), .A2(new_n14894_), .ZN(new_n14896_));
  AOI21_X1   g11851(.A1(new_n14896_), .A2(new_n12974_), .B(new_n3313_), .ZN(new_n14897_));
  XOR2_X1    g11852(.A1(new_n14897_), .A2(new_n12832_), .Z(new_n14898_));
  INV_X1     g11853(.I(new_n14852_), .ZN(new_n14899_));
  NOR2_X1    g11854(.A1(new_n14865_), .A2(new_n3111_), .ZN(new_n14900_));
  XOR2_X1    g11855(.A1(new_n14900_), .A2(new_n13309_), .Z(new_n14901_));
  NOR4_X1    g11856(.A1(new_n14901_), .A2(new_n3097_), .A3(new_n14899_), .A4(new_n14860_), .ZN(new_n14902_));
  NOR2_X1    g11857(.A1(new_n14365_), .A2(new_n3089_), .ZN(new_n14903_));
  XOR2_X1    g11858(.A1(new_n14903_), .A2(new_n14877_), .Z(new_n14904_));
  AOI22_X1   g11859(.A1(new_n14904_), .A2(new_n14874_), .B1(new_n14898_), .B2(new_n14902_), .ZN(new_n14905_));
  AOI21_X1   g11860(.A1(new_n13625_), .A2(pi0038), .B(new_n3290_), .ZN(new_n14906_));
  OAI22_X1   g11861(.A1(new_n14905_), .A2(new_n14893_), .B1(new_n3089_), .B2(new_n14906_), .ZN(new_n14907_));
  INV_X1     g11862(.I(new_n14907_), .ZN(new_n14908_));
  NAND2_X1   g11863(.A1(new_n14908_), .A2(new_n13613_), .ZN(new_n14909_));
  NOR2_X1    g11864(.A1(new_n3289_), .A2(new_n3089_), .ZN(new_n14910_));
  NOR2_X1    g11865(.A1(new_n14910_), .A2(pi0625), .ZN(new_n14911_));
  INV_X1     g11866(.I(new_n14911_), .ZN(new_n14912_));
  AOI21_X1   g11867(.A1(new_n14909_), .A2(pi1153), .B(new_n14912_), .ZN(new_n14913_));
  OAI21_X1   g11868(.A1(new_n14892_), .A2(new_n14913_), .B(new_n14081_), .ZN(new_n14914_));
  OAI21_X1   g11869(.A1(new_n14351_), .A2(new_n3089_), .B(pi0743), .ZN(new_n14915_));
  INV_X1     g11870(.I(new_n14915_), .ZN(new_n14916_));
  INV_X1     g11871(.I(new_n13405_), .ZN(new_n14917_));
  NAND4_X1   g11872(.A1(new_n13076_), .A2(pi0142), .A3(pi0743), .A4(new_n14917_), .ZN(new_n14918_));
  OR2_X2     g11873(.A1(new_n14918_), .A2(new_n14916_), .Z(new_n14919_));
  NAND2_X1   g11874(.A1(new_n14918_), .A2(new_n14916_), .ZN(new_n14920_));
  INV_X1     g11875(.I(pi0743), .ZN(new_n14921_));
  NOR2_X1    g11876(.A1(new_n14307_), .A2(new_n3089_), .ZN(new_n14922_));
  NOR2_X1    g11877(.A1(new_n14922_), .A2(new_n14921_), .ZN(new_n14923_));
  NAND3_X1   g11878(.A1(new_n14865_), .A2(pi0743), .A3(new_n13392_), .ZN(new_n14924_));
  XNOR2_X1   g11879(.A1(new_n14924_), .A2(new_n14923_), .ZN(new_n14925_));
  NAND3_X1   g11880(.A1(new_n14925_), .A2(pi0215), .A3(new_n5454_), .ZN(new_n14926_));
  XOR2_X1    g11881(.A1(new_n14924_), .A2(new_n14923_), .Z(new_n14927_));
  NAND3_X1   g11882(.A1(new_n14927_), .A2(pi0215), .A3(new_n13309_), .ZN(new_n14928_));
  AOI22_X1   g11883(.A1(new_n14926_), .A2(new_n14928_), .B1(new_n14919_), .B2(new_n14920_), .ZN(new_n14929_));
  NAND2_X1   g11884(.A1(new_n14370_), .A2(new_n14921_), .ZN(new_n14930_));
  NOR2_X1    g11885(.A1(new_n3089_), .A2(new_n14921_), .ZN(new_n14931_));
  INV_X1     g11886(.I(new_n14931_), .ZN(new_n14932_));
  NOR2_X1    g11887(.A1(new_n14320_), .A2(new_n14932_), .ZN(new_n14933_));
  AOI21_X1   g11888(.A1(new_n14933_), .A2(new_n14930_), .B(pi0142), .ZN(new_n14934_));
  NOR2_X1    g11889(.A1(new_n14934_), .A2(new_n13086_), .ZN(new_n14935_));
  INV_X1     g11890(.I(new_n14935_), .ZN(new_n14936_));
  NAND2_X1   g11891(.A1(new_n12980_), .A2(pi0743), .ZN(new_n14937_));
  NAND2_X1   g11892(.A1(new_n14325_), .A2(pi0142), .ZN(new_n14938_));
  NOR2_X1    g11893(.A1(new_n14321_), .A2(new_n3089_), .ZN(new_n14939_));
  NAND3_X1   g11894(.A1(new_n14377_), .A2(new_n14938_), .A3(new_n14939_), .ZN(new_n14940_));
  INV_X1     g11895(.I(new_n14938_), .ZN(new_n14941_));
  INV_X1     g11896(.I(new_n14939_), .ZN(new_n14942_));
  OAI21_X1   g11897(.A1(new_n14382_), .A2(new_n14942_), .B(new_n14941_), .ZN(new_n14943_));
  AOI21_X1   g11898(.A1(new_n14943_), .A2(new_n14940_), .B(new_n14932_), .ZN(new_n14944_));
  NAND2_X1   g11899(.A1(new_n14944_), .A2(new_n14937_), .ZN(new_n14945_));
  NOR3_X1    g11900(.A1(new_n14382_), .A2(new_n14942_), .A3(new_n14941_), .ZN(new_n14946_));
  AOI21_X1   g11901(.A1(new_n14377_), .A2(new_n14939_), .B(new_n14938_), .ZN(new_n14947_));
  OAI21_X1   g11902(.A1(new_n14946_), .A2(new_n14947_), .B(new_n14931_), .ZN(new_n14948_));
  NAND3_X1   g11903(.A1(new_n14948_), .A2(pi0743), .A3(new_n12980_), .ZN(new_n14949_));
  NAND3_X1   g11904(.A1(new_n14949_), .A2(new_n14945_), .A3(new_n5398_), .ZN(new_n14950_));
  NAND2_X1   g11905(.A1(new_n14950_), .A2(new_n12981_), .ZN(new_n14951_));
  NAND4_X1   g11906(.A1(new_n14949_), .A2(new_n14945_), .A3(new_n3092_), .A4(new_n5398_), .ZN(new_n14952_));
  AOI21_X1   g11907(.A1(new_n14951_), .A2(new_n14952_), .B(new_n14936_), .ZN(new_n14953_));
  AOI21_X1   g11908(.A1(pi0743), .A2(new_n13363_), .B(new_n14852_), .ZN(new_n14954_));
  INV_X1     g11909(.I(new_n14954_), .ZN(new_n14955_));
  NOR2_X1    g11910(.A1(new_n14955_), .A2(new_n3092_), .ZN(new_n14956_));
  OAI21_X1   g11911(.A1(new_n14953_), .A2(pi0223), .B(new_n14956_), .ZN(new_n14957_));
  AOI21_X1   g11912(.A1(new_n14927_), .A2(pi0223), .B(new_n13466_), .ZN(new_n14958_));
  NOR3_X1    g11913(.A1(new_n14925_), .A2(new_n3090_), .A3(new_n5398_), .ZN(new_n14959_));
  AOI21_X1   g11914(.A1(new_n14919_), .A2(new_n14920_), .B(new_n3098_), .ZN(new_n14960_));
  OAI21_X1   g11915(.A1(new_n14959_), .A2(new_n14958_), .B(new_n14960_), .ZN(new_n14961_));
  AOI21_X1   g11916(.A1(new_n14957_), .A2(new_n3097_), .B(new_n14961_), .ZN(new_n14962_));
  NAND2_X1   g11917(.A1(new_n14949_), .A2(new_n14945_), .ZN(new_n14963_));
  AOI21_X1   g11918(.A1(new_n14936_), .A2(new_n5455_), .B(new_n3313_), .ZN(new_n14964_));
  OAI21_X1   g11919(.A1(new_n14963_), .A2(new_n5455_), .B(new_n14964_), .ZN(new_n14965_));
  NAND2_X1   g11920(.A1(new_n14965_), .A2(new_n12832_), .ZN(new_n14966_));
  XOR2_X1    g11921(.A1(new_n14944_), .A2(new_n14937_), .Z(new_n14967_));
  NAND2_X1   g11922(.A1(new_n14967_), .A2(new_n5454_), .ZN(new_n14968_));
  NAND3_X1   g11923(.A1(new_n14968_), .A2(new_n12833_), .A3(new_n14964_), .ZN(new_n14969_));
  AOI21_X1   g11924(.A1(new_n14969_), .A2(new_n14966_), .B(new_n14955_), .ZN(new_n14970_));
  OAI21_X1   g11925(.A1(new_n14962_), .A2(new_n14929_), .B(new_n14970_), .ZN(new_n14971_));
  NAND2_X1   g11926(.A1(new_n13171_), .A2(new_n13172_), .ZN(new_n14972_));
  OAI22_X1   g11927(.A1(new_n14972_), .A2(pi0603), .B1(new_n13120_), .B2(new_n13122_), .ZN(new_n14973_));
  NAND2_X1   g11928(.A1(new_n14973_), .A2(pi0743), .ZN(new_n14974_));
  NAND2_X1   g11929(.A1(new_n14974_), .A2(new_n14931_), .ZN(new_n14975_));
  NOR2_X1    g11930(.A1(new_n14974_), .A2(new_n14931_), .ZN(new_n14976_));
  INV_X1     g11931(.I(new_n14976_), .ZN(new_n14977_));
  AOI21_X1   g11932(.A1(new_n14977_), .A2(new_n14975_), .B(new_n13173_), .ZN(new_n14978_));
  INV_X1     g11933(.I(new_n13145_), .ZN(new_n14979_));
  OAI21_X1   g11934(.A1(new_n14979_), .A2(new_n5794_), .B(new_n14336_), .ZN(new_n14980_));
  NOR2_X1    g11935(.A1(new_n14980_), .A2(new_n3089_), .ZN(new_n14981_));
  OR2_X2     g11936(.A1(new_n14336_), .A2(pi0743), .Z(new_n14982_));
  AOI22_X1   g11937(.A1(new_n13192_), .A2(new_n14982_), .B1(pi0142), .B2(new_n14336_), .ZN(new_n14983_));
  NAND3_X1   g11938(.A1(new_n14921_), .A2(pi0142), .A3(pi0299), .ZN(new_n14984_));
  NOR4_X1    g11939(.A1(new_n14981_), .A2(new_n13162_), .A3(new_n14983_), .A4(new_n14984_), .ZN(new_n14985_));
  OAI21_X1   g11940(.A1(new_n14978_), .A2(new_n3098_), .B(new_n14985_), .ZN(new_n14986_));
  INV_X1     g11941(.I(new_n14975_), .ZN(new_n14987_));
  OAI21_X1   g11942(.A1(new_n14987_), .A2(new_n14976_), .B(new_n13174_), .ZN(new_n14988_));
  INV_X1     g11943(.I(new_n14985_), .ZN(new_n14989_));
  NAND3_X1   g11944(.A1(new_n14988_), .A2(pi0299), .A3(new_n14989_), .ZN(new_n14990_));
  NAND2_X1   g11945(.A1(new_n14986_), .A2(new_n14990_), .ZN(new_n14991_));
  AOI21_X1   g11946(.A1(new_n14991_), .A2(new_n3183_), .B(pi0038), .ZN(new_n14992_));
  NOR2_X1    g11947(.A1(new_n14877_), .A2(new_n3259_), .ZN(new_n14993_));
  AOI21_X1   g11948(.A1(new_n3289_), .A2(new_n14993_), .B(pi0039), .ZN(new_n14994_));
  NAND2_X1   g11949(.A1(new_n13104_), .A2(pi0743), .ZN(new_n14995_));
  INV_X1     g11950(.I(new_n14995_), .ZN(new_n14996_));
  NOR4_X1    g11951(.A1(new_n3145_), .A2(pi0142), .A3(new_n9992_), .A4(new_n14996_), .ZN(new_n14997_));
  INV_X1     g11952(.I(new_n14997_), .ZN(new_n14998_));
  NOR2_X1    g11953(.A1(new_n14998_), .A2(new_n14994_), .ZN(new_n14999_));
  INV_X1     g11954(.I(new_n14999_), .ZN(new_n15000_));
  AOI21_X1   g11955(.A1(new_n14971_), .A2(new_n14992_), .B(new_n15000_), .ZN(new_n15001_));
  NOR2_X1    g11956(.A1(new_n15001_), .A2(new_n14430_), .ZN(new_n15002_));
  NAND2_X1   g11957(.A1(new_n13384_), .A2(pi0743), .ZN(new_n15003_));
  XOR2_X1    g11958(.A1(new_n15003_), .A2(new_n14932_), .Z(new_n15004_));
  NAND2_X1   g11959(.A1(new_n13500_), .A2(new_n14921_), .ZN(new_n15005_));
  AOI21_X1   g11960(.A1(new_n3089_), .A2(new_n13306_), .B(new_n15005_), .ZN(new_n15006_));
  AOI21_X1   g11961(.A1(new_n15004_), .A2(new_n15006_), .B(pi0142), .ZN(new_n15007_));
  NAND3_X1   g11962(.A1(new_n13537_), .A2(pi0735), .A3(new_n13539_), .ZN(new_n15008_));
  OAI22_X1   g11963(.A1(new_n15007_), .A2(new_n15008_), .B1(pi0735), .B2(new_n14963_), .ZN(new_n15009_));
  AOI21_X1   g11964(.A1(new_n13269_), .A2(new_n13241_), .B(new_n3089_), .ZN(new_n15010_));
  XOR2_X1    g11965(.A1(new_n15010_), .A2(new_n14931_), .Z(new_n15011_));
  AOI21_X1   g11966(.A1(new_n15011_), .A2(new_n13545_), .B(new_n14833_), .ZN(new_n15012_));
  NAND3_X1   g11967(.A1(new_n13457_), .A2(pi0142), .A3(pi0743), .ZN(new_n15013_));
  OR3_X2     g11968(.A1(new_n13457_), .A2(new_n14921_), .A3(new_n14931_), .Z(new_n15014_));
  NAND2_X1   g11969(.A1(new_n15014_), .A2(new_n15013_), .ZN(new_n15015_));
  NAND4_X1   g11970(.A1(new_n15015_), .A2(pi0735), .A3(new_n13507_), .A4(new_n14935_), .ZN(new_n15016_));
  XOR2_X1    g11971(.A1(new_n15016_), .A2(new_n15012_), .Z(new_n15017_));
  NOR2_X1    g11972(.A1(new_n14852_), .A2(new_n14833_), .ZN(new_n15018_));
  INV_X1     g11973(.I(new_n13463_), .ZN(new_n15019_));
  OAI21_X1   g11974(.A1(new_n15019_), .A2(new_n14998_), .B(new_n13324_), .ZN(new_n15020_));
  NAND4_X1   g11975(.A1(new_n14954_), .A2(pi0735), .A3(new_n12794_), .A4(new_n15020_), .ZN(new_n15021_));
  XOR2_X1    g11976(.A1(new_n15021_), .A2(new_n15018_), .Z(new_n15022_));
  NOR2_X1    g11977(.A1(new_n3312_), .A2(pi0215), .ZN(new_n15023_));
  INV_X1     g11978(.I(new_n15023_), .ZN(new_n15024_));
  OAI21_X1   g11979(.A1(new_n15017_), .A2(new_n15024_), .B(new_n5455_), .ZN(new_n15025_));
  AOI21_X1   g11980(.A1(new_n15025_), .A2(new_n15009_), .B(new_n5827_), .ZN(new_n15026_));
  NAND2_X1   g11981(.A1(new_n13564_), .A2(pi0142), .ZN(new_n15027_));
  XOR2_X1    g11982(.A1(new_n15027_), .A2(new_n14932_), .Z(new_n15028_));
  AOI21_X1   g11983(.A1(new_n15028_), .A2(new_n13342_), .B(new_n14833_), .ZN(new_n15029_));
  NAND2_X1   g11984(.A1(new_n14919_), .A2(new_n14920_), .ZN(new_n15030_));
  NAND2_X1   g11985(.A1(new_n13411_), .A2(pi0743), .ZN(new_n15031_));
  XOR2_X1    g11986(.A1(new_n15031_), .A2(new_n14931_), .Z(new_n15032_));
  NOR3_X1    g11987(.A1(new_n15032_), .A2(new_n14833_), .A3(new_n13475_), .ZN(new_n15033_));
  NAND2_X1   g11988(.A1(new_n15030_), .A2(new_n15033_), .ZN(new_n15034_));
  XNOR2_X1   g11989(.A1(new_n15029_), .A2(new_n15034_), .ZN(new_n15035_));
  NAND2_X1   g11990(.A1(new_n13572_), .A2(pi0142), .ZN(new_n15036_));
  XOR2_X1    g11991(.A1(new_n15036_), .A2(new_n14932_), .Z(new_n15037_));
  AOI21_X1   g11992(.A1(new_n15037_), .A2(new_n13348_), .B(new_n14833_), .ZN(new_n15038_));
  OAI21_X1   g11993(.A1(new_n13445_), .A2(new_n13400_), .B(pi0743), .ZN(new_n15039_));
  XOR2_X1    g11994(.A1(new_n15039_), .A2(new_n14931_), .Z(new_n15040_));
  NOR3_X1    g11995(.A1(new_n15040_), .A2(new_n14833_), .A3(new_n13488_), .ZN(new_n15041_));
  NAND2_X1   g11996(.A1(new_n14925_), .A2(new_n15041_), .ZN(new_n15042_));
  XOR2_X1    g11997(.A1(new_n15038_), .A2(new_n15042_), .Z(new_n15043_));
  AOI21_X1   g11998(.A1(new_n15043_), .A2(pi0215), .B(new_n13309_), .ZN(new_n15044_));
  XNOR2_X1   g11999(.A1(new_n15038_), .A2(new_n15042_), .ZN(new_n15045_));
  NOR3_X1    g12000(.A1(new_n15045_), .A2(new_n3111_), .A3(new_n5456_), .ZN(new_n15046_));
  OAI21_X1   g12001(.A1(new_n15046_), .A2(new_n15044_), .B(new_n15035_), .ZN(new_n15047_));
  NOR2_X1    g12002(.A1(new_n15026_), .A2(new_n15047_), .ZN(new_n15048_));
  INV_X1     g12003(.I(new_n13155_), .ZN(new_n15049_));
  NAND2_X1   g12004(.A1(new_n14980_), .A2(new_n3089_), .ZN(new_n15050_));
  NAND3_X1   g12005(.A1(new_n15050_), .A2(pi0680), .A3(new_n15049_), .ZN(new_n15051_));
  NOR2_X1    g12006(.A1(new_n13150_), .A2(new_n5375_), .ZN(new_n15052_));
  NOR3_X1    g12007(.A1(new_n13192_), .A2(pi0142), .A3(pi0743), .ZN(new_n15053_));
  OAI21_X1   g12008(.A1(new_n15049_), .A2(new_n5375_), .B(new_n13070_), .ZN(new_n15054_));
  NOR2_X1    g12009(.A1(new_n15054_), .A2(new_n15053_), .ZN(new_n15055_));
  OAI21_X1   g12010(.A1(new_n15052_), .A2(new_n15055_), .B(new_n14931_), .ZN(new_n15056_));
  NAND2_X1   g12011(.A1(new_n15056_), .A2(new_n15051_), .ZN(new_n15057_));
  NOR2_X1    g12012(.A1(new_n13174_), .A2(pi0142), .ZN(new_n15058_));
  NAND2_X1   g12013(.A1(new_n15058_), .A2(new_n14921_), .ZN(new_n15059_));
  AOI21_X1   g12014(.A1(new_n13159_), .A2(pi0680), .B(new_n13065_), .ZN(new_n15060_));
  NAND3_X1   g12015(.A1(new_n15059_), .A2(pi0299), .A3(new_n15060_), .ZN(new_n15061_));
  NOR3_X1    g12016(.A1(new_n13141_), .A2(new_n3089_), .A3(new_n5375_), .ZN(new_n15062_));
  INV_X1     g12017(.I(new_n15062_), .ZN(new_n15063_));
  AOI21_X1   g12018(.A1(new_n13137_), .A2(new_n15061_), .B(new_n15063_), .ZN(new_n15064_));
  AOI21_X1   g12019(.A1(new_n15057_), .A2(new_n15064_), .B(pi0743), .ZN(new_n15065_));
  INV_X1     g12020(.I(new_n13134_), .ZN(new_n15066_));
  NOR3_X1    g12021(.A1(new_n15058_), .A2(new_n5375_), .A3(new_n15066_), .ZN(new_n15067_));
  INV_X1     g12022(.I(new_n15067_), .ZN(new_n15068_));
  NOR2_X1    g12023(.A1(new_n15060_), .A2(pi0142), .ZN(new_n15069_));
  AOI21_X1   g12024(.A1(new_n15068_), .A2(new_n15069_), .B(new_n14973_), .ZN(new_n15070_));
  INV_X1     g12025(.I(new_n15070_), .ZN(new_n15071_));
  NOR4_X1    g12026(.A1(new_n15065_), .A2(new_n3183_), .A3(new_n14833_), .A4(new_n15071_), .ZN(new_n15072_));
  NOR2_X1    g12027(.A1(new_n15065_), .A2(new_n15071_), .ZN(new_n15073_));
  NOR3_X1    g12028(.A1(new_n15073_), .A2(pi0039), .A3(new_n14833_), .ZN(new_n15074_));
  NOR2_X1    g12029(.A1(new_n15074_), .A2(new_n15072_), .ZN(new_n15075_));
  AOI21_X1   g12030(.A1(new_n14988_), .A2(pi0299), .B(new_n14989_), .ZN(new_n15076_));
  NOR3_X1    g12031(.A1(new_n14978_), .A2(new_n3098_), .A3(new_n14985_), .ZN(new_n15077_));
  NOR2_X1    g12032(.A1(new_n15077_), .A2(new_n15076_), .ZN(new_n15078_));
  NOR2_X1    g12033(.A1(new_n15078_), .A2(new_n3259_), .ZN(new_n15079_));
  INV_X1     g12034(.I(new_n15079_), .ZN(new_n15080_));
  NOR2_X1    g12035(.A1(new_n15075_), .A2(new_n15080_), .ZN(new_n15081_));
  NOR2_X1    g12036(.A1(new_n15048_), .A2(new_n15081_), .ZN(new_n15082_));
  AND2_X2    g12037(.A1(new_n15022_), .A2(new_n3091_), .Z(new_n15083_));
  AOI21_X1   g12038(.A1(new_n15043_), .A2(pi0223), .B(new_n13466_), .ZN(new_n15084_));
  NOR3_X1    g12039(.A1(new_n15045_), .A2(new_n3090_), .A3(new_n5481_), .ZN(new_n15085_));
  NOR2_X1    g12040(.A1(new_n15085_), .A2(new_n15084_), .ZN(new_n15086_));
  NAND2_X1   g12041(.A1(new_n15035_), .A2(pi0299), .ZN(new_n15087_));
  OAI22_X1   g12042(.A1(new_n15086_), .A2(new_n15087_), .B1(pi0223), .B2(new_n15083_), .ZN(new_n15088_));
  NOR2_X1    g12043(.A1(new_n15009_), .A2(new_n5397_), .ZN(new_n15089_));
  XOR2_X1    g12044(.A1(new_n15089_), .A2(new_n12982_), .Z(new_n15090_));
  NOR2_X1    g12045(.A1(new_n15090_), .A2(new_n15017_), .ZN(new_n15091_));
  NAND2_X1   g12046(.A1(new_n15088_), .A2(new_n15091_), .ZN(new_n15092_));
  NOR3_X1    g12047(.A1(new_n14997_), .A2(pi0735), .A3(new_n13213_), .ZN(new_n15093_));
  NOR3_X1    g12048(.A1(new_n15093_), .A2(new_n14291_), .A3(new_n14994_), .ZN(new_n15094_));
  NAND3_X1   g12049(.A1(new_n15094_), .A2(new_n14910_), .A3(new_n14912_), .ZN(new_n15095_));
  NOR4_X1    g12050(.A1(new_n15082_), .A2(new_n15002_), .A3(new_n15092_), .A4(new_n15095_), .ZN(new_n15096_));
  AOI21_X1   g12051(.A1(new_n14914_), .A2(new_n15096_), .B(new_n13748_), .ZN(new_n15097_));
  INV_X1     g12052(.I(new_n3097_), .ZN(new_n15098_));
  INV_X1     g12053(.I(new_n14850_), .ZN(new_n15099_));
  OAI21_X1   g12054(.A1(new_n15099_), .A2(new_n14848_), .B(new_n14886_), .ZN(new_n15100_));
  INV_X1     g12055(.I(new_n14857_), .ZN(new_n15101_));
  AOI21_X1   g12056(.A1(new_n15100_), .A2(new_n3090_), .B(new_n15101_), .ZN(new_n15102_));
  OAI21_X1   g12057(.A1(new_n15102_), .A2(new_n15098_), .B(new_n14871_), .ZN(new_n15103_));
  INV_X1     g12058(.I(new_n14880_), .ZN(new_n15104_));
  INV_X1     g12059(.I(new_n14891_), .ZN(new_n15105_));
  AOI21_X1   g12060(.A1(new_n15103_), .A2(new_n15104_), .B(new_n15105_), .ZN(new_n15106_));
  NAND2_X1   g12061(.A1(new_n14908_), .A2(pi0625), .ZN(new_n15107_));
  AOI21_X1   g12062(.A1(new_n15107_), .A2(new_n13614_), .B(new_n14912_), .ZN(new_n15108_));
  INV_X1     g12063(.I(new_n15108_), .ZN(new_n15109_));
  AOI21_X1   g12064(.A1(new_n15106_), .A2(new_n15109_), .B(pi0608), .ZN(new_n15110_));
  OAI21_X1   g12065(.A1(new_n15082_), .A2(new_n15092_), .B(new_n15094_), .ZN(new_n15111_));
  NOR2_X1    g12066(.A1(new_n14910_), .A2(new_n13748_), .ZN(new_n15112_));
  NAND3_X1   g12067(.A1(new_n15096_), .A2(new_n15111_), .A3(new_n15112_), .ZN(new_n15113_));
  NOR3_X1    g12068(.A1(new_n15097_), .A2(new_n15110_), .A3(new_n15113_), .ZN(new_n15114_));
  INV_X1     g12069(.I(new_n14913_), .ZN(new_n15115_));
  AOI21_X1   g12070(.A1(new_n15106_), .A2(new_n15115_), .B(pi0608), .ZN(new_n15116_));
  INV_X1     g12071(.I(new_n15096_), .ZN(new_n15117_));
  OAI21_X1   g12072(.A1(new_n15116_), .A2(new_n15117_), .B(pi0778), .ZN(new_n15118_));
  NOR2_X1    g12073(.A1(new_n15113_), .A2(new_n15110_), .ZN(new_n15119_));
  NOR2_X1    g12074(.A1(new_n15118_), .A2(new_n15119_), .ZN(new_n15120_));
  NOR2_X1    g12075(.A1(new_n15120_), .A2(new_n15114_), .ZN(new_n15121_));
  AOI21_X1   g12076(.A1(new_n15106_), .A2(new_n15109_), .B(new_n13748_), .ZN(new_n15122_));
  NAND2_X1   g12077(.A1(new_n14892_), .A2(new_n15112_), .ZN(new_n15123_));
  NOR4_X1    g12078(.A1(new_n15122_), .A2(new_n15123_), .A3(new_n14892_), .A4(new_n14913_), .ZN(new_n15124_));
  NOR2_X1    g12079(.A1(new_n14892_), .A2(new_n14913_), .ZN(new_n15125_));
  OAI21_X1   g12080(.A1(new_n14892_), .A2(new_n15108_), .B(pi0778), .ZN(new_n15126_));
  NOR3_X1    g12081(.A1(new_n15106_), .A2(new_n13748_), .A3(new_n14910_), .ZN(new_n15127_));
  AOI21_X1   g12082(.A1(new_n15125_), .A2(new_n15127_), .B(new_n15126_), .ZN(new_n15128_));
  NOR2_X1    g12083(.A1(new_n15128_), .A2(new_n15124_), .ZN(new_n15129_));
  INV_X1     g12084(.I(new_n14910_), .ZN(new_n15130_));
  INV_X1     g12085(.I(new_n14929_), .ZN(new_n15131_));
  AOI21_X1   g12086(.A1(new_n14967_), .A2(new_n5398_), .B(new_n12982_), .ZN(new_n15132_));
  INV_X1     g12087(.I(new_n14952_), .ZN(new_n15133_));
  OAI21_X1   g12088(.A1(new_n15132_), .A2(new_n15133_), .B(new_n14935_), .ZN(new_n15134_));
  INV_X1     g12089(.I(new_n14956_), .ZN(new_n15135_));
  AOI21_X1   g12090(.A1(new_n15134_), .A2(new_n3090_), .B(new_n15135_), .ZN(new_n15136_));
  NAND3_X1   g12091(.A1(new_n14925_), .A2(pi0223), .A3(new_n5398_), .ZN(new_n15137_));
  NAND3_X1   g12092(.A1(new_n14927_), .A2(pi0223), .A3(new_n5397_), .ZN(new_n15138_));
  INV_X1     g12093(.I(new_n14960_), .ZN(new_n15139_));
  AOI21_X1   g12094(.A1(new_n15137_), .A2(new_n15138_), .B(new_n15139_), .ZN(new_n15140_));
  OAI21_X1   g12095(.A1(new_n15136_), .A2(new_n15098_), .B(new_n15140_), .ZN(new_n15141_));
  INV_X1     g12096(.I(new_n14970_), .ZN(new_n15142_));
  AOI21_X1   g12097(.A1(new_n15141_), .A2(new_n15131_), .B(new_n15142_), .ZN(new_n15143_));
  OAI21_X1   g12098(.A1(new_n15078_), .A2(pi0039), .B(new_n3259_), .ZN(new_n15144_));
  OAI21_X1   g12099(.A1(new_n15143_), .A2(new_n15144_), .B(new_n14999_), .ZN(new_n15145_));
  AOI21_X1   g12100(.A1(new_n15145_), .A2(new_n15130_), .B(new_n13775_), .ZN(new_n15146_));
  INV_X1     g12101(.I(new_n13780_), .ZN(new_n15147_));
  NOR2_X1    g12102(.A1(new_n14908_), .A2(new_n15147_), .ZN(new_n15148_));
  AOI21_X1   g12103(.A1(new_n15129_), .A2(new_n13784_), .B(pi0609), .ZN(new_n15149_));
  OAI21_X1   g12104(.A1(new_n15128_), .A2(new_n15124_), .B(pi0609), .ZN(new_n15150_));
  OAI21_X1   g12105(.A1(new_n15001_), .A2(new_n14910_), .B(new_n13776_), .ZN(new_n15151_));
  AOI21_X1   g12106(.A1(new_n14907_), .A2(new_n14467_), .B(pi0609), .ZN(new_n15152_));
  NOR2_X1    g12107(.A1(new_n15151_), .A2(new_n15152_), .ZN(new_n15153_));
  NOR2_X1    g12108(.A1(new_n15153_), .A2(new_n14465_), .ZN(new_n15154_));
  AOI21_X1   g12109(.A1(new_n15150_), .A2(new_n15154_), .B(pi0609), .ZN(new_n15155_));
  NOR4_X1    g12110(.A1(new_n15155_), .A2(new_n15149_), .A3(new_n15121_), .A4(new_n13801_), .ZN(new_n15156_));
  OAI21_X1   g12111(.A1(new_n15149_), .A2(new_n15121_), .B(pi0785), .ZN(new_n15157_));
  NOR3_X1    g12112(.A1(new_n15155_), .A2(new_n13801_), .A3(new_n15121_), .ZN(new_n15158_));
  NOR2_X1    g12113(.A1(new_n15158_), .A2(new_n15157_), .ZN(new_n15159_));
  NOR2_X1    g12114(.A1(new_n15159_), .A2(new_n15156_), .ZN(new_n15160_));
  OAI21_X1   g12115(.A1(new_n15146_), .A2(new_n15148_), .B(pi0609), .ZN(new_n15161_));
  AOI21_X1   g12116(.A1(new_n14907_), .A2(new_n13775_), .B(new_n13801_), .ZN(new_n15162_));
  NAND3_X1   g12117(.A1(new_n15153_), .A2(new_n15151_), .A3(new_n15162_), .ZN(new_n15163_));
  AOI21_X1   g12118(.A1(pi0785), .A2(new_n15161_), .B(new_n15163_), .ZN(new_n15164_));
  NAND2_X1   g12119(.A1(new_n15161_), .A2(pi0785), .ZN(new_n15165_));
  NAND2_X1   g12120(.A1(new_n15151_), .A2(new_n15162_), .ZN(new_n15166_));
  NOR3_X1    g12121(.A1(new_n15166_), .A2(new_n15151_), .A3(new_n15152_), .ZN(new_n15167_));
  NOR2_X1    g12122(.A1(new_n15165_), .A2(new_n15167_), .ZN(new_n15168_));
  NOR3_X1    g12123(.A1(new_n15164_), .A2(new_n15168_), .A3(new_n13816_), .ZN(new_n15169_));
  NOR2_X1    g12124(.A1(new_n15169_), .A2(new_n13819_), .ZN(new_n15170_));
  NAND2_X1   g12125(.A1(new_n15165_), .A2(new_n15167_), .ZN(new_n15171_));
  NAND3_X1   g12126(.A1(new_n15163_), .A2(pi0785), .A3(new_n15161_), .ZN(new_n15172_));
  NAND2_X1   g12127(.A1(new_n15171_), .A2(new_n15172_), .ZN(new_n15173_));
  NOR3_X1    g12128(.A1(new_n15173_), .A2(new_n13816_), .A3(new_n13818_), .ZN(new_n15174_));
  OAI21_X1   g12129(.A1(new_n15170_), .A2(new_n15174_), .B(new_n14908_), .ZN(new_n15175_));
  NOR2_X1    g12130(.A1(new_n14908_), .A2(new_n13805_), .ZN(new_n15176_));
  AOI21_X1   g12131(.A1(new_n15129_), .A2(new_n13805_), .B(new_n15176_), .ZN(new_n15177_));
  AOI21_X1   g12132(.A1(new_n15177_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n15178_));
  AOI21_X1   g12133(.A1(new_n15178_), .A2(new_n15175_), .B(pi0618), .ZN(new_n15179_));
  OAI21_X1   g12134(.A1(new_n15160_), .A2(new_n15179_), .B(pi0781), .ZN(new_n15180_));
  NOR2_X1    g12135(.A1(new_n15164_), .A2(new_n15168_), .ZN(new_n15181_));
  AOI21_X1   g12136(.A1(new_n15181_), .A2(pi1154), .B(new_n13819_), .ZN(new_n15182_));
  NAND4_X1   g12137(.A1(new_n15171_), .A2(new_n15172_), .A3(new_n13816_), .A4(pi1154), .ZN(new_n15183_));
  INV_X1     g12138(.I(new_n15183_), .ZN(new_n15184_));
  OAI21_X1   g12139(.A1(new_n15182_), .A2(new_n15184_), .B(new_n14908_), .ZN(new_n15185_));
  AOI21_X1   g12140(.A1(new_n15177_), .A2(pi0618), .B(new_n13837_), .ZN(new_n15186_));
  AOI21_X1   g12141(.A1(new_n15186_), .A2(new_n15185_), .B(pi0618), .ZN(new_n15187_));
  NOR3_X1    g12142(.A1(new_n15160_), .A2(new_n13855_), .A3(new_n15187_), .ZN(new_n15188_));
  XOR2_X1    g12143(.A1(new_n15188_), .A2(new_n15180_), .Z(new_n15189_));
  NOR4_X1    g12144(.A1(new_n15185_), .A2(new_n15175_), .A3(new_n13855_), .A4(new_n15181_), .ZN(new_n15190_));
  NAND2_X1   g12145(.A1(new_n15175_), .A2(pi0781), .ZN(new_n15191_));
  NAND2_X1   g12146(.A1(new_n15173_), .A2(pi0781), .ZN(new_n15192_));
  NOR2_X1    g12147(.A1(new_n15185_), .A2(new_n15192_), .ZN(new_n15193_));
  NOR2_X1    g12148(.A1(new_n15193_), .A2(new_n15191_), .ZN(new_n15194_));
  NOR2_X1    g12149(.A1(new_n15194_), .A2(new_n15190_), .ZN(new_n15195_));
  AOI21_X1   g12150(.A1(new_n15195_), .A2(pi0619), .B(new_n13904_), .ZN(new_n15196_));
  NOR4_X1    g12151(.A1(new_n15194_), .A2(new_n13860_), .A3(pi1159), .A4(new_n15190_), .ZN(new_n15197_));
  OAI21_X1   g12152(.A1(new_n15196_), .A2(new_n15197_), .B(new_n14908_), .ZN(new_n15198_));
  NAND2_X1   g12153(.A1(new_n14908_), .A2(new_n13879_), .ZN(new_n15199_));
  NAND2_X1   g12154(.A1(new_n15177_), .A2(new_n13880_), .ZN(new_n15200_));
  NAND2_X1   g12155(.A1(new_n15200_), .A2(new_n15199_), .ZN(new_n15201_));
  AOI21_X1   g12156(.A1(new_n15201_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n15202_));
  AOI21_X1   g12157(.A1(new_n15198_), .A2(new_n15202_), .B(pi0619), .ZN(new_n15203_));
  AOI21_X1   g12158(.A1(new_n15195_), .A2(pi1159), .B(new_n13904_), .ZN(new_n15204_));
  NAND3_X1   g12159(.A1(new_n15173_), .A2(pi0618), .A3(pi1154), .ZN(new_n15205_));
  NAND2_X1   g12160(.A1(new_n15169_), .A2(new_n13819_), .ZN(new_n15206_));
  AOI21_X1   g12161(.A1(new_n15206_), .A2(new_n15205_), .B(new_n14907_), .ZN(new_n15207_));
  NAND3_X1   g12162(.A1(new_n15171_), .A2(new_n15172_), .A3(pi1154), .ZN(new_n15208_));
  NAND2_X1   g12163(.A1(new_n15208_), .A2(new_n13818_), .ZN(new_n15209_));
  AOI21_X1   g12164(.A1(new_n15209_), .A2(new_n15183_), .B(new_n14907_), .ZN(new_n15210_));
  NAND4_X1   g12165(.A1(new_n15207_), .A2(new_n15210_), .A3(pi0781), .A4(new_n15173_), .ZN(new_n15211_));
  NAND3_X1   g12166(.A1(new_n15210_), .A2(pi0781), .A3(new_n15173_), .ZN(new_n15212_));
  NAND3_X1   g12167(.A1(new_n15212_), .A2(pi0781), .A3(new_n15175_), .ZN(new_n15213_));
  NAND4_X1   g12168(.A1(new_n15213_), .A2(new_n15211_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n15214_));
  INV_X1     g12169(.I(new_n15214_), .ZN(new_n15215_));
  OAI21_X1   g12170(.A1(new_n15204_), .A2(new_n15215_), .B(new_n14908_), .ZN(new_n15216_));
  INV_X1     g12171(.I(new_n13892_), .ZN(new_n15217_));
  AOI21_X1   g12172(.A1(new_n15201_), .A2(pi0619), .B(new_n15217_), .ZN(new_n15218_));
  AOI21_X1   g12173(.A1(new_n15216_), .A2(new_n15218_), .B(pi0619), .ZN(new_n15219_));
  NOR4_X1    g12174(.A1(new_n15189_), .A2(new_n13896_), .A3(new_n15203_), .A4(new_n15219_), .ZN(new_n15220_));
  OAI21_X1   g12175(.A1(new_n15189_), .A2(new_n15203_), .B(pi0789), .ZN(new_n15221_));
  NOR3_X1    g12176(.A1(new_n15189_), .A2(new_n13896_), .A3(new_n15219_), .ZN(new_n15222_));
  NOR2_X1    g12177(.A1(new_n15222_), .A2(new_n15221_), .ZN(new_n15223_));
  NOR2_X1    g12178(.A1(new_n15223_), .A2(new_n15220_), .ZN(new_n15224_));
  NOR4_X1    g12179(.A1(new_n15216_), .A2(new_n15198_), .A3(new_n13896_), .A4(new_n15195_), .ZN(new_n15225_));
  NAND2_X1   g12180(.A1(new_n15198_), .A2(pi0789), .ZN(new_n15226_));
  NOR2_X1    g12181(.A1(new_n15195_), .A2(new_n13896_), .ZN(new_n15227_));
  INV_X1     g12182(.I(new_n15227_), .ZN(new_n15228_));
  NOR2_X1    g12183(.A1(new_n15216_), .A2(new_n15228_), .ZN(new_n15229_));
  NOR2_X1    g12184(.A1(new_n15229_), .A2(new_n15226_), .ZN(new_n15230_));
  NOR2_X1    g12185(.A1(new_n15230_), .A2(new_n15225_), .ZN(new_n15231_));
  AOI21_X1   g12186(.A1(new_n15231_), .A2(pi1158), .B(new_n13954_), .ZN(new_n15232_));
  NAND2_X1   g12187(.A1(new_n15213_), .A2(new_n15211_), .ZN(new_n15233_));
  NAND3_X1   g12188(.A1(new_n15233_), .A2(pi0619), .A3(pi1159), .ZN(new_n15234_));
  INV_X1     g12189(.I(new_n15197_), .ZN(new_n15235_));
  AOI21_X1   g12190(.A1(new_n15235_), .A2(new_n15234_), .B(new_n14907_), .ZN(new_n15236_));
  NAND3_X1   g12191(.A1(new_n15233_), .A2(pi0619), .A3(pi1159), .ZN(new_n15237_));
  AOI21_X1   g12192(.A1(new_n15237_), .A2(new_n15214_), .B(new_n14907_), .ZN(new_n15238_));
  NAND4_X1   g12193(.A1(new_n15236_), .A2(new_n15238_), .A3(pi0789), .A4(new_n15233_), .ZN(new_n15239_));
  NAND2_X1   g12194(.A1(new_n15238_), .A2(new_n15227_), .ZN(new_n15240_));
  NAND3_X1   g12195(.A1(new_n15240_), .A2(pi0789), .A3(new_n15198_), .ZN(new_n15241_));
  NAND2_X1   g12196(.A1(new_n15241_), .A2(new_n15239_), .ZN(new_n15242_));
  NOR3_X1    g12197(.A1(new_n15242_), .A2(pi0626), .A3(new_n13929_), .ZN(new_n15243_));
  OAI21_X1   g12198(.A1(new_n15232_), .A2(new_n15243_), .B(new_n14908_), .ZN(new_n15244_));
  NAND2_X1   g12199(.A1(new_n14907_), .A2(new_n13918_), .ZN(new_n15245_));
  NAND3_X1   g12200(.A1(new_n15200_), .A2(new_n13919_), .A3(new_n15199_), .ZN(new_n15246_));
  NAND2_X1   g12201(.A1(new_n15246_), .A2(new_n15245_), .ZN(new_n15247_));
  AOI21_X1   g12202(.A1(new_n15247_), .A2(new_n13901_), .B(new_n13924_), .ZN(new_n15248_));
  NAND2_X1   g12203(.A1(new_n15244_), .A2(new_n15248_), .ZN(new_n15249_));
  NAND3_X1   g12204(.A1(new_n15242_), .A2(pi0626), .A3(pi1158), .ZN(new_n15251_));
  NAND4_X1   g12205(.A1(new_n15241_), .A2(pi0626), .A3(new_n13929_), .A4(new_n15239_), .ZN(new_n15252_));
  AOI21_X1   g12206(.A1(new_n15251_), .A2(new_n15252_), .B(new_n14907_), .ZN(new_n15253_));
  NOR3_X1    g12207(.A1(new_n15224_), .A2(new_n13901_), .A3(new_n13937_), .ZN(new_n15256_));
  AOI21_X1   g12208(.A1(new_n15249_), .A2(new_n13901_), .B(new_n15224_), .ZN(new_n15257_));
  INV_X1     g12209(.I(new_n14577_), .ZN(new_n15258_));
  NOR2_X1    g12210(.A1(new_n15224_), .A2(new_n15258_), .ZN(new_n15259_));
  NOR3_X1    g12211(.A1(new_n15257_), .A2(new_n13937_), .A3(new_n15259_), .ZN(new_n15260_));
  NOR2_X1    g12212(.A1(new_n15260_), .A2(new_n15256_), .ZN(new_n15261_));
  AOI21_X1   g12213(.A1(new_n15231_), .A2(pi0626), .B(new_n13954_), .ZN(new_n15262_));
  INV_X1     g12214(.I(new_n15252_), .ZN(new_n15263_));
  OAI21_X1   g12215(.A1(new_n15262_), .A2(new_n15263_), .B(new_n14908_), .ZN(new_n15264_));
  NOR4_X1    g12216(.A1(new_n15244_), .A2(new_n15264_), .A3(new_n13937_), .A4(new_n15231_), .ZN(new_n15265_));
  NAND2_X1   g12217(.A1(new_n15244_), .A2(pi0788), .ZN(new_n15266_));
  NOR3_X1    g12218(.A1(new_n15264_), .A2(new_n13937_), .A3(new_n15231_), .ZN(new_n15267_));
  NOR2_X1    g12219(.A1(new_n15267_), .A2(new_n15266_), .ZN(new_n15268_));
  NOR2_X1    g12220(.A1(new_n15268_), .A2(new_n15265_), .ZN(new_n15269_));
  INV_X1     g12221(.I(new_n13977_), .ZN(new_n15270_));
  AOI21_X1   g12222(.A1(new_n15246_), .A2(new_n15245_), .B(new_n13965_), .ZN(new_n15271_));
  NOR2_X1    g12223(.A1(new_n14908_), .A2(new_n13966_), .ZN(new_n15272_));
  NOR2_X1    g12224(.A1(new_n15271_), .A2(new_n15272_), .ZN(new_n15273_));
  AOI21_X1   g12225(.A1(new_n15273_), .A2(pi0628), .B(new_n13971_), .ZN(new_n15274_));
  NOR4_X1    g12226(.A1(new_n15271_), .A2(new_n13942_), .A3(pi1156), .A4(new_n15272_), .ZN(new_n15275_));
  OAI21_X1   g12227(.A1(new_n15274_), .A2(new_n15275_), .B(new_n14908_), .ZN(new_n15276_));
  INV_X1     g12228(.I(new_n15276_), .ZN(new_n15277_));
  NOR2_X1    g12229(.A1(new_n15277_), .A2(new_n15270_), .ZN(new_n15278_));
  AOI21_X1   g12230(.A1(new_n15269_), .A2(new_n15278_), .B(pi0628), .ZN(new_n15279_));
  NAND3_X1   g12231(.A1(new_n15242_), .A2(pi0626), .A3(pi1158), .ZN(new_n15280_));
  NAND3_X1   g12232(.A1(new_n15231_), .A2(new_n13901_), .A3(pi1158), .ZN(new_n15281_));
  AOI21_X1   g12233(.A1(new_n15281_), .A2(new_n15280_), .B(new_n14907_), .ZN(new_n15282_));
  NAND4_X1   g12234(.A1(new_n15282_), .A2(new_n15253_), .A3(pi0788), .A4(new_n15242_), .ZN(new_n15283_));
  NOR2_X1    g12235(.A1(new_n15231_), .A2(new_n13937_), .ZN(new_n15284_));
  NAND2_X1   g12236(.A1(new_n15253_), .A2(new_n15284_), .ZN(new_n15285_));
  NAND3_X1   g12237(.A1(new_n15285_), .A2(pi0788), .A3(new_n15244_), .ZN(new_n15286_));
  NAND2_X1   g12238(.A1(new_n15286_), .A2(new_n15283_), .ZN(new_n15287_));
  AOI21_X1   g12239(.A1(new_n15273_), .A2(pi1156), .B(new_n13971_), .ZN(new_n15288_));
  NAND3_X1   g12240(.A1(new_n15273_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n15289_));
  INV_X1     g12241(.I(new_n15289_), .ZN(new_n15290_));
  OAI21_X1   g12242(.A1(new_n15290_), .A2(new_n15288_), .B(new_n14908_), .ZN(new_n15291_));
  NOR4_X1    g12243(.A1(new_n15279_), .A2(new_n15261_), .A3(new_n13942_), .A4(new_n12777_), .ZN(new_n15294_));
  OAI21_X1   g12244(.A1(new_n15279_), .A2(new_n15261_), .B(pi0792), .ZN(new_n15295_));
  INV_X1     g12245(.I(new_n14606_), .ZN(new_n15296_));
  NOR2_X1    g12246(.A1(new_n15261_), .A2(new_n15296_), .ZN(new_n15297_));
  NOR2_X1    g12247(.A1(new_n15295_), .A2(new_n15297_), .ZN(new_n15298_));
  NOR2_X1    g12248(.A1(new_n15298_), .A2(new_n15294_), .ZN(new_n15299_));
  NOR2_X1    g12249(.A1(new_n14908_), .A2(new_n13994_), .ZN(new_n15300_));
  INV_X1     g12250(.I(new_n15300_), .ZN(new_n15301_));
  NAND3_X1   g12251(.A1(new_n15286_), .A2(new_n13994_), .A3(new_n15283_), .ZN(new_n15302_));
  NAND2_X1   g12252(.A1(new_n15302_), .A2(new_n15301_), .ZN(new_n15303_));
  NOR4_X1    g12253(.A1(new_n15291_), .A2(new_n12777_), .A3(new_n15273_), .A4(new_n15276_), .ZN(new_n15304_));
  NOR3_X1    g12254(.A1(new_n15291_), .A2(new_n12777_), .A3(new_n15273_), .ZN(new_n15305_));
  NOR3_X1    g12255(.A1(new_n15305_), .A2(new_n12777_), .A3(new_n15277_), .ZN(new_n15306_));
  NOR2_X1    g12256(.A1(new_n15306_), .A2(new_n15304_), .ZN(new_n15307_));
  AOI21_X1   g12257(.A1(new_n15307_), .A2(pi0647), .B(new_n14008_), .ZN(new_n15308_));
  INV_X1     g12258(.I(new_n15304_), .ZN(new_n15309_));
  INV_X1     g12259(.I(new_n15273_), .ZN(new_n15310_));
  INV_X1     g12260(.I(new_n15288_), .ZN(new_n15311_));
  NAND2_X1   g12261(.A1(new_n15311_), .A2(new_n15289_), .ZN(new_n15312_));
  NAND4_X1   g12262(.A1(new_n15312_), .A2(pi0792), .A3(new_n14908_), .A4(new_n15310_), .ZN(new_n15313_));
  NAND3_X1   g12263(.A1(new_n15313_), .A2(pi0792), .A3(new_n15276_), .ZN(new_n15314_));
  NAND2_X1   g12264(.A1(new_n15314_), .A2(new_n15309_), .ZN(new_n15315_));
  NOR3_X1    g12265(.A1(new_n15315_), .A2(new_n14005_), .A3(pi1157), .ZN(new_n15316_));
  OAI21_X1   g12266(.A1(new_n15308_), .A2(new_n15316_), .B(new_n14908_), .ZN(new_n15317_));
  NAND2_X1   g12267(.A1(new_n15317_), .A2(new_n14011_), .ZN(new_n15318_));
  INV_X1     g12268(.I(new_n15318_), .ZN(new_n15319_));
  AOI21_X1   g12269(.A1(new_n15319_), .A2(new_n15303_), .B(pi0647), .ZN(new_n15320_));
  NOR3_X1    g12270(.A1(new_n15268_), .A2(new_n13993_), .A3(new_n15265_), .ZN(new_n15321_));
  NOR3_X1    g12271(.A1(new_n15321_), .A2(new_n14005_), .A3(new_n15300_), .ZN(new_n15322_));
  AOI21_X1   g12272(.A1(new_n15307_), .A2(pi1157), .B(new_n14008_), .ZN(new_n15323_));
  NAND4_X1   g12273(.A1(new_n15314_), .A2(new_n15309_), .A3(new_n14005_), .A4(pi1157), .ZN(new_n15324_));
  INV_X1     g12274(.I(new_n15324_), .ZN(new_n15325_));
  OAI21_X1   g12275(.A1(new_n15323_), .A2(new_n15325_), .B(new_n14908_), .ZN(new_n15326_));
  NAND2_X1   g12276(.A1(new_n15326_), .A2(new_n14027_), .ZN(new_n15327_));
  OAI21_X1   g12277(.A1(new_n15322_), .A2(new_n15327_), .B(new_n14005_), .ZN(new_n15328_));
  INV_X1     g12278(.I(new_n15328_), .ZN(new_n15329_));
  NOR4_X1    g12279(.A1(new_n15299_), .A2(new_n12776_), .A3(new_n15320_), .A4(new_n15329_), .ZN(new_n15330_));
  INV_X1     g12280(.I(new_n15256_), .ZN(new_n15331_));
  OR2_X2     g12281(.A1(new_n15223_), .A2(new_n15220_), .Z(new_n15332_));
  INV_X1     g12282(.I(new_n15248_), .ZN(new_n15333_));
  OAI21_X1   g12283(.A1(new_n15282_), .A2(new_n15333_), .B(new_n13901_), .ZN(new_n15334_));
  AOI21_X1   g12284(.A1(new_n15332_), .A2(new_n15334_), .B(new_n13937_), .ZN(new_n15335_));
  INV_X1     g12285(.I(new_n15259_), .ZN(new_n15336_));
  NAND2_X1   g12286(.A1(new_n15335_), .A2(new_n15336_), .ZN(new_n15337_));
  NAND2_X1   g12287(.A1(new_n15337_), .A2(new_n15331_), .ZN(new_n15338_));
  INV_X1     g12288(.I(new_n15278_), .ZN(new_n15339_));
  OAI21_X1   g12289(.A1(new_n15287_), .A2(new_n15339_), .B(new_n13942_), .ZN(new_n15340_));
  NAND4_X1   g12290(.A1(new_n15338_), .A2(pi0628), .A3(pi0792), .A4(new_n15340_), .ZN(new_n15341_));
  AOI21_X1   g12291(.A1(new_n15338_), .A2(new_n15340_), .B(new_n12777_), .ZN(new_n15342_));
  NAND2_X1   g12292(.A1(new_n15338_), .A2(new_n14606_), .ZN(new_n15343_));
  NAND2_X1   g12293(.A1(new_n15342_), .A2(new_n15343_), .ZN(new_n15344_));
  AOI21_X1   g12294(.A1(new_n15344_), .A2(new_n15341_), .B(new_n15320_), .ZN(new_n15345_));
  NAND2_X1   g12295(.A1(new_n15328_), .A2(pi0787), .ZN(new_n15346_));
  AOI21_X1   g12296(.A1(new_n15341_), .A2(new_n15344_), .B(new_n15346_), .ZN(new_n15347_));
  NOR3_X1    g12297(.A1(new_n15347_), .A2(new_n15345_), .A3(new_n12776_), .ZN(new_n15348_));
  OAI21_X1   g12298(.A1(new_n15348_), .A2(new_n15330_), .B(new_n12775_), .ZN(new_n15349_));
  NAND2_X1   g12299(.A1(new_n15349_), .A2(new_n5787_), .ZN(new_n15350_));
  NAND2_X1   g12300(.A1(new_n15344_), .A2(new_n15341_), .ZN(new_n15351_));
  NOR2_X1    g12301(.A1(new_n15321_), .A2(new_n15300_), .ZN(new_n15352_));
  OAI21_X1   g12302(.A1(new_n15318_), .A2(new_n15352_), .B(new_n14005_), .ZN(new_n15353_));
  NAND4_X1   g12303(.A1(new_n15351_), .A2(pi0787), .A3(new_n15353_), .A4(new_n15328_), .ZN(new_n15354_));
  OAI21_X1   g12304(.A1(new_n15298_), .A2(new_n15294_), .B(new_n15353_), .ZN(new_n15355_));
  NAND3_X1   g12305(.A1(new_n15302_), .A2(pi0647), .A3(new_n15301_), .ZN(new_n15356_));
  NAND3_X1   g12306(.A1(new_n15356_), .A2(new_n14027_), .A3(new_n15326_), .ZN(new_n15357_));
  AOI21_X1   g12307(.A1(new_n15357_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n15358_));
  OAI21_X1   g12308(.A1(new_n15298_), .A2(new_n15294_), .B(new_n15358_), .ZN(new_n15359_));
  NAND3_X1   g12309(.A1(new_n15359_), .A2(new_n15355_), .A3(pi0787), .ZN(new_n15360_));
  NAND2_X1   g12310(.A1(new_n15360_), .A2(new_n15354_), .ZN(new_n15361_));
  NOR2_X1    g12311(.A1(new_n14907_), .A2(new_n14211_), .ZN(new_n15362_));
  AOI21_X1   g12312(.A1(new_n15352_), .A2(new_n14211_), .B(new_n15362_), .ZN(new_n15363_));
  OR3_X2     g12313(.A1(new_n15363_), .A2(new_n14204_), .A3(new_n14200_), .Z(new_n15364_));
  NAND3_X1   g12314(.A1(new_n15363_), .A2(pi0644), .A3(new_n14200_), .ZN(new_n15365_));
  AOI21_X1   g12315(.A1(new_n15364_), .A2(new_n15365_), .B(new_n14907_), .ZN(new_n15366_));
  NAND3_X1   g12316(.A1(new_n15315_), .A2(pi0647), .A3(pi1157), .ZN(new_n15367_));
  NAND3_X1   g12317(.A1(new_n15307_), .A2(pi0647), .A3(new_n14006_), .ZN(new_n15368_));
  AOI21_X1   g12318(.A1(new_n15368_), .A2(new_n15367_), .B(new_n14907_), .ZN(new_n15369_));
  NAND3_X1   g12319(.A1(new_n15315_), .A2(pi0647), .A3(pi1157), .ZN(new_n15370_));
  AOI21_X1   g12320(.A1(new_n15370_), .A2(new_n15324_), .B(new_n14907_), .ZN(new_n15371_));
  NAND4_X1   g12321(.A1(new_n15369_), .A2(new_n15371_), .A3(pi0787), .A4(new_n15315_), .ZN(new_n15372_));
  NOR2_X1    g12322(.A1(new_n15307_), .A2(new_n12776_), .ZN(new_n15373_));
  NAND2_X1   g12323(.A1(new_n15371_), .A2(new_n15373_), .ZN(new_n15374_));
  NAND3_X1   g12324(.A1(new_n15374_), .A2(pi0787), .A3(new_n15317_), .ZN(new_n15375_));
  NAND2_X1   g12325(.A1(new_n15375_), .A2(new_n15372_), .ZN(new_n15376_));
  NAND2_X1   g12326(.A1(new_n15376_), .A2(new_n14204_), .ZN(new_n15377_));
  NAND2_X1   g12327(.A1(new_n15377_), .A2(new_n14243_), .ZN(new_n15378_));
  OAI21_X1   g12328(.A1(new_n15366_), .A2(new_n15378_), .B(new_n14204_), .ZN(new_n15379_));
  AOI21_X1   g12329(.A1(new_n15361_), .A2(new_n15379_), .B(pi0790), .ZN(new_n15380_));
  INV_X1     g12330(.I(new_n15362_), .ZN(new_n15381_));
  NAND3_X1   g12331(.A1(new_n15302_), .A2(new_n14211_), .A3(new_n15301_), .ZN(new_n15382_));
  NAND3_X1   g12332(.A1(new_n15382_), .A2(pi0715), .A3(new_n15381_), .ZN(new_n15383_));
  XOR2_X1    g12333(.A1(new_n15383_), .A2(new_n14205_), .Z(new_n15384_));
  NOR2_X1    g12334(.A1(pi0715), .A2(pi1160), .ZN(new_n15385_));
  INV_X1     g12335(.I(new_n15385_), .ZN(new_n15386_));
  AOI21_X1   g12336(.A1(new_n15376_), .A2(pi0644), .B(new_n15386_), .ZN(new_n15387_));
  OAI21_X1   g12337(.A1(new_n15384_), .A2(new_n14907_), .B(new_n15387_), .ZN(new_n15388_));
  NAND2_X1   g12338(.A1(new_n5788_), .A2(new_n3089_), .ZN(new_n15389_));
  NOR2_X1    g12339(.A1(new_n9992_), .A2(new_n3089_), .ZN(new_n15390_));
  INV_X1     g12340(.I(new_n15390_), .ZN(new_n15391_));
  NOR2_X1    g12341(.A1(new_n14452_), .A2(new_n13748_), .ZN(new_n15392_));
  NOR2_X1    g12342(.A1(new_n14853_), .A2(new_n15392_), .ZN(new_n15393_));
  NOR2_X1    g12343(.A1(new_n15393_), .A2(new_n15390_), .ZN(new_n15394_));
  NOR2_X1    g12344(.A1(new_n13919_), .A2(new_n13966_), .ZN(new_n15395_));
  NAND3_X1   g12345(.A1(new_n15395_), .A2(new_n13803_), .A3(new_n13879_), .ZN(new_n15396_));
  NOR2_X1    g12346(.A1(new_n15396_), .A2(new_n15394_), .ZN(new_n15397_));
  NOR2_X1    g12347(.A1(new_n14006_), .A2(pi0647), .ZN(new_n15398_));
  NOR2_X1    g12348(.A1(new_n14005_), .A2(pi1157), .ZN(new_n15399_));
  NOR2_X1    g12349(.A1(new_n15398_), .A2(new_n15399_), .ZN(new_n15400_));
  NOR2_X1    g12350(.A1(new_n15400_), .A2(new_n12776_), .ZN(new_n15401_));
  INV_X1     g12351(.I(new_n15401_), .ZN(new_n15402_));
  NAND3_X1   g12352(.A1(new_n15397_), .A2(new_n14059_), .A3(new_n15402_), .ZN(new_n15403_));
  NAND2_X1   g12353(.A1(new_n15403_), .A2(new_n15391_), .ZN(new_n15404_));
  NOR2_X1    g12354(.A1(new_n14995_), .A2(new_n13775_), .ZN(new_n15405_));
  NOR2_X1    g12355(.A1(new_n15405_), .A2(new_n13801_), .ZN(new_n15406_));
  AOI21_X1   g12356(.A1(new_n15391_), .A2(new_n13778_), .B(new_n13766_), .ZN(new_n15407_));
  NAND2_X1   g12357(.A1(new_n15405_), .A2(new_n15407_), .ZN(new_n15408_));
  NAND3_X1   g12358(.A1(new_n15408_), .A2(pi0785), .A3(new_n15390_), .ZN(new_n15409_));
  XOR2_X1    g12359(.A1(new_n15409_), .A2(new_n15406_), .Z(new_n15410_));
  NAND2_X1   g12360(.A1(new_n15410_), .A2(pi0618), .ZN(new_n15411_));
  XOR2_X1    g12361(.A1(new_n15411_), .A2(new_n13819_), .Z(new_n15412_));
  NAND2_X1   g12362(.A1(new_n15412_), .A2(new_n15390_), .ZN(new_n15413_));
  NAND2_X1   g12363(.A1(new_n15413_), .A2(pi0781), .ZN(new_n15414_));
  NAND2_X1   g12364(.A1(new_n15410_), .A2(pi1154), .ZN(new_n15415_));
  XOR2_X1    g12365(.A1(new_n15415_), .A2(new_n13819_), .Z(new_n15416_));
  NAND2_X1   g12366(.A1(new_n15416_), .A2(new_n15390_), .ZN(new_n15417_));
  NOR3_X1    g12367(.A1(new_n15417_), .A2(new_n13855_), .A3(new_n15410_), .ZN(new_n15418_));
  XOR2_X1    g12368(.A1(new_n15418_), .A2(new_n15414_), .Z(new_n15419_));
  NAND2_X1   g12369(.A1(new_n15419_), .A2(pi0619), .ZN(new_n15420_));
  XOR2_X1    g12370(.A1(new_n15420_), .A2(new_n13904_), .Z(new_n15421_));
  NAND2_X1   g12371(.A1(new_n15421_), .A2(new_n15390_), .ZN(new_n15422_));
  NAND2_X1   g12372(.A1(new_n15422_), .A2(pi0789), .ZN(new_n15423_));
  NAND2_X1   g12373(.A1(new_n15419_), .A2(pi1159), .ZN(new_n15424_));
  XOR2_X1    g12374(.A1(new_n15424_), .A2(new_n13904_), .Z(new_n15425_));
  NAND2_X1   g12375(.A1(new_n15425_), .A2(new_n15390_), .ZN(new_n15426_));
  NOR3_X1    g12376(.A1(new_n15426_), .A2(new_n13896_), .A3(new_n15419_), .ZN(new_n15427_));
  XOR2_X1    g12377(.A1(new_n15427_), .A2(new_n15423_), .Z(new_n15428_));
  NOR2_X1    g12378(.A1(new_n15428_), .A2(pi0788), .ZN(new_n15429_));
  NAND2_X1   g12379(.A1(new_n15428_), .A2(new_n14153_), .ZN(new_n15430_));
  NAND2_X1   g12380(.A1(new_n14153_), .A2(new_n15390_), .ZN(new_n15431_));
  XOR2_X1    g12381(.A1(new_n15430_), .A2(new_n15431_), .Z(new_n15432_));
  AOI21_X1   g12382(.A1(new_n15432_), .A2(pi0788), .B(new_n15429_), .ZN(new_n15433_));
  INV_X1     g12383(.I(new_n15433_), .ZN(new_n15434_));
  NOR2_X1    g12384(.A1(new_n15434_), .A2(new_n13993_), .ZN(new_n15435_));
  AOI21_X1   g12385(.A1(new_n13993_), .A2(new_n15391_), .B(new_n15435_), .ZN(new_n15436_));
  NOR2_X1    g12386(.A1(new_n13879_), .A2(new_n13803_), .ZN(new_n15437_));
  NOR3_X1    g12387(.A1(new_n15393_), .A2(new_n15437_), .A3(new_n15390_), .ZN(new_n15438_));
  NAND2_X1   g12388(.A1(new_n14995_), .A2(new_n15391_), .ZN(new_n15439_));
  NAND4_X1   g12389(.A1(new_n15439_), .A2(new_n13220_), .A3(pi0735), .A4(new_n13748_), .ZN(new_n15440_));
  NAND3_X1   g12390(.A1(new_n15439_), .A2(new_n13220_), .A3(pi0735), .ZN(new_n15441_));
  NAND3_X1   g12391(.A1(new_n13220_), .A2(pi0625), .A3(pi0735), .ZN(new_n15442_));
  NAND2_X1   g12392(.A1(new_n15441_), .A2(new_n15442_), .ZN(new_n15443_));
  AOI21_X1   g12393(.A1(new_n15443_), .A2(new_n13614_), .B(new_n14081_), .ZN(new_n15444_));
  INV_X1     g12394(.I(new_n15442_), .ZN(new_n15445_));
  NOR2_X1    g12395(.A1(new_n13613_), .A2(new_n13614_), .ZN(new_n15446_));
  NOR2_X1    g12396(.A1(new_n15390_), .A2(pi1153), .ZN(new_n15447_));
  NAND2_X1   g12397(.A1(pi0608), .A2(pi0625), .ZN(new_n15448_));
  NOR4_X1    g12398(.A1(new_n14853_), .A2(new_n14995_), .A3(new_n15447_), .A4(new_n15448_), .ZN(new_n15449_));
  OAI21_X1   g12399(.A1(new_n15445_), .A2(new_n15446_), .B(new_n15449_), .ZN(new_n15450_));
  XOR2_X1    g12400(.A1(new_n15444_), .A2(new_n15450_), .Z(new_n15451_));
  OAI21_X1   g12401(.A1(new_n15451_), .A2(new_n13748_), .B(new_n15440_), .ZN(new_n15452_));
  NAND2_X1   g12402(.A1(new_n15452_), .A2(new_n13801_), .ZN(new_n15453_));
  NOR2_X1    g12403(.A1(new_n15452_), .A2(new_n13766_), .ZN(new_n15454_));
  XOR2_X1    g12404(.A1(new_n15454_), .A2(new_n14090_), .Z(new_n15455_));
  NAND4_X1   g12405(.A1(new_n15455_), .A2(new_n13783_), .A3(new_n15394_), .A4(new_n15408_), .ZN(new_n15456_));
  NOR2_X1    g12406(.A1(new_n15452_), .A2(new_n13778_), .ZN(new_n15457_));
  XOR2_X1    g12407(.A1(new_n15457_), .A2(new_n14694_), .Z(new_n15458_));
  INV_X1     g12408(.I(new_n15458_), .ZN(new_n15459_));
  NAND4_X1   g12409(.A1(new_n15456_), .A2(pi0785), .A3(new_n15394_), .A4(new_n15459_), .ZN(new_n15460_));
  NAND2_X1   g12410(.A1(new_n15460_), .A2(new_n15453_), .ZN(new_n15461_));
  NAND2_X1   g12411(.A1(new_n15461_), .A2(new_n13855_), .ZN(new_n15462_));
  AOI21_X1   g12412(.A1(new_n15393_), .A2(new_n13805_), .B(new_n15390_), .ZN(new_n15463_));
  NOR2_X1    g12413(.A1(new_n15461_), .A2(new_n13816_), .ZN(new_n15464_));
  XOR2_X1    g12414(.A1(new_n15464_), .A2(new_n13818_), .Z(new_n15465_));
  NAND2_X1   g12415(.A1(new_n15417_), .A2(new_n13823_), .ZN(new_n15466_));
  AOI21_X1   g12416(.A1(new_n15465_), .A2(new_n15463_), .B(new_n15466_), .ZN(new_n15467_));
  NAND2_X1   g12417(.A1(new_n15413_), .A2(new_n13823_), .ZN(new_n15468_));
  NOR2_X1    g12418(.A1(new_n15461_), .A2(new_n13817_), .ZN(new_n15469_));
  XOR2_X1    g12419(.A1(new_n15469_), .A2(new_n13819_), .Z(new_n15470_));
  NAND2_X1   g12420(.A1(new_n15463_), .A2(pi0781), .ZN(new_n15471_));
  NOR2_X1    g12421(.A1(new_n15470_), .A2(new_n15471_), .ZN(new_n15472_));
  OAI21_X1   g12422(.A1(new_n15467_), .A2(new_n15468_), .B(new_n15472_), .ZN(new_n15473_));
  NAND2_X1   g12423(.A1(new_n15473_), .A2(new_n15462_), .ZN(new_n15474_));
  NOR2_X1    g12424(.A1(new_n15474_), .A2(new_n13860_), .ZN(new_n15475_));
  XOR2_X1    g12425(.A1(new_n15475_), .A2(new_n13903_), .Z(new_n15476_));
  NAND2_X1   g12426(.A1(new_n15426_), .A2(new_n13884_), .ZN(new_n15477_));
  AOI21_X1   g12427(.A1(new_n15476_), .A2(new_n15438_), .B(new_n15477_), .ZN(new_n15478_));
  INV_X1     g12428(.I(new_n14143_), .ZN(new_n15479_));
  OAI21_X1   g12429(.A1(new_n15474_), .A2(new_n15479_), .B(new_n13896_), .ZN(new_n15480_));
  NOR2_X1    g12430(.A1(new_n15478_), .A2(new_n15480_), .ZN(new_n15481_));
  NOR2_X1    g12431(.A1(new_n15474_), .A2(new_n13868_), .ZN(new_n15482_));
  XOR2_X1    g12432(.A1(new_n15482_), .A2(new_n13903_), .Z(new_n15483_));
  NAND2_X1   g12433(.A1(new_n15483_), .A2(new_n15438_), .ZN(new_n15484_));
  NAND3_X1   g12434(.A1(new_n15484_), .A2(pi0648), .A3(new_n15422_), .ZN(new_n15485_));
  NOR3_X1    g12435(.A1(new_n13919_), .A2(new_n14162_), .A3(new_n15391_), .ZN(new_n15486_));
  AOI21_X1   g12436(.A1(new_n15486_), .A2(new_n13929_), .B(pi0641), .ZN(new_n15487_));
  OAI21_X1   g12437(.A1(new_n13929_), .A2(new_n15486_), .B(new_n15487_), .ZN(new_n15488_));
  AND2_X2    g12438(.A1(new_n15432_), .A2(new_n15488_), .Z(new_n15489_));
  OAI22_X1   g12439(.A1(new_n15481_), .A2(new_n15485_), .B1(new_n13937_), .B2(new_n15489_), .ZN(new_n15490_));
  NAND2_X1   g12440(.A1(new_n15490_), .A2(pi1156), .ZN(new_n15491_));
  XOR2_X1    g12441(.A1(new_n15491_), .A2(new_n13970_), .Z(new_n15492_));
  NOR2_X1    g12442(.A1(new_n15492_), .A2(new_n15433_), .ZN(new_n15493_));
  NAND2_X1   g12443(.A1(new_n15397_), .A2(new_n13942_), .ZN(new_n15494_));
  AND3_X2    g12444(.A1(new_n15494_), .A2(pi1156), .A3(new_n15391_), .Z(new_n15495_));
  OAI21_X1   g12445(.A1(new_n15493_), .A2(pi0629), .B(new_n15495_), .ZN(new_n15496_));
  NAND2_X1   g12446(.A1(new_n15490_), .A2(pi0628), .ZN(new_n15497_));
  XOR2_X1    g12447(.A1(new_n15497_), .A2(new_n13970_), .Z(new_n15498_));
  NOR2_X1    g12448(.A1(new_n15498_), .A2(new_n15433_), .ZN(new_n15499_));
  NAND2_X1   g12449(.A1(new_n15397_), .A2(pi0628), .ZN(new_n15500_));
  NAND4_X1   g12450(.A1(new_n15500_), .A2(pi0792), .A3(pi1156), .A4(new_n15391_), .ZN(new_n15501_));
  NOR2_X1    g12451(.A1(new_n15490_), .A2(new_n15501_), .ZN(new_n15502_));
  OAI21_X1   g12452(.A1(new_n15499_), .A2(pi0629), .B(new_n15502_), .ZN(new_n15503_));
  AOI21_X1   g12453(.A1(pi0792), .A2(new_n15496_), .B(new_n15503_), .ZN(new_n15504_));
  NAND3_X1   g12454(.A1(new_n15496_), .A2(new_n15503_), .A3(pi0792), .ZN(new_n15505_));
  INV_X1     g12455(.I(new_n15505_), .ZN(new_n15506_));
  NOR2_X1    g12456(.A1(new_n15506_), .A2(new_n15504_), .ZN(new_n15507_));
  AOI21_X1   g12457(.A1(new_n15507_), .A2(pi1157), .B(new_n14008_), .ZN(new_n15508_));
  INV_X1     g12458(.I(new_n15507_), .ZN(new_n15509_));
  NOR3_X1    g12459(.A1(new_n15509_), .A2(pi0647), .A3(new_n14006_), .ZN(new_n15510_));
  NOR2_X1    g12460(.A1(new_n15510_), .A2(new_n15508_), .ZN(new_n15511_));
  NOR2_X1    g12461(.A1(new_n15511_), .A2(new_n15436_), .ZN(new_n15512_));
  NAND2_X1   g12462(.A1(new_n15391_), .A2(new_n14006_), .ZN(new_n15513_));
  NAND4_X1   g12463(.A1(new_n15397_), .A2(pi0647), .A3(new_n14059_), .A4(new_n15513_), .ZN(new_n15514_));
  INV_X1     g12464(.I(new_n15514_), .ZN(new_n15515_));
  NOR2_X1    g12465(.A1(new_n15515_), .A2(new_n14010_), .ZN(new_n15516_));
  INV_X1     g12466(.I(new_n15516_), .ZN(new_n15517_));
  NOR2_X1    g12467(.A1(new_n15515_), .A2(pi0630), .ZN(new_n15518_));
  OAI21_X1   g12468(.A1(new_n15512_), .A2(new_n15517_), .B(new_n15518_), .ZN(new_n15519_));
  NOR2_X1    g12469(.A1(new_n15509_), .A2(new_n14005_), .ZN(new_n15520_));
  XOR2_X1    g12470(.A1(new_n15520_), .A2(new_n14007_), .Z(new_n15521_));
  NOR2_X1    g12471(.A1(new_n15436_), .A2(new_n12776_), .ZN(new_n15522_));
  NAND3_X1   g12472(.A1(new_n15519_), .A2(new_n15521_), .A3(new_n15522_), .ZN(new_n15523_));
  NAND2_X1   g12473(.A1(new_n15507_), .A2(new_n12776_), .ZN(new_n15524_));
  NAND2_X1   g12474(.A1(new_n15523_), .A2(new_n15524_), .ZN(new_n15525_));
  NAND3_X1   g12475(.A1(new_n15525_), .A2(pi0644), .A3(pi0715), .ZN(new_n15526_));
  NAND4_X1   g12476(.A1(new_n15523_), .A2(pi0644), .A3(new_n14200_), .A4(new_n15524_), .ZN(new_n15527_));
  AOI21_X1   g12477(.A1(new_n15526_), .A2(new_n15527_), .B(new_n15404_), .ZN(new_n15528_));
  NOR2_X1    g12478(.A1(new_n14211_), .A2(new_n15391_), .ZN(new_n15529_));
  AOI21_X1   g12479(.A1(new_n15436_), .A2(new_n14211_), .B(new_n15529_), .ZN(new_n15530_));
  NAND2_X1   g12480(.A1(new_n15530_), .A2(pi0715), .ZN(new_n15531_));
  XOR2_X1    g12481(.A1(new_n15531_), .A2(new_n14205_), .Z(new_n15532_));
  OAI21_X1   g12482(.A1(new_n15532_), .A2(new_n15391_), .B(new_n14203_), .ZN(new_n15533_));
  NAND2_X1   g12483(.A1(new_n15530_), .A2(pi0644), .ZN(new_n15534_));
  XOR2_X1    g12484(.A1(new_n15534_), .A2(new_n14217_), .Z(new_n15535_));
  AOI21_X1   g12485(.A1(new_n15535_), .A2(new_n15390_), .B(pi1160), .ZN(new_n15536_));
  OAI21_X1   g12486(.A1(new_n15528_), .A2(new_n15533_), .B(new_n15536_), .ZN(new_n15537_));
  NAND3_X1   g12487(.A1(new_n15525_), .A2(pi0644), .A3(pi0715), .ZN(new_n15538_));
  NAND4_X1   g12488(.A1(new_n15523_), .A2(new_n14204_), .A3(pi0715), .A4(new_n15524_), .ZN(new_n15539_));
  AOI21_X1   g12489(.A1(new_n15538_), .A2(new_n15539_), .B(new_n15404_), .ZN(new_n15540_));
  NAND4_X1   g12490(.A1(new_n15537_), .A2(pi0790), .A3(new_n15540_), .A4(pi0832), .ZN(new_n15541_));
  NAND2_X1   g12491(.A1(new_n15537_), .A2(new_n15540_), .ZN(new_n15542_));
  NAND3_X1   g12492(.A1(new_n15542_), .A2(new_n12775_), .A3(pi0832), .ZN(new_n15543_));
  NAND2_X1   g12493(.A1(new_n15543_), .A2(new_n15541_), .ZN(new_n15544_));
  NAND2_X1   g12494(.A1(pi0057), .A2(pi0142), .ZN(new_n15545_));
  AND3_X2    g12495(.A1(new_n15525_), .A2(new_n14799_), .A3(new_n15545_), .Z(new_n15546_));
  AOI22_X1   g12496(.A1(new_n15544_), .A2(new_n15546_), .B1(new_n5371_), .B2(new_n15389_), .ZN(new_n15547_));
  AOI21_X1   g12497(.A1(new_n15388_), .A2(new_n14204_), .B(new_n15547_), .ZN(new_n15548_));
  NAND2_X1   g12498(.A1(new_n15361_), .A2(new_n15548_), .ZN(new_n15549_));
  AOI21_X1   g12499(.A1(new_n15350_), .A2(new_n15380_), .B(new_n15549_), .ZN(po0299));
  NOR3_X1    g12500(.A1(new_n13632_), .A2(new_n3259_), .A3(new_n10708_), .ZN(new_n15551_));
  NAND4_X1   g12501(.A1(new_n13073_), .A2(new_n13096_), .A3(pi0038), .A4(new_n10708_), .ZN(new_n15552_));
  INV_X1     g12502(.I(new_n15552_), .ZN(new_n15553_));
  OAI21_X1   g12503(.A1(new_n15551_), .A2(new_n15553_), .B(new_n13624_), .ZN(new_n15554_));
  AOI21_X1   g12504(.A1(new_n5503_), .A2(new_n13310_), .B(new_n3259_), .ZN(new_n15555_));
  AOI21_X1   g12505(.A1(new_n14362_), .A2(new_n3259_), .B(new_n15555_), .ZN(new_n15556_));
  NOR2_X1    g12506(.A1(new_n14380_), .A2(new_n3183_), .ZN(new_n15557_));
  NAND2_X1   g12507(.A1(new_n14388_), .A2(pi0039), .ZN(new_n15558_));
  NOR3_X1    g12508(.A1(new_n15558_), .A2(new_n13180_), .A3(new_n15557_), .ZN(new_n15559_));
  NOR3_X1    g12509(.A1(new_n13180_), .A2(new_n3183_), .A3(new_n14387_), .ZN(new_n15560_));
  NOR3_X1    g12510(.A1(new_n15560_), .A2(new_n3183_), .A3(new_n14380_), .ZN(new_n15561_));
  NOR2_X1    g12511(.A1(new_n15561_), .A2(new_n15559_), .ZN(new_n15562_));
  NAND4_X1   g12512(.A1(new_n5492_), .A2(pi0038), .A3(pi0143), .A4(new_n13104_), .ZN(new_n15563_));
  OAI21_X1   g12513(.A1(pi0143), .A2(pi0774), .B(new_n15563_), .ZN(new_n15564_));
  AOI21_X1   g12514(.A1(new_n15556_), .A2(new_n15564_), .B(new_n3290_), .ZN(new_n15565_));
  INV_X1     g12515(.I(new_n15565_), .ZN(new_n15566_));
  AOI21_X1   g12516(.A1(new_n15554_), .A2(pi0774), .B(new_n15566_), .ZN(new_n15567_));
  NOR2_X1    g12517(.A1(new_n3289_), .A2(pi0143), .ZN(new_n15568_));
  NOR2_X1    g12518(.A1(new_n15567_), .A2(new_n15568_), .ZN(new_n15569_));
  NAND3_X1   g12519(.A1(new_n13097_), .A2(pi0038), .A3(pi0143), .ZN(new_n15570_));
  AOI21_X1   g12520(.A1(new_n15570_), .A2(new_n15552_), .B(new_n13625_), .ZN(new_n15571_));
  INV_X1     g12521(.I(pi0687), .ZN(new_n15572_));
  INV_X1     g12522(.I(pi0774), .ZN(new_n15573_));
  NAND2_X1   g12523(.A1(new_n15556_), .A2(new_n15564_), .ZN(new_n15574_));
  AOI21_X1   g12524(.A1(new_n15574_), .A2(new_n15572_), .B(new_n15573_), .ZN(new_n15575_));
  AOI21_X1   g12525(.A1(new_n15571_), .A2(new_n15575_), .B(new_n3290_), .ZN(new_n15576_));
  INV_X1     g12526(.I(new_n15576_), .ZN(new_n15577_));
  NAND2_X1   g12527(.A1(new_n14272_), .A2(new_n3183_), .ZN(new_n15578_));
  NAND2_X1   g12528(.A1(new_n15578_), .A2(pi0038), .ZN(new_n15579_));
  INV_X1     g12529(.I(new_n15579_), .ZN(new_n15580_));
  NOR2_X1    g12530(.A1(new_n13537_), .A2(new_n13586_), .ZN(new_n15581_));
  OAI21_X1   g12531(.A1(new_n13580_), .A2(new_n13583_), .B(new_n15581_), .ZN(new_n15582_));
  AOI21_X1   g12532(.A1(new_n15582_), .A2(pi0039), .B(new_n11324_), .ZN(new_n15583_));
  NOR3_X1    g12533(.A1(new_n13587_), .A2(new_n3183_), .A3(pi0299), .ZN(new_n15584_));
  OAI21_X1   g12534(.A1(new_n15584_), .A2(new_n15583_), .B(new_n13605_), .ZN(new_n15585_));
  NOR2_X1    g12535(.A1(new_n13109_), .A2(new_n13213_), .ZN(new_n15586_));
  INV_X1     g12536(.I(new_n15586_), .ZN(new_n15587_));
  NOR2_X1    g12537(.A1(new_n15587_), .A2(new_n3259_), .ZN(new_n15588_));
  INV_X1     g12538(.I(new_n15588_), .ZN(new_n15589_));
  NOR3_X1    g12539(.A1(new_n15585_), .A2(new_n15580_), .A3(new_n15589_), .ZN(new_n15590_));
  NAND3_X1   g12540(.A1(new_n13587_), .A2(pi0039), .A3(pi0299), .ZN(new_n15591_));
  NAND3_X1   g12541(.A1(new_n15582_), .A2(pi0039), .A3(new_n3098_), .ZN(new_n15592_));
  AOI21_X1   g12542(.A1(new_n15591_), .A2(new_n15592_), .B(new_n13577_), .ZN(new_n15593_));
  AOI21_X1   g12543(.A1(new_n15593_), .A2(new_n15588_), .B(new_n15579_), .ZN(new_n15594_));
  NOR2_X1    g12544(.A1(new_n15594_), .A2(new_n15590_), .ZN(new_n15595_));
  INV_X1     g12545(.I(new_n13511_), .ZN(new_n15596_));
  INV_X1     g12546(.I(new_n13520_), .ZN(new_n15597_));
  NOR2_X1    g12547(.A1(new_n13209_), .A2(new_n3183_), .ZN(new_n15598_));
  NOR2_X1    g12548(.A1(new_n3259_), .A2(pi0039), .ZN(new_n15599_));
  INV_X1     g12549(.I(new_n15599_), .ZN(new_n15600_));
  NOR2_X1    g12550(.A1(new_n13209_), .A2(new_n15600_), .ZN(new_n15601_));
  INV_X1     g12551(.I(new_n15601_), .ZN(new_n15602_));
  AOI21_X1   g12552(.A1(new_n13190_), .A2(new_n15598_), .B(new_n15602_), .ZN(new_n15603_));
  INV_X1     g12553(.I(new_n15598_), .ZN(new_n15604_));
  NOR4_X1    g12554(.A1(new_n13189_), .A2(new_n13187_), .A3(new_n15604_), .A4(new_n15601_), .ZN(new_n15605_));
  OAI21_X1   g12555(.A1(new_n15603_), .A2(new_n15605_), .B(pi0039), .ZN(new_n15606_));
  AOI21_X1   g12556(.A1(new_n15606_), .A2(new_n15596_), .B(new_n15597_), .ZN(new_n15607_));
  NOR2_X1    g12557(.A1(new_n15572_), .A2(pi0774), .ZN(new_n15608_));
  AOI21_X1   g12558(.A1(new_n15607_), .A2(new_n15608_), .B(pi0143), .ZN(new_n15609_));
  INV_X1     g12559(.I(new_n15609_), .ZN(new_n15610_));
  NAND3_X1   g12560(.A1(new_n13359_), .A2(pi0038), .A3(pi0039), .ZN(new_n15611_));
  INV_X1     g12561(.I(new_n13356_), .ZN(new_n15612_));
  NOR4_X1    g12562(.A1(new_n15612_), .A2(pi0038), .A3(new_n3183_), .A4(new_n13357_), .ZN(new_n15613_));
  INV_X1     g12563(.I(new_n15613_), .ZN(new_n15614_));
  AOI21_X1   g12564(.A1(new_n15614_), .A2(new_n15611_), .B(new_n13152_), .ZN(new_n15615_));
  AOI21_X1   g12565(.A1(new_n13198_), .A2(new_n3183_), .B(new_n3259_), .ZN(new_n15616_));
  INV_X1     g12566(.I(new_n15616_), .ZN(new_n15617_));
  AOI21_X1   g12567(.A1(new_n13434_), .A2(pi0039), .B(pi0299), .ZN(new_n15618_));
  NOR2_X1    g12568(.A1(new_n13452_), .A2(new_n15618_), .ZN(new_n15619_));
  NOR2_X1    g12569(.A1(new_n5504_), .A2(new_n13221_), .ZN(new_n15620_));
  INV_X1     g12570(.I(new_n15620_), .ZN(new_n15621_));
  NOR2_X1    g12571(.A1(new_n15621_), .A2(new_n3259_), .ZN(new_n15622_));
  NAND3_X1   g12572(.A1(new_n15619_), .A2(new_n15617_), .A3(new_n15622_), .ZN(new_n15623_));
  OAI21_X1   g12573(.A1(new_n13458_), .A2(new_n3183_), .B(new_n3098_), .ZN(new_n15624_));
  NAND2_X1   g12574(.A1(new_n13460_), .A2(new_n15624_), .ZN(new_n15625_));
  INV_X1     g12575(.I(new_n15622_), .ZN(new_n15626_));
  OAI21_X1   g12576(.A1(new_n15625_), .A2(new_n15626_), .B(new_n15616_), .ZN(new_n15627_));
  NAND2_X1   g12577(.A1(new_n15623_), .A2(new_n15627_), .ZN(new_n15628_));
  NOR3_X1    g12578(.A1(new_n14291_), .A2(new_n4368_), .A3(new_n13324_), .ZN(new_n15629_));
  INV_X1     g12579(.I(new_n15629_), .ZN(new_n15630_));
  AOI21_X1   g12580(.A1(new_n15630_), .A2(new_n15573_), .B(new_n10708_), .ZN(new_n15631_));
  NAND4_X1   g12581(.A1(new_n15610_), .A2(new_n15615_), .A3(new_n15628_), .A4(new_n15631_), .ZN(new_n15632_));
  NOR2_X1    g12582(.A1(new_n3290_), .A2(new_n10708_), .ZN(new_n15633_));
  INV_X1     g12583(.I(new_n15633_), .ZN(new_n15634_));
  AOI21_X1   g12584(.A1(new_n15632_), .A2(new_n15595_), .B(new_n15634_), .ZN(new_n15635_));
  NAND2_X1   g12585(.A1(new_n15635_), .A2(new_n15577_), .ZN(new_n15636_));
  NAND3_X1   g12586(.A1(new_n15593_), .A2(new_n15579_), .A3(new_n15588_), .ZN(new_n15637_));
  OAI21_X1   g12587(.A1(new_n15585_), .A2(new_n15589_), .B(new_n15580_), .ZN(new_n15638_));
  NAND2_X1   g12588(.A1(new_n15637_), .A2(new_n15638_), .ZN(new_n15639_));
  NOR3_X1    g12589(.A1(new_n15612_), .A2(new_n3183_), .A3(new_n13357_), .ZN(new_n15640_));
  NOR2_X1    g12590(.A1(new_n15640_), .A2(new_n4368_), .ZN(new_n15641_));
  OAI21_X1   g12591(.A1(new_n15641_), .A2(new_n15613_), .B(new_n14269_), .ZN(new_n15642_));
  NAND2_X1   g12592(.A1(new_n15628_), .A2(new_n15631_), .ZN(new_n15643_));
  NOR3_X1    g12593(.A1(new_n15643_), .A2(new_n15642_), .A3(new_n15609_), .ZN(new_n15644_));
  OAI21_X1   g12594(.A1(new_n15644_), .A2(new_n15639_), .B(new_n15633_), .ZN(new_n15645_));
  NAND2_X1   g12595(.A1(new_n15645_), .A2(new_n15576_), .ZN(new_n15646_));
  NAND3_X1   g12596(.A1(new_n15636_), .A2(new_n15646_), .A3(pi1153), .ZN(new_n15647_));
  NAND2_X1   g12597(.A1(new_n15647_), .A2(new_n13615_), .ZN(new_n15648_));
  NOR2_X1    g12598(.A1(new_n15645_), .A2(new_n15576_), .ZN(new_n15649_));
  NOR2_X1    g12599(.A1(new_n15635_), .A2(new_n15577_), .ZN(new_n15650_));
  NOR3_X1    g12600(.A1(new_n15650_), .A2(new_n15649_), .A3(new_n13614_), .ZN(new_n15651_));
  NAND2_X1   g12601(.A1(new_n15651_), .A2(new_n13620_), .ZN(new_n15652_));
  AOI21_X1   g12602(.A1(new_n15652_), .A2(new_n15648_), .B(new_n15569_), .ZN(new_n15653_));
  AOI21_X1   g12603(.A1(new_n13634_), .A2(new_n3289_), .B(pi0143), .ZN(new_n15654_));
  XOR2_X1    g12604(.A1(new_n14403_), .A2(new_n14401_), .Z(new_n15655_));
  NOR3_X1    g12605(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n10708_), .ZN(new_n15656_));
  NAND4_X1   g12606(.A1(new_n14421_), .A2(new_n14413_), .A3(new_n3259_), .A4(pi0143), .ZN(new_n15657_));
  INV_X1     g12607(.I(new_n15657_), .ZN(new_n15658_));
  OAI21_X1   g12608(.A1(new_n15656_), .A2(new_n15658_), .B(new_n15655_), .ZN(new_n15659_));
  NOR2_X1    g12609(.A1(new_n13721_), .A2(new_n15572_), .ZN(new_n15660_));
  OAI21_X1   g12610(.A1(new_n15660_), .A2(pi0143), .B(new_n13108_), .ZN(new_n15661_));
  INV_X1     g12611(.I(new_n15661_), .ZN(new_n15662_));
  AOI21_X1   g12612(.A1(new_n15659_), .A2(new_n15662_), .B(new_n3290_), .ZN(new_n15663_));
  NAND4_X1   g12613(.A1(new_n15571_), .A2(pi0143), .A3(new_n15572_), .A4(new_n3289_), .ZN(new_n15664_));
  NOR2_X1    g12614(.A1(new_n15663_), .A2(new_n15664_), .ZN(new_n15665_));
  NAND3_X1   g12615(.A1(new_n14422_), .A2(pi0038), .A3(pi0143), .ZN(new_n15666_));
  AOI21_X1   g12616(.A1(new_n15666_), .A2(new_n15657_), .B(new_n14404_), .ZN(new_n15667_));
  OAI21_X1   g12617(.A1(new_n15667_), .A2(new_n15661_), .B(new_n3289_), .ZN(new_n15668_));
  NOR4_X1    g12618(.A1(new_n15554_), .A2(new_n10708_), .A3(pi0687), .A4(new_n3290_), .ZN(new_n15669_));
  NOR2_X1    g12619(.A1(new_n15668_), .A2(new_n15669_), .ZN(new_n15670_));
  NOR3_X1    g12620(.A1(new_n15665_), .A2(new_n13613_), .A3(new_n15670_), .ZN(new_n15671_));
  NOR2_X1    g12621(.A1(new_n15671_), .A2(new_n13620_), .ZN(new_n15672_));
  XOR2_X1    g12622(.A1(new_n15668_), .A2(new_n15664_), .Z(new_n15673_));
  NOR3_X1    g12623(.A1(new_n15673_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n15674_));
  OAI21_X1   g12624(.A1(new_n15674_), .A2(new_n15672_), .B(new_n15654_), .ZN(new_n15675_));
  NAND2_X1   g12625(.A1(new_n15675_), .A2(pi0608), .ZN(new_n15676_));
  OAI21_X1   g12626(.A1(new_n15653_), .A2(new_n15676_), .B(pi0778), .ZN(new_n15677_));
  NOR2_X1    g12627(.A1(new_n15650_), .A2(new_n15649_), .ZN(new_n15678_));
  NAND3_X1   g12628(.A1(new_n15636_), .A2(new_n15646_), .A3(pi0625), .ZN(new_n15679_));
  NAND2_X1   g12629(.A1(new_n15679_), .A2(new_n13615_), .ZN(new_n15680_));
  NAND3_X1   g12630(.A1(new_n15678_), .A2(pi0625), .A3(new_n13620_), .ZN(new_n15681_));
  AOI21_X1   g12631(.A1(new_n15681_), .A2(new_n15680_), .B(new_n15569_), .ZN(new_n15682_));
  INV_X1     g12632(.I(new_n15654_), .ZN(new_n15683_));
  NAND3_X1   g12633(.A1(new_n15673_), .A2(pi0625), .A3(pi1153), .ZN(new_n15684_));
  NOR2_X1    g12634(.A1(new_n15665_), .A2(new_n15670_), .ZN(new_n15685_));
  NAND3_X1   g12635(.A1(new_n15685_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n15686_));
  AOI21_X1   g12636(.A1(new_n15684_), .A2(new_n15686_), .B(new_n15683_), .ZN(new_n15687_));
  NOR4_X1    g12637(.A1(new_n15682_), .A2(new_n13750_), .A3(new_n15678_), .A4(new_n15687_), .ZN(new_n15688_));
  XOR2_X1    g12638(.A1(new_n15688_), .A2(new_n15677_), .Z(new_n15689_));
  NOR2_X1    g12639(.A1(new_n15685_), .A2(new_n13748_), .ZN(new_n15690_));
  NAND2_X1   g12640(.A1(new_n15687_), .A2(new_n15690_), .ZN(new_n15691_));
  AOI21_X1   g12641(.A1(pi0778), .A2(new_n15675_), .B(new_n15691_), .ZN(new_n15692_));
  NAND3_X1   g12642(.A1(new_n15691_), .A2(pi0778), .A3(new_n15675_), .ZN(new_n15693_));
  INV_X1     g12643(.I(new_n15693_), .ZN(new_n15694_));
  NOR2_X1    g12644(.A1(new_n15694_), .A2(new_n15692_), .ZN(new_n15695_));
  NOR3_X1    g12645(.A1(new_n15567_), .A2(new_n13775_), .A3(new_n15568_), .ZN(new_n15696_));
  NOR2_X1    g12646(.A1(new_n15654_), .A2(new_n15147_), .ZN(new_n15697_));
  AOI21_X1   g12647(.A1(new_n15695_), .A2(new_n13784_), .B(pi0609), .ZN(new_n15699_));
  OAI21_X1   g12648(.A1(new_n15689_), .A2(new_n15699_), .B(pi0785), .ZN(new_n15700_));
  NAND2_X1   g12649(.A1(new_n15675_), .A2(pi0778), .ZN(new_n15701_));
  NAND3_X1   g12650(.A1(new_n15701_), .A2(new_n15687_), .A3(new_n15690_), .ZN(new_n15702_));
  AOI21_X1   g12651(.A1(new_n15702_), .A2(new_n15693_), .B(new_n13766_), .ZN(new_n15703_));
  OAI21_X1   g12652(.A1(new_n15571_), .A2(new_n15573_), .B(new_n15565_), .ZN(new_n15704_));
  INV_X1     g12653(.I(new_n15568_), .ZN(new_n15705_));
  NAND3_X1   g12654(.A1(new_n15704_), .A2(new_n13776_), .A3(new_n15705_), .ZN(new_n15706_));
  INV_X1     g12655(.I(new_n14467_), .ZN(new_n15707_));
  OAI21_X1   g12656(.A1(new_n15654_), .A2(new_n15707_), .B(new_n13766_), .ZN(new_n15708_));
  INV_X1     g12657(.I(new_n15708_), .ZN(new_n15709_));
  NOR2_X1    g12658(.A1(new_n15706_), .A2(new_n15709_), .ZN(new_n15710_));
  NOR2_X1    g12659(.A1(new_n15710_), .A2(new_n14465_), .ZN(new_n15711_));
  INV_X1     g12660(.I(new_n15711_), .ZN(new_n15712_));
  OAI21_X1   g12661(.A1(new_n15703_), .A2(new_n15712_), .B(new_n13766_), .ZN(new_n15713_));
  INV_X1     g12662(.I(new_n15713_), .ZN(new_n15714_));
  NOR3_X1    g12663(.A1(new_n15714_), .A2(new_n15689_), .A3(new_n13801_), .ZN(new_n15715_));
  NAND2_X1   g12664(.A1(new_n15715_), .A2(new_n15700_), .ZN(new_n15716_));
  NAND2_X1   g12665(.A1(new_n15688_), .A2(new_n15677_), .ZN(new_n15717_));
  NAND2_X1   g12666(.A1(new_n15704_), .A2(new_n15705_), .ZN(new_n15718_));
  NOR2_X1    g12667(.A1(new_n15651_), .A2(new_n13620_), .ZN(new_n15719_));
  NOR2_X1    g12668(.A1(new_n15647_), .A2(new_n13615_), .ZN(new_n15720_));
  OAI21_X1   g12669(.A1(new_n15719_), .A2(new_n15720_), .B(new_n15718_), .ZN(new_n15721_));
  INV_X1     g12670(.I(new_n15676_), .ZN(new_n15722_));
  AOI21_X1   g12671(.A1(new_n15722_), .A2(new_n15721_), .B(new_n13748_), .ZN(new_n15723_));
  AND2_X2    g12672(.A1(new_n15681_), .A2(new_n15680_), .Z(new_n15724_));
  NOR3_X1    g12673(.A1(new_n15687_), .A2(new_n13750_), .A3(new_n15678_), .ZN(new_n15725_));
  OAI21_X1   g12674(.A1(new_n15724_), .A2(new_n15569_), .B(new_n15725_), .ZN(new_n15726_));
  NAND2_X1   g12675(.A1(new_n15723_), .A2(new_n15726_), .ZN(new_n15727_));
  NAND2_X1   g12676(.A1(new_n15727_), .A2(new_n15717_), .ZN(new_n15728_));
  NAND2_X1   g12677(.A1(new_n15702_), .A2(new_n15693_), .ZN(new_n15729_));
  OAI21_X1   g12678(.A1(new_n15729_), .A2(new_n13785_), .B(new_n13766_), .ZN(new_n15730_));
  AOI21_X1   g12679(.A1(new_n15728_), .A2(new_n15730_), .B(new_n13801_), .ZN(new_n15731_));
  NAND3_X1   g12680(.A1(new_n15728_), .A2(new_n15713_), .A3(pi0785), .ZN(new_n15732_));
  NAND2_X1   g12681(.A1(new_n15731_), .A2(new_n15732_), .ZN(new_n15733_));
  NAND2_X1   g12682(.A1(new_n15716_), .A2(new_n15733_), .ZN(new_n15734_));
  INV_X1     g12683(.I(new_n15697_), .ZN(new_n15735_));
  AOI21_X1   g12684(.A1(new_n15706_), .A2(new_n15735_), .B(new_n13766_), .ZN(new_n15736_));
  NAND2_X1   g12685(.A1(new_n15654_), .A2(new_n13775_), .ZN(new_n15737_));
  OAI21_X1   g12686(.A1(new_n15569_), .A2(new_n13775_), .B(new_n15737_), .ZN(new_n15738_));
  NAND4_X1   g12687(.A1(new_n15738_), .A2(new_n15736_), .A3(new_n15710_), .A4(pi0785), .ZN(new_n15739_));
  NOR2_X1    g12688(.A1(new_n15736_), .A2(new_n13801_), .ZN(new_n15740_));
  NAND3_X1   g12689(.A1(new_n15738_), .A2(new_n15710_), .A3(pi0785), .ZN(new_n15741_));
  NAND2_X1   g12690(.A1(new_n15741_), .A2(new_n15740_), .ZN(new_n15742_));
  NAND2_X1   g12691(.A1(new_n15742_), .A2(new_n15739_), .ZN(new_n15743_));
  NAND3_X1   g12692(.A1(new_n15743_), .A2(pi0618), .A3(pi1154), .ZN(new_n15744_));
  OAI21_X1   g12693(.A1(new_n15696_), .A2(new_n15697_), .B(pi0609), .ZN(new_n15745_));
  NAND4_X1   g12694(.A1(new_n15708_), .A2(new_n15704_), .A3(new_n13776_), .A4(new_n15705_), .ZN(new_n15746_));
  INV_X1     g12695(.I(new_n15737_), .ZN(new_n15747_));
  AOI21_X1   g12696(.A1(new_n15718_), .A2(new_n13776_), .B(new_n15747_), .ZN(new_n15748_));
  NOR4_X1    g12697(.A1(new_n15745_), .A2(new_n13801_), .A3(new_n15748_), .A4(new_n15746_), .ZN(new_n15749_));
  NAND2_X1   g12698(.A1(new_n15745_), .A2(pi0785), .ZN(new_n15750_));
  NOR3_X1    g12699(.A1(new_n15748_), .A2(new_n13801_), .A3(new_n15746_), .ZN(new_n15751_));
  NOR2_X1    g12700(.A1(new_n15750_), .A2(new_n15751_), .ZN(new_n15752_));
  NOR4_X1    g12701(.A1(new_n15752_), .A2(new_n13816_), .A3(pi1154), .A4(new_n15749_), .ZN(new_n15753_));
  INV_X1     g12702(.I(new_n15753_), .ZN(new_n15754_));
  AOI21_X1   g12703(.A1(new_n15754_), .A2(new_n15744_), .B(new_n15683_), .ZN(new_n15755_));
  AOI21_X1   g12704(.A1(new_n15702_), .A2(new_n15693_), .B(new_n13803_), .ZN(new_n15756_));
  NOR2_X1    g12705(.A1(new_n15683_), .A2(new_n13805_), .ZN(new_n15757_));
  NOR2_X1    g12706(.A1(new_n15756_), .A2(new_n15757_), .ZN(new_n15758_));
  OAI21_X1   g12707(.A1(new_n15758_), .A2(pi0618), .B(new_n13824_), .ZN(new_n15759_));
  OAI21_X1   g12708(.A1(new_n15759_), .A2(new_n15755_), .B(new_n13816_), .ZN(new_n15760_));
  NOR2_X1    g12709(.A1(new_n15752_), .A2(new_n15749_), .ZN(new_n15761_));
  AOI21_X1   g12710(.A1(new_n15761_), .A2(pi1154), .B(new_n13819_), .ZN(new_n15762_));
  NAND4_X1   g12711(.A1(new_n15742_), .A2(new_n13816_), .A3(pi1154), .A4(new_n15739_), .ZN(new_n15763_));
  INV_X1     g12712(.I(new_n15763_), .ZN(new_n15764_));
  OAI21_X1   g12713(.A1(new_n15762_), .A2(new_n15764_), .B(new_n15654_), .ZN(new_n15765_));
  OAI21_X1   g12714(.A1(new_n15756_), .A2(new_n15757_), .B(pi0618), .ZN(new_n15766_));
  NAND3_X1   g12715(.A1(new_n15766_), .A2(new_n13836_), .A3(new_n15765_), .ZN(new_n15767_));
  NAND2_X1   g12716(.A1(new_n15767_), .A2(new_n13816_), .ZN(new_n15768_));
  NAND4_X1   g12717(.A1(new_n15734_), .A2(pi0781), .A3(new_n15760_), .A4(new_n15768_), .ZN(new_n15769_));
  NOR2_X1    g12718(.A1(new_n15731_), .A2(new_n15732_), .ZN(new_n15770_));
  NOR2_X1    g12719(.A1(new_n15715_), .A2(new_n15700_), .ZN(new_n15771_));
  OAI21_X1   g12720(.A1(new_n15771_), .A2(new_n15770_), .B(new_n15760_), .ZN(new_n15772_));
  AOI21_X1   g12721(.A1(new_n15767_), .A2(new_n13816_), .B(new_n13855_), .ZN(new_n15773_));
  OAI21_X1   g12722(.A1(new_n15771_), .A2(new_n15770_), .B(new_n15773_), .ZN(new_n15774_));
  NAND3_X1   g12723(.A1(new_n15772_), .A2(new_n15774_), .A3(pi0781), .ZN(new_n15775_));
  NAND2_X1   g12724(.A1(new_n15775_), .A2(new_n15769_), .ZN(new_n15776_));
  NAND3_X1   g12725(.A1(new_n15743_), .A2(pi0618), .A3(pi1154), .ZN(new_n15777_));
  AOI21_X1   g12726(.A1(new_n15777_), .A2(new_n15763_), .B(new_n15683_), .ZN(new_n15778_));
  NAND4_X1   g12727(.A1(new_n15755_), .A2(new_n15778_), .A3(pi0781), .A4(new_n15743_), .ZN(new_n15779_));
  AOI21_X1   g12728(.A1(new_n15761_), .A2(pi0618), .B(new_n13819_), .ZN(new_n15780_));
  OAI21_X1   g12729(.A1(new_n15780_), .A2(new_n15753_), .B(new_n15654_), .ZN(new_n15781_));
  NOR2_X1    g12730(.A1(new_n15761_), .A2(new_n13855_), .ZN(new_n15782_));
  NAND2_X1   g12731(.A1(new_n15778_), .A2(new_n15782_), .ZN(new_n15783_));
  NAND3_X1   g12732(.A1(new_n15783_), .A2(pi0781), .A3(new_n15781_), .ZN(new_n15784_));
  NAND2_X1   g12733(.A1(new_n15784_), .A2(new_n15779_), .ZN(new_n15785_));
  NAND3_X1   g12734(.A1(new_n15785_), .A2(pi0619), .A3(pi1159), .ZN(new_n15786_));
  NOR4_X1    g12735(.A1(new_n15765_), .A2(new_n15781_), .A3(new_n13855_), .A4(new_n15761_), .ZN(new_n15787_));
  NAND2_X1   g12736(.A1(new_n15781_), .A2(pi0781), .ZN(new_n15788_));
  INV_X1     g12737(.I(new_n15782_), .ZN(new_n15789_));
  NOR2_X1    g12738(.A1(new_n15765_), .A2(new_n15789_), .ZN(new_n15790_));
  NOR2_X1    g12739(.A1(new_n15790_), .A2(new_n15788_), .ZN(new_n15791_));
  NOR4_X1    g12740(.A1(new_n15791_), .A2(new_n13860_), .A3(pi1159), .A4(new_n15787_), .ZN(new_n15792_));
  INV_X1     g12741(.I(new_n15792_), .ZN(new_n15793_));
  AOI21_X1   g12742(.A1(new_n15793_), .A2(new_n15786_), .B(new_n15683_), .ZN(new_n15794_));
  NOR2_X1    g12743(.A1(new_n15654_), .A2(new_n13880_), .ZN(new_n15795_));
  AOI21_X1   g12744(.A1(new_n15758_), .A2(new_n13880_), .B(new_n15795_), .ZN(new_n15796_));
  NAND2_X1   g12745(.A1(new_n15796_), .A2(new_n13860_), .ZN(new_n15797_));
  NAND2_X1   g12746(.A1(new_n15797_), .A2(new_n13885_), .ZN(new_n15798_));
  OAI21_X1   g12747(.A1(new_n15794_), .A2(new_n15798_), .B(new_n13860_), .ZN(new_n15799_));
  NAND3_X1   g12748(.A1(new_n15785_), .A2(pi0619), .A3(pi1159), .ZN(new_n15800_));
  NAND4_X1   g12749(.A1(new_n15784_), .A2(new_n13860_), .A3(pi1159), .A4(new_n15779_), .ZN(new_n15801_));
  AOI21_X1   g12750(.A1(new_n15800_), .A2(new_n15801_), .B(new_n15683_), .ZN(new_n15802_));
  NAND2_X1   g12751(.A1(new_n15796_), .A2(pi0619), .ZN(new_n15803_));
  NAND2_X1   g12752(.A1(new_n15803_), .A2(new_n13892_), .ZN(new_n15804_));
  OAI21_X1   g12753(.A1(new_n15802_), .A2(new_n15804_), .B(new_n13860_), .ZN(new_n15805_));
  NAND4_X1   g12754(.A1(new_n15776_), .A2(pi0789), .A3(new_n15799_), .A4(new_n15805_), .ZN(new_n15806_));
  NAND2_X1   g12755(.A1(new_n15776_), .A2(new_n15799_), .ZN(new_n15807_));
  NAND3_X1   g12756(.A1(new_n15776_), .A2(pi0789), .A3(new_n15805_), .ZN(new_n15808_));
  NAND3_X1   g12757(.A1(new_n15808_), .A2(new_n15807_), .A3(pi0789), .ZN(new_n15809_));
  NAND2_X1   g12758(.A1(new_n15809_), .A2(new_n15806_), .ZN(new_n15810_));
  NAND4_X1   g12759(.A1(new_n15794_), .A2(new_n15802_), .A3(pi0789), .A4(new_n15785_), .ZN(new_n15811_));
  NOR2_X1    g12760(.A1(new_n15791_), .A2(new_n15787_), .ZN(new_n15812_));
  AOI21_X1   g12761(.A1(new_n15812_), .A2(pi0619), .B(new_n13904_), .ZN(new_n15813_));
  OAI21_X1   g12762(.A1(new_n15813_), .A2(new_n15792_), .B(new_n15654_), .ZN(new_n15814_));
  NOR2_X1    g12763(.A1(new_n15812_), .A2(new_n13896_), .ZN(new_n15815_));
  NAND2_X1   g12764(.A1(new_n15802_), .A2(new_n15815_), .ZN(new_n15816_));
  NAND3_X1   g12765(.A1(new_n15816_), .A2(pi0789), .A3(new_n15814_), .ZN(new_n15817_));
  NAND2_X1   g12766(.A1(new_n15817_), .A2(new_n15811_), .ZN(new_n15818_));
  NAND3_X1   g12767(.A1(new_n15818_), .A2(pi0626), .A3(pi1158), .ZN(new_n15819_));
  NAND4_X1   g12768(.A1(new_n15817_), .A2(new_n13901_), .A3(pi1158), .A4(new_n15811_), .ZN(new_n15820_));
  AOI21_X1   g12769(.A1(new_n15819_), .A2(new_n15820_), .B(new_n15683_), .ZN(new_n15821_));
  NOR2_X1    g12770(.A1(new_n15683_), .A2(new_n13919_), .ZN(new_n15822_));
  AOI21_X1   g12771(.A1(new_n15796_), .A2(new_n13919_), .B(new_n15822_), .ZN(new_n15823_));
  AOI21_X1   g12772(.A1(new_n15823_), .A2(new_n13901_), .B(new_n13924_), .ZN(new_n15824_));
  INV_X1     g12773(.I(new_n15824_), .ZN(new_n15825_));
  OAI21_X1   g12774(.A1(new_n15821_), .A2(new_n15825_), .B(new_n13901_), .ZN(new_n15826_));
  NAND3_X1   g12775(.A1(new_n15818_), .A2(pi0626), .A3(pi1158), .ZN(new_n15827_));
  NAND4_X1   g12776(.A1(new_n15817_), .A2(pi0626), .A3(new_n13929_), .A4(new_n15811_), .ZN(new_n15828_));
  AOI21_X1   g12777(.A1(new_n15827_), .A2(new_n15828_), .B(new_n15683_), .ZN(new_n15829_));
  NAND4_X1   g12778(.A1(new_n15826_), .A2(pi0626), .A3(new_n15810_), .A4(pi0788), .ZN(new_n15832_));
  NAND2_X1   g12779(.A1(new_n15826_), .A2(new_n15810_), .ZN(new_n15833_));
  NAND2_X1   g12780(.A1(new_n15810_), .A2(new_n14577_), .ZN(new_n15834_));
  NAND3_X1   g12781(.A1(new_n15833_), .A2(new_n15834_), .A3(pi0788), .ZN(new_n15835_));
  NAND2_X1   g12782(.A1(new_n15835_), .A2(new_n15832_), .ZN(new_n15836_));
  NAND4_X1   g12783(.A1(new_n15821_), .A2(new_n15829_), .A3(pi0788), .A4(new_n15818_), .ZN(new_n15837_));
  AOI21_X1   g12784(.A1(new_n15812_), .A2(pi1159), .B(new_n13904_), .ZN(new_n15838_));
  INV_X1     g12785(.I(new_n15801_), .ZN(new_n15839_));
  OAI21_X1   g12786(.A1(new_n15838_), .A2(new_n15839_), .B(new_n15654_), .ZN(new_n15840_));
  NOR4_X1    g12787(.A1(new_n15840_), .A2(new_n15814_), .A3(new_n13896_), .A4(new_n15812_), .ZN(new_n15841_));
  NAND2_X1   g12788(.A1(new_n15814_), .A2(pi0789), .ZN(new_n15842_));
  INV_X1     g12789(.I(new_n15815_), .ZN(new_n15843_));
  NOR2_X1    g12790(.A1(new_n15840_), .A2(new_n15843_), .ZN(new_n15844_));
  NOR2_X1    g12791(.A1(new_n15844_), .A2(new_n15842_), .ZN(new_n15845_));
  NOR2_X1    g12792(.A1(new_n15845_), .A2(new_n15841_), .ZN(new_n15846_));
  AOI21_X1   g12793(.A1(new_n15846_), .A2(pi1158), .B(new_n13954_), .ZN(new_n15847_));
  INV_X1     g12794(.I(new_n15820_), .ZN(new_n15848_));
  OAI21_X1   g12795(.A1(new_n15847_), .A2(new_n15848_), .B(new_n15654_), .ZN(new_n15849_));
  NAND2_X1   g12796(.A1(new_n15827_), .A2(new_n15828_), .ZN(new_n15850_));
  NOR2_X1    g12797(.A1(new_n15846_), .A2(new_n13937_), .ZN(new_n15851_));
  NAND3_X1   g12798(.A1(new_n15850_), .A2(new_n15654_), .A3(new_n15851_), .ZN(new_n15852_));
  NAND3_X1   g12799(.A1(new_n15852_), .A2(pi0788), .A3(new_n15849_), .ZN(new_n15853_));
  NAND2_X1   g12800(.A1(new_n15853_), .A2(new_n15837_), .ZN(new_n15854_));
  NOR2_X1    g12801(.A1(new_n15654_), .A2(new_n13966_), .ZN(new_n15855_));
  AOI21_X1   g12802(.A1(new_n15823_), .A2(new_n13966_), .B(new_n15855_), .ZN(new_n15856_));
  AOI21_X1   g12803(.A1(new_n15856_), .A2(pi0628), .B(new_n13971_), .ZN(new_n15857_));
  AND3_X2    g12804(.A1(new_n15856_), .A2(pi0628), .A3(new_n13969_), .Z(new_n15858_));
  OAI21_X1   g12805(.A1(new_n15858_), .A2(new_n15857_), .B(new_n15654_), .ZN(new_n15859_));
  NAND2_X1   g12806(.A1(new_n15859_), .A2(new_n13977_), .ZN(new_n15860_));
  OAI21_X1   g12807(.A1(new_n15854_), .A2(new_n15860_), .B(new_n13942_), .ZN(new_n15861_));
  AOI21_X1   g12808(.A1(new_n15836_), .A2(new_n15861_), .B(new_n12777_), .ZN(new_n15862_));
  AOI21_X1   g12809(.A1(new_n15856_), .A2(pi1156), .B(new_n13971_), .ZN(new_n15863_));
  AND3_X2    g12810(.A1(new_n15856_), .A2(pi1156), .A3(new_n13971_), .Z(new_n15864_));
  OAI21_X1   g12811(.A1(new_n15864_), .A2(new_n15863_), .B(new_n15654_), .ZN(new_n15865_));
  NAND2_X1   g12812(.A1(new_n15836_), .A2(new_n14606_), .ZN(new_n15868_));
  XOR2_X1    g12813(.A1(new_n15862_), .A2(new_n15868_), .Z(new_n15869_));
  NOR2_X1    g12814(.A1(new_n15654_), .A2(new_n13994_), .ZN(new_n15870_));
  INV_X1     g12815(.I(new_n15870_), .ZN(new_n15871_));
  NAND3_X1   g12816(.A1(new_n15853_), .A2(new_n13994_), .A3(new_n15837_), .ZN(new_n15872_));
  NAND2_X1   g12817(.A1(new_n15872_), .A2(new_n15871_), .ZN(new_n15873_));
  NOR4_X1    g12818(.A1(new_n15865_), .A2(new_n15859_), .A3(new_n12777_), .A4(new_n15856_), .ZN(new_n15874_));
  NAND2_X1   g12819(.A1(new_n15859_), .A2(pi0792), .ZN(new_n15875_));
  NOR3_X1    g12820(.A1(new_n15865_), .A2(new_n12777_), .A3(new_n15856_), .ZN(new_n15876_));
  NOR2_X1    g12821(.A1(new_n15876_), .A2(new_n15875_), .ZN(new_n15877_));
  NOR2_X1    g12822(.A1(new_n15877_), .A2(new_n15874_), .ZN(new_n15878_));
  NAND2_X1   g12823(.A1(new_n15878_), .A2(pi0647), .ZN(new_n15879_));
  NAND2_X1   g12824(.A1(new_n15879_), .A2(new_n14007_), .ZN(new_n15880_));
  NAND3_X1   g12825(.A1(new_n15878_), .A2(pi0647), .A3(new_n14006_), .ZN(new_n15881_));
  NAND2_X1   g12826(.A1(new_n15880_), .A2(new_n15881_), .ZN(new_n15882_));
  AOI21_X1   g12827(.A1(new_n15882_), .A2(new_n15654_), .B(new_n14012_), .ZN(new_n15883_));
  AOI21_X1   g12828(.A1(new_n15883_), .A2(new_n15873_), .B(pi0647), .ZN(new_n15884_));
  AOI21_X1   g12829(.A1(new_n15846_), .A2(pi0626), .B(new_n13954_), .ZN(new_n15885_));
  INV_X1     g12830(.I(new_n15828_), .ZN(new_n15886_));
  OAI21_X1   g12831(.A1(new_n15885_), .A2(new_n15886_), .B(new_n15654_), .ZN(new_n15887_));
  NOR4_X1    g12832(.A1(new_n15887_), .A2(new_n15849_), .A3(new_n13937_), .A4(new_n15846_), .ZN(new_n15888_));
  NAND2_X1   g12833(.A1(new_n15849_), .A2(pi0788), .ZN(new_n15889_));
  INV_X1     g12834(.I(new_n15851_), .ZN(new_n15890_));
  NOR2_X1    g12835(.A1(new_n15887_), .A2(new_n15890_), .ZN(new_n15891_));
  NOR2_X1    g12836(.A1(new_n15891_), .A2(new_n15889_), .ZN(new_n15892_));
  NOR3_X1    g12837(.A1(new_n15892_), .A2(new_n13993_), .A3(new_n15888_), .ZN(new_n15893_));
  NOR3_X1    g12838(.A1(new_n15893_), .A2(new_n14005_), .A3(new_n15870_), .ZN(new_n15894_));
  AOI21_X1   g12839(.A1(new_n15878_), .A2(pi1157), .B(new_n14008_), .ZN(new_n15895_));
  NOR4_X1    g12840(.A1(new_n15877_), .A2(pi0647), .A3(new_n14006_), .A4(new_n15874_), .ZN(new_n15896_));
  OAI21_X1   g12841(.A1(new_n15895_), .A2(new_n15896_), .B(new_n15654_), .ZN(new_n15897_));
  NAND2_X1   g12842(.A1(new_n15897_), .A2(new_n14027_), .ZN(new_n15898_));
  OAI21_X1   g12843(.A1(new_n15894_), .A2(new_n15898_), .B(new_n14005_), .ZN(new_n15899_));
  INV_X1     g12844(.I(new_n15899_), .ZN(new_n15900_));
  NOR4_X1    g12845(.A1(new_n15869_), .A2(new_n12776_), .A3(new_n15884_), .A4(new_n15900_), .ZN(new_n15901_));
  NAND4_X1   g12846(.A1(new_n15836_), .A2(new_n15861_), .A3(pi0628), .A4(pi0792), .ZN(new_n15902_));
  NAND2_X1   g12847(.A1(new_n15862_), .A2(new_n15868_), .ZN(new_n15903_));
  AOI21_X1   g12848(.A1(new_n15903_), .A2(new_n15902_), .B(new_n15884_), .ZN(new_n15904_));
  NAND2_X1   g12849(.A1(new_n15899_), .A2(pi0787), .ZN(new_n15905_));
  AOI21_X1   g12850(.A1(new_n15902_), .A2(new_n15903_), .B(new_n15905_), .ZN(new_n15906_));
  NOR3_X1    g12851(.A1(new_n15906_), .A2(new_n12776_), .A3(new_n15904_), .ZN(new_n15907_));
  OAI21_X1   g12852(.A1(new_n15907_), .A2(new_n15901_), .B(new_n12775_), .ZN(new_n15908_));
  NOR2_X1    g12853(.A1(new_n9992_), .A2(pi0143), .ZN(new_n15909_));
  NOR2_X1    g12854(.A1(new_n14652_), .A2(new_n15572_), .ZN(new_n15910_));
  INV_X1     g12855(.I(new_n15909_), .ZN(new_n15911_));
  OAI21_X1   g12856(.A1(new_n13219_), .A2(new_n15572_), .B(new_n15911_), .ZN(new_n15912_));
  NAND3_X1   g12857(.A1(new_n15912_), .A2(new_n15910_), .A3(new_n15909_), .ZN(new_n15913_));
  AOI21_X1   g12858(.A1(new_n13218_), .A2(pi0687), .B(new_n15909_), .ZN(new_n15914_));
  NOR3_X1    g12859(.A1(new_n15910_), .A2(new_n13614_), .A3(new_n15914_), .ZN(new_n15915_));
  XNOR2_X1   g12860(.A1(new_n15913_), .A2(new_n15915_), .ZN(new_n15916_));
  NAND2_X1   g12861(.A1(new_n15916_), .A2(pi0778), .ZN(new_n15917_));
  NAND2_X1   g12862(.A1(new_n15912_), .A2(new_n13748_), .ZN(new_n15918_));
  NAND2_X1   g12863(.A1(new_n15917_), .A2(new_n15918_), .ZN(new_n15919_));
  INV_X1     g12864(.I(new_n15919_), .ZN(new_n15920_));
  NOR2_X1    g12865(.A1(new_n15920_), .A2(new_n14048_), .ZN(new_n15921_));
  INV_X1     g12866(.I(new_n15921_), .ZN(new_n15922_));
  NOR2_X1    g12867(.A1(new_n15922_), .A2(new_n14051_), .ZN(new_n15923_));
  NAND2_X1   g12868(.A1(new_n15923_), .A2(new_n9992_), .ZN(new_n15924_));
  AOI21_X1   g12869(.A1(new_n15924_), .A2(new_n13966_), .B(new_n13919_), .ZN(new_n15925_));
  NAND2_X1   g12870(.A1(new_n15925_), .A2(new_n14061_), .ZN(new_n15926_));
  NAND2_X1   g12871(.A1(new_n15926_), .A2(pi0647), .ZN(new_n15927_));
  XOR2_X1    g12872(.A1(new_n15927_), .A2(new_n14008_), .Z(new_n15928_));
  NAND2_X1   g12873(.A1(new_n15928_), .A2(new_n15909_), .ZN(new_n15929_));
  NAND2_X1   g12874(.A1(new_n15929_), .A2(pi0787), .ZN(new_n15930_));
  NAND2_X1   g12875(.A1(new_n15926_), .A2(pi1157), .ZN(new_n15931_));
  XOR2_X1    g12876(.A1(new_n15931_), .A2(new_n14008_), .Z(new_n15932_));
  NAND2_X1   g12877(.A1(new_n15932_), .A2(new_n15909_), .ZN(new_n15933_));
  NOR3_X1    g12878(.A1(new_n15933_), .A2(new_n12776_), .A3(new_n15926_), .ZN(new_n15934_));
  XOR2_X1    g12879(.A1(new_n15934_), .A2(new_n15930_), .Z(new_n15935_));
  INV_X1     g12880(.I(new_n15923_), .ZN(new_n15936_));
  NAND2_X1   g12881(.A1(new_n15912_), .A2(new_n13103_), .ZN(new_n15937_));
  NOR2_X1    g12882(.A1(new_n15937_), .A2(new_n13613_), .ZN(new_n15938_));
  NAND2_X1   g12883(.A1(new_n15911_), .A2(new_n13614_), .ZN(new_n15939_));
  OAI21_X1   g12884(.A1(new_n15910_), .A2(new_n15939_), .B(pi0608), .ZN(new_n15940_));
  AOI21_X1   g12885(.A1(new_n13104_), .A2(new_n15573_), .B(new_n15909_), .ZN(new_n15941_));
  NOR2_X1    g12886(.A1(new_n15941_), .A2(pi1153), .ZN(new_n15942_));
  NAND2_X1   g12887(.A1(new_n15940_), .A2(new_n15942_), .ZN(new_n15943_));
  AOI21_X1   g12888(.A1(new_n15943_), .A2(new_n15938_), .B(new_n13748_), .ZN(new_n15944_));
  NOR2_X1    g12889(.A1(new_n15914_), .A2(new_n14082_), .ZN(new_n15945_));
  NAND3_X1   g12890(.A1(new_n15910_), .A2(new_n13614_), .A3(new_n15911_), .ZN(new_n15946_));
  OAI22_X1   g12891(.A1(new_n15946_), .A2(new_n15945_), .B1(new_n15937_), .B2(new_n13613_), .ZN(new_n15947_));
  NAND4_X1   g12892(.A1(new_n15947_), .A2(pi0778), .A3(new_n15937_), .A4(new_n15941_), .ZN(new_n15948_));
  XNOR2_X1   g12893(.A1(new_n15948_), .A2(new_n15944_), .ZN(new_n15949_));
  NAND2_X1   g12894(.A1(new_n15949_), .A2(new_n13801_), .ZN(new_n15950_));
  NOR2_X1    g12895(.A1(new_n15949_), .A2(new_n13778_), .ZN(new_n15951_));
  XOR2_X1    g12896(.A1(new_n15951_), .A2(new_n14694_), .Z(new_n15952_));
  NOR2_X1    g12897(.A1(new_n14096_), .A2(new_n15941_), .ZN(new_n15953_));
  AOI21_X1   g12898(.A1(new_n15953_), .A2(new_n14094_), .B(pi1155), .ZN(new_n15954_));
  NOR2_X1    g12899(.A1(new_n15954_), .A2(new_n13783_), .ZN(new_n15955_));
  OAI21_X1   g12900(.A1(new_n15952_), .A2(new_n15920_), .B(new_n15955_), .ZN(new_n15956_));
  AOI21_X1   g12901(.A1(new_n15941_), .A2(pi1155), .B(new_n9992_), .ZN(new_n15957_));
  NOR2_X1    g12902(.A1(new_n15957_), .A2(new_n14102_), .ZN(new_n15958_));
  NOR2_X1    g12903(.A1(new_n15958_), .A2(pi0660), .ZN(new_n15959_));
  NAND2_X1   g12904(.A1(new_n15956_), .A2(new_n15959_), .ZN(new_n15960_));
  NOR2_X1    g12905(.A1(new_n15949_), .A2(new_n13766_), .ZN(new_n15961_));
  XOR2_X1    g12906(.A1(new_n15961_), .A2(new_n14090_), .Z(new_n15962_));
  NAND4_X1   g12907(.A1(new_n15960_), .A2(pi0785), .A3(new_n15919_), .A4(new_n15962_), .ZN(new_n15963_));
  NAND2_X1   g12908(.A1(new_n15963_), .A2(new_n15950_), .ZN(new_n15964_));
  NAND2_X1   g12909(.A1(new_n15964_), .A2(new_n13855_), .ZN(new_n15965_));
  NOR2_X1    g12910(.A1(new_n15964_), .A2(new_n13816_), .ZN(new_n15966_));
  XOR2_X1    g12911(.A1(new_n15966_), .A2(new_n13818_), .Z(new_n15967_));
  NOR2_X1    g12912(.A1(new_n15954_), .A2(new_n13801_), .ZN(new_n15968_));
  NAND3_X1   g12913(.A1(new_n15958_), .A2(new_n15953_), .A3(pi0785), .ZN(new_n15969_));
  XOR2_X1    g12914(.A1(new_n15968_), .A2(new_n15969_), .Z(new_n15970_));
  NOR2_X1    g12915(.A1(new_n15970_), .A2(new_n13817_), .ZN(new_n15971_));
  OAI21_X1   g12916(.A1(new_n15971_), .A2(new_n9992_), .B(pi0618), .ZN(new_n15972_));
  NAND2_X1   g12917(.A1(new_n15972_), .A2(new_n13823_), .ZN(new_n15973_));
  AOI21_X1   g12918(.A1(new_n15967_), .A2(new_n15921_), .B(new_n15973_), .ZN(new_n15974_));
  OAI21_X1   g12919(.A1(new_n15971_), .A2(pi0618), .B(new_n9992_), .ZN(new_n15975_));
  NAND2_X1   g12920(.A1(new_n15975_), .A2(new_n13823_), .ZN(new_n15976_));
  NOR2_X1    g12921(.A1(new_n15964_), .A2(new_n13817_), .ZN(new_n15977_));
  XOR2_X1    g12922(.A1(new_n15977_), .A2(new_n13819_), .Z(new_n15978_));
  NOR3_X1    g12923(.A1(new_n15978_), .A2(new_n13855_), .A3(new_n15922_), .ZN(new_n15979_));
  OAI21_X1   g12924(.A1(new_n15974_), .A2(new_n15976_), .B(new_n15979_), .ZN(new_n15980_));
  NAND2_X1   g12925(.A1(new_n15980_), .A2(new_n15965_), .ZN(new_n15981_));
  NOR2_X1    g12926(.A1(new_n15981_), .A2(new_n13860_), .ZN(new_n15982_));
  XOR2_X1    g12927(.A1(new_n15982_), .A2(new_n13904_), .Z(new_n15983_));
  NOR2_X1    g12928(.A1(new_n15983_), .A2(new_n15936_), .ZN(new_n15984_));
  NAND2_X1   g12929(.A1(new_n15975_), .A2(pi0781), .ZN(new_n15985_));
  NOR3_X1    g12930(.A1(new_n15972_), .A2(new_n13855_), .A3(new_n15970_), .ZN(new_n15986_));
  XOR2_X1    g12931(.A1(new_n15986_), .A2(new_n15985_), .Z(new_n15987_));
  NAND2_X1   g12932(.A1(new_n15987_), .A2(pi1159), .ZN(new_n15988_));
  XOR2_X1    g12933(.A1(new_n15988_), .A2(new_n13904_), .Z(new_n15989_));
  NAND2_X1   g12934(.A1(new_n15989_), .A2(new_n15909_), .ZN(new_n15990_));
  NAND2_X1   g12935(.A1(new_n15990_), .A2(new_n13884_), .ZN(new_n15991_));
  INV_X1     g12936(.I(new_n15981_), .ZN(new_n15992_));
  AOI21_X1   g12937(.A1(new_n15992_), .A2(new_n14143_), .B(pi0789), .ZN(new_n15993_));
  OAI21_X1   g12938(.A1(new_n15984_), .A2(new_n15991_), .B(new_n15993_), .ZN(new_n15994_));
  NOR2_X1    g12939(.A1(new_n15981_), .A2(new_n13868_), .ZN(new_n15995_));
  XOR2_X1    g12940(.A1(new_n15995_), .A2(new_n13903_), .Z(new_n15996_));
  NAND2_X1   g12941(.A1(new_n15996_), .A2(new_n15923_), .ZN(new_n15997_));
  NAND2_X1   g12942(.A1(new_n15987_), .A2(pi0619), .ZN(new_n15998_));
  XOR2_X1    g12943(.A1(new_n15998_), .A2(new_n13904_), .Z(new_n15999_));
  NAND2_X1   g12944(.A1(new_n15999_), .A2(new_n15909_), .ZN(new_n16000_));
  NAND4_X1   g12945(.A1(new_n15994_), .A2(pi0648), .A3(new_n15997_), .A4(new_n16000_), .ZN(new_n16001_));
  NAND2_X1   g12946(.A1(new_n16000_), .A2(pi0789), .ZN(new_n16002_));
  NOR3_X1    g12947(.A1(new_n15990_), .A2(new_n13896_), .A3(new_n15987_), .ZN(new_n16003_));
  XOR2_X1    g12948(.A1(new_n16003_), .A2(new_n16002_), .Z(new_n16004_));
  NAND2_X1   g12949(.A1(new_n16004_), .A2(new_n14153_), .ZN(new_n16005_));
  NAND2_X1   g12950(.A1(new_n14153_), .A2(new_n15909_), .ZN(new_n16006_));
  XOR2_X1    g12951(.A1(new_n16005_), .A2(new_n16006_), .Z(new_n16007_));
  AOI21_X1   g12952(.A1(new_n15936_), .A2(new_n14162_), .B(new_n14164_), .ZN(new_n16008_));
  AOI21_X1   g12953(.A1(new_n16008_), .A2(new_n13929_), .B(pi0641), .ZN(new_n16009_));
  OAI21_X1   g12954(.A1(new_n13929_), .A2(new_n16008_), .B(new_n16009_), .ZN(new_n16010_));
  NAND2_X1   g12955(.A1(new_n16007_), .A2(new_n16010_), .ZN(new_n16011_));
  NAND2_X1   g12956(.A1(new_n16011_), .A2(pi0788), .ZN(new_n16012_));
  NAND2_X1   g12957(.A1(new_n16001_), .A2(new_n16012_), .ZN(new_n16013_));
  NOR2_X1    g12958(.A1(new_n16013_), .A2(pi0792), .ZN(new_n16014_));
  NAND2_X1   g12959(.A1(new_n16013_), .A2(pi1156), .ZN(new_n16015_));
  XOR2_X1    g12960(.A1(new_n16015_), .A2(new_n13971_), .Z(new_n16016_));
  NAND2_X1   g12961(.A1(new_n16007_), .A2(pi0788), .ZN(new_n16017_));
  OAI21_X1   g12962(.A1(pi0788), .A2(new_n16004_), .B(new_n16017_), .ZN(new_n16018_));
  OR2_X2     g12963(.A1(new_n15925_), .A2(new_n13977_), .Z(new_n16019_));
  NAND4_X1   g12964(.A1(new_n16016_), .A2(new_n14176_), .A3(new_n16018_), .A4(new_n16019_), .ZN(new_n16020_));
  NAND2_X1   g12965(.A1(new_n16013_), .A2(pi0628), .ZN(new_n16021_));
  XOR2_X1    g12966(.A1(new_n16021_), .A2(new_n13971_), .Z(new_n16022_));
  NAND4_X1   g12967(.A1(new_n16022_), .A2(new_n14181_), .A3(new_n16018_), .A4(new_n16019_), .ZN(new_n16023_));
  AOI21_X1   g12968(.A1(new_n16020_), .A2(new_n16023_), .B(new_n12777_), .ZN(new_n16024_));
  NOR2_X1    g12969(.A1(new_n16024_), .A2(new_n16014_), .ZN(new_n16025_));
  NOR2_X1    g12970(.A1(new_n16018_), .A2(new_n13993_), .ZN(new_n16026_));
  AOI21_X1   g12971(.A1(new_n13993_), .A2(new_n15911_), .B(new_n16026_), .ZN(new_n16027_));
  INV_X1     g12972(.I(new_n16027_), .ZN(new_n16028_));
  NAND2_X1   g12973(.A1(new_n16025_), .A2(pi1157), .ZN(new_n16029_));
  XOR2_X1    g12974(.A1(new_n16029_), .A2(new_n14008_), .Z(new_n16030_));
  NAND2_X1   g12975(.A1(new_n15929_), .A2(pi0630), .ZN(new_n16031_));
  AOI21_X1   g12976(.A1(new_n16030_), .A2(new_n16028_), .B(new_n16031_), .ZN(new_n16032_));
  NAND2_X1   g12977(.A1(new_n15933_), .A2(new_n14010_), .ZN(new_n16033_));
  NOR2_X1    g12978(.A1(new_n16032_), .A2(new_n16033_), .ZN(new_n16034_));
  NAND2_X1   g12979(.A1(new_n16025_), .A2(pi0647), .ZN(new_n16035_));
  XOR2_X1    g12980(.A1(new_n16035_), .A2(new_n14008_), .Z(new_n16036_));
  NAND3_X1   g12981(.A1(new_n16036_), .A2(pi0787), .A3(new_n16028_), .ZN(new_n16037_));
  OAI22_X1   g12982(.A1(new_n16034_), .A2(new_n16037_), .B1(pi0787), .B2(new_n16025_), .ZN(new_n16038_));
  NAND3_X1   g12983(.A1(new_n16038_), .A2(pi0644), .A3(pi0715), .ZN(new_n16039_));
  OR3_X2     g12984(.A1(new_n16038_), .A2(new_n14204_), .A3(new_n14205_), .Z(new_n16040_));
  AOI21_X1   g12985(.A1(new_n16040_), .A2(new_n16039_), .B(new_n15935_), .ZN(new_n16041_));
  NOR2_X1    g12986(.A1(new_n14211_), .A2(new_n15911_), .ZN(new_n16042_));
  AOI21_X1   g12987(.A1(new_n16027_), .A2(new_n14211_), .B(new_n16042_), .ZN(new_n16043_));
  NAND2_X1   g12988(.A1(new_n16043_), .A2(pi0715), .ZN(new_n16044_));
  XOR2_X1    g12989(.A1(new_n16044_), .A2(new_n14205_), .Z(new_n16045_));
  OAI21_X1   g12990(.A1(new_n16045_), .A2(new_n15911_), .B(new_n14203_), .ZN(new_n16046_));
  NAND2_X1   g12991(.A1(new_n16043_), .A2(pi0644), .ZN(new_n16047_));
  XOR2_X1    g12992(.A1(new_n16047_), .A2(new_n14217_), .Z(new_n16048_));
  AOI21_X1   g12993(.A1(new_n16048_), .A2(new_n15909_), .B(pi1160), .ZN(new_n16049_));
  OAI21_X1   g12994(.A1(new_n16041_), .A2(new_n16046_), .B(new_n16049_), .ZN(new_n16050_));
  NAND3_X1   g12995(.A1(new_n16038_), .A2(pi0644), .A3(pi0715), .ZN(new_n16051_));
  OR3_X2     g12996(.A1(new_n16038_), .A2(new_n14200_), .A3(new_n14205_), .Z(new_n16052_));
  AOI21_X1   g12997(.A1(new_n16052_), .A2(new_n16051_), .B(new_n15935_), .ZN(new_n16053_));
  NAND4_X1   g12998(.A1(new_n16050_), .A2(new_n16053_), .A3(pi0790), .A4(pi0832), .ZN(new_n16054_));
  NAND2_X1   g12999(.A1(new_n16050_), .A2(new_n16053_), .ZN(new_n16055_));
  NAND3_X1   g13000(.A1(new_n16055_), .A2(pi0832), .A3(new_n14801_), .ZN(new_n16056_));
  AOI21_X1   g13001(.A1(po1038), .A2(new_n10708_), .B(pi0832), .ZN(new_n16057_));
  NAND2_X1   g13002(.A1(new_n16038_), .A2(new_n16057_), .ZN(new_n16058_));
  AOI21_X1   g13003(.A1(new_n16056_), .A2(new_n16054_), .B(new_n16058_), .ZN(new_n16059_));
  AOI21_X1   g13004(.A1(new_n15908_), .A2(new_n7240_), .B(new_n16059_), .ZN(new_n16060_));
  NOR2_X1    g13005(.A1(new_n15907_), .A2(new_n15901_), .ZN(new_n16061_));
  AOI21_X1   g13006(.A1(new_n16061_), .A2(pi0715), .B(new_n14217_), .ZN(new_n16062_));
  NOR4_X1    g13007(.A1(new_n15907_), .A2(new_n15901_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n16063_));
  NOR2_X1    g13008(.A1(new_n16062_), .A2(new_n16063_), .ZN(new_n16064_));
  OAI21_X1   g13009(.A1(new_n12776_), .A2(new_n15904_), .B(new_n15906_), .ZN(new_n16065_));
  NOR2_X1    g13010(.A1(new_n15904_), .A2(new_n12776_), .ZN(new_n16066_));
  NAND2_X1   g13011(.A1(new_n15903_), .A2(new_n15902_), .ZN(new_n16067_));
  NAND3_X1   g13012(.A1(new_n16067_), .A2(pi0787), .A3(new_n15899_), .ZN(new_n16068_));
  NAND2_X1   g13013(.A1(new_n16066_), .A2(new_n16068_), .ZN(new_n16069_));
  NOR2_X1    g13014(.A1(new_n15873_), .A2(new_n14210_), .ZN(new_n16070_));
  AOI21_X1   g13015(.A1(new_n14210_), .A2(new_n15654_), .B(new_n16070_), .ZN(new_n16071_));
  OAI21_X1   g13016(.A1(new_n15683_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n16072_));
  NAND2_X1   g13017(.A1(new_n16071_), .A2(new_n16072_), .ZN(new_n16073_));
  AOI21_X1   g13018(.A1(new_n15882_), .A2(new_n15654_), .B(new_n12776_), .ZN(new_n16074_));
  NOR3_X1    g13019(.A1(new_n15897_), .A2(new_n12776_), .A3(new_n15878_), .ZN(new_n16075_));
  XNOR2_X1   g13020(.A1(new_n16074_), .A2(new_n16075_), .ZN(new_n16076_));
  AOI21_X1   g13021(.A1(new_n16073_), .A2(new_n14815_), .B(pi0644), .ZN(new_n16077_));
  AOI21_X1   g13022(.A1(new_n16065_), .A2(new_n16069_), .B(new_n16077_), .ZN(new_n16078_));
  AOI21_X1   g13023(.A1(new_n15683_), .A2(new_n14254_), .B(pi0644), .ZN(new_n16079_));
  NOR3_X1    g13024(.A1(new_n16076_), .A2(new_n16071_), .A3(new_n16079_), .ZN(new_n16080_));
  OAI21_X1   g13025(.A1(new_n16078_), .A2(pi0790), .B(new_n16080_), .ZN(new_n16081_));
  NOR3_X1    g13026(.A1(new_n16064_), .A2(new_n16060_), .A3(new_n16081_), .ZN(po0300));
  NAND2_X1   g13027(.A1(new_n14314_), .A2(new_n14329_), .ZN(new_n16083_));
  NAND3_X1   g13028(.A1(new_n14344_), .A2(new_n14339_), .A3(new_n14347_), .ZN(new_n16084_));
  NAND2_X1   g13029(.A1(new_n16084_), .A2(new_n16083_), .ZN(new_n16085_));
  NOR3_X1    g13030(.A1(new_n16085_), .A2(new_n12986_), .A3(new_n12992_), .ZN(new_n16086_));
  NAND3_X1   g13031(.A1(new_n12977_), .A2(new_n16086_), .A3(pi0758), .ZN(new_n16087_));
  NAND4_X1   g13032(.A1(new_n13093_), .A2(new_n13088_), .A3(new_n16083_), .A4(new_n16084_), .ZN(new_n16088_));
  NAND3_X1   g13033(.A1(new_n13085_), .A2(new_n16088_), .A3(pi0758), .ZN(new_n16089_));
  INV_X1     g13034(.I(pi0758), .ZN(new_n16090_));
  NOR3_X1    g13035(.A1(new_n14338_), .A2(new_n3183_), .A3(new_n16090_), .ZN(new_n16091_));
  NOR3_X1    g13036(.A1(new_n14356_), .A2(pi0039), .A3(new_n16090_), .ZN(new_n16092_));
  NOR2_X1    g13037(.A1(new_n14298_), .A2(new_n7969_), .ZN(new_n16093_));
  OAI21_X1   g13038(.A1(new_n16092_), .A2(new_n16091_), .B(new_n16093_), .ZN(new_n16094_));
  AOI22_X1   g13039(.A1(new_n16087_), .A2(new_n16089_), .B1(new_n3183_), .B2(new_n16094_), .ZN(new_n16095_));
  AOI21_X1   g13040(.A1(new_n13203_), .A2(pi0758), .B(new_n3259_), .ZN(new_n16096_));
  XOR2_X1    g13041(.A1(new_n13723_), .A2(new_n16096_), .Z(new_n16097_));
  NAND2_X1   g13042(.A1(new_n16097_), .A2(pi0144), .ZN(new_n16098_));
  NOR2_X1    g13043(.A1(new_n16098_), .A2(new_n3259_), .ZN(new_n16099_));
  NOR2_X1    g13044(.A1(new_n16090_), .A2(pi0144), .ZN(new_n16100_));
  INV_X1     g13045(.I(new_n16100_), .ZN(new_n16101_));
  NOR2_X1    g13046(.A1(new_n15562_), .A2(new_n16101_), .ZN(new_n16102_));
  OAI21_X1   g13047(.A1(new_n16095_), .A2(new_n16099_), .B(new_n16102_), .ZN(new_n16103_));
  NOR2_X1    g13048(.A1(new_n3289_), .A2(pi0144), .ZN(new_n16104_));
  INV_X1     g13049(.I(new_n16104_), .ZN(new_n16105_));
  OAI21_X1   g13050(.A1(new_n16103_), .A2(new_n3290_), .B(new_n16105_), .ZN(new_n16106_));
  NOR3_X1    g13051(.A1(new_n13085_), .A2(new_n16088_), .A3(new_n16090_), .ZN(new_n16107_));
  NOR3_X1    g13052(.A1(new_n12977_), .A2(new_n16086_), .A3(new_n16090_), .ZN(new_n16108_));
  NAND2_X1   g13053(.A1(new_n16094_), .A2(new_n3183_), .ZN(new_n16109_));
  OAI21_X1   g13054(.A1(new_n16107_), .A2(new_n16108_), .B(new_n16109_), .ZN(new_n16110_));
  INV_X1     g13055(.I(new_n16099_), .ZN(new_n16111_));
  NAND4_X1   g13056(.A1(new_n13194_), .A2(pi0039), .A3(new_n14388_), .A4(new_n14380_), .ZN(new_n16112_));
  OAI21_X1   g13057(.A1(new_n15558_), .A2(new_n13180_), .B(new_n15557_), .ZN(new_n16113_));
  NAND2_X1   g13058(.A1(new_n16113_), .A2(new_n16112_), .ZN(new_n16114_));
  NAND2_X1   g13059(.A1(new_n16114_), .A2(new_n16100_), .ZN(new_n16115_));
  AOI21_X1   g13060(.A1(new_n16110_), .A2(new_n16111_), .B(new_n16115_), .ZN(new_n16116_));
  NOR2_X1    g13061(.A1(new_n7969_), .A2(new_n16090_), .ZN(new_n16117_));
  NOR2_X1    g13062(.A1(new_n14270_), .A2(new_n7969_), .ZN(new_n16118_));
  XNOR2_X1   g13063(.A1(new_n16118_), .A2(new_n16117_), .ZN(new_n16119_));
  OAI21_X1   g13064(.A1(new_n16119_), .A2(new_n13152_), .B(new_n3211_), .ZN(new_n16120_));
  NAND3_X1   g13065(.A1(new_n13198_), .A2(pi0144), .A3(pi0758), .ZN(new_n16121_));
  NAND3_X1   g13066(.A1(new_n13200_), .A2(new_n7969_), .A3(pi0758), .ZN(new_n16122_));
  AOI21_X1   g13067(.A1(new_n16122_), .A2(new_n16121_), .B(new_n13191_), .ZN(new_n16123_));
  NAND2_X1   g13068(.A1(new_n3289_), .A2(pi0736), .ZN(new_n16124_));
  NOR2_X1    g13069(.A1(new_n15629_), .A2(new_n16124_), .ZN(new_n16125_));
  AOI22_X1   g13070(.A1(new_n16120_), .A2(new_n16123_), .B1(new_n16098_), .B2(new_n16125_), .ZN(new_n16126_));
  NAND3_X1   g13071(.A1(new_n15596_), .A2(new_n7969_), .A3(new_n16090_), .ZN(new_n16127_));
  NOR2_X1    g13072(.A1(new_n15597_), .A2(new_n3183_), .ZN(new_n16128_));
  AOI21_X1   g13073(.A1(new_n16127_), .A2(new_n16128_), .B(pi0144), .ZN(new_n16129_));
  NOR3_X1    g13074(.A1(new_n16129_), .A2(pi0758), .A3(new_n13461_), .ZN(new_n16130_));
  AOI21_X1   g13075(.A1(new_n16130_), .A2(new_n13359_), .B(pi0144), .ZN(new_n16131_));
  NAND3_X1   g13076(.A1(new_n14284_), .A2(pi0144), .A3(new_n3290_), .ZN(new_n16132_));
  NOR3_X1    g13077(.A1(new_n16126_), .A2(new_n16131_), .A3(new_n16132_), .ZN(new_n16133_));
  OAI21_X1   g13078(.A1(new_n16133_), .A2(new_n16116_), .B(pi0736), .ZN(new_n16134_));
  AOI21_X1   g13079(.A1(new_n16134_), .A2(pi1153), .B(new_n13620_), .ZN(new_n16135_));
  INV_X1     g13080(.I(pi0736), .ZN(new_n16136_));
  INV_X1     g13081(.I(new_n16126_), .ZN(new_n16137_));
  NOR2_X1    g13082(.A1(new_n16131_), .A2(new_n16132_), .ZN(new_n16138_));
  NAND2_X1   g13083(.A1(new_n16137_), .A2(new_n16138_), .ZN(new_n16139_));
  AOI21_X1   g13084(.A1(new_n16139_), .A2(new_n16103_), .B(new_n16136_), .ZN(new_n16140_));
  NOR3_X1    g13085(.A1(new_n16140_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n16141_));
  OAI21_X1   g13086(.A1(new_n16141_), .A2(new_n16135_), .B(new_n16106_), .ZN(new_n16142_));
  NAND3_X1   g13087(.A1(new_n14422_), .A2(pi0038), .A3(pi0144), .ZN(new_n16143_));
  NAND3_X1   g13088(.A1(new_n14424_), .A2(new_n3259_), .A3(pi0144), .ZN(new_n16144_));
  AOI21_X1   g13089(.A1(new_n16144_), .A2(new_n16143_), .B(new_n14404_), .ZN(new_n16145_));
  NOR2_X1    g13090(.A1(new_n13206_), .A2(new_n3259_), .ZN(new_n16146_));
  NOR3_X1    g13091(.A1(new_n13109_), .A2(new_n3259_), .A3(new_n16146_), .ZN(new_n16147_));
  NOR3_X1    g13092(.A1(new_n13108_), .A2(new_n3259_), .A3(new_n13206_), .ZN(new_n16148_));
  NOR2_X1    g13093(.A1(new_n16147_), .A2(new_n16148_), .ZN(new_n16149_));
  OAI21_X1   g13094(.A1(new_n16145_), .A2(new_n16124_), .B(new_n7969_), .ZN(new_n16150_));
  AND2_X2    g13095(.A1(new_n16150_), .A2(new_n14428_), .Z(new_n16151_));
  NAND2_X1   g13096(.A1(new_n13627_), .A2(pi0144), .ZN(new_n16152_));
  NAND2_X1   g13097(.A1(new_n16152_), .A2(pi0625), .ZN(new_n16153_));
  XOR2_X1    g13098(.A1(new_n16153_), .A2(new_n13620_), .Z(new_n16154_));
  AOI21_X1   g13099(.A1(new_n16151_), .A2(new_n16154_), .B(new_n14081_), .ZN(new_n16155_));
  NAND2_X1   g13100(.A1(new_n16142_), .A2(new_n16155_), .ZN(new_n16156_));
  AOI21_X1   g13101(.A1(new_n16116_), .A2(new_n3289_), .B(new_n16104_), .ZN(new_n16157_));
  NAND3_X1   g13102(.A1(new_n16140_), .A2(pi0625), .A3(pi1153), .ZN(new_n16158_));
  NAND3_X1   g13103(.A1(new_n16134_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n16159_));
  AOI21_X1   g13104(.A1(new_n16158_), .A2(new_n16159_), .B(new_n16157_), .ZN(new_n16160_));
  NAND2_X1   g13105(.A1(new_n16152_), .A2(pi1153), .ZN(new_n16161_));
  XOR2_X1    g13106(.A1(new_n16161_), .A2(new_n13620_), .Z(new_n16162_));
  NAND2_X1   g13107(.A1(new_n16151_), .A2(new_n16162_), .ZN(new_n16163_));
  NAND3_X1   g13108(.A1(new_n16140_), .A2(new_n16163_), .A3(new_n13749_), .ZN(new_n16164_));
  OR2_X2     g13109(.A1(new_n16160_), .A2(new_n16164_), .Z(new_n16165_));
  AOI21_X1   g13110(.A1(pi0778), .A2(new_n16156_), .B(new_n16165_), .ZN(new_n16166_));
  INV_X1     g13111(.I(new_n16156_), .ZN(new_n16167_));
  NOR2_X1    g13112(.A1(new_n16160_), .A2(new_n16164_), .ZN(new_n16168_));
  NOR3_X1    g13113(.A1(new_n16167_), .A2(new_n16168_), .A3(new_n13748_), .ZN(new_n16169_));
  NOR2_X1    g13114(.A1(new_n16166_), .A2(new_n16169_), .ZN(new_n16170_));
  AOI21_X1   g13115(.A1(new_n16151_), .A2(new_n16154_), .B(new_n13748_), .ZN(new_n16171_));
  NAND3_X1   g13116(.A1(new_n16151_), .A2(new_n16162_), .A3(pi0778), .ZN(new_n16172_));
  XOR2_X1    g13117(.A1(new_n16171_), .A2(new_n16172_), .Z(new_n16173_));
  NAND3_X1   g13118(.A1(new_n13627_), .A2(pi0144), .A3(new_n13775_), .ZN(new_n16174_));
  OAI21_X1   g13119(.A1(new_n16106_), .A2(new_n13775_), .B(new_n16174_), .ZN(new_n16175_));
  NAND3_X1   g13120(.A1(new_n16175_), .A2(pi0609), .A3(pi1155), .ZN(new_n16176_));
  INV_X1     g13121(.I(new_n16174_), .ZN(new_n16177_));
  AOI21_X1   g13122(.A1(new_n13776_), .A2(new_n16157_), .B(new_n16177_), .ZN(new_n16178_));
  NAND3_X1   g13123(.A1(new_n16178_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n16179_));
  AOI21_X1   g13124(.A1(new_n16179_), .A2(new_n16176_), .B(new_n16152_), .ZN(new_n16180_));
  NOR2_X1    g13125(.A1(new_n16180_), .A2(new_n13785_), .ZN(new_n16181_));
  AOI21_X1   g13126(.A1(new_n16173_), .A2(new_n16181_), .B(pi0609), .ZN(new_n16182_));
  OAI21_X1   g13127(.A1(new_n16170_), .A2(new_n16182_), .B(pi0785), .ZN(new_n16183_));
  OAI21_X1   g13128(.A1(new_n16167_), .A2(new_n13748_), .B(new_n16168_), .ZN(new_n16184_));
  NAND3_X1   g13129(.A1(new_n16165_), .A2(new_n16156_), .A3(pi0778), .ZN(new_n16185_));
  NAND2_X1   g13130(.A1(new_n16184_), .A2(new_n16185_), .ZN(new_n16186_));
  NOR2_X1    g13131(.A1(new_n16173_), .A2(new_n13766_), .ZN(new_n16187_));
  INV_X1     g13132(.I(new_n16152_), .ZN(new_n16188_));
  AOI21_X1   g13133(.A1(new_n16178_), .A2(pi1155), .B(new_n14694_), .ZN(new_n16189_));
  NOR3_X1    g13134(.A1(new_n16175_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n16190_));
  OAI21_X1   g13135(.A1(new_n16189_), .A2(new_n16190_), .B(new_n16188_), .ZN(new_n16191_));
  NAND2_X1   g13136(.A1(new_n16191_), .A2(new_n13793_), .ZN(new_n16192_));
  OAI21_X1   g13137(.A1(new_n16187_), .A2(new_n16192_), .B(new_n13766_), .ZN(new_n16193_));
  NAND3_X1   g13138(.A1(new_n16186_), .A2(pi0785), .A3(new_n16193_), .ZN(new_n16194_));
  XOR2_X1    g13139(.A1(new_n16183_), .A2(new_n16194_), .Z(new_n16195_));
  NAND3_X1   g13140(.A1(new_n16175_), .A2(pi0609), .A3(pi1155), .ZN(new_n16196_));
  NAND2_X1   g13141(.A1(new_n16157_), .A2(new_n13776_), .ZN(new_n16197_));
  NAND4_X1   g13142(.A1(new_n16197_), .A2(new_n13766_), .A3(pi1155), .A4(new_n16174_), .ZN(new_n16198_));
  AOI21_X1   g13143(.A1(new_n16196_), .A2(new_n16198_), .B(new_n16152_), .ZN(new_n16199_));
  NAND4_X1   g13144(.A1(new_n16180_), .A2(pi0785), .A3(new_n16199_), .A4(new_n16175_), .ZN(new_n16200_));
  INV_X1     g13145(.I(new_n16200_), .ZN(new_n16201_));
  AOI21_X1   g13146(.A1(new_n16178_), .A2(pi0609), .B(new_n14694_), .ZN(new_n16202_));
  NOR3_X1    g13147(.A1(new_n16175_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n16203_));
  OAI21_X1   g13148(.A1(new_n16202_), .A2(new_n16203_), .B(new_n16188_), .ZN(new_n16204_));
  NAND2_X1   g13149(.A1(new_n16204_), .A2(pi0785), .ZN(new_n16205_));
  NOR3_X1    g13150(.A1(new_n16191_), .A2(new_n13801_), .A3(new_n16178_), .ZN(new_n16206_));
  NOR2_X1    g13151(.A1(new_n16206_), .A2(new_n16205_), .ZN(new_n16207_));
  NOR2_X1    g13152(.A1(new_n16207_), .A2(new_n16201_), .ZN(new_n16208_));
  AOI21_X1   g13153(.A1(new_n16208_), .A2(pi0618), .B(new_n13819_), .ZN(new_n16209_));
  NOR2_X1    g13154(.A1(new_n16178_), .A2(new_n13801_), .ZN(new_n16210_));
  NAND2_X1   g13155(.A1(new_n16199_), .A2(new_n16210_), .ZN(new_n16211_));
  NAND3_X1   g13156(.A1(new_n16211_), .A2(pi0785), .A3(new_n16204_), .ZN(new_n16212_));
  NAND4_X1   g13157(.A1(new_n16212_), .A2(pi0618), .A3(new_n16200_), .A4(new_n13817_), .ZN(new_n16213_));
  INV_X1     g13158(.I(new_n16213_), .ZN(new_n16214_));
  OAI21_X1   g13159(.A1(new_n16209_), .A2(new_n16214_), .B(new_n16188_), .ZN(new_n16215_));
  NAND2_X1   g13160(.A1(new_n16188_), .A2(new_n13803_), .ZN(new_n16216_));
  NAND2_X1   g13161(.A1(new_n16173_), .A2(new_n13805_), .ZN(new_n16217_));
  NAND2_X1   g13162(.A1(new_n16217_), .A2(new_n16216_), .ZN(new_n16218_));
  INV_X1     g13163(.I(new_n16218_), .ZN(new_n16219_));
  NAND2_X1   g13164(.A1(new_n16219_), .A2(new_n13816_), .ZN(new_n16220_));
  NAND3_X1   g13165(.A1(new_n16220_), .A2(new_n13824_), .A3(new_n16215_), .ZN(new_n16221_));
  NAND2_X1   g13166(.A1(new_n16221_), .A2(new_n13816_), .ZN(new_n16222_));
  NAND2_X1   g13167(.A1(new_n16212_), .A2(new_n16200_), .ZN(new_n16223_));
  NAND3_X1   g13168(.A1(new_n16223_), .A2(pi0618), .A3(pi1154), .ZN(new_n16224_));
  NAND4_X1   g13169(.A1(new_n16212_), .A2(new_n13816_), .A3(new_n16200_), .A4(pi1154), .ZN(new_n16225_));
  AOI21_X1   g13170(.A1(new_n16224_), .A2(new_n16225_), .B(new_n16152_), .ZN(new_n16226_));
  OAI21_X1   g13171(.A1(new_n16218_), .A2(new_n13816_), .B(new_n13836_), .ZN(new_n16227_));
  OAI21_X1   g13172(.A1(new_n16227_), .A2(new_n16226_), .B(new_n13816_), .ZN(new_n16228_));
  NAND4_X1   g13173(.A1(new_n16195_), .A2(new_n16228_), .A3(new_n16222_), .A4(pi0781), .ZN(new_n16229_));
  NAND2_X1   g13174(.A1(new_n16195_), .A2(new_n16222_), .ZN(new_n16230_));
  NAND3_X1   g13175(.A1(new_n16195_), .A2(new_n16228_), .A3(pi0781), .ZN(new_n16231_));
  NAND3_X1   g13176(.A1(new_n16231_), .A2(new_n16230_), .A3(pi0781), .ZN(new_n16232_));
  NAND2_X1   g13177(.A1(new_n16232_), .A2(new_n16229_), .ZN(new_n16233_));
  NAND3_X1   g13178(.A1(new_n16223_), .A2(pi0618), .A3(pi1154), .ZN(new_n16234_));
  AOI21_X1   g13179(.A1(new_n16234_), .A2(new_n16213_), .B(new_n16152_), .ZN(new_n16235_));
  NAND4_X1   g13180(.A1(new_n16235_), .A2(new_n16226_), .A3(pi0781), .A4(new_n16223_), .ZN(new_n16236_));
  NOR2_X1    g13181(.A1(new_n16208_), .A2(new_n13855_), .ZN(new_n16237_));
  NAND2_X1   g13182(.A1(new_n16226_), .A2(new_n16237_), .ZN(new_n16238_));
  NAND3_X1   g13183(.A1(new_n16238_), .A2(pi0781), .A3(new_n16215_), .ZN(new_n16239_));
  NAND2_X1   g13184(.A1(new_n16239_), .A2(new_n16236_), .ZN(new_n16240_));
  NAND3_X1   g13185(.A1(new_n16240_), .A2(pi0619), .A3(pi1159), .ZN(new_n16241_));
  NAND4_X1   g13186(.A1(new_n16239_), .A2(pi0619), .A3(new_n13868_), .A4(new_n16236_), .ZN(new_n16242_));
  AOI21_X1   g13187(.A1(new_n16241_), .A2(new_n16242_), .B(new_n16152_), .ZN(new_n16243_));
  NOR2_X1    g13188(.A1(new_n16188_), .A2(new_n13880_), .ZN(new_n16244_));
  AOI21_X1   g13189(.A1(new_n16219_), .A2(new_n13880_), .B(new_n16244_), .ZN(new_n16245_));
  OAI21_X1   g13190(.A1(new_n16245_), .A2(pi0619), .B(new_n13885_), .ZN(new_n16246_));
  OAI21_X1   g13191(.A1(new_n16243_), .A2(new_n16246_), .B(new_n13860_), .ZN(new_n16247_));
  NAND3_X1   g13192(.A1(new_n16240_), .A2(pi0619), .A3(pi1159), .ZN(new_n16248_));
  NAND4_X1   g13193(.A1(new_n16239_), .A2(new_n13860_), .A3(pi1159), .A4(new_n16236_), .ZN(new_n16249_));
  AOI21_X1   g13194(.A1(new_n16248_), .A2(new_n16249_), .B(new_n16152_), .ZN(new_n16250_));
  OAI21_X1   g13195(.A1(new_n16245_), .A2(new_n13860_), .B(new_n13892_), .ZN(new_n16251_));
  OAI21_X1   g13196(.A1(new_n16250_), .A2(new_n16251_), .B(new_n13860_), .ZN(new_n16252_));
  NAND4_X1   g13197(.A1(new_n16233_), .A2(new_n16247_), .A3(new_n16252_), .A4(pi0789), .ZN(new_n16253_));
  NAND2_X1   g13198(.A1(new_n16233_), .A2(new_n16247_), .ZN(new_n16254_));
  NAND3_X1   g13199(.A1(new_n16233_), .A2(new_n16252_), .A3(pi0789), .ZN(new_n16255_));
  NAND3_X1   g13200(.A1(new_n16255_), .A2(new_n16254_), .A3(pi0789), .ZN(new_n16256_));
  NAND2_X1   g13201(.A1(new_n16256_), .A2(new_n16253_), .ZN(new_n16257_));
  NAND4_X1   g13202(.A1(new_n16243_), .A2(new_n16250_), .A3(pi0789), .A4(new_n16240_), .ZN(new_n16258_));
  INV_X1     g13203(.I(new_n16243_), .ZN(new_n16259_));
  AOI21_X1   g13204(.A1(new_n16239_), .A2(new_n16236_), .B(new_n13896_), .ZN(new_n16260_));
  NAND2_X1   g13205(.A1(new_n16250_), .A2(new_n16260_), .ZN(new_n16261_));
  NAND3_X1   g13206(.A1(new_n16261_), .A2(new_n16259_), .A3(pi0789), .ZN(new_n16262_));
  NAND2_X1   g13207(.A1(new_n16262_), .A2(new_n16258_), .ZN(new_n16263_));
  NAND3_X1   g13208(.A1(new_n16263_), .A2(pi0626), .A3(pi1158), .ZN(new_n16264_));
  NAND4_X1   g13209(.A1(new_n16262_), .A2(new_n13901_), .A3(pi1158), .A4(new_n16258_), .ZN(new_n16265_));
  AOI21_X1   g13210(.A1(new_n16264_), .A2(new_n16265_), .B(new_n16152_), .ZN(new_n16266_));
  NOR2_X1    g13211(.A1(new_n16152_), .A2(new_n13919_), .ZN(new_n16267_));
  AOI21_X1   g13212(.A1(new_n16245_), .A2(new_n13919_), .B(new_n16267_), .ZN(new_n16268_));
  OAI21_X1   g13213(.A1(new_n16268_), .A2(pi0626), .B(new_n13923_), .ZN(new_n16269_));
  OAI21_X1   g13214(.A1(new_n16266_), .A2(new_n16269_), .B(new_n13901_), .ZN(new_n16270_));
  NAND3_X1   g13215(.A1(new_n16263_), .A2(pi0626), .A3(pi1158), .ZN(new_n16271_));
  NAND4_X1   g13216(.A1(new_n16262_), .A2(pi0626), .A3(new_n13929_), .A4(new_n16258_), .ZN(new_n16272_));
  AOI21_X1   g13217(.A1(new_n16271_), .A2(new_n16272_), .B(new_n16152_), .ZN(new_n16273_));
  NAND4_X1   g13218(.A1(new_n16270_), .A2(new_n16257_), .A3(pi0626), .A4(pi0788), .ZN(new_n16276_));
  AOI21_X1   g13219(.A1(new_n16270_), .A2(new_n16257_), .B(new_n13937_), .ZN(new_n16277_));
  NAND2_X1   g13220(.A1(new_n16257_), .A2(new_n14577_), .ZN(new_n16278_));
  NAND2_X1   g13221(.A1(new_n16277_), .A2(new_n16278_), .ZN(new_n16279_));
  NAND2_X1   g13222(.A1(new_n16279_), .A2(new_n16276_), .ZN(new_n16280_));
  NAND4_X1   g13223(.A1(new_n16266_), .A2(new_n16273_), .A3(pi0788), .A4(new_n16263_), .ZN(new_n16281_));
  NOR2_X1    g13224(.A1(new_n16266_), .A2(new_n13937_), .ZN(new_n16282_));
  NAND2_X1   g13225(.A1(new_n16271_), .A2(new_n16272_), .ZN(new_n16283_));
  AOI21_X1   g13226(.A1(new_n16262_), .A2(new_n16258_), .B(new_n13937_), .ZN(new_n16284_));
  NAND3_X1   g13227(.A1(new_n16283_), .A2(new_n16188_), .A3(new_n16284_), .ZN(new_n16285_));
  NAND2_X1   g13228(.A1(new_n16282_), .A2(new_n16285_), .ZN(new_n16286_));
  NAND2_X1   g13229(.A1(new_n16286_), .A2(new_n16281_), .ZN(new_n16287_));
  NOR2_X1    g13230(.A1(new_n16188_), .A2(new_n13966_), .ZN(new_n16288_));
  AOI21_X1   g13231(.A1(new_n16268_), .A2(new_n13966_), .B(new_n16288_), .ZN(new_n16289_));
  AOI21_X1   g13232(.A1(new_n16289_), .A2(pi0628), .B(new_n13971_), .ZN(new_n16290_));
  INV_X1     g13233(.I(new_n16289_), .ZN(new_n16291_));
  NOR3_X1    g13234(.A1(new_n16291_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n16292_));
  OAI21_X1   g13235(.A1(new_n16292_), .A2(new_n16290_), .B(new_n16188_), .ZN(new_n16293_));
  INV_X1     g13236(.I(new_n16293_), .ZN(new_n16294_));
  NOR2_X1    g13237(.A1(new_n16294_), .A2(new_n15270_), .ZN(new_n16295_));
  INV_X1     g13238(.I(new_n16295_), .ZN(new_n16296_));
  OAI21_X1   g13239(.A1(new_n16287_), .A2(new_n16296_), .B(new_n13942_), .ZN(new_n16297_));
  AOI21_X1   g13240(.A1(new_n16280_), .A2(new_n16297_), .B(new_n12777_), .ZN(new_n16298_));
  AOI21_X1   g13241(.A1(new_n16289_), .A2(pi1156), .B(new_n13971_), .ZN(new_n16299_));
  NOR3_X1    g13242(.A1(new_n16291_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n16300_));
  OAI21_X1   g13243(.A1(new_n16300_), .A2(new_n16299_), .B(new_n16188_), .ZN(new_n16301_));
  NAND2_X1   g13244(.A1(new_n16280_), .A2(new_n14606_), .ZN(new_n16304_));
  NOR2_X1    g13245(.A1(new_n16298_), .A2(new_n16304_), .ZN(new_n16305_));
  XOR2_X1    g13246(.A1(new_n16277_), .A2(new_n16278_), .Z(new_n16306_));
  XOR2_X1    g13247(.A1(new_n16282_), .A2(new_n16285_), .Z(new_n16307_));
  AOI21_X1   g13248(.A1(new_n16307_), .A2(new_n16295_), .B(pi0628), .ZN(new_n16308_));
  OAI21_X1   g13249(.A1(new_n16306_), .A2(new_n16308_), .B(pi0792), .ZN(new_n16309_));
  NOR2_X1    g13250(.A1(new_n16306_), .A2(new_n15296_), .ZN(new_n16310_));
  NOR2_X1    g13251(.A1(new_n16309_), .A2(new_n16310_), .ZN(new_n16311_));
  NOR2_X1    g13252(.A1(new_n16311_), .A2(new_n16305_), .ZN(new_n16312_));
  NOR2_X1    g13253(.A1(new_n16188_), .A2(new_n13994_), .ZN(new_n16313_));
  AOI21_X1   g13254(.A1(new_n16287_), .A2(new_n13994_), .B(new_n16313_), .ZN(new_n16314_));
  NAND2_X1   g13255(.A1(new_n16293_), .A2(pi0792), .ZN(new_n16315_));
  NOR3_X1    g13256(.A1(new_n16301_), .A2(new_n12777_), .A3(new_n16289_), .ZN(new_n16316_));
  NAND2_X1   g13257(.A1(new_n16316_), .A2(new_n16315_), .ZN(new_n16317_));
  NOR2_X1    g13258(.A1(new_n16316_), .A2(new_n16315_), .ZN(new_n16318_));
  INV_X1     g13259(.I(new_n16318_), .ZN(new_n16319_));
  NAND2_X1   g13260(.A1(new_n16319_), .A2(new_n16317_), .ZN(new_n16320_));
  NAND3_X1   g13261(.A1(new_n16320_), .A2(pi0647), .A3(pi1157), .ZN(new_n16321_));
  INV_X1     g13262(.I(new_n16320_), .ZN(new_n16322_));
  NAND3_X1   g13263(.A1(new_n16322_), .A2(pi0647), .A3(new_n14008_), .ZN(new_n16323_));
  AOI21_X1   g13264(.A1(new_n16323_), .A2(new_n16321_), .B(new_n16152_), .ZN(new_n16324_));
  NOR2_X1    g13265(.A1(new_n16324_), .A2(new_n14012_), .ZN(new_n16325_));
  AOI21_X1   g13266(.A1(new_n16325_), .A2(new_n16314_), .B(pi0647), .ZN(new_n16326_));
  INV_X1     g13267(.I(new_n16313_), .ZN(new_n16327_));
  OAI21_X1   g13268(.A1(new_n16307_), .A2(new_n13993_), .B(new_n16327_), .ZN(new_n16328_));
  INV_X1     g13269(.I(new_n14027_), .ZN(new_n16329_));
  NAND3_X1   g13270(.A1(new_n16320_), .A2(pi0647), .A3(pi1157), .ZN(new_n16330_));
  NAND4_X1   g13271(.A1(new_n16319_), .A2(new_n14005_), .A3(pi1157), .A4(new_n16317_), .ZN(new_n16331_));
  AOI21_X1   g13272(.A1(new_n16330_), .A2(new_n16331_), .B(new_n16152_), .ZN(new_n16332_));
  NOR2_X1    g13273(.A1(new_n16332_), .A2(new_n16329_), .ZN(new_n16333_));
  INV_X1     g13274(.I(new_n16333_), .ZN(new_n16334_));
  AOI21_X1   g13275(.A1(new_n16328_), .A2(pi0647), .B(new_n16334_), .ZN(new_n16335_));
  NOR2_X1    g13276(.A1(new_n16335_), .A2(pi0647), .ZN(new_n16336_));
  NOR4_X1    g13277(.A1(new_n16312_), .A2(new_n12776_), .A3(new_n16326_), .A4(new_n16336_), .ZN(new_n16337_));
  NAND2_X1   g13278(.A1(new_n16309_), .A2(new_n16310_), .ZN(new_n16338_));
  NAND2_X1   g13279(.A1(new_n16298_), .A2(new_n16304_), .ZN(new_n16339_));
  AOI21_X1   g13280(.A1(new_n16338_), .A2(new_n16339_), .B(new_n16326_), .ZN(new_n16340_));
  OAI21_X1   g13281(.A1(new_n16335_), .A2(pi0647), .B(pi0787), .ZN(new_n16341_));
  AOI21_X1   g13282(.A1(new_n16338_), .A2(new_n16339_), .B(new_n16341_), .ZN(new_n16342_));
  NOR3_X1    g13283(.A1(new_n16342_), .A2(new_n12776_), .A3(new_n16340_), .ZN(new_n16343_));
  OAI21_X1   g13284(.A1(new_n16343_), .A2(new_n16337_), .B(new_n12775_), .ZN(new_n16344_));
  NAND2_X1   g13285(.A1(new_n16344_), .A2(new_n5787_), .ZN(new_n16345_));
  NAND2_X1   g13286(.A1(new_n16338_), .A2(new_n16339_), .ZN(new_n16346_));
  INV_X1     g13287(.I(new_n16326_), .ZN(new_n16347_));
  INV_X1     g13288(.I(new_n16336_), .ZN(new_n16348_));
  NAND4_X1   g13289(.A1(new_n16346_), .A2(new_n16348_), .A3(pi0787), .A4(new_n16347_), .ZN(new_n16349_));
  OAI21_X1   g13290(.A1(new_n16311_), .A2(new_n16305_), .B(new_n16347_), .ZN(new_n16350_));
  OAI21_X1   g13291(.A1(new_n16314_), .A2(new_n14005_), .B(new_n16333_), .ZN(new_n16351_));
  AOI21_X1   g13292(.A1(new_n16351_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n16352_));
  OAI21_X1   g13293(.A1(new_n16311_), .A2(new_n16305_), .B(new_n16352_), .ZN(new_n16353_));
  NAND3_X1   g13294(.A1(new_n16350_), .A2(new_n16353_), .A3(pi0787), .ZN(new_n16354_));
  NAND2_X1   g13295(.A1(new_n16354_), .A2(new_n16349_), .ZN(new_n16355_));
  NAND2_X1   g13296(.A1(new_n16188_), .A2(new_n14210_), .ZN(new_n16356_));
  OAI21_X1   g13297(.A1(new_n16328_), .A2(new_n14210_), .B(new_n16356_), .ZN(new_n16357_));
  INV_X1     g13298(.I(new_n16357_), .ZN(new_n16358_));
  NAND4_X1   g13299(.A1(new_n16324_), .A2(pi0787), .A3(new_n16332_), .A4(new_n16320_), .ZN(new_n16359_));
  NOR2_X1    g13300(.A1(new_n16324_), .A2(new_n12776_), .ZN(new_n16360_));
  NAND3_X1   g13301(.A1(new_n16332_), .A2(pi0787), .A3(new_n16320_), .ZN(new_n16361_));
  NAND2_X1   g13302(.A1(new_n16360_), .A2(new_n16361_), .ZN(new_n16362_));
  NAND2_X1   g13303(.A1(new_n16362_), .A2(new_n16359_), .ZN(new_n16363_));
  NAND2_X1   g13304(.A1(pi0644), .A2(pi0715), .ZN(new_n16365_));
  OAI21_X1   g13305(.A1(new_n16358_), .A2(new_n16365_), .B(new_n14204_), .ZN(new_n16366_));
  AOI21_X1   g13306(.A1(new_n16355_), .A2(new_n16366_), .B(pi0790), .ZN(new_n16367_));
  NAND2_X1   g13307(.A1(new_n16363_), .A2(pi0644), .ZN(new_n16368_));
  NOR2_X1    g13308(.A1(new_n14204_), .A2(pi0715), .ZN(new_n16369_));
  NAND3_X1   g13309(.A1(new_n16368_), .A2(new_n16357_), .A3(new_n16369_), .ZN(new_n16370_));
  NAND2_X1   g13310(.A1(new_n5788_), .A2(new_n7969_), .ZN(new_n16371_));
  INV_X1     g13311(.I(new_n14142_), .ZN(new_n16372_));
  NOR2_X1    g13312(.A1(new_n13778_), .A2(pi0609), .ZN(new_n16373_));
  NOR2_X1    g13313(.A1(new_n13766_), .A2(pi1155), .ZN(new_n16374_));
  OAI21_X1   g13314(.A1(new_n16373_), .A2(new_n16374_), .B(pi0785), .ZN(new_n16375_));
  INV_X1     g13315(.I(new_n16375_), .ZN(new_n16376_));
  NOR2_X1    g13316(.A1(new_n13105_), .A2(new_n16090_), .ZN(new_n16377_));
  INV_X1     g13317(.I(new_n16377_), .ZN(new_n16378_));
  NOR2_X1    g13318(.A1(new_n16378_), .A2(new_n16376_), .ZN(new_n16379_));
  INV_X1     g13319(.I(new_n16379_), .ZN(new_n16380_));
  XNOR2_X1   g13320(.A1(pi0618), .A2(pi1154), .ZN(new_n16381_));
  NOR2_X1    g13321(.A1(new_n16381_), .A2(new_n13855_), .ZN(new_n16382_));
  NOR2_X1    g13322(.A1(new_n13775_), .A2(new_n16382_), .ZN(new_n16383_));
  INV_X1     g13323(.I(new_n16383_), .ZN(new_n16384_));
  OAI21_X1   g13324(.A1(new_n16384_), .A2(pi1159), .B(new_n13860_), .ZN(new_n16385_));
  AOI21_X1   g13325(.A1(pi1159), .A2(new_n16384_), .B(new_n16385_), .ZN(new_n16386_));
  NOR2_X1    g13326(.A1(new_n16386_), .A2(new_n13896_), .ZN(new_n16387_));
  INV_X1     g13327(.I(new_n16387_), .ZN(new_n16388_));
  NOR2_X1    g13328(.A1(new_n16388_), .A2(new_n16380_), .ZN(new_n16389_));
  NAND2_X1   g13329(.A1(new_n16389_), .A2(new_n16372_), .ZN(new_n16390_));
  NOR2_X1    g13330(.A1(new_n16390_), .A2(new_n13993_), .ZN(new_n16391_));
  NOR2_X1    g13331(.A1(new_n9992_), .A2(new_n7969_), .ZN(new_n16392_));
  INV_X1     g13332(.I(new_n16392_), .ZN(new_n16393_));
  NAND2_X1   g13333(.A1(new_n16393_), .A2(new_n14200_), .ZN(new_n16394_));
  NAND4_X1   g13334(.A1(new_n16391_), .A2(pi0644), .A3(new_n14211_), .A4(new_n16394_), .ZN(new_n16395_));
  NOR3_X1    g13335(.A1(new_n13219_), .A2(new_n13613_), .A3(new_n16136_), .ZN(new_n16396_));
  INV_X1     g13336(.I(new_n16396_), .ZN(new_n16397_));
  NOR2_X1    g13337(.A1(new_n16392_), .A2(new_n13614_), .ZN(new_n16398_));
  AOI21_X1   g13338(.A1(new_n16397_), .A2(new_n16398_), .B(new_n13748_), .ZN(new_n16399_));
  AOI21_X1   g13339(.A1(new_n13218_), .A2(pi0736), .B(new_n16392_), .ZN(new_n16400_));
  NOR2_X1    g13340(.A1(new_n16396_), .A2(new_n16400_), .ZN(new_n16401_));
  NOR2_X1    g13341(.A1(new_n16401_), .A2(pi1153), .ZN(new_n16402_));
  NAND3_X1   g13342(.A1(new_n16402_), .A2(pi0778), .A3(new_n16400_), .ZN(new_n16403_));
  NOR2_X1    g13343(.A1(new_n16403_), .A2(new_n16399_), .ZN(new_n16404_));
  NAND2_X1   g13344(.A1(new_n16403_), .A2(new_n16399_), .ZN(new_n16405_));
  INV_X1     g13345(.I(new_n16405_), .ZN(new_n16406_));
  NOR2_X1    g13346(.A1(new_n16406_), .A2(new_n16404_), .ZN(new_n16407_));
  NOR2_X1    g13347(.A1(new_n16407_), .A2(new_n15396_), .ZN(new_n16408_));
  INV_X1     g13348(.I(new_n16408_), .ZN(new_n16409_));
  NOR2_X1    g13349(.A1(new_n16409_), .A2(new_n14058_), .ZN(new_n16410_));
  AOI21_X1   g13350(.A1(new_n16410_), .A2(new_n15402_), .B(new_n16392_), .ZN(new_n16411_));
  OAI21_X1   g13351(.A1(new_n16410_), .A2(pi0630), .B(pi0647), .ZN(new_n16412_));
  NAND2_X1   g13352(.A1(new_n16412_), .A2(pi1157), .ZN(new_n16413_));
  NAND3_X1   g13353(.A1(new_n16391_), .A2(pi0630), .A3(pi1157), .ZN(new_n16415_));
  XNOR2_X1   g13354(.A1(new_n16413_), .A2(new_n16415_), .ZN(new_n16416_));
  XNOR2_X1   g13355(.A1(pi0630), .A2(pi0647), .ZN(new_n16417_));
  NAND2_X1   g13356(.A1(new_n15400_), .A2(new_n16417_), .ZN(new_n16418_));
  NAND2_X1   g13357(.A1(new_n16418_), .A2(pi0787), .ZN(new_n16419_));
  NOR2_X1    g13358(.A1(new_n13942_), .A2(pi0629), .ZN(new_n16420_));
  NOR2_X1    g13359(.A1(new_n13976_), .A2(pi0628), .ZN(new_n16421_));
  NOR4_X1    g13360(.A1(new_n13990_), .A2(new_n13991_), .A3(new_n16420_), .A4(new_n16421_), .ZN(new_n16422_));
  NOR2_X1    g13361(.A1(new_n16422_), .A2(new_n12777_), .ZN(new_n16423_));
  INV_X1     g13362(.I(new_n16423_), .ZN(new_n16424_));
  INV_X1     g13363(.I(new_n16390_), .ZN(new_n16425_));
  NAND2_X1   g13364(.A1(new_n16390_), .A2(new_n13942_), .ZN(new_n16426_));
  AOI22_X1   g13365(.A1(new_n16426_), .A2(new_n16408_), .B1(new_n16425_), .B2(pi0629), .ZN(new_n16427_));
  NAND2_X1   g13366(.A1(new_n16390_), .A2(new_n15270_), .ZN(new_n16428_));
  NAND4_X1   g13367(.A1(new_n16428_), .A2(pi0628), .A3(new_n16409_), .A4(new_n16392_), .ZN(new_n16429_));
  AOI21_X1   g13368(.A1(new_n13969_), .A2(new_n16429_), .B(new_n16427_), .ZN(new_n16430_));
  OAI21_X1   g13369(.A1(new_n16430_), .A2(new_n16424_), .B(new_n16419_), .ZN(new_n16431_));
  INV_X1     g13370(.I(new_n16407_), .ZN(new_n16432_));
  NAND2_X1   g13371(.A1(new_n13880_), .A2(new_n16393_), .ZN(new_n16433_));
  OAI21_X1   g13372(.A1(new_n16432_), .A2(new_n16433_), .B(new_n13803_), .ZN(new_n16434_));
  NAND2_X1   g13373(.A1(new_n13220_), .A2(pi0625), .ZN(new_n16435_));
  NAND2_X1   g13374(.A1(new_n16392_), .A2(pi1153), .ZN(new_n16436_));
  NOR4_X1    g13375(.A1(new_n16435_), .A2(new_n16378_), .A3(new_n16136_), .A4(new_n16436_), .ZN(new_n16437_));
  NOR3_X1    g13376(.A1(new_n16437_), .A2(new_n16402_), .A3(new_n14081_), .ZN(new_n16438_));
  NOR2_X1    g13377(.A1(new_n16438_), .A2(new_n13748_), .ZN(new_n16439_));
  NAND2_X1   g13378(.A1(new_n16439_), .A2(new_n13801_), .ZN(new_n16440_));
  NOR2_X1    g13379(.A1(new_n16439_), .A2(new_n13778_), .ZN(new_n16441_));
  XOR2_X1    g13380(.A1(new_n16441_), .A2(new_n14090_), .Z(new_n16442_));
  NAND2_X1   g13381(.A1(new_n16442_), .A2(new_n16432_), .ZN(new_n16443_));
  INV_X1     g13382(.I(new_n13779_), .ZN(new_n16444_));
  AOI21_X1   g13383(.A1(new_n13778_), .A2(new_n16393_), .B(new_n16444_), .ZN(new_n16445_));
  AOI21_X1   g13384(.A1(new_n16445_), .A2(new_n16377_), .B(new_n13783_), .ZN(new_n16446_));
  OAI21_X1   g13385(.A1(pi1155), .A2(new_n16392_), .B(new_n14101_), .ZN(new_n16447_));
  OAI21_X1   g13386(.A1(new_n16447_), .A2(new_n16378_), .B(new_n13783_), .ZN(new_n16448_));
  AOI21_X1   g13387(.A1(new_n16443_), .A2(new_n16446_), .B(new_n16448_), .ZN(new_n16449_));
  NOR2_X1    g13388(.A1(new_n16439_), .A2(new_n13766_), .ZN(new_n16450_));
  XOR2_X1    g13389(.A1(new_n16450_), .A2(new_n14090_), .Z(new_n16451_));
  NAND3_X1   g13390(.A1(new_n16451_), .A2(pi0785), .A3(new_n16432_), .ZN(new_n16452_));
  OAI21_X1   g13391(.A1(new_n16449_), .A2(new_n16452_), .B(new_n16440_), .ZN(new_n16453_));
  NAND2_X1   g13392(.A1(new_n16453_), .A2(new_n13855_), .ZN(new_n16454_));
  AOI21_X1   g13393(.A1(new_n16432_), .A2(new_n13805_), .B(new_n16392_), .ZN(new_n16455_));
  INV_X1     g13394(.I(new_n16455_), .ZN(new_n16456_));
  NOR2_X1    g13395(.A1(new_n16453_), .A2(new_n13817_), .ZN(new_n16457_));
  XOR2_X1    g13396(.A1(new_n16457_), .A2(new_n13819_), .Z(new_n16458_));
  NOR2_X1    g13397(.A1(new_n16392_), .A2(pi1154), .ZN(new_n16459_));
  NAND2_X1   g13398(.A1(new_n13776_), .A2(new_n13816_), .ZN(new_n16460_));
  NOR2_X1    g13399(.A1(new_n16460_), .A2(new_n16459_), .ZN(new_n16461_));
  AOI21_X1   g13400(.A1(new_n16379_), .A2(new_n16461_), .B(new_n13823_), .ZN(new_n16462_));
  OAI21_X1   g13401(.A1(new_n16458_), .A2(new_n16456_), .B(new_n16462_), .ZN(new_n16463_));
  NAND2_X1   g13402(.A1(new_n13776_), .A2(pi0618), .ZN(new_n16464_));
  NOR2_X1    g13403(.A1(new_n16464_), .A2(new_n16459_), .ZN(new_n16465_));
  AOI21_X1   g13404(.A1(new_n16379_), .A2(new_n16465_), .B(pi0627), .ZN(new_n16466_));
  NAND2_X1   g13405(.A1(new_n16463_), .A2(new_n16466_), .ZN(new_n16467_));
  NOR2_X1    g13406(.A1(new_n16453_), .A2(new_n13816_), .ZN(new_n16468_));
  XOR2_X1    g13407(.A1(new_n16468_), .A2(new_n13818_), .Z(new_n16469_));
  NAND4_X1   g13408(.A1(new_n16467_), .A2(pi0781), .A3(new_n16455_), .A4(new_n16469_), .ZN(new_n16470_));
  NAND2_X1   g13409(.A1(new_n16470_), .A2(new_n16454_), .ZN(new_n16471_));
  NOR2_X1    g13410(.A1(new_n16471_), .A2(new_n13868_), .ZN(new_n16472_));
  XOR2_X1    g13411(.A1(new_n16472_), .A2(new_n13904_), .Z(new_n16473_));
  NOR2_X1    g13412(.A1(pi0648), .A2(pi0789), .ZN(new_n16474_));
  OAI21_X1   g13413(.A1(new_n16473_), .A2(new_n16434_), .B(new_n16474_), .ZN(new_n16475_));
  NAND3_X1   g13414(.A1(new_n13775_), .A2(new_n16382_), .A3(pi0619), .ZN(new_n16476_));
  NOR2_X1    g13415(.A1(new_n16380_), .A2(new_n16476_), .ZN(new_n16477_));
  INV_X1     g13416(.I(new_n16477_), .ZN(new_n16478_));
  NAND4_X1   g13417(.A1(new_n16475_), .A2(new_n13868_), .A3(new_n16393_), .A4(new_n16478_), .ZN(new_n16479_));
  NOR2_X1    g13418(.A1(new_n16392_), .A2(new_n13868_), .ZN(new_n16480_));
  AOI21_X1   g13419(.A1(new_n16478_), .A2(new_n16480_), .B(pi0648), .ZN(new_n16481_));
  NAND2_X1   g13420(.A1(new_n16479_), .A2(new_n16481_), .ZN(new_n16482_));
  NOR2_X1    g13421(.A1(new_n16471_), .A2(new_n13860_), .ZN(new_n16483_));
  XOR2_X1    g13422(.A1(new_n16483_), .A2(new_n13904_), .Z(new_n16484_));
  OAI21_X1   g13423(.A1(new_n13919_), .A2(new_n16392_), .B(new_n16434_), .ZN(new_n16485_));
  OAI21_X1   g13424(.A1(new_n16393_), .A2(new_n13929_), .B(new_n13901_), .ZN(new_n16486_));
  NAND2_X1   g13425(.A1(new_n16389_), .A2(new_n16486_), .ZN(new_n16487_));
  NOR2_X1    g13426(.A1(new_n13937_), .A2(pi0641), .ZN(new_n16488_));
  AOI21_X1   g13427(.A1(new_n16487_), .A2(new_n16488_), .B(new_n14140_), .ZN(new_n16489_));
  NOR4_X1    g13428(.A1(new_n16484_), .A2(new_n16434_), .A3(new_n16485_), .A4(new_n16489_), .ZN(new_n16490_));
  NAND2_X1   g13429(.A1(new_n16482_), .A2(new_n16490_), .ZN(new_n16491_));
  NAND2_X1   g13430(.A1(new_n16471_), .A2(new_n13896_), .ZN(new_n16492_));
  NAND4_X1   g13431(.A1(new_n13901_), .A2(new_n13937_), .A3(pi0641), .A4(pi1158), .ZN(new_n16494_));
  NOR2_X1    g13432(.A1(new_n16485_), .A2(new_n16494_), .ZN(new_n16495_));
  NAND2_X1   g13433(.A1(new_n16492_), .A2(new_n16495_), .ZN(new_n16496_));
  NAND2_X1   g13434(.A1(new_n16430_), .A2(pi0792), .ZN(new_n16497_));
  NOR2_X1    g13435(.A1(new_n16392_), .A2(new_n12776_), .ZN(new_n16498_));
  NAND4_X1   g13436(.A1(new_n16491_), .A2(new_n16496_), .A3(new_n16497_), .A4(new_n16498_), .ZN(new_n16499_));
  OAI21_X1   g13437(.A1(new_n16416_), .A2(new_n16431_), .B(new_n16499_), .ZN(new_n16500_));
  NOR2_X1    g13438(.A1(new_n16500_), .A2(new_n14204_), .ZN(new_n16501_));
  XOR2_X1    g13439(.A1(new_n16501_), .A2(new_n14205_), .Z(new_n16502_));
  NAND4_X1   g13440(.A1(new_n16502_), .A2(new_n14203_), .A3(new_n16395_), .A4(new_n16411_), .ZN(new_n16503_));
  INV_X1     g13441(.I(new_n16411_), .ZN(new_n16504_));
  NOR2_X1    g13442(.A1(new_n16500_), .A2(new_n14200_), .ZN(new_n16505_));
  XOR2_X1    g13443(.A1(new_n16505_), .A2(new_n14217_), .Z(new_n16506_));
  NOR2_X1    g13444(.A1(new_n16506_), .A2(new_n16504_), .ZN(new_n16507_));
  AOI21_X1   g13445(.A1(new_n16503_), .A2(new_n16507_), .B(new_n14799_), .ZN(new_n16508_));
  XOR2_X1    g13446(.A1(new_n16508_), .A2(new_n14800_), .Z(new_n16509_));
  NAND2_X1   g13447(.A1(pi0057), .A2(pi0144), .ZN(new_n16510_));
  AND3_X2    g13448(.A1(new_n16500_), .A2(new_n14799_), .A3(new_n16510_), .Z(new_n16511_));
  AOI22_X1   g13449(.A1(new_n16509_), .A2(new_n16511_), .B1(new_n5371_), .B2(new_n16371_), .ZN(new_n16512_));
  AOI21_X1   g13450(.A1(new_n16370_), .A2(new_n14204_), .B(new_n16512_), .ZN(new_n16513_));
  NAND2_X1   g13451(.A1(new_n16355_), .A2(new_n16513_), .ZN(new_n16514_));
  AOI21_X1   g13452(.A1(new_n16345_), .A2(new_n16367_), .B(new_n16514_), .ZN(po0301));
  NOR2_X1    g13453(.A1(new_n9992_), .A2(pi0145), .ZN(new_n16516_));
  INV_X1     g13454(.I(pi0767), .ZN(new_n16517_));
  AOI21_X1   g13455(.A1(new_n13104_), .A2(new_n16517_), .B(new_n16516_), .ZN(new_n16518_));
  NOR2_X1    g13456(.A1(new_n14096_), .A2(new_n16518_), .ZN(new_n16519_));
  AOI21_X1   g13457(.A1(new_n16519_), .A2(new_n14094_), .B(pi1155), .ZN(new_n16520_));
  NOR2_X1    g13458(.A1(new_n16520_), .A2(new_n13801_), .ZN(new_n16521_));
  NAND2_X1   g13459(.A1(new_n16518_), .A2(pi1155), .ZN(new_n16522_));
  AOI21_X1   g13460(.A1(new_n16522_), .A2(new_n2723_), .B(new_n14102_), .ZN(new_n16523_));
  NAND3_X1   g13461(.A1(new_n16523_), .A2(pi0785), .A3(new_n16519_), .ZN(new_n16524_));
  XOR2_X1    g13462(.A1(new_n16521_), .A2(new_n16524_), .Z(new_n16525_));
  NOR2_X1    g13463(.A1(new_n16525_), .A2(new_n13817_), .ZN(new_n16526_));
  OAI21_X1   g13464(.A1(new_n16526_), .A2(pi0618), .B(new_n9992_), .ZN(new_n16527_));
  NAND2_X1   g13465(.A1(new_n16527_), .A2(pi0781), .ZN(new_n16528_));
  OAI21_X1   g13466(.A1(new_n16526_), .A2(new_n9992_), .B(pi0618), .ZN(new_n16529_));
  NOR3_X1    g13467(.A1(new_n16529_), .A2(new_n13855_), .A3(new_n16525_), .ZN(new_n16530_));
  XOR2_X1    g13468(.A1(new_n16530_), .A2(new_n16528_), .Z(new_n16531_));
  NAND2_X1   g13469(.A1(new_n16531_), .A2(pi0619), .ZN(new_n16532_));
  XOR2_X1    g13470(.A1(new_n16532_), .A2(new_n13904_), .Z(new_n16533_));
  NAND2_X1   g13471(.A1(new_n16533_), .A2(new_n16516_), .ZN(new_n16534_));
  NAND2_X1   g13472(.A1(new_n16534_), .A2(pi0789), .ZN(new_n16535_));
  INV_X1     g13473(.I(new_n16516_), .ZN(new_n16536_));
  NAND2_X1   g13474(.A1(new_n16531_), .A2(pi1159), .ZN(new_n16537_));
  XOR2_X1    g13475(.A1(new_n16537_), .A2(new_n13903_), .Z(new_n16538_));
  NOR2_X1    g13476(.A1(new_n16538_), .A2(new_n16536_), .ZN(new_n16539_));
  INV_X1     g13477(.I(new_n16539_), .ZN(new_n16540_));
  NOR3_X1    g13478(.A1(new_n16540_), .A2(new_n13896_), .A3(new_n16531_), .ZN(new_n16541_));
  XOR2_X1    g13479(.A1(new_n16541_), .A2(new_n16535_), .Z(new_n16542_));
  NAND2_X1   g13480(.A1(new_n16542_), .A2(new_n14153_), .ZN(new_n16543_));
  NAND2_X1   g13481(.A1(new_n14153_), .A2(new_n16516_), .ZN(new_n16544_));
  XOR2_X1    g13482(.A1(new_n16543_), .A2(new_n16544_), .Z(new_n16545_));
  INV_X1     g13483(.I(new_n14055_), .ZN(new_n16546_));
  NOR3_X1    g13484(.A1(new_n16546_), .A2(pi1156), .A3(new_n14181_), .ZN(new_n16547_));
  OR2_X2     g13485(.A1(new_n16542_), .A2(pi0788), .Z(new_n16548_));
  NAND2_X1   g13486(.A1(new_n16545_), .A2(pi0788), .ZN(new_n16549_));
  INV_X1     g13487(.I(pi0698), .ZN(new_n16550_));
  AOI21_X1   g13488(.A1(new_n13218_), .A2(new_n16550_), .B(new_n16516_), .ZN(new_n16551_));
  INV_X1     g13489(.I(new_n16551_), .ZN(new_n16552_));
  NOR3_X1    g13490(.A1(new_n13219_), .A2(pi0625), .A3(pi0698), .ZN(new_n16553_));
  NAND3_X1   g13491(.A1(new_n16552_), .A2(new_n16553_), .A3(new_n16516_), .ZN(new_n16554_));
  NOR3_X1    g13492(.A1(new_n16553_), .A2(new_n13614_), .A3(new_n16551_), .ZN(new_n16555_));
  XOR2_X1    g13493(.A1(new_n16554_), .A2(new_n16555_), .Z(new_n16556_));
  NAND2_X1   g13494(.A1(new_n16552_), .A2(new_n13748_), .ZN(new_n16557_));
  OAI21_X1   g13495(.A1(new_n16556_), .A2(new_n13748_), .B(new_n16557_), .ZN(new_n16558_));
  NAND2_X1   g13496(.A1(new_n16558_), .A2(new_n14049_), .ZN(new_n16559_));
  NOR2_X1    g13497(.A1(new_n16559_), .A2(new_n14051_), .ZN(new_n16560_));
  NAND2_X1   g13498(.A1(new_n16560_), .A2(new_n9992_), .ZN(new_n16561_));
  AOI21_X1   g13499(.A1(new_n16561_), .A2(new_n13966_), .B(new_n13919_), .ZN(new_n16562_));
  INV_X1     g13500(.I(new_n16562_), .ZN(new_n16563_));
  AOI21_X1   g13501(.A1(new_n16549_), .A2(new_n16548_), .B(new_n16563_), .ZN(new_n16564_));
  NOR2_X1    g13502(.A1(new_n16564_), .A2(new_n16547_), .ZN(new_n16565_));
  INV_X1     g13503(.I(new_n14176_), .ZN(new_n16566_));
  INV_X1     g13504(.I(new_n14056_), .ZN(new_n16567_));
  NOR2_X1    g13505(.A1(new_n16567_), .A2(new_n13969_), .ZN(new_n16568_));
  AOI21_X1   g13506(.A1(new_n16568_), .A2(new_n16566_), .B(new_n12777_), .ZN(new_n16569_));
  INV_X1     g13507(.I(new_n16569_), .ZN(new_n16570_));
  NOR2_X1    g13508(.A1(new_n16564_), .A2(new_n16570_), .ZN(new_n16571_));
  NOR2_X1    g13509(.A1(new_n13976_), .A2(new_n12777_), .ZN(new_n16572_));
  XNOR2_X1   g13510(.A1(new_n16571_), .A2(new_n16572_), .ZN(new_n16573_));
  INV_X1     g13511(.I(new_n16419_), .ZN(new_n16574_));
  NOR3_X1    g13512(.A1(new_n14005_), .A2(pi0630), .A3(pi1157), .ZN(new_n16575_));
  AOI21_X1   g13513(.A1(pi0630), .A2(new_n15398_), .B(new_n16575_), .ZN(new_n16576_));
  AND3_X2    g13514(.A1(new_n16549_), .A2(new_n13994_), .A3(new_n16548_), .Z(new_n16577_));
  AOI21_X1   g13515(.A1(new_n13993_), .A2(new_n16536_), .B(new_n16577_), .ZN(new_n16578_));
  NOR2_X1    g13516(.A1(new_n16536_), .A2(pi0647), .ZN(new_n16579_));
  NOR2_X1    g13517(.A1(new_n16563_), .A2(new_n14060_), .ZN(new_n16580_));
  AOI21_X1   g13518(.A1(new_n16580_), .A2(pi0647), .B(new_n16579_), .ZN(new_n16581_));
  NAND2_X1   g13519(.A1(new_n16581_), .A2(pi0630), .ZN(new_n16582_));
  NOR2_X1    g13520(.A1(new_n16580_), .A2(new_n14005_), .ZN(new_n16583_));
  XOR2_X1    g13521(.A1(new_n16583_), .A2(new_n14007_), .Z(new_n16584_));
  NAND2_X1   g13522(.A1(new_n16584_), .A2(new_n16516_), .ZN(new_n16585_));
  NOR2_X1    g13523(.A1(new_n16585_), .A2(new_n14012_), .ZN(new_n16586_));
  XOR2_X1    g13524(.A1(new_n16586_), .A2(new_n16582_), .Z(new_n16587_));
  OAI21_X1   g13525(.A1(new_n12776_), .A2(new_n16587_), .B(new_n16578_), .ZN(new_n16588_));
  AOI21_X1   g13526(.A1(new_n16588_), .A2(new_n16576_), .B(new_n16574_), .ZN(new_n16589_));
  OAI21_X1   g13527(.A1(new_n16573_), .A2(new_n16565_), .B(new_n16589_), .ZN(new_n16590_));
  NOR3_X1    g13528(.A1(new_n16551_), .A2(new_n13613_), .A3(new_n13203_), .ZN(new_n16591_));
  INV_X1     g13529(.I(new_n16518_), .ZN(new_n16592_));
  NOR2_X1    g13530(.A1(new_n16516_), .A2(pi1153), .ZN(new_n16593_));
  INV_X1     g13531(.I(new_n16593_), .ZN(new_n16594_));
  OAI21_X1   g13532(.A1(new_n16553_), .A2(new_n16594_), .B(pi0608), .ZN(new_n16595_));
  NAND3_X1   g13533(.A1(new_n16595_), .A2(new_n13614_), .A3(new_n16592_), .ZN(new_n16596_));
  AOI21_X1   g13534(.A1(new_n16596_), .A2(new_n16591_), .B(new_n13748_), .ZN(new_n16597_));
  NOR2_X1    g13535(.A1(new_n16551_), .A2(new_n13203_), .ZN(new_n16598_));
  NAND2_X1   g13536(.A1(new_n16553_), .A2(new_n16593_), .ZN(new_n16599_));
  AOI21_X1   g13537(.A1(new_n14083_), .A2(new_n16552_), .B(new_n16599_), .ZN(new_n16600_));
  NOR2_X1    g13538(.A1(new_n16600_), .A2(new_n16591_), .ZN(new_n16601_));
  NOR4_X1    g13539(.A1(new_n16601_), .A2(new_n13748_), .A3(new_n16592_), .A4(new_n16598_), .ZN(new_n16602_));
  XOR2_X1    g13540(.A1(new_n16602_), .A2(new_n16597_), .Z(new_n16603_));
  NAND2_X1   g13541(.A1(new_n16603_), .A2(new_n13801_), .ZN(new_n16604_));
  NOR2_X1    g13542(.A1(new_n16603_), .A2(new_n13778_), .ZN(new_n16605_));
  XOR2_X1    g13543(.A1(new_n16605_), .A2(new_n14090_), .Z(new_n16606_));
  NAND2_X1   g13544(.A1(new_n16606_), .A2(new_n16558_), .ZN(new_n16607_));
  NOR2_X1    g13545(.A1(new_n16520_), .A2(new_n13783_), .ZN(new_n16608_));
  NAND2_X1   g13546(.A1(new_n16607_), .A2(new_n16608_), .ZN(new_n16609_));
  NOR2_X1    g13547(.A1(new_n16523_), .A2(pi0660), .ZN(new_n16610_));
  NAND2_X1   g13548(.A1(new_n16609_), .A2(new_n16610_), .ZN(new_n16611_));
  NOR2_X1    g13549(.A1(new_n16603_), .A2(new_n13766_), .ZN(new_n16612_));
  XOR2_X1    g13550(.A1(new_n16612_), .A2(new_n14090_), .Z(new_n16613_));
  NAND4_X1   g13551(.A1(new_n16611_), .A2(pi0785), .A3(new_n16558_), .A4(new_n16613_), .ZN(new_n16614_));
  NAND2_X1   g13552(.A1(new_n16614_), .A2(new_n16604_), .ZN(new_n16615_));
  NAND2_X1   g13553(.A1(new_n16615_), .A2(new_n13855_), .ZN(new_n16616_));
  INV_X1     g13554(.I(new_n16559_), .ZN(new_n16617_));
  NOR2_X1    g13555(.A1(new_n16615_), .A2(new_n13816_), .ZN(new_n16618_));
  XOR2_X1    g13556(.A1(new_n16618_), .A2(new_n13818_), .Z(new_n16619_));
  NAND2_X1   g13557(.A1(new_n16529_), .A2(new_n13823_), .ZN(new_n16620_));
  AOI21_X1   g13558(.A1(new_n16619_), .A2(new_n16617_), .B(new_n16620_), .ZN(new_n16621_));
  NAND2_X1   g13559(.A1(new_n16527_), .A2(new_n13823_), .ZN(new_n16622_));
  NOR2_X1    g13560(.A1(new_n16615_), .A2(new_n13817_), .ZN(new_n16623_));
  XOR2_X1    g13561(.A1(new_n16623_), .A2(new_n13819_), .Z(new_n16624_));
  NOR3_X1    g13562(.A1(new_n16624_), .A2(new_n13855_), .A3(new_n16559_), .ZN(new_n16625_));
  OAI21_X1   g13563(.A1(new_n16621_), .A2(new_n16622_), .B(new_n16625_), .ZN(new_n16626_));
  NAND2_X1   g13564(.A1(new_n16626_), .A2(new_n16616_), .ZN(new_n16627_));
  NOR2_X1    g13565(.A1(new_n16627_), .A2(new_n13860_), .ZN(new_n16628_));
  XOR2_X1    g13566(.A1(new_n16628_), .A2(new_n13903_), .Z(new_n16629_));
  NAND2_X1   g13567(.A1(new_n16540_), .A2(new_n13884_), .ZN(new_n16630_));
  AOI21_X1   g13568(.A1(new_n16629_), .A2(new_n16560_), .B(new_n16630_), .ZN(new_n16631_));
  OAI21_X1   g13569(.A1(new_n16627_), .A2(new_n15479_), .B(new_n13896_), .ZN(new_n16632_));
  NOR2_X1    g13570(.A1(new_n16631_), .A2(new_n16632_), .ZN(new_n16633_));
  NOR2_X1    g13571(.A1(new_n16627_), .A2(new_n13868_), .ZN(new_n16634_));
  XOR2_X1    g13572(.A1(new_n16634_), .A2(new_n13903_), .Z(new_n16635_));
  NAND2_X1   g13573(.A1(new_n16635_), .A2(new_n16560_), .ZN(new_n16636_));
  NAND4_X1   g13574(.A1(new_n16636_), .A2(pi0648), .A3(new_n16423_), .A4(new_n16534_), .ZN(new_n16637_));
  OAI21_X1   g13575(.A1(new_n16633_), .A2(new_n16637_), .B(new_n13937_), .ZN(new_n16638_));
  INV_X1     g13576(.I(new_n14162_), .ZN(new_n16639_));
  NOR2_X1    g13577(.A1(new_n16560_), .A2(new_n16639_), .ZN(new_n16640_));
  NOR2_X1    g13578(.A1(new_n16640_), .A2(new_n14164_), .ZN(new_n16641_));
  AOI21_X1   g13579(.A1(new_n16641_), .A2(new_n13929_), .B(pi0641), .ZN(new_n16642_));
  OAI21_X1   g13580(.A1(new_n13929_), .A2(new_n16641_), .B(new_n16642_), .ZN(new_n16643_));
  NAND4_X1   g13581(.A1(new_n16590_), .A2(new_n16545_), .A3(new_n16638_), .A4(new_n16643_), .ZN(new_n16644_));
  AOI21_X1   g13582(.A1(new_n16581_), .A2(pi1157), .B(new_n12776_), .ZN(new_n16645_));
  AOI22_X1   g13583(.A1(new_n16585_), .A2(new_n16645_), .B1(new_n12776_), .B2(new_n16580_), .ZN(new_n16646_));
  NAND2_X1   g13584(.A1(new_n16644_), .A2(pi0644), .ZN(new_n16647_));
  XOR2_X1    g13585(.A1(new_n16647_), .A2(new_n14205_), .Z(new_n16648_));
  NOR2_X1    g13586(.A1(new_n16648_), .A2(new_n16646_), .ZN(new_n16649_));
  NOR2_X1    g13587(.A1(new_n16578_), .A2(new_n14210_), .ZN(new_n16650_));
  AOI21_X1   g13588(.A1(new_n14210_), .A2(new_n16536_), .B(new_n16650_), .ZN(new_n16651_));
  NAND2_X1   g13589(.A1(new_n16651_), .A2(pi0715), .ZN(new_n16652_));
  XOR2_X1    g13590(.A1(new_n16652_), .A2(new_n14205_), .Z(new_n16653_));
  OAI21_X1   g13591(.A1(new_n16653_), .A2(new_n16536_), .B(new_n14203_), .ZN(new_n16654_));
  NAND2_X1   g13592(.A1(new_n16651_), .A2(pi0644), .ZN(new_n16655_));
  XOR2_X1    g13593(.A1(new_n16655_), .A2(new_n14217_), .Z(new_n16656_));
  AOI21_X1   g13594(.A1(new_n16656_), .A2(new_n16516_), .B(pi1160), .ZN(new_n16657_));
  OAI21_X1   g13595(.A1(new_n16649_), .A2(new_n16654_), .B(new_n16657_), .ZN(new_n16658_));
  NAND2_X1   g13596(.A1(new_n16644_), .A2(pi0715), .ZN(new_n16659_));
  XOR2_X1    g13597(.A1(new_n16659_), .A2(new_n14205_), .Z(new_n16660_));
  NOR2_X1    g13598(.A1(new_n16660_), .A2(new_n16646_), .ZN(new_n16661_));
  AOI21_X1   g13599(.A1(new_n16658_), .A2(new_n16661_), .B(new_n14799_), .ZN(new_n16662_));
  XOR2_X1    g13600(.A1(new_n16662_), .A2(new_n14801_), .Z(new_n16663_));
  NOR2_X1    g13601(.A1(new_n16663_), .A2(new_n16644_), .ZN(new_n16664_));
  NOR2_X1    g13602(.A1(new_n14428_), .A2(pi0145), .ZN(new_n16665_));
  NOR2_X1    g13603(.A1(new_n16665_), .A2(new_n13994_), .ZN(new_n16666_));
  NAND2_X1   g13604(.A1(new_n13109_), .A2(new_n5641_), .ZN(new_n16667_));
  NAND2_X1   g13605(.A1(new_n16667_), .A2(pi0038), .ZN(new_n16668_));
  NOR4_X1    g13606(.A1(new_n15562_), .A2(new_n5641_), .A3(new_n16517_), .A4(new_n14362_), .ZN(new_n16669_));
  NOR4_X1    g13607(.A1(new_n13107_), .A2(new_n3259_), .A3(new_n5641_), .A4(pi0767), .ZN(new_n16670_));
  OAI21_X1   g13608(.A1(new_n16669_), .A2(new_n13097_), .B(new_n16670_), .ZN(new_n16671_));
  XOR2_X1    g13609(.A1(new_n16671_), .A2(new_n16668_), .Z(new_n16672_));
  NOR2_X1    g13610(.A1(new_n3289_), .A2(pi0145), .ZN(new_n16673_));
  AOI21_X1   g13611(.A1(new_n16672_), .A2(new_n3289_), .B(new_n16673_), .ZN(new_n16674_));
  NAND2_X1   g13612(.A1(new_n16674_), .A2(new_n13776_), .ZN(new_n16675_));
  OAI21_X1   g13613(.A1(new_n15147_), .A2(new_n16665_), .B(new_n16675_), .ZN(new_n16676_));
  NAND2_X1   g13614(.A1(new_n16676_), .A2(pi0609), .ZN(new_n16677_));
  NAND2_X1   g13615(.A1(new_n16677_), .A2(pi0785), .ZN(new_n16678_));
  INV_X1     g13616(.I(new_n16674_), .ZN(new_n16679_));
  INV_X1     g13617(.I(new_n16665_), .ZN(new_n16680_));
  NOR2_X1    g13618(.A1(new_n16680_), .A2(new_n13776_), .ZN(new_n16681_));
  AOI21_X1   g13619(.A1(new_n16679_), .A2(new_n13776_), .B(new_n16681_), .ZN(new_n16682_));
  AOI21_X1   g13620(.A1(new_n16680_), .A2(new_n14467_), .B(pi0609), .ZN(new_n16683_));
  NOR2_X1    g13621(.A1(new_n16675_), .A2(new_n16683_), .ZN(new_n16684_));
  INV_X1     g13622(.I(new_n16684_), .ZN(new_n16685_));
  NOR3_X1    g13623(.A1(new_n16685_), .A2(new_n13801_), .A3(new_n16682_), .ZN(new_n16686_));
  XOR2_X1    g13624(.A1(new_n16678_), .A2(new_n16686_), .Z(new_n16687_));
  NOR2_X1    g13625(.A1(new_n16687_), .A2(pi0781), .ZN(new_n16688_));
  INV_X1     g13626(.I(new_n16381_), .ZN(new_n16689_));
  XNOR2_X1   g13627(.A1(new_n16678_), .A2(new_n16686_), .ZN(new_n16690_));
  NAND3_X1   g13628(.A1(new_n16690_), .A2(new_n16689_), .A3(new_n16665_), .ZN(new_n16691_));
  NAND3_X1   g13629(.A1(new_n16687_), .A2(new_n16689_), .A3(new_n16680_), .ZN(new_n16692_));
  NAND2_X1   g13630(.A1(new_n16691_), .A2(new_n16692_), .ZN(new_n16693_));
  AOI21_X1   g13631(.A1(new_n16693_), .A2(pi0781), .B(new_n16688_), .ZN(new_n16694_));
  NOR2_X1    g13632(.A1(new_n16694_), .A2(pi0789), .ZN(new_n16695_));
  XNOR2_X1   g13633(.A1(pi0619), .A2(pi1159), .ZN(new_n16696_));
  INV_X1     g13634(.I(new_n16696_), .ZN(new_n16697_));
  NAND2_X1   g13635(.A1(new_n16694_), .A2(new_n16697_), .ZN(new_n16698_));
  NAND2_X1   g13636(.A1(new_n16665_), .A2(new_n16697_), .ZN(new_n16699_));
  XOR2_X1    g13637(.A1(new_n16698_), .A2(new_n16699_), .Z(new_n16700_));
  AOI21_X1   g13638(.A1(new_n16700_), .A2(pi0789), .B(new_n16695_), .ZN(new_n16701_));
  NOR2_X1    g13639(.A1(new_n16701_), .A2(pi0788), .ZN(new_n16702_));
  OR3_X2     g13640(.A1(new_n16701_), .A2(new_n14141_), .A3(new_n16680_), .Z(new_n16703_));
  NAND3_X1   g13641(.A1(new_n16701_), .A2(new_n14153_), .A3(new_n16680_), .ZN(new_n16704_));
  AOI21_X1   g13642(.A1(new_n16703_), .A2(new_n16704_), .B(new_n13937_), .ZN(new_n16705_));
  NOR3_X1    g13643(.A1(new_n16705_), .A2(new_n16702_), .A3(new_n13993_), .ZN(new_n16706_));
  OAI21_X1   g13644(.A1(new_n16706_), .A2(new_n16666_), .B(new_n14211_), .ZN(new_n16707_));
  NOR2_X1    g13645(.A1(new_n16665_), .A2(new_n14211_), .ZN(new_n16708_));
  INV_X1     g13646(.I(new_n16708_), .ZN(new_n16709_));
  AOI21_X1   g13647(.A1(new_n16680_), .A2(new_n14254_), .B(pi0644), .ZN(new_n16710_));
  AOI21_X1   g13648(.A1(new_n16707_), .A2(new_n16709_), .B(new_n16710_), .ZN(new_n16711_));
  INV_X1     g13649(.I(new_n16711_), .ZN(new_n16712_));
  NAND2_X1   g13650(.A1(new_n16667_), .A2(new_n13720_), .ZN(new_n16713_));
  NOR2_X1    g13651(.A1(new_n3290_), .A2(new_n3259_), .ZN(new_n16714_));
  INV_X1     g13652(.I(new_n16714_), .ZN(new_n16715_));
  NAND2_X1   g13653(.A1(new_n16715_), .A2(new_n5641_), .ZN(new_n16716_));
  NAND4_X1   g13654(.A1(new_n15655_), .A2(new_n16550_), .A3(new_n16713_), .A4(new_n16716_), .ZN(new_n16717_));
  AOI21_X1   g13655(.A1(new_n16717_), .A2(new_n14424_), .B(new_n5641_), .ZN(new_n16718_));
  NAND2_X1   g13656(.A1(new_n16665_), .A2(new_n16718_), .ZN(new_n16719_));
  NAND2_X1   g13657(.A1(new_n16719_), .A2(new_n3290_), .ZN(new_n16720_));
  NAND2_X1   g13658(.A1(new_n16720_), .A2(pi0698), .ZN(new_n16721_));
  NAND2_X1   g13659(.A1(new_n16721_), .A2(pi0625), .ZN(new_n16722_));
  XOR2_X1    g13660(.A1(new_n16722_), .A2(new_n13620_), .Z(new_n16723_));
  NAND2_X1   g13661(.A1(new_n16723_), .A2(new_n16665_), .ZN(new_n16724_));
  NAND2_X1   g13662(.A1(new_n16724_), .A2(pi0778), .ZN(new_n16725_));
  NAND2_X1   g13663(.A1(new_n16721_), .A2(pi1153), .ZN(new_n16726_));
  XOR2_X1    g13664(.A1(new_n16726_), .A2(new_n13620_), .Z(new_n16727_));
  NAND2_X1   g13665(.A1(new_n16727_), .A2(new_n16665_), .ZN(new_n16728_));
  NOR3_X1    g13666(.A1(new_n16728_), .A2(new_n13748_), .A3(new_n16721_), .ZN(new_n16729_));
  XNOR2_X1   g13667(.A1(new_n16729_), .A2(new_n16725_), .ZN(new_n16730_));
  INV_X1     g13668(.I(new_n16730_), .ZN(new_n16731_));
  INV_X1     g13669(.I(new_n16672_), .ZN(new_n16732_));
  NOR2_X1    g13670(.A1(new_n5641_), .A2(new_n16517_), .ZN(new_n16733_));
  NOR2_X1    g13671(.A1(new_n13453_), .A2(new_n5641_), .ZN(new_n16734_));
  XOR2_X1    g13672(.A1(new_n16734_), .A2(new_n16733_), .Z(new_n16735_));
  NAND2_X1   g13673(.A1(new_n16735_), .A2(new_n13521_), .ZN(new_n16736_));
  NAND3_X1   g13674(.A1(new_n14270_), .A2(pi0145), .A3(pi0767), .ZN(new_n16737_));
  NAND3_X1   g13675(.A1(new_n14272_), .A2(new_n5641_), .A3(pi0767), .ZN(new_n16738_));
  AOI21_X1   g13676(.A1(new_n16737_), .A2(new_n16738_), .B(new_n13152_), .ZN(new_n16739_));
  NAND3_X1   g13677(.A1(new_n13198_), .A2(pi0145), .A3(pi0767), .ZN(new_n16740_));
  NAND3_X1   g13678(.A1(new_n13200_), .A2(pi0145), .A3(new_n16517_), .ZN(new_n16741_));
  AOI21_X1   g13679(.A1(new_n16741_), .A2(new_n16740_), .B(new_n13191_), .ZN(new_n16742_));
  OAI21_X1   g13680(.A1(new_n16739_), .A2(new_n3262_), .B(new_n16742_), .ZN(new_n16743_));
  NAND3_X1   g13681(.A1(new_n16736_), .A2(new_n3183_), .A3(new_n16743_), .ZN(new_n16744_));
  NOR2_X1    g13682(.A1(new_n14284_), .A2(new_n16517_), .ZN(new_n16745_));
  XOR2_X1    g13683(.A1(new_n16745_), .A2(new_n16733_), .Z(new_n16746_));
  NAND3_X1   g13684(.A1(new_n16744_), .A2(new_n16746_), .A3(new_n13359_), .ZN(new_n16747_));
  NAND3_X1   g13685(.A1(new_n16747_), .A2(new_n16550_), .A3(new_n3290_), .ZN(new_n16748_));
  OAI21_X1   g13686(.A1(new_n15587_), .A2(new_n5641_), .B(new_n16517_), .ZN(new_n16749_));
  NAND2_X1   g13687(.A1(new_n16749_), .A2(new_n13209_), .ZN(new_n16750_));
  INV_X1     g13688(.I(new_n13220_), .ZN(new_n16751_));
  OAI21_X1   g13689(.A1(new_n16751_), .A2(new_n5641_), .B(new_n13105_), .ZN(new_n16752_));
  NAND4_X1   g13690(.A1(new_n5503_), .A2(new_n16752_), .A3(new_n3290_), .A4(new_n16733_), .ZN(new_n16753_));
  AOI21_X1   g13691(.A1(new_n16750_), .A2(new_n3259_), .B(new_n16753_), .ZN(new_n16754_));
  NAND2_X1   g13692(.A1(new_n16748_), .A2(new_n16754_), .ZN(new_n16755_));
  AOI21_X1   g13693(.A1(new_n16755_), .A2(new_n16550_), .B(new_n16732_), .ZN(new_n16756_));
  NAND3_X1   g13694(.A1(new_n16756_), .A2(pi0625), .A3(pi1153), .ZN(new_n16757_));
  NOR2_X1    g13695(.A1(new_n16756_), .A2(new_n13613_), .ZN(new_n16758_));
  NAND2_X1   g13696(.A1(new_n16758_), .A2(new_n13620_), .ZN(new_n16759_));
  NAND2_X1   g13697(.A1(new_n16759_), .A2(new_n16757_), .ZN(new_n16760_));
  NAND2_X1   g13698(.A1(new_n16728_), .A2(new_n14081_), .ZN(new_n16761_));
  AOI21_X1   g13699(.A1(new_n16760_), .A2(new_n16679_), .B(new_n16761_), .ZN(new_n16762_));
  NOR2_X1    g13700(.A1(new_n16756_), .A2(new_n13614_), .ZN(new_n16763_));
  NOR2_X1    g13701(.A1(new_n16763_), .A2(new_n13620_), .ZN(new_n16764_));
  NOR3_X1    g13702(.A1(new_n16756_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n16765_));
  OAI21_X1   g13703(.A1(new_n16764_), .A2(new_n16765_), .B(new_n16679_), .ZN(new_n16766_));
  NAND2_X1   g13704(.A1(new_n16766_), .A2(new_n14081_), .ZN(new_n16767_));
  NOR2_X1    g13705(.A1(new_n16724_), .A2(new_n13748_), .ZN(new_n16768_));
  OAI21_X1   g13706(.A1(new_n16767_), .A2(new_n16762_), .B(new_n16768_), .ZN(new_n16769_));
  NOR2_X1    g13707(.A1(new_n16756_), .A2(pi0778), .ZN(new_n16770_));
  INV_X1     g13708(.I(new_n16770_), .ZN(new_n16771_));
  NAND2_X1   g13709(.A1(new_n16769_), .A2(new_n16771_), .ZN(new_n16772_));
  NAND3_X1   g13710(.A1(new_n16772_), .A2(pi0609), .A3(pi1155), .ZN(new_n16773_));
  NAND4_X1   g13711(.A1(new_n16769_), .A2(new_n13766_), .A3(pi1155), .A4(new_n16771_), .ZN(new_n16774_));
  AOI21_X1   g13712(.A1(new_n16773_), .A2(new_n16774_), .B(new_n16731_), .ZN(new_n16775_));
  NAND2_X1   g13713(.A1(new_n16677_), .A2(pi0660), .ZN(new_n16776_));
  OAI21_X1   g13714(.A1(new_n16775_), .A2(new_n16776_), .B(pi0785), .ZN(new_n16777_));
  NAND3_X1   g13715(.A1(new_n16769_), .A2(pi0609), .A3(new_n16771_), .ZN(new_n16778_));
  XOR2_X1    g13716(.A1(new_n16778_), .A2(new_n14694_), .Z(new_n16779_));
  NOR2_X1    g13717(.A1(new_n13801_), .A2(pi0660), .ZN(new_n16780_));
  NAND3_X1   g13718(.A1(new_n16772_), .A2(new_n16685_), .A3(new_n16780_), .ZN(new_n16781_));
  AOI21_X1   g13719(.A1(new_n16779_), .A2(new_n16730_), .B(new_n16781_), .ZN(new_n16782_));
  NAND2_X1   g13720(.A1(new_n16782_), .A2(new_n16777_), .ZN(new_n16783_));
  INV_X1     g13721(.I(new_n16783_), .ZN(new_n16784_));
  NOR2_X1    g13722(.A1(new_n16782_), .A2(new_n16777_), .ZN(new_n16785_));
  NOR2_X1    g13723(.A1(new_n16680_), .A2(new_n13805_), .ZN(new_n16786_));
  AOI21_X1   g13724(.A1(new_n16730_), .A2(new_n13805_), .B(new_n16786_), .ZN(new_n16787_));
  OAI21_X1   g13725(.A1(new_n16680_), .A2(new_n13816_), .B(new_n13877_), .ZN(new_n16788_));
  AOI21_X1   g13726(.A1(new_n16687_), .A2(new_n16788_), .B(new_n13819_), .ZN(new_n16789_));
  AOI21_X1   g13727(.A1(new_n16787_), .A2(new_n16789_), .B(pi0618), .ZN(new_n16790_));
  INV_X1     g13728(.I(new_n16790_), .ZN(new_n16791_));
  OAI21_X1   g13729(.A1(new_n16784_), .A2(new_n16785_), .B(new_n16791_), .ZN(new_n16792_));
  AOI21_X1   g13730(.A1(new_n16680_), .A2(new_n13824_), .B(pi0618), .ZN(new_n16793_));
  NOR3_X1    g13731(.A1(new_n16687_), .A2(pi1154), .A3(new_n16793_), .ZN(new_n16794_));
  OAI21_X1   g13732(.A1(new_n16787_), .A2(new_n13816_), .B(new_n16794_), .ZN(new_n16795_));
  INV_X1     g13733(.I(new_n16795_), .ZN(new_n16796_));
  NOR2_X1    g13734(.A1(new_n16796_), .A2(pi0618), .ZN(new_n16797_));
  NOR2_X1    g13735(.A1(new_n16797_), .A2(new_n13855_), .ZN(new_n16798_));
  OAI21_X1   g13736(.A1(new_n16784_), .A2(new_n16785_), .B(new_n16798_), .ZN(new_n16799_));
  AOI21_X1   g13737(.A1(pi0781), .A2(new_n16792_), .B(new_n16799_), .ZN(new_n16800_));
  INV_X1     g13738(.I(new_n16785_), .ZN(new_n16801_));
  AOI21_X1   g13739(.A1(new_n16801_), .A2(new_n16783_), .B(new_n16790_), .ZN(new_n16802_));
  INV_X1     g13740(.I(new_n16798_), .ZN(new_n16803_));
  AOI21_X1   g13741(.A1(new_n16801_), .A2(new_n16783_), .B(new_n16803_), .ZN(new_n16804_));
  NOR3_X1    g13742(.A1(new_n16802_), .A2(new_n16804_), .A3(new_n13855_), .ZN(new_n16805_));
  OAI21_X1   g13743(.A1(new_n16800_), .A2(new_n16805_), .B(new_n13896_), .ZN(new_n16806_));
  NAND2_X1   g13744(.A1(new_n16806_), .A2(new_n14143_), .ZN(new_n16807_));
  OAI21_X1   g13745(.A1(new_n13855_), .A2(new_n16802_), .B(new_n16804_), .ZN(new_n16808_));
  NAND3_X1   g13746(.A1(new_n16792_), .A2(new_n16799_), .A3(pi0781), .ZN(new_n16809_));
  NAND2_X1   g13747(.A1(new_n16808_), .A2(new_n16809_), .ZN(new_n16810_));
  INV_X1     g13748(.I(new_n16787_), .ZN(new_n16811_));
  NOR2_X1    g13749(.A1(new_n16811_), .A2(new_n13879_), .ZN(new_n16812_));
  AOI21_X1   g13750(.A1(new_n13879_), .A2(new_n16680_), .B(new_n16812_), .ZN(new_n16813_));
  INV_X1     g13751(.I(new_n16813_), .ZN(new_n16814_));
  NOR2_X1    g13752(.A1(new_n16814_), .A2(new_n13860_), .ZN(new_n16815_));
  AOI21_X1   g13753(.A1(new_n16680_), .A2(new_n13885_), .B(pi0619), .ZN(new_n16816_));
  OR3_X2     g13754(.A1(new_n16694_), .A2(pi1159), .A3(new_n16816_), .Z(new_n16817_));
  OAI21_X1   g13755(.A1(new_n16815_), .A2(new_n16817_), .B(new_n13860_), .ZN(new_n16818_));
  AOI21_X1   g13756(.A1(new_n16810_), .A2(new_n16818_), .B(pi0789), .ZN(new_n16819_));
  OAI21_X1   g13757(.A1(new_n16680_), .A2(new_n13860_), .B(new_n13916_), .ZN(new_n16820_));
  AOI21_X1   g13758(.A1(new_n16694_), .A2(new_n16820_), .B(new_n13904_), .ZN(new_n16821_));
  AOI21_X1   g13759(.A1(new_n16814_), .A2(new_n16821_), .B(pi0619), .ZN(new_n16822_));
  AOI21_X1   g13760(.A1(new_n16808_), .A2(new_n16809_), .B(new_n16822_), .ZN(new_n16823_));
  INV_X1     g13761(.I(new_n16823_), .ZN(new_n16824_));
  AOI21_X1   g13762(.A1(new_n16807_), .A2(new_n16819_), .B(new_n16824_), .ZN(new_n16825_));
  INV_X1     g13763(.I(new_n16705_), .ZN(new_n16826_));
  NAND2_X1   g13764(.A1(new_n16813_), .A2(new_n16639_), .ZN(new_n16827_));
  NOR2_X1    g13765(.A1(new_n13919_), .A2(new_n14162_), .ZN(new_n16828_));
  INV_X1     g13766(.I(new_n16828_), .ZN(new_n16829_));
  XOR2_X1    g13767(.A1(new_n16827_), .A2(new_n16829_), .Z(new_n16830_));
  NAND2_X1   g13768(.A1(new_n16830_), .A2(new_n16665_), .ZN(new_n16831_));
  OAI21_X1   g13769(.A1(new_n16831_), .A2(pi1158), .B(new_n13922_), .ZN(new_n16832_));
  AOI21_X1   g13770(.A1(pi1158), .A2(new_n16831_), .B(new_n16832_), .ZN(new_n16833_));
  NOR2_X1    g13771(.A1(new_n16833_), .A2(new_n16826_), .ZN(new_n16834_));
  OAI21_X1   g13772(.A1(new_n16825_), .A2(new_n16423_), .B(new_n16834_), .ZN(new_n16835_));
  NOR2_X1    g13773(.A1(new_n16706_), .A2(new_n16666_), .ZN(new_n16836_));
  INV_X1     g13774(.I(new_n16836_), .ZN(new_n16837_));
  NAND4_X1   g13775(.A1(new_n16787_), .A2(new_n13880_), .A3(new_n15395_), .A4(new_n16665_), .ZN(new_n16838_));
  INV_X1     g13776(.I(new_n15395_), .ZN(new_n16839_));
  NOR4_X1    g13777(.A1(new_n16787_), .A2(new_n13879_), .A3(new_n16839_), .A4(new_n16665_), .ZN(new_n16840_));
  INV_X1     g13778(.I(new_n16840_), .ZN(new_n16841_));
  NAND2_X1   g13779(.A1(new_n16841_), .A2(new_n16838_), .ZN(new_n16842_));
  NAND3_X1   g13780(.A1(new_n16842_), .A2(pi0628), .A3(pi1156), .ZN(new_n16843_));
  NOR3_X1    g13781(.A1(new_n16842_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n16844_));
  INV_X1     g13782(.I(new_n16844_), .ZN(new_n16845_));
  AOI21_X1   g13783(.A1(new_n16845_), .A2(new_n16843_), .B(new_n16680_), .ZN(new_n16846_));
  NAND3_X1   g13784(.A1(new_n16842_), .A2(pi0628), .A3(pi1156), .ZN(new_n16847_));
  NAND4_X1   g13785(.A1(new_n16841_), .A2(new_n13942_), .A3(pi1156), .A4(new_n16838_), .ZN(new_n16848_));
  AOI21_X1   g13786(.A1(new_n16847_), .A2(new_n16848_), .B(new_n16680_), .ZN(new_n16849_));
  NAND4_X1   g13787(.A1(new_n16846_), .A2(pi0792), .A3(new_n16842_), .A4(new_n16849_), .ZN(new_n16850_));
  INV_X1     g13788(.I(new_n16843_), .ZN(new_n16851_));
  OAI21_X1   g13789(.A1(new_n16851_), .A2(new_n16844_), .B(new_n16665_), .ZN(new_n16852_));
  NAND3_X1   g13790(.A1(new_n16849_), .A2(pi0792), .A3(new_n16842_), .ZN(new_n16853_));
  NAND3_X1   g13791(.A1(new_n16853_), .A2(pi0792), .A3(new_n16852_), .ZN(new_n16854_));
  AOI21_X1   g13792(.A1(new_n16854_), .A2(new_n16850_), .B(pi0647), .ZN(new_n16855_));
  NOR2_X1    g13793(.A1(new_n16680_), .A2(new_n14005_), .ZN(new_n16856_));
  OAI21_X1   g13794(.A1(new_n16855_), .A2(new_n16856_), .B(new_n14011_), .ZN(new_n16857_));
  NAND2_X1   g13795(.A1(new_n16854_), .A2(new_n16850_), .ZN(new_n16858_));
  AOI21_X1   g13796(.A1(new_n16665_), .A2(new_n14005_), .B(new_n14006_), .ZN(new_n16859_));
  INV_X1     g13797(.I(new_n16859_), .ZN(new_n16860_));
  AOI21_X1   g13798(.A1(new_n16858_), .A2(pi0647), .B(new_n16860_), .ZN(new_n16861_));
  NAND3_X1   g13799(.A1(new_n16857_), .A2(new_n16861_), .A3(new_n14010_), .ZN(new_n16862_));
  NOR2_X1    g13800(.A1(new_n16855_), .A2(new_n16856_), .ZN(new_n16863_));
  NOR3_X1    g13801(.A1(new_n16863_), .A2(new_n14010_), .A3(new_n14006_), .ZN(new_n16864_));
  INV_X1     g13802(.I(new_n16864_), .ZN(new_n16865_));
  AOI21_X1   g13803(.A1(new_n16865_), .A2(new_n16862_), .B(new_n12776_), .ZN(new_n16866_));
  INV_X1     g13804(.I(new_n16576_), .ZN(new_n16867_));
  NOR2_X1    g13805(.A1(new_n16419_), .A2(new_n16867_), .ZN(new_n16868_));
  OAI21_X1   g13806(.A1(new_n16866_), .A2(new_n16837_), .B(new_n16868_), .ZN(new_n16869_));
  NAND2_X1   g13807(.A1(new_n16869_), .A2(new_n16835_), .ZN(new_n16870_));
  INV_X1     g13808(.I(new_n16702_), .ZN(new_n16871_));
  INV_X1     g13809(.I(new_n13985_), .ZN(new_n16872_));
  NOR2_X1    g13810(.A1(new_n16872_), .A2(new_n13942_), .ZN(new_n16873_));
  AOI21_X1   g13811(.A1(new_n13942_), .A2(new_n13977_), .B(new_n16873_), .ZN(new_n16874_));
  INV_X1     g13812(.I(new_n16874_), .ZN(new_n16875_));
  NOR2_X1    g13813(.A1(new_n16846_), .A2(new_n13976_), .ZN(new_n16876_));
  NOR2_X1    g13814(.A1(new_n16849_), .A2(pi0629), .ZN(new_n16877_));
  OAI21_X1   g13815(.A1(new_n16876_), .A2(new_n16877_), .B(pi0792), .ZN(new_n16878_));
  AOI22_X1   g13816(.A1(new_n16826_), .A2(new_n16871_), .B1(new_n16875_), .B2(new_n16878_), .ZN(new_n16879_));
  NAND3_X1   g13817(.A1(new_n16870_), .A2(pi0790), .A3(new_n16879_), .ZN(new_n16880_));
  AOI21_X1   g13818(.A1(new_n16880_), .A2(new_n14204_), .B(new_n16712_), .ZN(new_n16881_));
  NAND4_X1   g13819(.A1(new_n16870_), .A2(pi0644), .A3(pi0715), .A4(new_n16879_), .ZN(new_n16882_));
  AOI21_X1   g13820(.A1(new_n16810_), .A2(new_n13896_), .B(new_n15479_), .ZN(new_n16883_));
  OAI21_X1   g13821(.A1(new_n16800_), .A2(new_n16805_), .B(new_n16818_), .ZN(new_n16884_));
  NAND2_X1   g13822(.A1(new_n16884_), .A2(new_n13896_), .ZN(new_n16885_));
  OAI21_X1   g13823(.A1(new_n16885_), .A2(new_n16883_), .B(new_n16823_), .ZN(new_n16886_));
  INV_X1     g13824(.I(new_n16834_), .ZN(new_n16887_));
  AOI21_X1   g13825(.A1(new_n16886_), .A2(new_n16424_), .B(new_n16887_), .ZN(new_n16888_));
  INV_X1     g13826(.I(new_n16862_), .ZN(new_n16889_));
  OAI21_X1   g13827(.A1(new_n16889_), .A2(new_n16864_), .B(pi0787), .ZN(new_n16890_));
  INV_X1     g13828(.I(new_n16868_), .ZN(new_n16891_));
  AOI21_X1   g13829(.A1(new_n16890_), .A2(new_n16836_), .B(new_n16891_), .ZN(new_n16892_));
  OAI21_X1   g13830(.A1(new_n16892_), .A2(new_n16888_), .B(new_n16879_), .ZN(new_n16893_));
  NAND3_X1   g13831(.A1(new_n16893_), .A2(pi0644), .A3(new_n14200_), .ZN(new_n16894_));
  AOI21_X1   g13832(.A1(new_n14006_), .A2(new_n16863_), .B(new_n16861_), .ZN(new_n16895_));
  NOR2_X1    g13833(.A1(new_n16895_), .A2(new_n12776_), .ZN(new_n16896_));
  NOR2_X1    g13834(.A1(new_n16858_), .A2(pi0787), .ZN(new_n16897_));
  AOI21_X1   g13835(.A1(new_n16837_), .A2(new_n14211_), .B(new_n16708_), .ZN(new_n16898_));
  NOR2_X1    g13836(.A1(new_n14243_), .A2(pi0644), .ZN(new_n16899_));
  AOI21_X1   g13837(.A1(new_n16711_), .A2(pi0715), .B(pi0644), .ZN(new_n16900_));
  OAI21_X1   g13838(.A1(new_n16896_), .A2(new_n16897_), .B(pi0790), .ZN(new_n16901_));
  OAI22_X1   g13839(.A1(new_n16901_), .A2(new_n16900_), .B1(new_n16898_), .B2(new_n16899_), .ZN(new_n16902_));
  OAI21_X1   g13840(.A1(new_n16896_), .A2(new_n16897_), .B(new_n16902_), .ZN(new_n16903_));
  AOI21_X1   g13841(.A1(new_n16894_), .A2(new_n16882_), .B(new_n16903_), .ZN(new_n16904_));
  OAI21_X1   g13842(.A1(new_n16904_), .A2(new_n16881_), .B(new_n7240_), .ZN(new_n16905_));
  AOI21_X1   g13843(.A1(po1038), .A2(new_n5641_), .B(pi0832), .ZN(new_n16906_));
  AOI21_X1   g13844(.A1(new_n16905_), .A2(new_n16906_), .B(new_n16664_), .ZN(po0302));
  NOR4_X1    g13845(.A1(new_n14833_), .A2(new_n14921_), .A3(new_n5741_), .A4(new_n5800_), .ZN(new_n16908_));
  NOR2_X1    g13846(.A1(new_n14921_), .A2(new_n5741_), .ZN(new_n16909_));
  NOR3_X1    g13847(.A1(new_n16909_), .A2(pi0735), .A3(new_n5800_), .ZN(new_n16910_));
  NOR2_X1    g13848(.A1(new_n16910_), .A2(new_n16908_), .ZN(new_n16911_));
  NAND2_X1   g13849(.A1(new_n16911_), .A2(pi0832), .ZN(new_n16912_));
  NOR2_X1    g13850(.A1(new_n2723_), .A2(new_n14799_), .ZN(new_n16913_));
  XOR2_X1    g13851(.A1(new_n16912_), .A2(new_n16913_), .Z(new_n16914_));
  INV_X1     g13852(.I(new_n16911_), .ZN(new_n16915_));
  NOR2_X1    g13853(.A1(new_n12784_), .A2(pi0146), .ZN(new_n16916_));
  AOI21_X1   g13854(.A1(new_n12784_), .A2(new_n16915_), .B(new_n16916_), .ZN(new_n16917_));
  INV_X1     g13855(.I(new_n16917_), .ZN(new_n16918_));
  AOI21_X1   g13856(.A1(new_n13086_), .A2(new_n5452_), .B(new_n14833_), .ZN(new_n16919_));
  NOR2_X1    g13857(.A1(new_n5451_), .A2(pi0907), .ZN(new_n16920_));
  INV_X1     g13858(.I(new_n16920_), .ZN(new_n16921_));
  NAND2_X1   g13859(.A1(new_n16921_), .A2(pi0146), .ZN(new_n16922_));
  NOR4_X1    g13860(.A1(new_n12974_), .A2(pi0743), .A3(new_n5800_), .A4(new_n16922_), .ZN(new_n16923_));
  NOR2_X1    g13861(.A1(new_n16919_), .A2(new_n16923_), .ZN(new_n16924_));
  NAND3_X1   g13862(.A1(new_n12980_), .A2(pi0146), .A3(new_n16920_), .ZN(new_n16925_));
  OAI21_X1   g13863(.A1(new_n16924_), .A2(new_n16925_), .B(new_n3312_), .ZN(new_n16926_));
  XOR2_X1    g13864(.A1(new_n16926_), .A2(new_n12833_), .Z(new_n16927_));
  NAND2_X1   g13865(.A1(new_n16927_), .A2(new_n16918_), .ZN(new_n16928_));
  NAND2_X1   g13866(.A1(new_n13078_), .A2(new_n16911_), .ZN(new_n16929_));
  NAND2_X1   g13867(.A1(new_n13078_), .A2(new_n5398_), .ZN(new_n16930_));
  XOR2_X1    g13868(.A1(new_n16929_), .A2(new_n16930_), .Z(new_n16931_));
  AOI21_X1   g13869(.A1(new_n16931_), .A2(pi0146), .B(new_n3512_), .ZN(new_n16932_));
  NOR2_X1    g13870(.A1(new_n16915_), .A2(new_n5397_), .ZN(new_n16933_));
  XOR2_X1    g13871(.A1(new_n13091_), .A2(new_n16933_), .Z(new_n16934_));
  NOR3_X1    g13872(.A1(new_n16932_), .A2(new_n2847_), .A3(new_n16934_), .ZN(new_n16935_));
  OAI21_X1   g13873(.A1(new_n16917_), .A2(new_n3092_), .B(new_n3090_), .ZN(new_n16936_));
  NOR3_X1    g13874(.A1(new_n13086_), .A2(new_n5397_), .A3(new_n16911_), .ZN(new_n16937_));
  NOR3_X1    g13875(.A1(new_n13086_), .A2(new_n5398_), .A3(new_n16915_), .ZN(new_n16938_));
  OAI21_X1   g13876(.A1(new_n16937_), .A2(new_n16938_), .B(pi0146), .ZN(new_n16939_));
  NAND2_X1   g13877(.A1(new_n12973_), .A2(new_n5398_), .ZN(new_n16940_));
  XNOR2_X1   g13878(.A1(new_n16940_), .A2(new_n16933_), .ZN(new_n16941_));
  NAND2_X1   g13879(.A1(new_n16941_), .A2(pi0146), .ZN(new_n16942_));
  NAND2_X1   g13880(.A1(new_n3092_), .A2(pi0299), .ZN(new_n16943_));
  AOI21_X1   g13881(.A1(new_n16942_), .A2(new_n16939_), .B(new_n16943_), .ZN(new_n16944_));
  OAI21_X1   g13882(.A1(new_n16935_), .A2(new_n16936_), .B(new_n16944_), .ZN(new_n16945_));
  NAND2_X1   g13883(.A1(new_n16929_), .A2(pi0215), .ZN(new_n16946_));
  NAND3_X1   g13884(.A1(new_n16946_), .A2(new_n2847_), .A3(new_n13081_), .ZN(new_n16947_));
  NAND2_X1   g13885(.A1(new_n16911_), .A2(pi0299), .ZN(new_n16948_));
  XOR2_X1    g13886(.A1(new_n13069_), .A2(new_n16948_), .Z(new_n16949_));
  AOI21_X1   g13887(.A1(new_n16949_), .A2(pi0146), .B(new_n3212_), .ZN(new_n16950_));
  NAND2_X1   g13888(.A1(new_n13162_), .A2(new_n16911_), .ZN(new_n16951_));
  XOR2_X1    g13889(.A1(new_n13163_), .A2(new_n16951_), .Z(new_n16952_));
  NOR3_X1    g13890(.A1(new_n5504_), .A2(new_n2847_), .A3(new_n2723_), .ZN(new_n16954_));
  NAND2_X1   g13891(.A1(new_n16952_), .A2(new_n16954_), .ZN(new_n16955_));
  OAI21_X1   g13892(.A1(new_n16955_), .A2(new_n16950_), .B(new_n3183_), .ZN(new_n16956_));
  NAND3_X1   g13893(.A1(new_n16956_), .A2(new_n13080_), .A3(new_n16947_), .ZN(new_n16957_));
  AOI21_X1   g13894(.A1(new_n16945_), .A2(new_n16928_), .B(new_n16957_), .ZN(new_n16958_));
  OAI21_X1   g13895(.A1(new_n8297_), .A2(pi0146), .B(new_n14799_), .ZN(new_n16959_));
  OAI22_X1   g13896(.A1(new_n16958_), .A2(new_n16959_), .B1(new_n2847_), .B2(new_n16914_), .ZN(po0303));
  INV_X1     g13897(.I(new_n16913_), .ZN(new_n16961_));
  INV_X1     g13898(.I(pi0726), .ZN(new_n16962_));
  NAND2_X1   g13899(.A1(pi0770), .A2(pi0907), .ZN(new_n16963_));
  NAND3_X1   g13900(.A1(new_n16963_), .A2(new_n16962_), .A3(pi0947), .ZN(new_n16964_));
  NAND4_X1   g13901(.A1(pi0726), .A2(pi0770), .A3(pi0907), .A4(pi0947), .ZN(new_n16965_));
  NAND3_X1   g13902(.A1(new_n16964_), .A2(pi0832), .A3(new_n16965_), .ZN(new_n16966_));
  XOR2_X1    g13903(.A1(new_n16966_), .A2(new_n16961_), .Z(new_n16967_));
  NOR2_X1    g13904(.A1(new_n5741_), .A2(pi0947), .ZN(new_n16968_));
  INV_X1     g13905(.I(new_n16968_), .ZN(new_n16969_));
  NOR2_X1    g13906(.A1(new_n14298_), .A2(new_n16969_), .ZN(new_n16970_));
  AOI21_X1   g13907(.A1(new_n12986_), .A2(new_n12988_), .B(new_n12991_), .ZN(new_n16971_));
  AOI21_X1   g13908(.A1(new_n16971_), .A2(new_n16968_), .B(pi0299), .ZN(new_n16972_));
  INV_X1     g13909(.I(new_n16972_), .ZN(new_n16973_));
  NOR2_X1    g13910(.A1(new_n13086_), .A2(new_n16969_), .ZN(new_n16974_));
  NOR2_X1    g13911(.A1(new_n16974_), .A2(new_n3312_), .ZN(new_n16975_));
  NOR2_X1    g13912(.A1(new_n16975_), .A2(new_n3111_), .ZN(new_n16976_));
  NOR2_X1    g13913(.A1(new_n12935_), .A2(new_n16969_), .ZN(new_n16977_));
  NOR2_X1    g13914(.A1(new_n12809_), .A2(new_n16969_), .ZN(new_n16978_));
  NOR2_X1    g13915(.A1(new_n16978_), .A2(new_n3313_), .ZN(new_n16979_));
  NAND3_X1   g13916(.A1(new_n16977_), .A2(pi0215), .A3(new_n16979_), .ZN(new_n16980_));
  XOR2_X1    g13917(.A1(new_n16976_), .A2(new_n16980_), .Z(new_n16981_));
  NAND2_X1   g13918(.A1(new_n16981_), .A2(pi0299), .ZN(new_n16982_));
  NAND2_X1   g13919(.A1(new_n16982_), .A2(new_n16973_), .ZN(new_n16983_));
  NOR2_X1    g13920(.A1(new_n16983_), .A2(new_n3183_), .ZN(new_n16984_));
  AOI21_X1   g13921(.A1(new_n3183_), .A2(new_n16970_), .B(new_n16984_), .ZN(new_n16985_));
  NOR2_X1    g13922(.A1(new_n3259_), .A2(new_n9530_), .ZN(new_n16986_));
  NOR2_X1    g13923(.A1(new_n16968_), .A2(new_n3183_), .ZN(new_n16987_));
  NOR2_X1    g13924(.A1(new_n16968_), .A2(new_n3098_), .ZN(new_n16988_));
  NOR2_X1    g13925(.A1(new_n13086_), .A2(new_n5800_), .ZN(new_n16989_));
  AOI21_X1   g13926(.A1(new_n13086_), .A2(new_n5451_), .B(new_n5453_), .ZN(new_n16990_));
  OAI21_X1   g13927(.A1(new_n5451_), .A2(new_n12973_), .B(new_n16990_), .ZN(new_n16991_));
  INV_X1     g13928(.I(new_n16991_), .ZN(new_n16992_));
  NOR2_X1    g13929(.A1(new_n16992_), .A2(new_n16989_), .ZN(new_n16993_));
  NOR2_X1    g13930(.A1(new_n16993_), .A2(new_n3312_), .ZN(new_n16994_));
  NOR2_X1    g13931(.A1(new_n16994_), .A2(new_n3111_), .ZN(new_n16995_));
  INV_X1     g13932(.I(new_n13343_), .ZN(new_n16996_));
  NOR2_X1    g13933(.A1(new_n16996_), .A2(new_n16968_), .ZN(new_n16997_));
  NAND3_X1   g13934(.A1(new_n13080_), .A2(pi0215), .A3(new_n16997_), .ZN(new_n16998_));
  XOR2_X1    g13935(.A1(new_n16995_), .A2(new_n16998_), .Z(new_n16999_));
  INV_X1     g13936(.I(new_n16999_), .ZN(new_n17000_));
  NOR3_X1    g13937(.A1(new_n12935_), .A2(new_n3111_), .A3(new_n5800_), .ZN(new_n17001_));
  NOR2_X1    g13938(.A1(new_n17000_), .A2(new_n17001_), .ZN(new_n17002_));
  INV_X1     g13939(.I(new_n16971_), .ZN(new_n17003_));
  NOR2_X1    g13940(.A1(new_n17003_), .A2(new_n3098_), .ZN(new_n17004_));
  NAND2_X1   g13941(.A1(new_n17002_), .A2(new_n17004_), .ZN(new_n17005_));
  NOR2_X1    g13942(.A1(new_n17005_), .A2(new_n16988_), .ZN(new_n17006_));
  NAND2_X1   g13943(.A1(new_n17005_), .A2(new_n16988_), .ZN(new_n17007_));
  INV_X1     g13944(.I(new_n17007_), .ZN(new_n17008_));
  NOR2_X1    g13945(.A1(new_n17008_), .A2(new_n17006_), .ZN(new_n17009_));
  NOR2_X1    g13946(.A1(new_n17009_), .A2(new_n13071_), .ZN(new_n17010_));
  INV_X1     g13947(.I(new_n17010_), .ZN(new_n17011_));
  NOR2_X1    g13948(.A1(new_n17011_), .A2(new_n16987_), .ZN(new_n17012_));
  NAND2_X1   g13949(.A1(new_n17011_), .A2(new_n16987_), .ZN(new_n17013_));
  INV_X1     g13950(.I(new_n17013_), .ZN(new_n17014_));
  NOR2_X1    g13951(.A1(new_n17014_), .A2(new_n17012_), .ZN(new_n17015_));
  NAND2_X1   g13952(.A1(new_n17015_), .A2(pi0147), .ZN(new_n17016_));
  XOR2_X1    g13953(.A1(new_n17016_), .A2(new_n16986_), .Z(new_n17017_));
  NOR2_X1    g13954(.A1(new_n17017_), .A2(new_n16985_), .ZN(new_n17018_));
  INV_X1     g13955(.I(pi0770), .ZN(new_n17019_));
  NAND2_X1   g13956(.A1(new_n16962_), .A2(new_n17019_), .ZN(new_n17020_));
  AOI21_X1   g13957(.A1(new_n13108_), .A2(new_n16968_), .B(new_n3259_), .ZN(new_n17021_));
  INV_X1     g13958(.I(new_n17021_), .ZN(new_n17022_));
  AOI21_X1   g13959(.A1(new_n9530_), .A2(new_n13109_), .B(new_n17022_), .ZN(new_n17023_));
  OAI21_X1   g13960(.A1(new_n17018_), .A2(new_n17020_), .B(new_n17023_), .ZN(new_n17024_));
  NOR2_X1    g13961(.A1(new_n13109_), .A2(new_n5452_), .ZN(new_n17025_));
  NOR2_X1    g13962(.A1(new_n17025_), .A2(new_n3259_), .ZN(new_n17026_));
  NOR2_X1    g13963(.A1(new_n13625_), .A2(new_n5453_), .ZN(new_n17027_));
  INV_X1     g13964(.I(new_n17027_), .ZN(new_n17028_));
  NAND2_X1   g13965(.A1(new_n17028_), .A2(new_n9530_), .ZN(new_n17029_));
  AOI21_X1   g13966(.A1(new_n17029_), .A2(new_n17026_), .B(pi0770), .ZN(new_n17030_));
  NOR2_X1    g13967(.A1(new_n14298_), .A2(new_n5452_), .ZN(new_n17031_));
  NAND2_X1   g13968(.A1(new_n17031_), .A2(new_n3183_), .ZN(new_n17032_));
  NOR2_X1    g13969(.A1(new_n12942_), .A2(new_n3111_), .ZN(new_n17033_));
  INV_X1     g13970(.I(new_n17033_), .ZN(new_n17034_));
  NAND2_X1   g13971(.A1(new_n17034_), .A2(pi0299), .ZN(new_n17035_));
  NOR2_X1    g13972(.A1(new_n17003_), .A2(new_n5452_), .ZN(new_n17036_));
  NOR2_X1    g13973(.A1(new_n12839_), .A2(new_n12834_), .ZN(new_n17037_));
  NAND2_X1   g13974(.A1(new_n12784_), .A2(new_n5453_), .ZN(new_n17038_));
  NOR3_X1    g13975(.A1(new_n17037_), .A2(new_n3098_), .A3(new_n17038_), .ZN(new_n17039_));
  NAND2_X1   g13976(.A1(new_n17036_), .A2(new_n17039_), .ZN(new_n17040_));
  XNOR2_X1   g13977(.A1(new_n17040_), .A2(new_n17035_), .ZN(new_n17041_));
  INV_X1     g13978(.I(new_n17041_), .ZN(new_n17042_));
  OAI21_X1   g13979(.A1(new_n17042_), .A2(new_n3183_), .B(new_n17032_), .ZN(new_n17043_));
  NOR2_X1    g13980(.A1(new_n14874_), .A2(new_n3183_), .ZN(new_n17044_));
  NOR2_X1    g13981(.A1(new_n12990_), .A2(new_n12989_), .ZN(new_n17045_));
  NOR2_X1    g13982(.A1(new_n17045_), .A2(pi0947), .ZN(new_n17046_));
  NOR2_X1    g13983(.A1(new_n17046_), .A2(new_n3090_), .ZN(new_n17047_));
  INV_X1     g13984(.I(new_n17047_), .ZN(new_n17048_));
  NAND2_X1   g13985(.A1(new_n12987_), .A2(new_n3160_), .ZN(new_n17049_));
  NAND2_X1   g13986(.A1(new_n12986_), .A2(new_n17049_), .ZN(new_n17050_));
  AOI21_X1   g13987(.A1(new_n17050_), .A2(new_n5452_), .B(pi0223), .ZN(new_n17051_));
  INV_X1     g13988(.I(new_n17045_), .ZN(new_n17052_));
  AOI21_X1   g13989(.A1(new_n17052_), .A2(new_n16969_), .B(new_n3090_), .ZN(new_n17053_));
  NOR3_X1    g13990(.A1(new_n17051_), .A2(pi0299), .A3(new_n17053_), .ZN(new_n17054_));
  NOR2_X1    g13991(.A1(new_n17054_), .A2(new_n17048_), .ZN(new_n17055_));
  AOI21_X1   g13992(.A1(pi0299), .A2(new_n17055_), .B(new_n17000_), .ZN(new_n17056_));
  NOR2_X1    g13993(.A1(new_n17056_), .A2(new_n5800_), .ZN(new_n17057_));
  INV_X1     g13994(.I(new_n17057_), .ZN(new_n17058_));
  NOR3_X1    g13995(.A1(new_n17058_), .A2(new_n3183_), .A3(new_n5453_), .ZN(new_n17059_));
  XNOR2_X1   g13996(.A1(new_n17059_), .A2(new_n17044_), .ZN(new_n17060_));
  NAND2_X1   g13997(.A1(new_n17060_), .A2(pi0147), .ZN(new_n17061_));
  XNOR2_X1   g13998(.A1(new_n17061_), .A2(new_n16986_), .ZN(new_n17062_));
  NAND2_X1   g13999(.A1(new_n17062_), .A2(new_n17043_), .ZN(new_n17063_));
  AOI21_X1   g14000(.A1(new_n17024_), .A2(new_n17030_), .B(new_n17063_), .ZN(new_n17064_));
  NOR3_X1    g14001(.A1(new_n13625_), .A2(new_n3259_), .A3(pi0947), .ZN(new_n17065_));
  AOI21_X1   g14002(.A1(new_n14874_), .A2(new_n5800_), .B(pi0039), .ZN(new_n17066_));
  NOR2_X1    g14003(.A1(new_n3098_), .A2(pi0947), .ZN(new_n17067_));
  OAI21_X1   g14004(.A1(new_n13086_), .A2(new_n16969_), .B(new_n16991_), .ZN(new_n17068_));
  NAND2_X1   g14005(.A1(new_n17068_), .A2(new_n3313_), .ZN(new_n17069_));
  NAND2_X1   g14006(.A1(new_n17069_), .A2(new_n3111_), .ZN(new_n17070_));
  INV_X1     g14007(.I(new_n17070_), .ZN(new_n17071_));
  NOR2_X1    g14008(.A1(new_n13080_), .A2(new_n3111_), .ZN(new_n17072_));
  INV_X1     g14009(.I(new_n17072_), .ZN(new_n17073_));
  NOR2_X1    g14010(.A1(new_n17073_), .A2(new_n16977_), .ZN(new_n17074_));
  NAND2_X1   g14011(.A1(new_n17071_), .A2(new_n17074_), .ZN(new_n17075_));
  AOI21_X1   g14012(.A1(new_n17075_), .A2(new_n16996_), .B(new_n5800_), .ZN(new_n17076_));
  NAND2_X1   g14013(.A1(new_n17076_), .A2(new_n17004_), .ZN(new_n17077_));
  XOR2_X1    g14014(.A1(new_n17077_), .A2(new_n17067_), .Z(new_n17078_));
  AOI21_X1   g14015(.A1(new_n17078_), .A2(pi0039), .B(new_n17066_), .ZN(new_n17079_));
  AND2_X2    g14016(.A1(new_n17079_), .A2(new_n3259_), .Z(new_n17080_));
  NOR2_X1    g14017(.A1(new_n17080_), .A2(new_n17065_), .ZN(new_n17081_));
  NAND3_X1   g14018(.A1(new_n17081_), .A2(pi0147), .A3(pi0770), .ZN(new_n17082_));
  OR3_X2     g14019(.A1(new_n17081_), .A2(pi0147), .A3(new_n17019_), .Z(new_n17083_));
  AOI21_X1   g14020(.A1(new_n13624_), .A2(pi0947), .B(new_n3259_), .ZN(new_n17084_));
  AOI21_X1   g14021(.A1(new_n14874_), .A2(pi0947), .B(pi0039), .ZN(new_n17085_));
  INV_X1     g14022(.I(new_n17085_), .ZN(new_n17086_));
  AOI21_X1   g14023(.A1(new_n16971_), .A2(pi0947), .B(pi0299), .ZN(new_n17087_));
  NOR2_X1    g14024(.A1(new_n12809_), .A2(new_n5800_), .ZN(new_n17088_));
  NOR2_X1    g14025(.A1(new_n17088_), .A2(new_n3313_), .ZN(new_n17089_));
  NOR2_X1    g14026(.A1(new_n17089_), .A2(pi0215), .ZN(new_n17090_));
  OAI21_X1   g14027(.A1(new_n16989_), .A2(new_n3312_), .B(new_n17090_), .ZN(new_n17091_));
  INV_X1     g14028(.I(new_n17091_), .ZN(new_n17092_));
  NOR2_X1    g14029(.A1(new_n17001_), .A2(new_n3098_), .ZN(new_n17093_));
  INV_X1     g14030(.I(new_n17093_), .ZN(new_n17094_));
  NOR2_X1    g14031(.A1(new_n17094_), .A2(new_n17092_), .ZN(new_n17095_));
  NOR2_X1    g14032(.A1(new_n17087_), .A2(new_n17095_), .ZN(new_n17096_));
  OAI21_X1   g14033(.A1(new_n17096_), .A2(new_n3183_), .B(new_n17086_), .ZN(new_n17097_));
  AOI21_X1   g14034(.A1(new_n17097_), .A2(new_n3259_), .B(new_n17084_), .ZN(new_n17098_));
  INV_X1     g14035(.I(new_n17098_), .ZN(new_n17099_));
  NAND3_X1   g14036(.A1(new_n17099_), .A2(new_n9530_), .A3(new_n16962_), .ZN(new_n17100_));
  NAND3_X1   g14037(.A1(new_n17100_), .A2(pi0770), .A3(new_n13634_), .ZN(new_n17101_));
  AOI21_X1   g14038(.A1(new_n17083_), .A2(new_n17082_), .B(new_n17101_), .ZN(new_n17102_));
  OAI21_X1   g14039(.A1(new_n17064_), .A2(new_n8297_), .B(new_n17102_), .ZN(new_n17103_));
  AOI21_X1   g14040(.A1(new_n8345_), .A2(new_n9530_), .B(pi0832), .ZN(new_n17104_));
  AOI22_X1   g14041(.A1(new_n17103_), .A2(new_n17104_), .B1(pi0147), .B2(new_n16967_), .ZN(po0304));
  NAND2_X1   g14042(.A1(new_n16971_), .A2(new_n3098_), .ZN(new_n17106_));
  OAI21_X1   g14043(.A1(new_n16981_), .A2(new_n3098_), .B(new_n17106_), .ZN(new_n17107_));
  OAI21_X1   g14044(.A1(new_n17107_), .A2(new_n4329_), .B(new_n14263_), .ZN(new_n17108_));
  OAI21_X1   g14045(.A1(new_n17009_), .A2(new_n17108_), .B(new_n3098_), .ZN(new_n17109_));
  NAND2_X1   g14046(.A1(new_n17109_), .A2(pi0148), .ZN(new_n17110_));
  NOR2_X1    g14047(.A1(new_n5800_), .A2(pi0749), .ZN(new_n17111_));
  OAI21_X1   g14048(.A1(new_n14874_), .A2(pi0148), .B(new_n15599_), .ZN(new_n17112_));
  OAI21_X1   g14049(.A1(new_n5452_), .A2(new_n14298_), .B(new_n17112_), .ZN(new_n17113_));
  AOI21_X1   g14050(.A1(new_n17113_), .A2(new_n17111_), .B(pi0039), .ZN(new_n17114_));
  NOR3_X1    g14051(.A1(new_n17058_), .A2(new_n4329_), .A3(new_n14263_), .ZN(new_n17115_));
  NOR3_X1    g14052(.A1(new_n17057_), .A2(pi0148), .A3(new_n14263_), .ZN(new_n17116_));
  OAI21_X1   g14053(.A1(new_n17115_), .A2(new_n17116_), .B(new_n17042_), .ZN(new_n17117_));
  AOI21_X1   g14054(.A1(new_n17110_), .A2(new_n17114_), .B(new_n17117_), .ZN(new_n17118_));
  NAND3_X1   g14055(.A1(new_n13108_), .A2(pi0148), .A3(new_n17111_), .ZN(new_n17119_));
  XOR2_X1    g14056(.A1(new_n17025_), .A2(new_n17119_), .Z(new_n17120_));
  NOR2_X1    g14057(.A1(new_n17120_), .A2(new_n3259_), .ZN(new_n17121_));
  OAI21_X1   g14058(.A1(new_n17118_), .A2(pi0706), .B(new_n17121_), .ZN(new_n17122_));
  NOR2_X1    g14059(.A1(new_n3290_), .A2(new_n5788_), .ZN(new_n17123_));
  INV_X1     g14060(.I(new_n17123_), .ZN(new_n17124_));
  NOR2_X1    g14061(.A1(new_n17076_), .A2(new_n3098_), .ZN(new_n17125_));
  XOR2_X1    g14062(.A1(new_n17125_), .A2(new_n12666_), .Z(new_n17126_));
  INV_X1     g14063(.I(new_n14366_), .ZN(new_n17127_));
  AOI21_X1   g14064(.A1(new_n17087_), .A2(pi0749), .B(pi0148), .ZN(new_n17128_));
  OAI21_X1   g14065(.A1(new_n14263_), .A2(new_n5800_), .B(new_n17112_), .ZN(new_n17129_));
  NAND3_X1   g14066(.A1(new_n3183_), .A2(new_n4329_), .A3(new_n14263_), .ZN(new_n17130_));
  NAND3_X1   g14067(.A1(new_n17129_), .A2(new_n14874_), .A3(new_n17130_), .ZN(new_n17131_));
  OAI22_X1   g14068(.A1(new_n17127_), .A2(new_n17131_), .B1(new_n17128_), .B2(new_n17003_), .ZN(new_n17132_));
  NOR2_X1    g14069(.A1(new_n17092_), .A2(new_n17001_), .ZN(new_n17133_));
  NOR2_X1    g14070(.A1(new_n14263_), .A2(new_n5800_), .ZN(new_n17134_));
  NOR2_X1    g14071(.A1(new_n13109_), .A2(new_n17134_), .ZN(new_n17135_));
  NAND2_X1   g14072(.A1(pi0038), .A2(pi0706), .ZN(new_n17136_));
  OAI21_X1   g14073(.A1(new_n17135_), .A2(new_n17136_), .B(new_n4329_), .ZN(new_n17137_));
  NAND2_X1   g14074(.A1(new_n17124_), .A2(new_n4329_), .ZN(new_n17138_));
  NOR2_X1    g14075(.A1(new_n17134_), .A2(new_n9992_), .ZN(new_n17139_));
  NAND2_X1   g14076(.A1(new_n16968_), .A2(pi0706), .ZN(new_n17140_));
  OAI21_X1   g14077(.A1(new_n17139_), .A2(new_n17140_), .B(new_n14799_), .ZN(new_n17141_));
  NOR4_X1    g14078(.A1(new_n2723_), .A2(pi0057), .A3(new_n4329_), .A4(pi0832), .ZN(new_n17142_));
  AOI22_X1   g14079(.A1(new_n17138_), .A2(new_n5371_), .B1(new_n17141_), .B2(new_n17142_), .ZN(new_n17143_));
  NOR2_X1    g14080(.A1(new_n13625_), .A2(new_n17143_), .ZN(new_n17144_));
  AND3_X2    g14081(.A1(new_n17133_), .A2(new_n17137_), .A3(new_n17144_), .Z(new_n17145_));
  NAND3_X1   g14082(.A1(new_n17126_), .A2(new_n17132_), .A3(new_n17145_), .ZN(new_n17146_));
  AOI21_X1   g14083(.A1(new_n17122_), .A2(new_n17124_), .B(new_n17146_), .ZN(po0305));
  INV_X1     g14084(.I(pi0725), .ZN(new_n17148_));
  NOR2_X1    g14085(.A1(new_n5800_), .A2(pi0755), .ZN(new_n17149_));
  NOR2_X1    g14086(.A1(new_n14298_), .A2(new_n17149_), .ZN(new_n17150_));
  XOR2_X1    g14087(.A1(new_n17150_), .A2(new_n13094_), .Z(new_n17151_));
  NAND2_X1   g14088(.A1(new_n17151_), .A2(pi0149), .ZN(new_n17152_));
  INV_X1     g14089(.I(pi0755), .ZN(new_n17153_));
  NOR3_X1    g14090(.A1(new_n17058_), .A2(new_n7475_), .A3(new_n17153_), .ZN(new_n17154_));
  NOR3_X1    g14091(.A1(new_n17057_), .A2(new_n7475_), .A3(pi0755), .ZN(new_n17155_));
  OAI21_X1   g14092(.A1(new_n17154_), .A2(new_n17155_), .B(new_n17042_), .ZN(new_n17156_));
  NOR2_X1    g14093(.A1(new_n17002_), .A2(new_n3098_), .ZN(new_n17157_));
  INV_X1     g14094(.I(new_n17157_), .ZN(new_n17158_));
  NAND2_X1   g14095(.A1(new_n17003_), .A2(new_n3098_), .ZN(new_n17159_));
  OAI21_X1   g14096(.A1(new_n17159_), .A2(pi0755), .B(new_n16968_), .ZN(new_n17160_));
  NOR3_X1    g14097(.A1(new_n17158_), .A2(new_n7475_), .A3(new_n17160_), .ZN(new_n17161_));
  NOR3_X1    g14098(.A1(new_n17157_), .A2(pi0149), .A3(new_n17160_), .ZN(new_n17162_));
  OAI21_X1   g14099(.A1(new_n17161_), .A2(new_n17162_), .B(new_n17107_), .ZN(new_n17163_));
  NAND3_X1   g14100(.A1(new_n17156_), .A2(new_n3262_), .A3(new_n17163_), .ZN(new_n17164_));
  NAND2_X1   g14101(.A1(new_n17164_), .A2(new_n17152_), .ZN(new_n17165_));
  AOI21_X1   g14102(.A1(new_n17165_), .A2(new_n16970_), .B(new_n17148_), .ZN(new_n17166_));
  INV_X1     g14103(.I(new_n17095_), .ZN(new_n17167_));
  NAND4_X1   g14104(.A1(new_n17076_), .A2(new_n7475_), .A3(new_n3098_), .A4(new_n17167_), .ZN(new_n17168_));
  NAND2_X1   g14105(.A1(new_n3183_), .A2(new_n7475_), .ZN(new_n17169_));
  AOI21_X1   g14106(.A1(new_n14366_), .A2(new_n17169_), .B(pi0755), .ZN(new_n17170_));
  OAI21_X1   g14107(.A1(pi0149), .A2(new_n16971_), .B(new_n17087_), .ZN(new_n17171_));
  AOI21_X1   g14108(.A1(new_n17168_), .A2(new_n17170_), .B(new_n17171_), .ZN(new_n17172_));
  NOR2_X1    g14109(.A1(new_n13624_), .A2(new_n7475_), .ZN(new_n17173_));
  OAI21_X1   g14110(.A1(new_n13109_), .A2(new_n17149_), .B(pi0038), .ZN(new_n17174_));
  OAI21_X1   g14111(.A1(new_n17173_), .A2(new_n17174_), .B(new_n3259_), .ZN(new_n17175_));
  AOI21_X1   g14112(.A1(new_n12794_), .A2(new_n5453_), .B(pi0039), .ZN(new_n17176_));
  NOR3_X1    g14113(.A1(new_n17176_), .A2(new_n17153_), .A3(new_n5800_), .ZN(new_n17177_));
  NOR2_X1    g14114(.A1(new_n17177_), .A2(pi0038), .ZN(new_n17178_));
  NAND2_X1   g14115(.A1(pi0149), .A2(pi0725), .ZN(new_n17179_));
  NOR4_X1    g14116(.A1(new_n17152_), .A2(new_n13109_), .A3(new_n17178_), .A4(new_n17179_), .ZN(new_n17180_));
  OAI21_X1   g14117(.A1(new_n17172_), .A2(new_n17175_), .B(new_n17180_), .ZN(new_n17181_));
  OAI21_X1   g14118(.A1(new_n17166_), .A2(new_n17181_), .B(new_n8297_), .ZN(new_n17182_));
  AOI21_X1   g14119(.A1(new_n17166_), .A2(new_n17181_), .B(new_n17182_), .ZN(new_n17183_));
  NOR2_X1    g14120(.A1(new_n8345_), .A2(new_n14799_), .ZN(new_n17184_));
  XOR2_X1    g14121(.A1(new_n17183_), .A2(new_n17184_), .Z(new_n17185_));
  AOI21_X1   g14122(.A1(new_n17148_), .A2(new_n16968_), .B(new_n17149_), .ZN(new_n17186_));
  NOR2_X1    g14123(.A1(new_n17186_), .A2(new_n14799_), .ZN(new_n17187_));
  XOR2_X1    g14124(.A1(new_n17187_), .A2(new_n16913_), .Z(new_n17188_));
  OAI21_X1   g14125(.A1(new_n17185_), .A2(new_n17188_), .B(pi0149), .ZN(po0306));
  NOR2_X1    g14126(.A1(pi0150), .A2(pi0751), .ZN(new_n17190_));
  NAND3_X1   g14127(.A1(new_n17066_), .A2(pi0751), .A3(new_n14874_), .ZN(new_n17191_));
  INV_X1     g14128(.I(pi0751), .ZN(new_n17192_));
  NAND3_X1   g14129(.A1(new_n17066_), .A2(new_n17192_), .A3(new_n14298_), .ZN(new_n17193_));
  NAND2_X1   g14130(.A1(new_n17191_), .A2(new_n17193_), .ZN(new_n17194_));
  AOI21_X1   g14131(.A1(new_n17194_), .A2(pi0150), .B(pi0038), .ZN(new_n17195_));
  NOR4_X1    g14132(.A1(new_n17195_), .A2(new_n3183_), .A3(new_n17127_), .A4(new_n17190_), .ZN(new_n17196_));
  NOR2_X1    g14133(.A1(new_n5800_), .A2(pi0751), .ZN(new_n17197_));
  OAI21_X1   g14134(.A1(new_n13109_), .A2(new_n17197_), .B(pi0038), .ZN(new_n17198_));
  AOI21_X1   g14135(.A1(new_n13625_), .A2(pi0150), .B(new_n17198_), .ZN(new_n17199_));
  OAI21_X1   g14136(.A1(new_n17196_), .A2(pi0701), .B(new_n17199_), .ZN(new_n17200_));
  NAND2_X1   g14137(.A1(pi0751), .A2(pi0947), .ZN(new_n17201_));
  OAI21_X1   g14138(.A1(new_n17176_), .A2(new_n17201_), .B(new_n3259_), .ZN(new_n17202_));
  NOR2_X1    g14139(.A1(new_n13109_), .A2(new_n10629_), .ZN(new_n17203_));
  AOI21_X1   g14140(.A1(new_n17203_), .A2(new_n17202_), .B(pi0701), .ZN(new_n17204_));
  NAND2_X1   g14141(.A1(new_n17200_), .A2(new_n17204_), .ZN(new_n17205_));
  NOR2_X1    g14142(.A1(new_n10629_), .A2(new_n17192_), .ZN(new_n17206_));
  NOR2_X1    g14143(.A1(new_n17057_), .A2(new_n10629_), .ZN(new_n17207_));
  XNOR2_X1   g14144(.A1(new_n17207_), .A2(new_n17206_), .ZN(new_n17208_));
  NAND2_X1   g14145(.A1(new_n17009_), .A2(pi0751), .ZN(new_n17209_));
  XOR2_X1    g14146(.A1(new_n17209_), .A2(new_n17206_), .Z(new_n17210_));
  OAI22_X1   g14147(.A1(new_n17210_), .A2(new_n16983_), .B1(new_n17041_), .B2(new_n17208_), .ZN(new_n17211_));
  NAND2_X1   g14148(.A1(new_n17211_), .A2(pi0039), .ZN(new_n17212_));
  NAND3_X1   g14149(.A1(new_n14874_), .A2(pi0751), .A3(pi0947), .ZN(new_n17213_));
  NAND3_X1   g14150(.A1(new_n14874_), .A2(new_n17192_), .A3(new_n5800_), .ZN(new_n17214_));
  AOI21_X1   g14151(.A1(new_n17213_), .A2(new_n17214_), .B(new_n5741_), .ZN(new_n17215_));
  NOR2_X1    g14152(.A1(new_n14298_), .A2(new_n10629_), .ZN(new_n17216_));
  OAI21_X1   g14153(.A1(new_n17215_), .A2(pi0039), .B(new_n17216_), .ZN(new_n17217_));
  NAND4_X1   g14154(.A1(new_n17212_), .A2(new_n3259_), .A3(new_n17205_), .A4(new_n17217_), .ZN(new_n17218_));
  NAND2_X1   g14155(.A1(new_n17218_), .A2(new_n8297_), .ZN(new_n17219_));
  XNOR2_X1   g14156(.A1(new_n17219_), .A2(new_n17184_), .ZN(new_n17220_));
  NOR2_X1    g14157(.A1(new_n5800_), .A2(pi0701), .ZN(new_n17221_));
  OAI21_X1   g14158(.A1(new_n5741_), .A2(new_n17201_), .B(new_n17221_), .ZN(new_n17222_));
  NAND4_X1   g14159(.A1(pi0701), .A2(pi0751), .A3(pi0907), .A4(pi0947), .ZN(new_n17223_));
  NAND3_X1   g14160(.A1(new_n17222_), .A2(pi0832), .A3(new_n17223_), .ZN(new_n17224_));
  XOR2_X1    g14161(.A1(new_n17224_), .A2(new_n16961_), .Z(new_n17225_));
  OAI21_X1   g14162(.A1(new_n17220_), .A2(new_n17225_), .B(pi0150), .ZN(po0307));
  INV_X1     g14163(.I(pi0723), .ZN(new_n17227_));
  NOR2_X1    g14164(.A1(new_n14298_), .A2(pi0745), .ZN(new_n17228_));
  NOR3_X1    g14165(.A1(new_n14298_), .A2(new_n3538_), .A3(new_n5800_), .ZN(new_n17229_));
  XNOR2_X1   g14166(.A1(new_n17229_), .A2(new_n17228_), .ZN(new_n17230_));
  AOI21_X1   g14167(.A1(new_n14365_), .A2(pi0151), .B(pi0745), .ZN(new_n17231_));
  NAND2_X1   g14168(.A1(new_n13081_), .A2(new_n3538_), .ZN(new_n17232_));
  OAI21_X1   g14169(.A1(new_n16977_), .A2(new_n17232_), .B(new_n13080_), .ZN(new_n17233_));
  NOR2_X1    g14170(.A1(new_n16977_), .A2(new_n3111_), .ZN(new_n17234_));
  NAND2_X1   g14171(.A1(new_n17233_), .A2(new_n17234_), .ZN(new_n17235_));
  NAND2_X1   g14172(.A1(new_n17235_), .A2(new_n3098_), .ZN(new_n17236_));
  NOR2_X1    g14173(.A1(new_n16991_), .A2(new_n3313_), .ZN(new_n17237_));
  INV_X1     g14174(.I(new_n17237_), .ZN(new_n17238_));
  AOI21_X1   g14175(.A1(new_n17238_), .A2(new_n3538_), .B(new_n12831_), .ZN(new_n17239_));
  AOI21_X1   g14176(.A1(new_n17239_), .A2(new_n17089_), .B(pi0151), .ZN(new_n17240_));
  NOR3_X1    g14177(.A1(new_n17240_), .A2(new_n12809_), .A3(new_n17070_), .ZN(new_n17241_));
  AOI21_X1   g14178(.A1(new_n17241_), .A2(new_n17236_), .B(pi0745), .ZN(new_n17242_));
  OAI21_X1   g14179(.A1(new_n13085_), .A2(new_n17231_), .B(new_n17242_), .ZN(new_n17243_));
  AOI21_X1   g14180(.A1(new_n17243_), .A2(new_n17087_), .B(new_n3183_), .ZN(new_n17244_));
  XOR2_X1    g14181(.A1(new_n17244_), .A2(new_n4368_), .Z(new_n17245_));
  OAI21_X1   g14182(.A1(new_n17245_), .A2(new_n17230_), .B(new_n17227_), .ZN(new_n17246_));
  NAND2_X1   g14183(.A1(new_n13625_), .A2(pi0151), .ZN(new_n17247_));
  OAI21_X1   g14184(.A1(pi0745), .A2(new_n5800_), .B(new_n13108_), .ZN(new_n17248_));
  NAND4_X1   g14185(.A1(new_n17246_), .A2(pi0038), .A3(new_n17247_), .A4(new_n17248_), .ZN(new_n17249_));
  NAND2_X1   g14186(.A1(pi0745), .A2(pi0947), .ZN(new_n17250_));
  OAI21_X1   g14187(.A1(new_n17176_), .A2(new_n17250_), .B(new_n3259_), .ZN(new_n17251_));
  NOR2_X1    g14188(.A1(new_n13109_), .A2(new_n3538_), .ZN(new_n17252_));
  AOI21_X1   g14189(.A1(new_n17252_), .A2(new_n17251_), .B(pi0723), .ZN(new_n17253_));
  NAND2_X1   g14190(.A1(new_n17249_), .A2(new_n17253_), .ZN(new_n17254_));
  NOR2_X1    g14191(.A1(new_n16970_), .A2(pi0039), .ZN(new_n17255_));
  INV_X1     g14192(.I(new_n17255_), .ZN(new_n17256_));
  INV_X1     g14193(.I(new_n16979_), .ZN(new_n17257_));
  AOI21_X1   g14194(.A1(new_n3538_), .A2(new_n12809_), .B(new_n17257_), .ZN(new_n17258_));
  AOI21_X1   g14195(.A1(new_n17258_), .A2(new_n17038_), .B(new_n3111_), .ZN(new_n17259_));
  INV_X1     g14196(.I(new_n17239_), .ZN(new_n17260_));
  NOR3_X1    g14197(.A1(new_n17260_), .A2(new_n3111_), .A3(new_n17233_), .ZN(new_n17261_));
  XNOR2_X1   g14198(.A1(new_n17261_), .A2(new_n17259_), .ZN(new_n17262_));
  INV_X1     g14199(.I(new_n17036_), .ZN(new_n17263_));
  NAND2_X1   g14200(.A1(new_n17263_), .A2(pi0151), .ZN(new_n17264_));
  NAND3_X1   g14201(.A1(new_n17264_), .A2(pi0745), .A3(new_n17055_), .ZN(new_n17265_));
  AOI21_X1   g14202(.A1(new_n3098_), .A2(new_n17265_), .B(new_n17262_), .ZN(new_n17266_));
  AOI21_X1   g14203(.A1(new_n16972_), .A2(pi0745), .B(pi0151), .ZN(new_n17267_));
  INV_X1     g14204(.I(new_n17001_), .ZN(new_n17268_));
  NAND3_X1   g14205(.A1(new_n16994_), .A2(pi0215), .A3(new_n17258_), .ZN(new_n17269_));
  OAI22_X1   g14206(.A1(new_n17269_), .A2(new_n17260_), .B1(new_n3098_), .B2(new_n17268_), .ZN(new_n17270_));
  NOR2_X1    g14207(.A1(new_n3259_), .A2(new_n3111_), .ZN(new_n17271_));
  NAND4_X1   g14208(.A1(new_n17270_), .A2(new_n16971_), .A3(new_n17233_), .A4(new_n17271_), .ZN(new_n17272_));
  NOR2_X1    g14209(.A1(new_n17272_), .A2(new_n17267_), .ZN(new_n17273_));
  OAI21_X1   g14210(.A1(new_n17266_), .A2(pi0039), .B(new_n17273_), .ZN(new_n17274_));
  AOI21_X1   g14211(.A1(new_n17274_), .A2(new_n17230_), .B(new_n17256_), .ZN(new_n17275_));
  AOI21_X1   g14212(.A1(new_n17254_), .A2(new_n17275_), .B(new_n8345_), .ZN(new_n17276_));
  XOR2_X1    g14213(.A1(new_n17276_), .A2(new_n17184_), .Z(new_n17277_));
  NOR2_X1    g14214(.A1(new_n5800_), .A2(pi0723), .ZN(new_n17278_));
  OAI21_X1   g14215(.A1(new_n5741_), .A2(new_n17250_), .B(new_n17278_), .ZN(new_n17279_));
  NAND4_X1   g14216(.A1(pi0723), .A2(pi0745), .A3(pi0907), .A4(pi0947), .ZN(new_n17280_));
  NAND3_X1   g14217(.A1(new_n17279_), .A2(pi0832), .A3(new_n17280_), .ZN(new_n17281_));
  XOR2_X1    g14218(.A1(new_n17281_), .A2(new_n16961_), .Z(new_n17282_));
  OAI21_X1   g14219(.A1(new_n17277_), .A2(new_n17282_), .B(pi0151), .ZN(po0308));
  INV_X1     g14220(.I(new_n16975_), .ZN(new_n17284_));
  AOI21_X1   g14221(.A1(new_n16993_), .A2(pi0152), .B(new_n17284_), .ZN(new_n17285_));
  NOR2_X1    g14222(.A1(new_n12784_), .A2(new_n5158_), .ZN(new_n17286_));
  NAND2_X1   g14223(.A1(new_n17038_), .A2(new_n13446_), .ZN(new_n17287_));
  NAND2_X1   g14224(.A1(new_n17287_), .A2(new_n17286_), .ZN(new_n17288_));
  NOR3_X1    g14225(.A1(new_n17285_), .A2(new_n16997_), .A3(new_n17288_), .ZN(new_n17289_));
  NOR3_X1    g14226(.A1(new_n17289_), .A2(pi0299), .A3(pi0759), .ZN(new_n17290_));
  AOI21_X1   g14227(.A1(new_n5158_), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n17291_));
  NAND2_X1   g14228(.A1(new_n17034_), .A2(new_n16969_), .ZN(new_n17292_));
  NAND2_X1   g14229(.A1(new_n17291_), .A2(new_n17292_), .ZN(new_n17293_));
  INV_X1     g14230(.I(new_n17053_), .ZN(new_n17294_));
  AOI21_X1   g14231(.A1(new_n5158_), .A2(new_n17045_), .B(new_n17294_), .ZN(new_n17295_));
  NOR2_X1    g14232(.A1(new_n17295_), .A2(pi0299), .ZN(new_n17296_));
  OAI21_X1   g14233(.A1(new_n17290_), .A2(new_n17293_), .B(new_n17296_), .ZN(new_n17297_));
  OAI21_X1   g14234(.A1(new_n5398_), .A2(new_n13086_), .B(new_n16940_), .ZN(new_n17298_));
  NAND3_X1   g14235(.A1(new_n17298_), .A2(new_n3091_), .A3(new_n16968_), .ZN(new_n17299_));
  NAND3_X1   g14236(.A1(new_n17298_), .A2(new_n3092_), .A3(new_n16969_), .ZN(new_n17300_));
  NAND2_X1   g14237(.A1(new_n17299_), .A2(new_n17300_), .ZN(new_n17301_));
  NAND3_X1   g14238(.A1(new_n17301_), .A2(pi0152), .A3(pi0223), .ZN(new_n17302_));
  OR2_X2     g14239(.A1(new_n16978_), .A2(new_n17286_), .Z(new_n17303_));
  AOI21_X1   g14240(.A1(new_n17302_), .A2(new_n3092_), .B(new_n17303_), .ZN(new_n17304_));
  AOI21_X1   g14241(.A1(new_n17297_), .A2(new_n17304_), .B(pi0039), .ZN(new_n17305_));
  NOR2_X1    g14242(.A1(new_n17048_), .A2(new_n3098_), .ZN(new_n17306_));
  INV_X1     g14243(.I(new_n17306_), .ZN(new_n17307_));
  AOI21_X1   g14244(.A1(new_n17307_), .A2(new_n5158_), .B(new_n17045_), .ZN(new_n17308_));
  INV_X1     g14245(.I(pi0759), .ZN(new_n17309_));
  NAND3_X1   g14246(.A1(new_n17298_), .A2(pi0947), .A3(new_n3091_), .ZN(new_n17310_));
  NAND3_X1   g14247(.A1(new_n17298_), .A2(new_n5800_), .A3(new_n3092_), .ZN(new_n17311_));
  NAND2_X1   g14248(.A1(new_n17310_), .A2(new_n17311_), .ZN(new_n17312_));
  NAND2_X1   g14249(.A1(new_n17312_), .A2(pi0152), .ZN(new_n17313_));
  NAND2_X1   g14250(.A1(new_n17038_), .A2(new_n3091_), .ZN(new_n17314_));
  OAI21_X1   g14251(.A1(new_n17314_), .A2(new_n17286_), .B(new_n3090_), .ZN(new_n17315_));
  AOI21_X1   g14252(.A1(new_n17298_), .A2(new_n5453_), .B(new_n3091_), .ZN(new_n17316_));
  NAND2_X1   g14253(.A1(new_n17316_), .A2(new_n17315_), .ZN(new_n17317_));
  OAI21_X1   g14254(.A1(new_n17313_), .A2(new_n17317_), .B(new_n17309_), .ZN(new_n17318_));
  INV_X1     g14255(.I(new_n17295_), .ZN(new_n17319_));
  AOI21_X1   g14256(.A1(new_n17285_), .A2(new_n12831_), .B(new_n17288_), .ZN(new_n17320_));
  NOR4_X1    g14257(.A1(new_n17320_), .A2(new_n17319_), .A3(new_n3098_), .A4(new_n17291_), .ZN(new_n17321_));
  OAI21_X1   g14258(.A1(new_n17318_), .A2(new_n17308_), .B(new_n17321_), .ZN(new_n17322_));
  OAI21_X1   g14259(.A1(new_n17305_), .A2(new_n17322_), .B(new_n3259_), .ZN(new_n17323_));
  NOR2_X1    g14260(.A1(new_n17309_), .A2(new_n5800_), .ZN(new_n17324_));
  NOR2_X1    g14261(.A1(new_n14298_), .A2(new_n17324_), .ZN(new_n17325_));
  XOR2_X1    g14262(.A1(new_n17325_), .A2(new_n13094_), .Z(new_n17326_));
  INV_X1     g14263(.I(pi0696), .ZN(new_n17327_));
  AND4_X2    g14264(.A1(pi0152), .A2(new_n17326_), .A3(new_n13624_), .A4(new_n16970_), .Z(new_n17330_));
  AND2_X2    g14265(.A1(new_n17285_), .A2(new_n12974_), .Z(new_n17331_));
  OAI21_X1   g14266(.A1(new_n17069_), .A2(new_n5800_), .B(new_n3111_), .ZN(new_n17332_));
  NOR3_X1    g14267(.A1(new_n17088_), .A2(new_n17286_), .A3(new_n3313_), .ZN(new_n17333_));
  OAI21_X1   g14268(.A1(new_n17331_), .A2(new_n17332_), .B(new_n17333_), .ZN(new_n17334_));
  NAND2_X1   g14269(.A1(new_n17334_), .A2(new_n17094_), .ZN(new_n17335_));
  INV_X1     g14270(.I(new_n17074_), .ZN(new_n17336_));
  NOR2_X1    g14271(.A1(new_n17336_), .A2(new_n5158_), .ZN(new_n17337_));
  AOI21_X1   g14272(.A1(new_n17335_), .A2(new_n17337_), .B(pi0759), .ZN(new_n17338_));
  OAI21_X1   g14273(.A1(new_n17313_), .A2(new_n3090_), .B(new_n3092_), .ZN(new_n17339_));
  AOI21_X1   g14274(.A1(new_n17326_), .A2(pi0152), .B(pi0038), .ZN(new_n17340_));
  OAI21_X1   g14275(.A1(new_n14291_), .A2(new_n16968_), .B(new_n3211_), .ZN(new_n17341_));
  NAND3_X1   g14276(.A1(new_n17341_), .A2(pi0696), .A3(new_n17324_), .ZN(new_n17342_));
  NAND2_X1   g14277(.A1(new_n17342_), .A2(new_n5158_), .ZN(new_n17343_));
  NAND3_X1   g14278(.A1(new_n3183_), .A2(new_n5158_), .A3(new_n17309_), .ZN(new_n17344_));
  NAND3_X1   g14279(.A1(new_n17343_), .A2(new_n13108_), .A3(new_n17344_), .ZN(new_n17345_));
  NOR4_X1    g14280(.A1(new_n17340_), .A2(new_n17088_), .A3(new_n17286_), .A4(new_n17345_), .ZN(new_n17346_));
  NAND4_X1   g14281(.A1(new_n17346_), .A2(new_n17339_), .A3(new_n14366_), .A4(new_n17308_), .ZN(new_n17347_));
  OAI21_X1   g14282(.A1(new_n17338_), .A2(new_n17347_), .B(new_n8297_), .ZN(new_n17348_));
  AOI21_X1   g14283(.A1(new_n17323_), .A2(new_n17330_), .B(new_n17348_), .ZN(new_n17349_));
  XNOR2_X1   g14284(.A1(new_n17349_), .A2(new_n17184_), .ZN(new_n17350_));
  NOR2_X1    g14285(.A1(new_n17324_), .A2(new_n9992_), .ZN(new_n17351_));
  NOR3_X1    g14286(.A1(new_n17351_), .A2(new_n17327_), .A3(new_n16969_), .ZN(new_n17352_));
  OAI21_X1   g14287(.A1(new_n9992_), .A2(pi0152), .B(pi0832), .ZN(new_n17353_));
  OAI22_X1   g14288(.A1(new_n17350_), .A2(new_n5158_), .B1(new_n17352_), .B2(new_n17353_), .ZN(po0309));
  INV_X1     g14289(.I(pi0766), .ZN(new_n17355_));
  NAND2_X1   g14290(.A1(new_n14299_), .A2(new_n17355_), .ZN(new_n17356_));
  AOI22_X1   g14291(.A1(new_n17086_), .A2(new_n17356_), .B1(new_n2837_), .B2(new_n14298_), .ZN(new_n17357_));
  NOR3_X1    g14292(.A1(new_n16993_), .A2(new_n3312_), .A3(new_n17257_), .ZN(new_n17358_));
  NOR2_X1    g14293(.A1(new_n17358_), .A2(pi0153), .ZN(new_n17359_));
  AOI21_X1   g14294(.A1(pi0153), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n17360_));
  NOR2_X1    g14295(.A1(new_n17360_), .A2(new_n17034_), .ZN(new_n17361_));
  NAND2_X1   g14296(.A1(new_n17268_), .A2(pi0215), .ZN(new_n17362_));
  OAI22_X1   g14297(.A1(new_n17359_), .A2(new_n12809_), .B1(new_n17361_), .B2(new_n17362_), .ZN(new_n17363_));
  NOR2_X1    g14298(.A1(new_n16971_), .A2(pi0153), .ZN(new_n17364_));
  OAI21_X1   g14299(.A1(new_n16973_), .A2(new_n17364_), .B(new_n17355_), .ZN(new_n17365_));
  AOI21_X1   g14300(.A1(new_n17238_), .A2(new_n2837_), .B(new_n12831_), .ZN(new_n17366_));
  NAND4_X1   g14301(.A1(new_n17363_), .A2(pi0299), .A3(new_n17365_), .A4(new_n17366_), .ZN(new_n17367_));
  INV_X1     g14302(.I(new_n17055_), .ZN(new_n17368_));
  INV_X1     g14303(.I(new_n17366_), .ZN(new_n17369_));
  INV_X1     g14304(.I(new_n17089_), .ZN(new_n17370_));
  AOI21_X1   g14305(.A1(new_n2837_), .A2(new_n12809_), .B(new_n17370_), .ZN(new_n17371_));
  NAND2_X1   g14306(.A1(new_n17371_), .A2(pi0215), .ZN(new_n17372_));
  NAND2_X1   g14307(.A1(new_n17372_), .A2(new_n5741_), .ZN(new_n17373_));
  AOI22_X1   g14308(.A1(new_n17360_), .A2(pi0299), .B1(new_n12784_), .B2(new_n17373_), .ZN(new_n17374_));
  NOR3_X1    g14309(.A1(new_n17368_), .A2(new_n17369_), .A3(new_n17374_), .ZN(new_n17375_));
  NOR3_X1    g14310(.A1(new_n17263_), .A2(new_n3259_), .A3(new_n17355_), .ZN(new_n17376_));
  OAI21_X1   g14311(.A1(new_n17375_), .A2(pi0153), .B(new_n17376_), .ZN(new_n17377_));
  AOI21_X1   g14312(.A1(new_n3183_), .A2(new_n17367_), .B(new_n17377_), .ZN(new_n17378_));
  OAI21_X1   g14313(.A1(new_n17378_), .A2(new_n17357_), .B(new_n16970_), .ZN(new_n17379_));
  NOR2_X1    g14314(.A1(new_n17336_), .A2(new_n3098_), .ZN(new_n17380_));
  NOR2_X1    g14315(.A1(new_n13081_), .A2(new_n17355_), .ZN(new_n17381_));
  OAI21_X1   g14316(.A1(new_n17380_), .A2(pi0153), .B(new_n17381_), .ZN(new_n17382_));
  NAND2_X1   g14317(.A1(new_n17382_), .A2(new_n17070_), .ZN(new_n17383_));
  INV_X1     g14318(.I(new_n17087_), .ZN(new_n17384_));
  NOR3_X1    g14319(.A1(new_n17369_), .A2(new_n17384_), .A3(new_n17371_), .ZN(new_n17385_));
  AOI21_X1   g14320(.A1(new_n17383_), .A2(new_n17385_), .B(pi0153), .ZN(new_n17386_));
  NAND2_X1   g14321(.A1(new_n3183_), .A2(new_n2837_), .ZN(new_n17387_));
  OAI22_X1   g14322(.A1(new_n17357_), .A2(pi0038), .B1(pi0766), .B2(new_n17387_), .ZN(new_n17388_));
  OR3_X2     g14323(.A1(new_n17388_), .A2(new_n17127_), .A3(new_n17003_), .Z(new_n17389_));
  NOR2_X1    g14324(.A1(new_n17123_), .A2(pi0700), .ZN(new_n17390_));
  OAI21_X1   g14325(.A1(new_n17386_), .A2(new_n17389_), .B(new_n17390_), .ZN(new_n17391_));
  INV_X1     g14326(.I(pi0700), .ZN(new_n17392_));
  AOI21_X1   g14327(.A1(pi0766), .A2(pi0947), .B(new_n2723_), .ZN(new_n17393_));
  AOI21_X1   g14328(.A1(new_n5503_), .A2(new_n17393_), .B(pi0038), .ZN(new_n17394_));
  NOR4_X1    g14329(.A1(new_n13625_), .A2(new_n2837_), .A3(new_n17392_), .A4(new_n17394_), .ZN(new_n17395_));
  NAND2_X1   g14330(.A1(new_n17391_), .A2(new_n17395_), .ZN(new_n17396_));
  NOR3_X1    g14331(.A1(new_n17176_), .A2(new_n17355_), .A3(new_n5800_), .ZN(new_n17397_));
  NOR2_X1    g14332(.A1(new_n16969_), .A2(pi0832), .ZN(new_n17401_));
  NAND2_X1   g14333(.A1(new_n5371_), .A2(pi0153), .ZN(new_n17402_));
  NOR2_X1    g14334(.A1(new_n13109_), .A2(new_n17402_), .ZN(new_n17403_));
  OAI21_X1   g14335(.A1(new_n17397_), .A2(pi0038), .B(new_n17403_), .ZN(new_n17404_));
  AOI21_X1   g14336(.A1(new_n17379_), .A2(new_n17396_), .B(new_n17404_), .ZN(po0310));
  NAND2_X1   g14337(.A1(new_n17078_), .A2(pi0039), .ZN(new_n17406_));
  XOR2_X1    g14338(.A1(new_n17406_), .A2(new_n3404_), .Z(new_n17407_));
  NAND3_X1   g14339(.A1(new_n17407_), .A2(new_n17085_), .A3(new_n17096_), .ZN(new_n17408_));
  INV_X1     g14340(.I(pi0742), .ZN(new_n17409_));
  OAI21_X1   g14341(.A1(pi0154), .A2(new_n13624_), .B(new_n17084_), .ZN(new_n17410_));
  AOI21_X1   g14342(.A1(new_n17410_), .A2(new_n17409_), .B(new_n3259_), .ZN(new_n17411_));
  NAND2_X1   g14343(.A1(new_n14874_), .A2(new_n17411_), .ZN(new_n17412_));
  AOI21_X1   g14344(.A1(new_n17408_), .A2(new_n3336_), .B(new_n17412_), .ZN(new_n17413_));
  INV_X1     g14345(.I(pi0704), .ZN(new_n17414_));
  NAND2_X1   g14346(.A1(new_n17414_), .A2(new_n17409_), .ZN(new_n17415_));
  OAI21_X1   g14347(.A1(new_n13634_), .A2(new_n17415_), .B(pi0154), .ZN(new_n17416_));
  OAI21_X1   g14348(.A1(new_n17413_), .A2(new_n17416_), .B(new_n8297_), .ZN(new_n17417_));
  NAND2_X1   g14349(.A1(pi0742), .A2(pi0907), .ZN(new_n17418_));
  NAND3_X1   g14350(.A1(new_n17418_), .A2(new_n17414_), .A3(pi0947), .ZN(new_n17419_));
  NAND4_X1   g14351(.A1(pi0704), .A2(pi0742), .A3(pi0907), .A4(pi0947), .ZN(new_n17420_));
  NAND3_X1   g14352(.A1(new_n17419_), .A2(pi0832), .A3(new_n17420_), .ZN(new_n17421_));
  XOR2_X1    g14353(.A1(new_n17421_), .A2(new_n16961_), .Z(new_n17422_));
  NOR2_X1    g14354(.A1(new_n3336_), .A2(pi0832), .ZN(new_n17423_));
  NAND2_X1   g14355(.A1(new_n17422_), .A2(new_n17423_), .ZN(new_n17424_));
  OAI21_X1   g14356(.A1(pi0154), .A2(new_n14874_), .B(new_n17255_), .ZN(new_n17425_));
  INV_X1     g14357(.I(new_n16983_), .ZN(new_n17426_));
  NAND2_X1   g14358(.A1(new_n17009_), .A2(pi0039), .ZN(new_n17427_));
  XOR2_X1    g14359(.A1(new_n17427_), .A2(new_n3404_), .Z(new_n17428_));
  OAI21_X1   g14360(.A1(new_n17022_), .A2(new_n17409_), .B(new_n3336_), .ZN(new_n17429_));
  AOI22_X1   g14361(.A1(new_n17428_), .A2(new_n17426_), .B1(new_n13723_), .B2(new_n17429_), .ZN(new_n17430_));
  OAI21_X1   g14362(.A1(new_n17430_), .A2(new_n17425_), .B(new_n17414_), .ZN(new_n17431_));
  NOR2_X1    g14363(.A1(new_n17057_), .A2(new_n3183_), .ZN(new_n17432_));
  XOR2_X1    g14364(.A1(new_n17432_), .A2(new_n3404_), .Z(new_n17433_));
  NAND2_X1   g14365(.A1(new_n17042_), .A2(pi0038), .ZN(new_n17434_));
  OAI21_X1   g14366(.A1(new_n17433_), .A2(new_n17434_), .B(new_n17425_), .ZN(new_n17435_));
  NAND2_X1   g14367(.A1(new_n17026_), .A2(pi0742), .ZN(new_n17436_));
  AOI21_X1   g14368(.A1(new_n17436_), .A2(new_n3336_), .B(new_n13109_), .ZN(new_n17437_));
  NAND4_X1   g14369(.A1(new_n17431_), .A2(new_n17031_), .A3(new_n17435_), .A4(new_n17437_), .ZN(new_n17438_));
  AOI21_X1   g14370(.A1(new_n17417_), .A2(new_n17424_), .B(new_n17438_), .ZN(po0311));
  INV_X1     g14371(.I(pi0686), .ZN(new_n17440_));
  NAND2_X1   g14372(.A1(pi0757), .A2(pi0907), .ZN(new_n17441_));
  NAND3_X1   g14373(.A1(new_n17441_), .A2(new_n17440_), .A3(pi0947), .ZN(new_n17442_));
  NAND4_X1   g14374(.A1(pi0686), .A2(pi0757), .A3(pi0907), .A4(pi0947), .ZN(new_n17443_));
  NAND3_X1   g14375(.A1(new_n17442_), .A2(pi0832), .A3(new_n17443_), .ZN(new_n17444_));
  XOR2_X1    g14376(.A1(new_n17444_), .A2(new_n16961_), .Z(new_n17445_));
  INV_X1     g14377(.I(pi0757), .ZN(new_n17446_));
  NAND2_X1   g14378(.A1(new_n8297_), .A2(pi0686), .ZN(new_n17447_));
  AOI21_X1   g14379(.A1(new_n17099_), .A2(new_n17447_), .B(new_n17446_), .ZN(new_n17448_));
  NOR2_X1    g14380(.A1(new_n17440_), .A2(new_n17446_), .ZN(new_n17449_));
  NOR2_X1    g14381(.A1(new_n16968_), .A2(new_n3259_), .ZN(new_n17450_));
  OAI21_X1   g14382(.A1(new_n17014_), .A2(new_n17012_), .B(new_n13723_), .ZN(new_n17451_));
  XOR2_X1    g14383(.A1(new_n17451_), .A2(new_n17450_), .Z(new_n17452_));
  NAND2_X1   g14384(.A1(new_n17452_), .A2(pi0757), .ZN(new_n17453_));
  XOR2_X1    g14385(.A1(new_n17453_), .A2(new_n17449_), .Z(new_n17454_));
  NOR2_X1    g14386(.A1(new_n17081_), .A2(new_n17440_), .ZN(new_n17455_));
  XNOR2_X1   g14387(.A1(new_n17455_), .A2(new_n17449_), .ZN(new_n17456_));
  NOR2_X1    g14388(.A1(new_n17060_), .A2(pi0038), .ZN(new_n17457_));
  NOR2_X1    g14389(.A1(new_n17027_), .A2(new_n3259_), .ZN(new_n17458_));
  NOR2_X1    g14390(.A1(new_n17457_), .A2(new_n17458_), .ZN(new_n17459_));
  NAND2_X1   g14391(.A1(new_n8345_), .A2(new_n8020_), .ZN(new_n17460_));
  NAND3_X1   g14392(.A1(new_n13634_), .A2(pi0155), .A3(new_n17460_), .ZN(new_n17461_));
  NOR4_X1    g14393(.A1(new_n17454_), .A2(new_n17456_), .A3(new_n17459_), .A4(new_n17461_), .ZN(new_n17462_));
  AOI21_X1   g14394(.A1(new_n16985_), .A2(new_n3259_), .B(new_n17021_), .ZN(new_n17463_));
  INV_X1     g14395(.I(new_n17463_), .ZN(new_n17464_));
  INV_X1     g14396(.I(new_n17026_), .ZN(new_n17465_));
  OAI21_X1   g14397(.A1(new_n17043_), .A2(pi0038), .B(new_n17465_), .ZN(new_n17466_));
  NAND2_X1   g14398(.A1(new_n17466_), .A2(pi0757), .ZN(new_n17467_));
  XOR2_X1    g14399(.A1(new_n17467_), .A2(new_n17449_), .Z(new_n17468_));
  NOR2_X1    g14400(.A1(new_n17468_), .A2(new_n17464_), .ZN(new_n17469_));
  OAI21_X1   g14401(.A1(new_n17462_), .A2(new_n17448_), .B(new_n17469_), .ZN(new_n17470_));
  AOI22_X1   g14402(.A1(new_n17470_), .A2(new_n14799_), .B1(pi0155), .B2(new_n17445_), .ZN(po0312));
  INV_X1     g14403(.I(new_n17459_), .ZN(new_n17472_));
  NAND2_X1   g14404(.A1(new_n17452_), .A2(pi0741), .ZN(new_n17473_));
  INV_X1     g14405(.I(pi0724), .ZN(new_n17474_));
  INV_X1     g14406(.I(pi0741), .ZN(new_n17475_));
  NOR2_X1    g14407(.A1(new_n17474_), .A2(new_n17475_), .ZN(new_n17476_));
  XNOR2_X1   g14408(.A1(new_n17473_), .A2(new_n17476_), .ZN(new_n17477_));
  NAND2_X1   g14409(.A1(new_n17466_), .A2(pi0741), .ZN(new_n17478_));
  XNOR2_X1   g14410(.A1(new_n17478_), .A2(new_n17476_), .ZN(new_n17479_));
  NAND2_X1   g14411(.A1(new_n17099_), .A2(new_n17474_), .ZN(new_n17480_));
  AOI21_X1   g14412(.A1(new_n17479_), .A2(new_n17463_), .B(new_n17480_), .ZN(new_n17481_));
  NAND2_X1   g14413(.A1(pi0741), .A2(pi0907), .ZN(new_n17482_));
  NAND3_X1   g14414(.A1(new_n17482_), .A2(new_n17474_), .A3(pi0947), .ZN(new_n17483_));
  NAND4_X1   g14415(.A1(pi0724), .A2(pi0741), .A3(pi0907), .A4(pi0947), .ZN(new_n17484_));
  NAND3_X1   g14416(.A1(new_n17483_), .A2(pi0832), .A3(new_n17484_), .ZN(new_n17485_));
  XOR2_X1    g14417(.A1(new_n17485_), .A2(new_n16961_), .Z(new_n17486_));
  NOR2_X1    g14418(.A1(new_n9505_), .A2(new_n17475_), .ZN(new_n17487_));
  NAND2_X1   g14419(.A1(new_n17486_), .A2(new_n17487_), .ZN(new_n17488_));
  OAI21_X1   g14420(.A1(new_n17481_), .A2(new_n17488_), .B(new_n9505_), .ZN(new_n17489_));
  NOR2_X1    g14421(.A1(new_n17081_), .A2(new_n17474_), .ZN(new_n17490_));
  XOR2_X1    g14422(.A1(new_n17490_), .A2(new_n17476_), .Z(new_n17491_));
  NAND2_X1   g14423(.A1(new_n17491_), .A2(new_n13634_), .ZN(new_n17492_));
  NAND3_X1   g14424(.A1(new_n17492_), .A2(new_n8297_), .A3(new_n17489_), .ZN(new_n17493_));
  AOI21_X1   g14425(.A1(new_n17477_), .A2(new_n17472_), .B(new_n17493_), .ZN(po0313));
  INV_X1     g14426(.I(pi0688), .ZN(new_n17495_));
  NOR2_X1    g14427(.A1(new_n5800_), .A2(pi0760), .ZN(new_n17496_));
  NOR2_X1    g14428(.A1(new_n14298_), .A2(new_n17496_), .ZN(new_n17497_));
  XOR2_X1    g14429(.A1(new_n17497_), .A2(new_n13094_), .Z(new_n17498_));
  NAND2_X1   g14430(.A1(new_n17498_), .A2(pi0157), .ZN(new_n17499_));
  INV_X1     g14431(.I(pi0760), .ZN(new_n17500_));
  NOR3_X1    g14432(.A1(new_n17009_), .A2(new_n10692_), .A3(new_n17500_), .ZN(new_n17501_));
  NOR4_X1    g14433(.A1(new_n17008_), .A2(pi0157), .A3(new_n17500_), .A4(new_n17006_), .ZN(new_n17502_));
  OAI21_X1   g14434(.A1(new_n17501_), .A2(new_n17502_), .B(new_n17057_), .ZN(new_n17503_));
  NOR3_X1    g14435(.A1(new_n17041_), .A2(new_n10692_), .A3(new_n17500_), .ZN(new_n17504_));
  NOR3_X1    g14436(.A1(new_n17042_), .A2(new_n10692_), .A3(pi0760), .ZN(new_n17505_));
  OAI21_X1   g14437(.A1(new_n17505_), .A2(new_n17504_), .B(new_n17426_), .ZN(new_n17506_));
  NAND3_X1   g14438(.A1(new_n17503_), .A2(new_n3262_), .A3(new_n17506_), .ZN(new_n17507_));
  NAND2_X1   g14439(.A1(new_n17507_), .A2(new_n17499_), .ZN(new_n17508_));
  AOI21_X1   g14440(.A1(new_n17508_), .A2(new_n16970_), .B(new_n17495_), .ZN(new_n17509_));
  NAND4_X1   g14441(.A1(new_n17076_), .A2(new_n10692_), .A3(new_n3098_), .A4(new_n17167_), .ZN(new_n17510_));
  NAND2_X1   g14442(.A1(new_n3183_), .A2(new_n10692_), .ZN(new_n17511_));
  AOI21_X1   g14443(.A1(new_n14366_), .A2(new_n17511_), .B(pi0760), .ZN(new_n17512_));
  OAI21_X1   g14444(.A1(pi0157), .A2(new_n16971_), .B(new_n17087_), .ZN(new_n17513_));
  AOI21_X1   g14445(.A1(new_n17510_), .A2(new_n17512_), .B(new_n17513_), .ZN(new_n17514_));
  NOR2_X1    g14446(.A1(new_n13624_), .A2(new_n10692_), .ZN(new_n17515_));
  OAI21_X1   g14447(.A1(new_n13109_), .A2(new_n17496_), .B(pi0038), .ZN(new_n17516_));
  OAI21_X1   g14448(.A1(new_n17515_), .A2(new_n17516_), .B(new_n3259_), .ZN(new_n17517_));
  NOR3_X1    g14449(.A1(new_n17176_), .A2(new_n17500_), .A3(new_n5800_), .ZN(new_n17518_));
  NOR2_X1    g14450(.A1(new_n17518_), .A2(pi0038), .ZN(new_n17519_));
  NAND2_X1   g14451(.A1(pi0157), .A2(pi0688), .ZN(new_n17520_));
  NOR4_X1    g14452(.A1(new_n17499_), .A2(new_n13109_), .A3(new_n17519_), .A4(new_n17520_), .ZN(new_n17521_));
  OAI21_X1   g14453(.A1(new_n17514_), .A2(new_n17517_), .B(new_n17521_), .ZN(new_n17522_));
  OAI21_X1   g14454(.A1(new_n17509_), .A2(new_n17522_), .B(new_n8297_), .ZN(new_n17523_));
  AOI21_X1   g14455(.A1(new_n17509_), .A2(new_n17522_), .B(new_n17523_), .ZN(new_n17524_));
  XOR2_X1    g14456(.A1(new_n17524_), .A2(new_n17184_), .Z(new_n17525_));
  AOI21_X1   g14457(.A1(new_n17495_), .A2(new_n16968_), .B(new_n17496_), .ZN(new_n17526_));
  NOR2_X1    g14458(.A1(new_n17526_), .A2(new_n14799_), .ZN(new_n17527_));
  XOR2_X1    g14459(.A1(new_n17527_), .A2(new_n16913_), .Z(new_n17528_));
  OAI21_X1   g14460(.A1(new_n17525_), .A2(new_n17528_), .B(pi0157), .ZN(po0314));
  NOR2_X1    g14461(.A1(pi0158), .A2(pi0753), .ZN(new_n17530_));
  NAND3_X1   g14462(.A1(new_n17066_), .A2(pi0753), .A3(new_n14874_), .ZN(new_n17531_));
  INV_X1     g14463(.I(pi0753), .ZN(new_n17532_));
  NAND3_X1   g14464(.A1(new_n17066_), .A2(new_n17532_), .A3(new_n14298_), .ZN(new_n17533_));
  NAND2_X1   g14465(.A1(new_n17531_), .A2(new_n17533_), .ZN(new_n17534_));
  AOI21_X1   g14466(.A1(new_n17534_), .A2(pi0158), .B(pi0038), .ZN(new_n17535_));
  NOR4_X1    g14467(.A1(new_n17535_), .A2(new_n3183_), .A3(new_n17127_), .A4(new_n17530_), .ZN(new_n17536_));
  NOR2_X1    g14468(.A1(new_n5800_), .A2(pi0753), .ZN(new_n17537_));
  OAI21_X1   g14469(.A1(new_n13109_), .A2(new_n17537_), .B(pi0038), .ZN(new_n17538_));
  AOI21_X1   g14470(.A1(new_n13625_), .A2(pi0158), .B(new_n17538_), .ZN(new_n17539_));
  OAI21_X1   g14471(.A1(new_n17536_), .A2(pi0702), .B(new_n17539_), .ZN(new_n17540_));
  NAND2_X1   g14472(.A1(pi0753), .A2(pi0947), .ZN(new_n17541_));
  OAI21_X1   g14473(.A1(new_n17176_), .A2(new_n17541_), .B(new_n3259_), .ZN(new_n17542_));
  NOR2_X1    g14474(.A1(new_n13109_), .A2(new_n5661_), .ZN(new_n17543_));
  AOI21_X1   g14475(.A1(new_n17543_), .A2(new_n17542_), .B(pi0702), .ZN(new_n17544_));
  NAND2_X1   g14476(.A1(new_n17540_), .A2(new_n17544_), .ZN(new_n17545_));
  NOR2_X1    g14477(.A1(new_n5661_), .A2(new_n17532_), .ZN(new_n17546_));
  NOR2_X1    g14478(.A1(new_n17057_), .A2(new_n5661_), .ZN(new_n17547_));
  XNOR2_X1   g14479(.A1(new_n17547_), .A2(new_n17546_), .ZN(new_n17548_));
  NAND2_X1   g14480(.A1(new_n17009_), .A2(pi0753), .ZN(new_n17549_));
  XOR2_X1    g14481(.A1(new_n17549_), .A2(new_n17546_), .Z(new_n17550_));
  OAI22_X1   g14482(.A1(new_n17550_), .A2(new_n16983_), .B1(new_n17041_), .B2(new_n17548_), .ZN(new_n17551_));
  NAND2_X1   g14483(.A1(new_n17551_), .A2(pi0039), .ZN(new_n17552_));
  NAND3_X1   g14484(.A1(new_n14874_), .A2(pi0753), .A3(pi0947), .ZN(new_n17553_));
  NAND3_X1   g14485(.A1(new_n14874_), .A2(new_n17532_), .A3(new_n5800_), .ZN(new_n17554_));
  AOI21_X1   g14486(.A1(new_n17553_), .A2(new_n17554_), .B(new_n5741_), .ZN(new_n17555_));
  NOR2_X1    g14487(.A1(new_n14298_), .A2(new_n5661_), .ZN(new_n17556_));
  OAI21_X1   g14488(.A1(new_n17555_), .A2(pi0039), .B(new_n17556_), .ZN(new_n17557_));
  NAND4_X1   g14489(.A1(new_n17552_), .A2(new_n3259_), .A3(new_n17545_), .A4(new_n17557_), .ZN(new_n17558_));
  NAND2_X1   g14490(.A1(new_n17558_), .A2(new_n8297_), .ZN(new_n17559_));
  XNOR2_X1   g14491(.A1(new_n17559_), .A2(new_n17184_), .ZN(new_n17560_));
  NOR2_X1    g14492(.A1(new_n5800_), .A2(pi0702), .ZN(new_n17561_));
  OAI21_X1   g14493(.A1(new_n5741_), .A2(new_n17541_), .B(new_n17561_), .ZN(new_n17562_));
  NAND4_X1   g14494(.A1(pi0702), .A2(pi0753), .A3(pi0907), .A4(pi0947), .ZN(new_n17563_));
  NAND3_X1   g14495(.A1(new_n17562_), .A2(pi0832), .A3(new_n17563_), .ZN(new_n17564_));
  XOR2_X1    g14496(.A1(new_n17564_), .A2(new_n16961_), .Z(new_n17565_));
  OAI21_X1   g14497(.A1(new_n17560_), .A2(new_n17565_), .B(pi0158), .ZN(po0315));
  NOR2_X1    g14498(.A1(pi0159), .A2(pi0754), .ZN(new_n17567_));
  NAND3_X1   g14499(.A1(new_n17066_), .A2(pi0754), .A3(new_n14874_), .ZN(new_n17568_));
  INV_X1     g14500(.I(pi0754), .ZN(new_n17569_));
  NAND3_X1   g14501(.A1(new_n17066_), .A2(new_n17569_), .A3(new_n14298_), .ZN(new_n17570_));
  NAND2_X1   g14502(.A1(new_n17568_), .A2(new_n17570_), .ZN(new_n17571_));
  AOI21_X1   g14503(.A1(new_n17571_), .A2(pi0159), .B(pi0038), .ZN(new_n17572_));
  NOR4_X1    g14504(.A1(new_n17572_), .A2(new_n3183_), .A3(new_n17127_), .A4(new_n17567_), .ZN(new_n17573_));
  NOR2_X1    g14505(.A1(new_n5800_), .A2(pi0754), .ZN(new_n17574_));
  OAI21_X1   g14506(.A1(new_n13109_), .A2(new_n17574_), .B(pi0038), .ZN(new_n17575_));
  AOI21_X1   g14507(.A1(new_n13625_), .A2(pi0159), .B(new_n17575_), .ZN(new_n17576_));
  OAI21_X1   g14508(.A1(new_n17573_), .A2(pi0709), .B(new_n17576_), .ZN(new_n17577_));
  NAND2_X1   g14509(.A1(pi0754), .A2(pi0947), .ZN(new_n17578_));
  OAI21_X1   g14510(.A1(new_n17176_), .A2(new_n17578_), .B(new_n3259_), .ZN(new_n17579_));
  NOR2_X1    g14511(.A1(new_n13109_), .A2(new_n5662_), .ZN(new_n17580_));
  AOI21_X1   g14512(.A1(new_n17580_), .A2(new_n17579_), .B(pi0709), .ZN(new_n17581_));
  NAND2_X1   g14513(.A1(new_n17577_), .A2(new_n17581_), .ZN(new_n17582_));
  NOR2_X1    g14514(.A1(new_n5662_), .A2(new_n17569_), .ZN(new_n17583_));
  NOR2_X1    g14515(.A1(new_n17057_), .A2(new_n5662_), .ZN(new_n17584_));
  XNOR2_X1   g14516(.A1(new_n17584_), .A2(new_n17583_), .ZN(new_n17585_));
  NAND2_X1   g14517(.A1(new_n17009_), .A2(pi0754), .ZN(new_n17586_));
  XOR2_X1    g14518(.A1(new_n17586_), .A2(new_n17583_), .Z(new_n17587_));
  OAI22_X1   g14519(.A1(new_n17587_), .A2(new_n16983_), .B1(new_n17041_), .B2(new_n17585_), .ZN(new_n17588_));
  NAND2_X1   g14520(.A1(new_n17588_), .A2(pi0039), .ZN(new_n17589_));
  NAND3_X1   g14521(.A1(new_n14874_), .A2(pi0754), .A3(pi0947), .ZN(new_n17590_));
  NAND3_X1   g14522(.A1(new_n14874_), .A2(new_n17569_), .A3(new_n5800_), .ZN(new_n17591_));
  AOI21_X1   g14523(.A1(new_n17590_), .A2(new_n17591_), .B(new_n5741_), .ZN(new_n17592_));
  NOR2_X1    g14524(.A1(new_n14298_), .A2(new_n5662_), .ZN(new_n17593_));
  OAI21_X1   g14525(.A1(new_n17592_), .A2(pi0039), .B(new_n17593_), .ZN(new_n17594_));
  NAND4_X1   g14526(.A1(new_n17589_), .A2(new_n3259_), .A3(new_n17582_), .A4(new_n17594_), .ZN(new_n17595_));
  NAND2_X1   g14527(.A1(new_n17595_), .A2(new_n8297_), .ZN(new_n17596_));
  XNOR2_X1   g14528(.A1(new_n17596_), .A2(new_n17184_), .ZN(new_n17597_));
  NOR2_X1    g14529(.A1(new_n5800_), .A2(pi0709), .ZN(new_n17598_));
  OAI21_X1   g14530(.A1(new_n5741_), .A2(new_n17578_), .B(new_n17598_), .ZN(new_n17599_));
  NAND4_X1   g14531(.A1(pi0709), .A2(pi0754), .A3(pi0907), .A4(pi0947), .ZN(new_n17600_));
  NAND3_X1   g14532(.A1(new_n17599_), .A2(pi0832), .A3(new_n17600_), .ZN(new_n17601_));
  XOR2_X1    g14533(.A1(new_n17601_), .A2(new_n16961_), .Z(new_n17602_));
  OAI21_X1   g14534(.A1(new_n17597_), .A2(new_n17602_), .B(pi0159), .ZN(po0316));
  INV_X1     g14535(.I(pi0734), .ZN(new_n17604_));
  NOR2_X1    g14536(.A1(new_n5800_), .A2(pi0756), .ZN(new_n17605_));
  NOR2_X1    g14537(.A1(new_n14298_), .A2(new_n17605_), .ZN(new_n17606_));
  XOR2_X1    g14538(.A1(new_n17606_), .A2(new_n13094_), .Z(new_n17607_));
  NAND2_X1   g14539(.A1(new_n17607_), .A2(pi0160), .ZN(new_n17608_));
  INV_X1     g14540(.I(pi0756), .ZN(new_n17609_));
  NOR3_X1    g14541(.A1(new_n17058_), .A2(new_n5664_), .A3(new_n17609_), .ZN(new_n17610_));
  NOR3_X1    g14542(.A1(new_n17057_), .A2(new_n5664_), .A3(pi0756), .ZN(new_n17611_));
  OAI21_X1   g14543(.A1(new_n17610_), .A2(new_n17611_), .B(new_n17042_), .ZN(new_n17612_));
  OAI21_X1   g14544(.A1(new_n17159_), .A2(pi0756), .B(new_n16968_), .ZN(new_n17613_));
  NOR3_X1    g14545(.A1(new_n17158_), .A2(new_n5664_), .A3(new_n17613_), .ZN(new_n17614_));
  NOR3_X1    g14546(.A1(new_n17157_), .A2(pi0160), .A3(new_n17613_), .ZN(new_n17615_));
  OAI21_X1   g14547(.A1(new_n17614_), .A2(new_n17615_), .B(new_n17107_), .ZN(new_n17616_));
  NAND3_X1   g14548(.A1(new_n17612_), .A2(new_n3262_), .A3(new_n17616_), .ZN(new_n17617_));
  NAND2_X1   g14549(.A1(new_n17617_), .A2(new_n17608_), .ZN(new_n17618_));
  AOI21_X1   g14550(.A1(new_n17618_), .A2(new_n16970_), .B(new_n17604_), .ZN(new_n17619_));
  NOR3_X1    g14551(.A1(new_n17125_), .A2(new_n5664_), .A3(new_n3098_), .ZN(new_n17620_));
  NOR3_X1    g14552(.A1(new_n17076_), .A2(pi0160), .A3(new_n3098_), .ZN(new_n17621_));
  OAI21_X1   g14553(.A1(new_n17620_), .A2(new_n17621_), .B(new_n17133_), .ZN(new_n17622_));
  NAND2_X1   g14554(.A1(new_n3183_), .A2(new_n5664_), .ZN(new_n17623_));
  AOI21_X1   g14555(.A1(new_n14366_), .A2(new_n17623_), .B(pi0756), .ZN(new_n17624_));
  OAI21_X1   g14556(.A1(pi0160), .A2(new_n16971_), .B(new_n17087_), .ZN(new_n17625_));
  AOI21_X1   g14557(.A1(new_n17622_), .A2(new_n17624_), .B(new_n17625_), .ZN(new_n17626_));
  NOR2_X1    g14558(.A1(new_n13624_), .A2(new_n5664_), .ZN(new_n17627_));
  OAI21_X1   g14559(.A1(new_n13109_), .A2(new_n17605_), .B(pi0038), .ZN(new_n17628_));
  OAI21_X1   g14560(.A1(new_n17627_), .A2(new_n17628_), .B(new_n3259_), .ZN(new_n17629_));
  NOR3_X1    g14561(.A1(new_n17176_), .A2(new_n17609_), .A3(new_n5800_), .ZN(new_n17630_));
  NOR2_X1    g14562(.A1(new_n17630_), .A2(pi0038), .ZN(new_n17631_));
  NAND2_X1   g14563(.A1(pi0160), .A2(pi0734), .ZN(new_n17632_));
  NOR4_X1    g14564(.A1(new_n17608_), .A2(new_n13109_), .A3(new_n17631_), .A4(new_n17632_), .ZN(new_n17633_));
  OAI21_X1   g14565(.A1(new_n17626_), .A2(new_n17629_), .B(new_n17633_), .ZN(new_n17634_));
  OAI21_X1   g14566(.A1(new_n17619_), .A2(new_n17634_), .B(new_n8297_), .ZN(new_n17635_));
  AOI21_X1   g14567(.A1(new_n17619_), .A2(new_n17634_), .B(new_n17635_), .ZN(new_n17636_));
  XOR2_X1    g14568(.A1(new_n17636_), .A2(new_n17184_), .Z(new_n17637_));
  AOI21_X1   g14569(.A1(new_n17604_), .A2(new_n16968_), .B(new_n17605_), .ZN(new_n17638_));
  NOR2_X1    g14570(.A1(new_n17638_), .A2(new_n14799_), .ZN(new_n17639_));
  XOR2_X1    g14571(.A1(new_n17639_), .A2(new_n16913_), .Z(new_n17640_));
  OAI21_X1   g14572(.A1(new_n17637_), .A2(new_n17640_), .B(pi0160), .ZN(po0317));
  AOI21_X1   g14573(.A1(new_n16993_), .A2(pi0161), .B(new_n17284_), .ZN(new_n17642_));
  NOR2_X1    g14574(.A1(new_n12784_), .A2(new_n4981_), .ZN(new_n17643_));
  NAND2_X1   g14575(.A1(new_n17287_), .A2(new_n17643_), .ZN(new_n17644_));
  NOR3_X1    g14576(.A1(new_n17642_), .A2(new_n16997_), .A3(new_n17644_), .ZN(new_n17645_));
  NOR3_X1    g14577(.A1(new_n17645_), .A2(pi0299), .A3(pi0758), .ZN(new_n17646_));
  AOI21_X1   g14578(.A1(new_n4981_), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n17647_));
  NAND2_X1   g14579(.A1(new_n17647_), .A2(new_n17292_), .ZN(new_n17648_));
  AOI21_X1   g14580(.A1(new_n4981_), .A2(new_n17045_), .B(new_n17294_), .ZN(new_n17649_));
  NOR2_X1    g14581(.A1(new_n17649_), .A2(pi0299), .ZN(new_n17650_));
  OAI21_X1   g14582(.A1(new_n17646_), .A2(new_n17648_), .B(new_n17650_), .ZN(new_n17651_));
  OAI21_X1   g14583(.A1(new_n16978_), .A2(new_n17643_), .B(new_n3091_), .ZN(new_n17652_));
  NAND2_X1   g14584(.A1(new_n17301_), .A2(pi0161), .ZN(new_n17653_));
  AOI21_X1   g14585(.A1(new_n17653_), .A2(new_n17652_), .B(pi0223), .ZN(new_n17654_));
  AOI21_X1   g14586(.A1(new_n17651_), .A2(new_n17654_), .B(pi0039), .ZN(new_n17655_));
  AOI21_X1   g14587(.A1(new_n17307_), .A2(new_n4981_), .B(new_n17045_), .ZN(new_n17656_));
  NAND2_X1   g14588(.A1(new_n17312_), .A2(pi0161), .ZN(new_n17657_));
  OAI21_X1   g14589(.A1(new_n17314_), .A2(new_n17643_), .B(new_n3090_), .ZN(new_n17658_));
  NAND2_X1   g14590(.A1(new_n17316_), .A2(new_n17658_), .ZN(new_n17659_));
  OAI21_X1   g14591(.A1(new_n17657_), .A2(new_n17659_), .B(new_n16090_), .ZN(new_n17660_));
  INV_X1     g14592(.I(new_n17649_), .ZN(new_n17661_));
  AOI21_X1   g14593(.A1(new_n17642_), .A2(new_n12831_), .B(new_n17644_), .ZN(new_n17662_));
  NOR4_X1    g14594(.A1(new_n17662_), .A2(new_n17661_), .A3(new_n3098_), .A4(new_n17647_), .ZN(new_n17663_));
  OAI21_X1   g14595(.A1(new_n17660_), .A2(new_n17656_), .B(new_n17663_), .ZN(new_n17664_));
  OAI21_X1   g14596(.A1(new_n17655_), .A2(new_n17664_), .B(new_n3259_), .ZN(new_n17665_));
  NOR2_X1    g14597(.A1(new_n16090_), .A2(new_n5800_), .ZN(new_n17666_));
  NOR2_X1    g14598(.A1(new_n14298_), .A2(new_n17666_), .ZN(new_n17667_));
  XOR2_X1    g14599(.A1(new_n17667_), .A2(new_n13094_), .Z(new_n17668_));
  AND4_X2    g14600(.A1(pi0161), .A2(new_n17668_), .A3(new_n13624_), .A4(new_n16970_), .Z(new_n17671_));
  AND2_X2    g14601(.A1(new_n17642_), .A2(new_n12974_), .Z(new_n17672_));
  NOR3_X1    g14602(.A1(new_n17088_), .A2(new_n17643_), .A3(new_n3313_), .ZN(new_n17673_));
  OAI21_X1   g14603(.A1(new_n17672_), .A2(new_n17332_), .B(new_n17673_), .ZN(new_n17674_));
  NAND2_X1   g14604(.A1(new_n17674_), .A2(new_n17094_), .ZN(new_n17675_));
  NOR2_X1    g14605(.A1(new_n17336_), .A2(new_n4981_), .ZN(new_n17676_));
  AOI21_X1   g14606(.A1(new_n17675_), .A2(new_n17676_), .B(pi0758), .ZN(new_n17677_));
  OAI21_X1   g14607(.A1(new_n17657_), .A2(new_n3090_), .B(new_n3092_), .ZN(new_n17678_));
  AOI21_X1   g14608(.A1(new_n17668_), .A2(pi0161), .B(pi0038), .ZN(new_n17679_));
  NAND3_X1   g14609(.A1(new_n17341_), .A2(pi0736), .A3(new_n17666_), .ZN(new_n17680_));
  NAND2_X1   g14610(.A1(new_n17680_), .A2(new_n4981_), .ZN(new_n17681_));
  NAND3_X1   g14611(.A1(new_n3183_), .A2(new_n4981_), .A3(new_n16090_), .ZN(new_n17682_));
  NAND3_X1   g14612(.A1(new_n17681_), .A2(new_n13108_), .A3(new_n17682_), .ZN(new_n17683_));
  NOR4_X1    g14613(.A1(new_n17679_), .A2(new_n17088_), .A3(new_n17643_), .A4(new_n17683_), .ZN(new_n17684_));
  NAND4_X1   g14614(.A1(new_n17684_), .A2(new_n17678_), .A3(new_n14366_), .A4(new_n17656_), .ZN(new_n17685_));
  OAI21_X1   g14615(.A1(new_n17677_), .A2(new_n17685_), .B(new_n8297_), .ZN(new_n17686_));
  AOI21_X1   g14616(.A1(new_n17665_), .A2(new_n17671_), .B(new_n17686_), .ZN(new_n17687_));
  XNOR2_X1   g14617(.A1(new_n17687_), .A2(new_n17184_), .ZN(new_n17688_));
  NOR2_X1    g14618(.A1(new_n17666_), .A2(new_n9992_), .ZN(new_n17689_));
  NOR3_X1    g14619(.A1(new_n17689_), .A2(new_n16136_), .A3(new_n16969_), .ZN(new_n17690_));
  OAI21_X1   g14620(.A1(new_n9992_), .A2(pi0161), .B(pi0832), .ZN(new_n17691_));
  OAI22_X1   g14621(.A1(new_n17688_), .A2(new_n4981_), .B1(new_n17690_), .B2(new_n17691_), .ZN(po0318));
  NOR2_X1    g14622(.A1(new_n5800_), .A2(pi0761), .ZN(new_n17693_));
  NOR2_X1    g14623(.A1(new_n14298_), .A2(new_n17693_), .ZN(new_n17694_));
  XOR2_X1    g14624(.A1(new_n17694_), .A2(new_n13094_), .Z(new_n17695_));
  NAND2_X1   g14625(.A1(new_n17695_), .A2(pi0162), .ZN(new_n17696_));
  NOR3_X1    g14626(.A1(new_n17058_), .A2(new_n8108_), .A3(new_n13099_), .ZN(new_n17697_));
  NOR3_X1    g14627(.A1(new_n17057_), .A2(new_n8108_), .A3(pi0761), .ZN(new_n17698_));
  OAI21_X1   g14628(.A1(new_n17697_), .A2(new_n17698_), .B(new_n17042_), .ZN(new_n17699_));
  OAI21_X1   g14629(.A1(new_n17107_), .A2(new_n8108_), .B(pi0761), .ZN(new_n17700_));
  OAI21_X1   g14630(.A1(new_n17009_), .A2(new_n17700_), .B(new_n3098_), .ZN(new_n17701_));
  NAND2_X1   g14631(.A1(new_n17701_), .A2(pi0162), .ZN(new_n17702_));
  NAND3_X1   g14632(.A1(new_n17702_), .A2(new_n3262_), .A3(new_n17699_), .ZN(new_n17703_));
  NAND2_X1   g14633(.A1(new_n17703_), .A2(new_n17696_), .ZN(new_n17704_));
  AOI21_X1   g14634(.A1(new_n17704_), .A2(new_n16970_), .B(new_n13226_), .ZN(new_n17705_));
  NOR2_X1    g14635(.A1(new_n8108_), .A2(new_n13099_), .ZN(new_n17706_));
  NAND2_X1   g14636(.A1(new_n17106_), .A2(pi0761), .ZN(new_n17707_));
  AOI21_X1   g14637(.A1(new_n17076_), .A2(pi0299), .B(new_n17707_), .ZN(new_n17708_));
  XOR2_X1    g14638(.A1(new_n17708_), .A2(new_n17706_), .Z(new_n17709_));
  AOI21_X1   g14639(.A1(new_n17709_), .A2(new_n14366_), .B(pi0039), .ZN(new_n17710_));
  NAND2_X1   g14640(.A1(pi0162), .A2(pi0299), .ZN(new_n17711_));
  OAI21_X1   g14641(.A1(new_n17133_), .A2(new_n17711_), .B(new_n5800_), .ZN(new_n17712_));
  NOR2_X1    g14642(.A1(new_n17712_), .A2(new_n16971_), .ZN(new_n17713_));
  NOR4_X1    g14643(.A1(new_n17710_), .A2(new_n3098_), .A3(new_n13099_), .A4(new_n17713_), .ZN(new_n17714_));
  NOR2_X1    g14644(.A1(new_n13624_), .A2(new_n8108_), .ZN(new_n17715_));
  OAI21_X1   g14645(.A1(new_n13109_), .A2(new_n17693_), .B(pi0038), .ZN(new_n17716_));
  OAI21_X1   g14646(.A1(new_n17715_), .A2(new_n17716_), .B(new_n3259_), .ZN(new_n17717_));
  NOR3_X1    g14647(.A1(new_n17176_), .A2(new_n13099_), .A3(new_n5800_), .ZN(new_n17718_));
  NOR2_X1    g14648(.A1(new_n17718_), .A2(pi0038), .ZN(new_n17719_));
  NAND2_X1   g14649(.A1(pi0162), .A2(pi0738), .ZN(new_n17720_));
  NOR4_X1    g14650(.A1(new_n17696_), .A2(new_n13109_), .A3(new_n17719_), .A4(new_n17720_), .ZN(new_n17721_));
  OAI21_X1   g14651(.A1(new_n17714_), .A2(new_n17717_), .B(new_n17721_), .ZN(new_n17722_));
  OAI21_X1   g14652(.A1(new_n17705_), .A2(new_n17722_), .B(new_n8297_), .ZN(new_n17723_));
  AOI21_X1   g14653(.A1(new_n17705_), .A2(new_n17722_), .B(new_n17723_), .ZN(new_n17724_));
  XOR2_X1    g14654(.A1(new_n17724_), .A2(new_n17184_), .Z(new_n17725_));
  AOI21_X1   g14655(.A1(new_n13226_), .A2(new_n16968_), .B(new_n17693_), .ZN(new_n17726_));
  NOR2_X1    g14656(.A1(new_n17726_), .A2(new_n14799_), .ZN(new_n17727_));
  XOR2_X1    g14657(.A1(new_n17727_), .A2(new_n16913_), .Z(new_n17728_));
  OAI21_X1   g14658(.A1(new_n17725_), .A2(new_n17728_), .B(pi0162), .ZN(po0319));
  INV_X1     g14659(.I(pi0737), .ZN(new_n17730_));
  NOR2_X1    g14660(.A1(new_n5800_), .A2(pi0777), .ZN(new_n17731_));
  NOR2_X1    g14661(.A1(new_n14298_), .A2(new_n17731_), .ZN(new_n17732_));
  XOR2_X1    g14662(.A1(new_n17732_), .A2(new_n13094_), .Z(new_n17733_));
  NAND2_X1   g14663(.A1(new_n17733_), .A2(pi0163), .ZN(new_n17734_));
  INV_X1     g14664(.I(pi0777), .ZN(new_n17735_));
  NOR3_X1    g14665(.A1(new_n17058_), .A2(new_n9456_), .A3(new_n17735_), .ZN(new_n17736_));
  NOR3_X1    g14666(.A1(new_n17057_), .A2(new_n9456_), .A3(pi0777), .ZN(new_n17737_));
  OAI21_X1   g14667(.A1(new_n17736_), .A2(new_n17737_), .B(new_n17042_), .ZN(new_n17738_));
  OAI21_X1   g14668(.A1(new_n17159_), .A2(pi0777), .B(new_n16968_), .ZN(new_n17739_));
  NOR3_X1    g14669(.A1(new_n17158_), .A2(new_n9456_), .A3(new_n17739_), .ZN(new_n17740_));
  NOR3_X1    g14670(.A1(new_n17157_), .A2(pi0163), .A3(new_n17739_), .ZN(new_n17741_));
  OAI21_X1   g14671(.A1(new_n17740_), .A2(new_n17741_), .B(new_n17107_), .ZN(new_n17742_));
  NAND3_X1   g14672(.A1(new_n17738_), .A2(new_n3262_), .A3(new_n17742_), .ZN(new_n17743_));
  NAND2_X1   g14673(.A1(new_n17743_), .A2(new_n17734_), .ZN(new_n17744_));
  AOI21_X1   g14674(.A1(new_n17744_), .A2(new_n16970_), .B(new_n17730_), .ZN(new_n17745_));
  NAND4_X1   g14675(.A1(new_n17076_), .A2(new_n9456_), .A3(new_n3098_), .A4(new_n17167_), .ZN(new_n17746_));
  NAND2_X1   g14676(.A1(new_n3183_), .A2(new_n9456_), .ZN(new_n17747_));
  AOI21_X1   g14677(.A1(new_n14366_), .A2(new_n17747_), .B(pi0777), .ZN(new_n17748_));
  OAI21_X1   g14678(.A1(pi0163), .A2(new_n16971_), .B(new_n17087_), .ZN(new_n17749_));
  AOI21_X1   g14679(.A1(new_n17746_), .A2(new_n17748_), .B(new_n17749_), .ZN(new_n17750_));
  NOR2_X1    g14680(.A1(new_n13624_), .A2(new_n9456_), .ZN(new_n17751_));
  OAI21_X1   g14681(.A1(new_n13109_), .A2(new_n17731_), .B(pi0038), .ZN(new_n17752_));
  OAI21_X1   g14682(.A1(new_n17751_), .A2(new_n17752_), .B(new_n3259_), .ZN(new_n17753_));
  NOR3_X1    g14683(.A1(new_n17176_), .A2(new_n17735_), .A3(new_n5800_), .ZN(new_n17754_));
  NOR2_X1    g14684(.A1(new_n17754_), .A2(pi0038), .ZN(new_n17755_));
  NAND2_X1   g14685(.A1(pi0163), .A2(pi0737), .ZN(new_n17756_));
  NOR4_X1    g14686(.A1(new_n17734_), .A2(new_n13109_), .A3(new_n17755_), .A4(new_n17756_), .ZN(new_n17757_));
  OAI21_X1   g14687(.A1(new_n17750_), .A2(new_n17753_), .B(new_n17757_), .ZN(new_n17758_));
  OAI21_X1   g14688(.A1(new_n17745_), .A2(new_n17758_), .B(new_n8297_), .ZN(new_n17759_));
  AOI21_X1   g14689(.A1(new_n17745_), .A2(new_n17758_), .B(new_n17759_), .ZN(new_n17760_));
  XOR2_X1    g14690(.A1(new_n17760_), .A2(new_n17184_), .Z(new_n17761_));
  AOI21_X1   g14691(.A1(new_n17730_), .A2(new_n16968_), .B(new_n17731_), .ZN(new_n17762_));
  NOR2_X1    g14692(.A1(new_n17762_), .A2(new_n14799_), .ZN(new_n17763_));
  XOR2_X1    g14693(.A1(new_n17763_), .A2(new_n16913_), .Z(new_n17764_));
  OAI21_X1   g14694(.A1(new_n17761_), .A2(new_n17764_), .B(pi0163), .ZN(po0320));
  NAND2_X1   g14695(.A1(new_n17060_), .A2(pi0164), .ZN(new_n17766_));
  NAND2_X1   g14696(.A1(pi0038), .A2(pi0164), .ZN(new_n17767_));
  XOR2_X1    g14697(.A1(new_n17766_), .A2(new_n17767_), .Z(new_n17768_));
  INV_X1     g14698(.I(pi0752), .ZN(new_n17769_));
  OAI21_X1   g14699(.A1(new_n17022_), .A2(new_n17769_), .B(new_n7491_), .ZN(new_n17770_));
  NAND4_X1   g14700(.A1(new_n17768_), .A2(new_n13108_), .A3(new_n17043_), .A4(new_n17770_), .ZN(new_n17771_));
  INV_X1     g14701(.I(new_n16985_), .ZN(new_n17772_));
  NAND2_X1   g14702(.A1(new_n17015_), .A2(pi0164), .ZN(new_n17773_));
  XOR2_X1    g14703(.A1(new_n17773_), .A2(new_n17767_), .Z(new_n17774_));
  OAI21_X1   g14704(.A1(new_n17465_), .A2(new_n17769_), .B(new_n7491_), .ZN(new_n17775_));
  NAND4_X1   g14705(.A1(new_n17774_), .A2(new_n17772_), .A3(new_n17027_), .A4(new_n17775_), .ZN(new_n17776_));
  INV_X1     g14706(.I(pi0703), .ZN(new_n17777_));
  NAND2_X1   g14707(.A1(new_n17777_), .A2(pi0164), .ZN(new_n17778_));
  AOI21_X1   g14708(.A1(new_n13634_), .A2(pi0752), .B(new_n17778_), .ZN(new_n17779_));
  OAI21_X1   g14709(.A1(new_n17779_), .A2(new_n17098_), .B(pi0752), .ZN(new_n17780_));
  AOI21_X1   g14710(.A1(new_n17776_), .A2(new_n17771_), .B(new_n17780_), .ZN(new_n17781_));
  INV_X1     g14711(.I(new_n17065_), .ZN(new_n17782_));
  NOR4_X1    g14712(.A1(new_n17782_), .A2(new_n7491_), .A3(new_n17777_), .A4(new_n17769_), .ZN(new_n17783_));
  NOR3_X1    g14713(.A1(new_n17781_), .A2(new_n8345_), .A3(new_n17783_), .ZN(new_n17784_));
  XOR2_X1    g14714(.A1(new_n17784_), .A2(new_n17184_), .Z(new_n17785_));
  NAND2_X1   g14715(.A1(pi0752), .A2(pi0907), .ZN(new_n17786_));
  NAND3_X1   g14716(.A1(new_n17786_), .A2(new_n17777_), .A3(pi0947), .ZN(new_n17787_));
  NAND4_X1   g14717(.A1(pi0703), .A2(pi0752), .A3(pi0907), .A4(pi0947), .ZN(new_n17788_));
  NAND3_X1   g14718(.A1(new_n17787_), .A2(pi0832), .A3(new_n17788_), .ZN(new_n17789_));
  XOR2_X1    g14719(.A1(new_n17789_), .A2(new_n16961_), .Z(new_n17790_));
  OAI21_X1   g14720(.A1(new_n17785_), .A2(new_n17790_), .B(pi0164), .ZN(po0321));
  NAND2_X1   g14721(.A1(new_n17060_), .A2(pi0165), .ZN(new_n17792_));
  NAND2_X1   g14722(.A1(pi0038), .A2(pi0165), .ZN(new_n17793_));
  XOR2_X1    g14723(.A1(new_n17792_), .A2(new_n17793_), .Z(new_n17794_));
  OAI21_X1   g14724(.A1(new_n17022_), .A2(new_n15573_), .B(new_n10640_), .ZN(new_n17795_));
  NAND4_X1   g14725(.A1(new_n17794_), .A2(new_n13108_), .A3(new_n17043_), .A4(new_n17795_), .ZN(new_n17796_));
  NAND2_X1   g14726(.A1(new_n17015_), .A2(pi0165), .ZN(new_n17797_));
  XOR2_X1    g14727(.A1(new_n17797_), .A2(new_n17793_), .Z(new_n17798_));
  OAI21_X1   g14728(.A1(new_n17465_), .A2(new_n15573_), .B(new_n10640_), .ZN(new_n17799_));
  NAND4_X1   g14729(.A1(new_n17798_), .A2(new_n17772_), .A3(new_n17027_), .A4(new_n17799_), .ZN(new_n17800_));
  NAND2_X1   g14730(.A1(new_n15572_), .A2(pi0165), .ZN(new_n17801_));
  AOI21_X1   g14731(.A1(new_n13634_), .A2(pi0774), .B(new_n17801_), .ZN(new_n17802_));
  OAI21_X1   g14732(.A1(new_n17802_), .A2(new_n17098_), .B(pi0774), .ZN(new_n17803_));
  AOI21_X1   g14733(.A1(new_n17800_), .A2(new_n17796_), .B(new_n17803_), .ZN(new_n17804_));
  NOR4_X1    g14734(.A1(new_n17782_), .A2(new_n10640_), .A3(new_n15572_), .A4(new_n15573_), .ZN(new_n17805_));
  NOR3_X1    g14735(.A1(new_n17804_), .A2(new_n8345_), .A3(new_n17805_), .ZN(new_n17806_));
  XOR2_X1    g14736(.A1(new_n17806_), .A2(new_n17184_), .Z(new_n17807_));
  NAND2_X1   g14737(.A1(pi0774), .A2(pi0907), .ZN(new_n17808_));
  NAND3_X1   g14738(.A1(new_n17808_), .A2(new_n15572_), .A3(pi0947), .ZN(new_n17809_));
  NAND4_X1   g14739(.A1(pi0687), .A2(pi0774), .A3(pi0907), .A4(pi0947), .ZN(new_n17810_));
  NAND3_X1   g14740(.A1(new_n17809_), .A2(pi0832), .A3(new_n17810_), .ZN(new_n17811_));
  XOR2_X1    g14741(.A1(new_n17811_), .A2(new_n16961_), .Z(new_n17812_));
  OAI21_X1   g14742(.A1(new_n17807_), .A2(new_n17812_), .B(pi0165), .ZN(po0322));
  AOI21_X1   g14743(.A1(new_n16993_), .A2(pi0166), .B(new_n17284_), .ZN(new_n17814_));
  INV_X1     g14744(.I(new_n16997_), .ZN(new_n17815_));
  AOI21_X1   g14745(.A1(new_n4808_), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n17816_));
  AND2_X2    g14746(.A1(new_n17816_), .A2(pi0299), .Z(new_n17817_));
  OAI21_X1   g14747(.A1(new_n17817_), .A2(new_n16968_), .B(new_n17033_), .ZN(new_n17818_));
  NOR2_X1    g14748(.A1(new_n12784_), .A2(pi0166), .ZN(new_n17819_));
  AOI21_X1   g14749(.A1(new_n5452_), .A2(new_n12784_), .B(new_n17819_), .ZN(new_n17820_));
  OAI21_X1   g14750(.A1(new_n17820_), .A2(new_n3313_), .B(new_n3111_), .ZN(new_n17821_));
  NAND3_X1   g14751(.A1(new_n17818_), .A2(new_n17815_), .A3(new_n17821_), .ZN(new_n17822_));
  NOR2_X1    g14752(.A1(pi0039), .A2(pi0772), .ZN(new_n17823_));
  INV_X1     g14753(.I(new_n17823_), .ZN(new_n17824_));
  AOI21_X1   g14754(.A1(new_n17822_), .A2(new_n17814_), .B(new_n17824_), .ZN(new_n17825_));
  OAI21_X1   g14755(.A1(new_n4808_), .A2(new_n3090_), .B(new_n17045_), .ZN(new_n17826_));
  NAND2_X1   g14756(.A1(new_n17826_), .A2(new_n5452_), .ZN(new_n17827_));
  NAND2_X1   g14757(.A1(new_n17827_), .A2(new_n3098_), .ZN(new_n17828_));
  NOR2_X1    g14758(.A1(new_n17820_), .A2(new_n3092_), .ZN(new_n17829_));
  NOR2_X1    g14759(.A1(new_n17829_), .A2(pi0223), .ZN(new_n17830_));
  AOI21_X1   g14760(.A1(new_n17088_), .A2(new_n3091_), .B(new_n4808_), .ZN(new_n17831_));
  NAND4_X1   g14761(.A1(new_n17301_), .A2(new_n17828_), .A3(new_n17830_), .A4(new_n17831_), .ZN(new_n17832_));
  OAI21_X1   g14762(.A1(new_n17306_), .A2(pi0166), .B(new_n17052_), .ZN(new_n17833_));
  NAND2_X1   g14763(.A1(new_n17833_), .A2(new_n17827_), .ZN(new_n17834_));
  NAND3_X1   g14764(.A1(new_n17316_), .A2(new_n16968_), .A3(new_n17298_), .ZN(new_n17835_));
  INV_X1     g14765(.I(new_n17298_), .ZN(new_n17836_));
  NAND3_X1   g14766(.A1(new_n17316_), .A2(new_n16969_), .A3(new_n17836_), .ZN(new_n17837_));
  NAND2_X1   g14767(.A1(new_n17830_), .A2(pi0166), .ZN(new_n17838_));
  AOI21_X1   g14768(.A1(new_n17837_), .A2(new_n17835_), .B(new_n17838_), .ZN(new_n17839_));
  AOI21_X1   g14769(.A1(new_n17834_), .A2(new_n17839_), .B(pi0772), .ZN(new_n17840_));
  OAI21_X1   g14770(.A1(new_n17825_), .A2(new_n17832_), .B(new_n17840_), .ZN(new_n17841_));
  AOI21_X1   g14771(.A1(new_n17814_), .A2(new_n12831_), .B(new_n17821_), .ZN(new_n17842_));
  NOR3_X1    g14772(.A1(new_n17842_), .A2(new_n3098_), .A3(new_n17816_), .ZN(new_n17843_));
  AOI21_X1   g14773(.A1(new_n17841_), .A2(new_n17843_), .B(pi0038), .ZN(new_n17844_));
  INV_X1     g14774(.I(pi0772), .ZN(new_n17845_));
  NOR2_X1    g14775(.A1(new_n17845_), .A2(new_n5800_), .ZN(new_n17846_));
  NAND3_X1   g14776(.A1(new_n14874_), .A2(pi0039), .A3(new_n17846_), .ZN(new_n17847_));
  OR3_X2     g14777(.A1(new_n14298_), .A2(pi0039), .A3(new_n17846_), .Z(new_n17848_));
  AOI21_X1   g14778(.A1(new_n17847_), .A2(new_n17848_), .B(new_n4808_), .ZN(new_n17849_));
  AND2_X2    g14779(.A1(new_n17814_), .A2(new_n12974_), .Z(new_n17850_));
  AOI21_X1   g14780(.A1(new_n5800_), .A2(new_n12784_), .B(new_n17819_), .ZN(new_n17851_));
  NOR2_X1    g14781(.A1(new_n17851_), .A2(new_n3313_), .ZN(new_n17852_));
  OAI21_X1   g14782(.A1(new_n17850_), .A2(new_n17332_), .B(new_n17852_), .ZN(new_n17853_));
  NAND2_X1   g14783(.A1(new_n17074_), .A2(pi0166), .ZN(new_n17854_));
  AOI21_X1   g14784(.A1(new_n17853_), .A2(new_n17094_), .B(new_n17854_), .ZN(new_n17855_));
  AOI21_X1   g14785(.A1(new_n4808_), .A2(new_n17823_), .B(new_n17127_), .ZN(new_n17856_));
  NOR3_X1    g14786(.A1(new_n17855_), .A2(pi0772), .A3(new_n17856_), .ZN(new_n17857_));
  INV_X1     g14787(.I(new_n17851_), .ZN(new_n17858_));
  OAI22_X1   g14788(.A1(new_n17833_), .A2(new_n3090_), .B1(new_n3092_), .B2(new_n17858_), .ZN(new_n17859_));
  NAND3_X1   g14789(.A1(new_n17859_), .A2(pi0166), .A3(new_n17312_), .ZN(new_n17860_));
  NOR2_X1    g14790(.A1(new_n13109_), .A2(new_n17846_), .ZN(new_n17861_));
  NAND2_X1   g14791(.A1(pi0038), .A2(pi0727), .ZN(new_n17862_));
  OAI21_X1   g14792(.A1(new_n17861_), .A2(new_n17862_), .B(new_n4808_), .ZN(new_n17863_));
  AOI21_X1   g14793(.A1(new_n17863_), .A2(new_n13624_), .B(pi0038), .ZN(new_n17864_));
  OAI21_X1   g14794(.A1(new_n17857_), .A2(new_n17860_), .B(new_n17864_), .ZN(new_n17865_));
  INV_X1     g14795(.I(pi0727), .ZN(new_n17866_));
  NOR4_X1    g14796(.A1(new_n14291_), .A2(pi0039), .A3(new_n16968_), .A4(new_n17846_), .ZN(new_n17867_));
  NOR2_X1    g14797(.A1(new_n17867_), .A2(pi0038), .ZN(new_n17868_));
  NAND2_X1   g14798(.A1(new_n13108_), .A2(pi0166), .ZN(new_n17869_));
  OAI21_X1   g14799(.A1(new_n17868_), .A2(new_n17869_), .B(new_n17866_), .ZN(new_n17870_));
  AOI21_X1   g14800(.A1(new_n17865_), .A2(new_n17849_), .B(new_n17870_), .ZN(new_n17871_));
  NAND2_X1   g14801(.A1(new_n17849_), .A2(new_n16970_), .ZN(new_n17872_));
  NOR3_X1    g14802(.A1(new_n17871_), .A2(new_n17844_), .A3(new_n17872_), .ZN(new_n17873_));
  NOR2_X1    g14803(.A1(new_n17873_), .A2(new_n8345_), .ZN(new_n17874_));
  XNOR2_X1   g14804(.A1(new_n17874_), .A2(new_n17184_), .ZN(new_n17875_));
  NOR2_X1    g14805(.A1(new_n17846_), .A2(new_n9992_), .ZN(new_n17876_));
  NOR3_X1    g14806(.A1(new_n17876_), .A2(new_n17866_), .A3(new_n16969_), .ZN(new_n17877_));
  OAI21_X1   g14807(.A1(new_n9992_), .A2(pi0166), .B(pi0832), .ZN(new_n17878_));
  OAI22_X1   g14808(.A1(new_n17875_), .A2(new_n4808_), .B1(new_n17877_), .B2(new_n17878_), .ZN(po0323));
  INV_X1     g14809(.I(pi0705), .ZN(new_n17880_));
  INV_X1     g14810(.I(pi0768), .ZN(new_n17881_));
  NAND2_X1   g14811(.A1(pi0038), .A2(pi0167), .ZN(new_n17882_));
  NAND2_X1   g14812(.A1(new_n17060_), .A2(pi0167), .ZN(new_n17883_));
  XOR2_X1    g14813(.A1(new_n17883_), .A2(new_n17882_), .Z(new_n17884_));
  NAND2_X1   g14814(.A1(new_n17884_), .A2(new_n17043_), .ZN(new_n17885_));
  NAND3_X1   g14815(.A1(new_n17885_), .A2(new_n17880_), .A3(new_n17881_), .ZN(new_n17886_));
  AOI21_X1   g14816(.A1(new_n17028_), .A2(new_n8029_), .B(new_n17465_), .ZN(new_n17887_));
  NOR2_X1    g14817(.A1(new_n13108_), .A2(pi0167), .ZN(new_n17888_));
  OAI21_X1   g14818(.A1(new_n17022_), .A2(new_n17888_), .B(new_n17881_), .ZN(new_n17889_));
  AOI21_X1   g14819(.A1(new_n17886_), .A2(new_n17887_), .B(new_n17889_), .ZN(new_n17890_));
  NOR2_X1    g14820(.A1(new_n17084_), .A2(new_n17881_), .ZN(new_n17891_));
  NOR2_X1    g14821(.A1(new_n17891_), .A2(pi0167), .ZN(new_n17892_));
  NOR3_X1    g14822(.A1(new_n13632_), .A2(new_n3259_), .A3(new_n17881_), .ZN(new_n17893_));
  NOR3_X1    g14823(.A1(new_n13097_), .A2(pi0038), .A3(new_n17881_), .ZN(new_n17894_));
  OAI21_X1   g14824(.A1(new_n17893_), .A2(new_n17894_), .B(new_n13624_), .ZN(new_n17895_));
  NOR2_X1    g14825(.A1(new_n17895_), .A2(pi0167), .ZN(new_n17896_));
  NAND2_X1   g14826(.A1(new_n8297_), .A2(new_n17880_), .ZN(new_n17897_));
  OAI22_X1   g14827(.A1(new_n17896_), .A2(new_n17897_), .B1(new_n13625_), .B2(new_n17892_), .ZN(new_n17898_));
  NOR2_X1    g14828(.A1(new_n17079_), .A2(new_n8029_), .ZN(new_n17899_));
  XOR2_X1    g14829(.A1(new_n17899_), .A2(new_n17882_), .Z(new_n17900_));
  NOR2_X1    g14830(.A1(new_n17900_), .A2(new_n17097_), .ZN(new_n17901_));
  NAND2_X1   g14831(.A1(pi0768), .A2(pi0907), .ZN(new_n17902_));
  NAND3_X1   g14832(.A1(new_n17902_), .A2(new_n17880_), .A3(pi0947), .ZN(new_n17903_));
  NAND4_X1   g14833(.A1(pi0705), .A2(pi0768), .A3(pi0907), .A4(pi0947), .ZN(new_n17904_));
  NAND3_X1   g14834(.A1(new_n17903_), .A2(pi0832), .A3(new_n17904_), .ZN(new_n17905_));
  XOR2_X1    g14835(.A1(new_n17905_), .A2(new_n16961_), .Z(new_n17906_));
  NOR2_X1    g14836(.A1(new_n8029_), .A2(pi0832), .ZN(new_n17907_));
  AOI22_X1   g14837(.A1(new_n17901_), .A2(new_n17898_), .B1(new_n17906_), .B2(new_n17907_), .ZN(new_n17908_));
  NAND2_X1   g14838(.A1(new_n17015_), .A2(pi0167), .ZN(new_n17909_));
  XNOR2_X1   g14839(.A1(new_n17909_), .A2(new_n17882_), .ZN(new_n17910_));
  NOR4_X1    g14840(.A1(new_n17890_), .A2(new_n16985_), .A3(new_n17908_), .A4(new_n17910_), .ZN(po0324));
  INV_X1     g14841(.I(pi0763), .ZN(new_n17912_));
  NAND2_X1   g14842(.A1(new_n14299_), .A2(new_n17912_), .ZN(new_n17913_));
  AOI22_X1   g14843(.A1(new_n17086_), .A2(new_n17913_), .B1(new_n4635_), .B2(new_n14298_), .ZN(new_n17914_));
  NOR2_X1    g14844(.A1(new_n17358_), .A2(pi0168), .ZN(new_n17915_));
  AOI21_X1   g14845(.A1(pi0168), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n17916_));
  NOR2_X1    g14846(.A1(new_n17916_), .A2(new_n17034_), .ZN(new_n17917_));
  OAI22_X1   g14847(.A1(new_n17915_), .A2(new_n12809_), .B1(new_n17917_), .B2(new_n17362_), .ZN(new_n17918_));
  NOR2_X1    g14848(.A1(new_n16971_), .A2(pi0168), .ZN(new_n17919_));
  OAI21_X1   g14849(.A1(new_n16973_), .A2(new_n17919_), .B(new_n17912_), .ZN(new_n17920_));
  AOI21_X1   g14850(.A1(new_n17238_), .A2(new_n4635_), .B(new_n12831_), .ZN(new_n17921_));
  NAND4_X1   g14851(.A1(new_n17918_), .A2(pi0299), .A3(new_n17920_), .A4(new_n17921_), .ZN(new_n17922_));
  INV_X1     g14852(.I(new_n17921_), .ZN(new_n17923_));
  AOI21_X1   g14853(.A1(new_n4635_), .A2(new_n12809_), .B(new_n17370_), .ZN(new_n17924_));
  NAND2_X1   g14854(.A1(new_n17924_), .A2(pi0215), .ZN(new_n17925_));
  NAND2_X1   g14855(.A1(new_n17925_), .A2(new_n5741_), .ZN(new_n17926_));
  AOI22_X1   g14856(.A1(new_n17916_), .A2(pi0299), .B1(new_n12784_), .B2(new_n17926_), .ZN(new_n17927_));
  NOR3_X1    g14857(.A1(new_n17368_), .A2(new_n17923_), .A3(new_n17927_), .ZN(new_n17928_));
  NOR3_X1    g14858(.A1(new_n17263_), .A2(new_n3259_), .A3(new_n17912_), .ZN(new_n17929_));
  OAI21_X1   g14859(.A1(new_n17928_), .A2(pi0168), .B(new_n17929_), .ZN(new_n17930_));
  AOI21_X1   g14860(.A1(new_n3183_), .A2(new_n17922_), .B(new_n17930_), .ZN(new_n17931_));
  OAI21_X1   g14861(.A1(new_n17931_), .A2(new_n17914_), .B(new_n16970_), .ZN(new_n17932_));
  NOR2_X1    g14862(.A1(new_n13081_), .A2(new_n17912_), .ZN(new_n17933_));
  OAI21_X1   g14863(.A1(new_n17380_), .A2(pi0168), .B(new_n17933_), .ZN(new_n17934_));
  NAND2_X1   g14864(.A1(new_n17934_), .A2(new_n17070_), .ZN(new_n17935_));
  NOR3_X1    g14865(.A1(new_n17923_), .A2(new_n17384_), .A3(new_n17924_), .ZN(new_n17936_));
  AOI21_X1   g14866(.A1(new_n17935_), .A2(new_n17936_), .B(pi0168), .ZN(new_n17937_));
  NAND2_X1   g14867(.A1(new_n3183_), .A2(new_n4635_), .ZN(new_n17938_));
  OAI22_X1   g14868(.A1(new_n17914_), .A2(pi0038), .B1(pi0763), .B2(new_n17938_), .ZN(new_n17939_));
  OR3_X2     g14869(.A1(new_n17939_), .A2(new_n17127_), .A3(new_n17003_), .Z(new_n17940_));
  NOR2_X1    g14870(.A1(new_n17123_), .A2(pi0699), .ZN(new_n17941_));
  OAI21_X1   g14871(.A1(new_n17937_), .A2(new_n17940_), .B(new_n17941_), .ZN(new_n17942_));
  INV_X1     g14872(.I(pi0699), .ZN(new_n17943_));
  AOI21_X1   g14873(.A1(pi0763), .A2(pi0947), .B(new_n2723_), .ZN(new_n17944_));
  AOI21_X1   g14874(.A1(new_n5503_), .A2(new_n17944_), .B(pi0038), .ZN(new_n17945_));
  NOR4_X1    g14875(.A1(new_n13625_), .A2(new_n4635_), .A3(new_n17943_), .A4(new_n17945_), .ZN(new_n17946_));
  NAND2_X1   g14876(.A1(new_n17942_), .A2(new_n17946_), .ZN(new_n17947_));
  NOR3_X1    g14877(.A1(new_n17176_), .A2(new_n17912_), .A3(new_n5800_), .ZN(new_n17948_));
  NAND2_X1   g14878(.A1(new_n5371_), .A2(pi0168), .ZN(new_n17952_));
  NOR2_X1    g14879(.A1(new_n13109_), .A2(new_n17952_), .ZN(new_n17953_));
  OAI21_X1   g14880(.A1(new_n17948_), .A2(pi0038), .B(new_n17953_), .ZN(new_n17954_));
  AOI21_X1   g14881(.A1(new_n17932_), .A2(new_n17947_), .B(new_n17954_), .ZN(po0325));
  INV_X1     g14882(.I(pi0746), .ZN(new_n17956_));
  NAND2_X1   g14883(.A1(new_n14299_), .A2(new_n17956_), .ZN(new_n17957_));
  AOI22_X1   g14884(.A1(new_n17086_), .A2(new_n17957_), .B1(new_n4474_), .B2(new_n14298_), .ZN(new_n17958_));
  NOR2_X1    g14885(.A1(new_n17358_), .A2(pi0169), .ZN(new_n17959_));
  AOI21_X1   g14886(.A1(pi0169), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n17960_));
  NOR2_X1    g14887(.A1(new_n17960_), .A2(new_n17034_), .ZN(new_n17961_));
  OAI22_X1   g14888(.A1(new_n17959_), .A2(new_n12809_), .B1(new_n17961_), .B2(new_n17362_), .ZN(new_n17962_));
  NOR2_X1    g14889(.A1(new_n16971_), .A2(pi0169), .ZN(new_n17963_));
  OAI21_X1   g14890(.A1(new_n16973_), .A2(new_n17963_), .B(new_n17956_), .ZN(new_n17964_));
  AOI21_X1   g14891(.A1(new_n17238_), .A2(new_n4474_), .B(new_n12831_), .ZN(new_n17965_));
  NAND4_X1   g14892(.A1(new_n17962_), .A2(pi0299), .A3(new_n17964_), .A4(new_n17965_), .ZN(new_n17966_));
  INV_X1     g14893(.I(new_n17965_), .ZN(new_n17967_));
  AOI21_X1   g14894(.A1(new_n4474_), .A2(new_n12809_), .B(new_n17370_), .ZN(new_n17968_));
  NAND2_X1   g14895(.A1(new_n17968_), .A2(pi0215), .ZN(new_n17969_));
  NAND2_X1   g14896(.A1(new_n17969_), .A2(new_n5741_), .ZN(new_n17970_));
  AOI22_X1   g14897(.A1(new_n17960_), .A2(pi0299), .B1(new_n12784_), .B2(new_n17970_), .ZN(new_n17971_));
  NOR3_X1    g14898(.A1(new_n17368_), .A2(new_n17967_), .A3(new_n17971_), .ZN(new_n17972_));
  NOR3_X1    g14899(.A1(new_n17263_), .A2(new_n3259_), .A3(new_n17956_), .ZN(new_n17973_));
  OAI21_X1   g14900(.A1(new_n17972_), .A2(pi0169), .B(new_n17973_), .ZN(new_n17974_));
  AOI21_X1   g14901(.A1(new_n3183_), .A2(new_n17966_), .B(new_n17974_), .ZN(new_n17975_));
  OAI21_X1   g14902(.A1(new_n17975_), .A2(new_n17958_), .B(new_n16970_), .ZN(new_n17976_));
  NOR2_X1    g14903(.A1(new_n13081_), .A2(new_n17956_), .ZN(new_n17977_));
  OAI21_X1   g14904(.A1(new_n17380_), .A2(pi0169), .B(new_n17977_), .ZN(new_n17978_));
  NAND2_X1   g14905(.A1(new_n17978_), .A2(new_n17070_), .ZN(new_n17979_));
  NOR3_X1    g14906(.A1(new_n17967_), .A2(new_n17384_), .A3(new_n17968_), .ZN(new_n17980_));
  AOI21_X1   g14907(.A1(new_n17979_), .A2(new_n17980_), .B(pi0169), .ZN(new_n17981_));
  NAND2_X1   g14908(.A1(new_n3183_), .A2(new_n4474_), .ZN(new_n17982_));
  OAI22_X1   g14909(.A1(new_n17958_), .A2(pi0038), .B1(pi0746), .B2(new_n17982_), .ZN(new_n17983_));
  OR3_X2     g14910(.A1(new_n17983_), .A2(new_n17127_), .A3(new_n17003_), .Z(new_n17984_));
  NOR2_X1    g14911(.A1(new_n17123_), .A2(pi0729), .ZN(new_n17985_));
  OAI21_X1   g14912(.A1(new_n17981_), .A2(new_n17984_), .B(new_n17985_), .ZN(new_n17986_));
  INV_X1     g14913(.I(pi0729), .ZN(new_n17987_));
  AOI21_X1   g14914(.A1(pi0746), .A2(pi0947), .B(new_n2723_), .ZN(new_n17988_));
  AOI21_X1   g14915(.A1(new_n5503_), .A2(new_n17988_), .B(pi0038), .ZN(new_n17989_));
  NOR4_X1    g14916(.A1(new_n13625_), .A2(new_n4474_), .A3(new_n17987_), .A4(new_n17989_), .ZN(new_n17990_));
  NAND2_X1   g14917(.A1(new_n17986_), .A2(new_n17990_), .ZN(new_n17991_));
  NOR3_X1    g14918(.A1(new_n17176_), .A2(new_n17956_), .A3(new_n5800_), .ZN(new_n17992_));
  NAND2_X1   g14919(.A1(new_n5371_), .A2(pi0169), .ZN(new_n17996_));
  NOR2_X1    g14920(.A1(new_n13109_), .A2(new_n17996_), .ZN(new_n17997_));
  OAI21_X1   g14921(.A1(new_n17992_), .A2(pi0038), .B(new_n17997_), .ZN(new_n17998_));
  AOI21_X1   g14922(.A1(new_n17976_), .A2(new_n17991_), .B(new_n17998_), .ZN(po0326));
  INV_X1     g14923(.I(pi0748), .ZN(new_n18000_));
  OAI21_X1   g14924(.A1(new_n17022_), .A2(new_n18000_), .B(new_n4150_), .ZN(new_n18001_));
  NAND2_X1   g14925(.A1(new_n18001_), .A2(new_n13108_), .ZN(new_n18002_));
  OR2_X2     g14926(.A1(new_n17084_), .A2(new_n18000_), .Z(new_n18003_));
  AOI21_X1   g14927(.A1(new_n18003_), .A2(new_n4150_), .B(new_n13625_), .ZN(new_n18004_));
  NOR3_X1    g14928(.A1(new_n13634_), .A2(pi0730), .A3(pi0748), .ZN(new_n18005_));
  NOR3_X1    g14929(.A1(new_n18005_), .A2(new_n4150_), .A3(new_n17124_), .ZN(new_n18006_));
  NAND3_X1   g14930(.A1(new_n16971_), .A2(pi0299), .A3(pi0947), .ZN(new_n18007_));
  NAND3_X1   g14931(.A1(new_n16971_), .A2(new_n3098_), .A3(new_n5800_), .ZN(new_n18008_));
  AOI21_X1   g14932(.A1(new_n18007_), .A2(new_n18008_), .B(new_n4150_), .ZN(new_n18009_));
  OAI21_X1   g14933(.A1(pi0170), .A2(new_n12784_), .B(new_n17089_), .ZN(new_n18010_));
  OAI21_X1   g14934(.A1(new_n17380_), .A2(pi0170), .B(new_n12942_), .ZN(new_n18011_));
  AOI21_X1   g14935(.A1(new_n17238_), .A2(new_n4150_), .B(new_n12831_), .ZN(new_n18012_));
  NOR2_X1    g14936(.A1(new_n17071_), .A2(new_n18012_), .ZN(new_n18013_));
  AOI21_X1   g14937(.A1(new_n18011_), .A2(new_n18013_), .B(new_n18010_), .ZN(new_n18014_));
  OAI21_X1   g14938(.A1(new_n18014_), .A2(new_n18009_), .B(new_n3262_), .ZN(new_n18015_));
  AOI21_X1   g14939(.A1(pi0170), .A2(new_n17263_), .B(new_n17368_), .ZN(new_n18016_));
  NOR2_X1    g14940(.A1(new_n14874_), .A2(pi0170), .ZN(new_n18017_));
  OAI21_X1   g14941(.A1(new_n18017_), .A2(new_n17031_), .B(new_n3183_), .ZN(new_n18018_));
  INV_X1     g14942(.I(new_n18012_), .ZN(new_n18019_));
  INV_X1     g14943(.I(new_n18017_), .ZN(new_n18020_));
  OAI21_X1   g14944(.A1(new_n18010_), .A2(new_n3111_), .B(new_n5741_), .ZN(new_n18021_));
  AOI21_X1   g14945(.A1(pi0170), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n18022_));
  AOI22_X1   g14946(.A1(new_n18022_), .A2(pi0299), .B1(new_n12784_), .B2(new_n18021_), .ZN(new_n18023_));
  OAI21_X1   g14947(.A1(new_n17465_), .A2(new_n18000_), .B(new_n4150_), .ZN(new_n18024_));
  INV_X1     g14948(.I(pi0730), .ZN(new_n18025_));
  NOR2_X1    g14949(.A1(new_n13109_), .A2(new_n18025_), .ZN(new_n18026_));
  AOI21_X1   g14950(.A1(new_n18024_), .A2(new_n18026_), .B(pi0038), .ZN(new_n18027_));
  NOR4_X1    g14951(.A1(new_n18023_), .A2(new_n18019_), .A3(new_n18020_), .A4(new_n18027_), .ZN(new_n18028_));
  OAI21_X1   g14952(.A1(new_n18016_), .A2(new_n18018_), .B(new_n18028_), .ZN(new_n18029_));
  AOI21_X1   g14953(.A1(new_n17086_), .A2(new_n18015_), .B(new_n18029_), .ZN(new_n18030_));
  OAI21_X1   g14954(.A1(new_n18004_), .A2(new_n18006_), .B(new_n18030_), .ZN(new_n18031_));
  NOR3_X1    g14955(.A1(new_n17003_), .A2(new_n3098_), .A3(new_n16969_), .ZN(new_n18032_));
  NOR3_X1    g14956(.A1(new_n17003_), .A2(pi0299), .A3(new_n16968_), .ZN(new_n18033_));
  NOR2_X1    g14957(.A1(new_n3183_), .A2(new_n4150_), .ZN(new_n18034_));
  OAI21_X1   g14958(.A1(new_n18032_), .A2(new_n18033_), .B(new_n18034_), .ZN(new_n18035_));
  NOR2_X1    g14959(.A1(new_n17358_), .A2(pi0170), .ZN(new_n18036_));
  NOR2_X1    g14960(.A1(new_n18022_), .A2(new_n17034_), .ZN(new_n18037_));
  OAI22_X1   g14961(.A1(new_n18036_), .A2(new_n12809_), .B1(new_n18037_), .B2(new_n17362_), .ZN(new_n18038_));
  NAND3_X1   g14962(.A1(new_n18038_), .A2(pi0038), .A3(new_n18012_), .ZN(new_n18039_));
  AOI21_X1   g14963(.A1(new_n18035_), .A2(new_n3098_), .B(new_n18039_), .ZN(new_n18040_));
  NAND2_X1   g14964(.A1(new_n17124_), .A2(new_n4150_), .ZN(new_n18041_));
  NOR2_X1    g14965(.A1(new_n9992_), .A2(new_n4150_), .ZN(new_n18042_));
  OAI21_X1   g14966(.A1(new_n18000_), .A2(new_n5800_), .B(new_n16913_), .ZN(new_n18043_));
  OAI21_X1   g14967(.A1(new_n18043_), .A2(new_n18042_), .B(new_n18025_), .ZN(new_n18044_));
  INV_X1     g14968(.I(new_n17401_), .ZN(new_n18045_));
  AOI21_X1   g14969(.A1(pi0057), .A2(pi0170), .B(new_n18045_), .ZN(new_n18046_));
  AOI22_X1   g14970(.A1(new_n18041_), .A2(new_n5371_), .B1(new_n18044_), .B2(new_n18046_), .ZN(new_n18047_));
  NOR2_X1    g14971(.A1(new_n18020_), .A2(new_n18047_), .ZN(new_n18048_));
  OAI21_X1   g14972(.A1(new_n18040_), .A2(new_n17255_), .B(new_n18048_), .ZN(new_n18049_));
  AOI21_X1   g14973(.A1(new_n18031_), .A2(new_n18002_), .B(new_n18049_), .ZN(po0327));
  INV_X1     g14974(.I(pi0764), .ZN(new_n18051_));
  NAND2_X1   g14975(.A1(new_n14299_), .A2(new_n18051_), .ZN(new_n18052_));
  AOI22_X1   g14976(.A1(new_n17086_), .A2(new_n18052_), .B1(new_n3989_), .B2(new_n14298_), .ZN(new_n18053_));
  NOR2_X1    g14977(.A1(new_n17358_), .A2(pi0171), .ZN(new_n18054_));
  AOI21_X1   g14978(.A1(pi0171), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n18055_));
  NOR2_X1    g14979(.A1(new_n18055_), .A2(new_n17034_), .ZN(new_n18056_));
  OAI22_X1   g14980(.A1(new_n18054_), .A2(new_n12809_), .B1(new_n18056_), .B2(new_n17362_), .ZN(new_n18057_));
  NOR2_X1    g14981(.A1(new_n16971_), .A2(pi0171), .ZN(new_n18058_));
  OAI21_X1   g14982(.A1(new_n16973_), .A2(new_n18058_), .B(new_n18051_), .ZN(new_n18059_));
  AOI21_X1   g14983(.A1(new_n17238_), .A2(new_n3989_), .B(new_n12831_), .ZN(new_n18060_));
  NAND4_X1   g14984(.A1(new_n18057_), .A2(pi0299), .A3(new_n18059_), .A4(new_n18060_), .ZN(new_n18061_));
  INV_X1     g14985(.I(new_n18060_), .ZN(new_n18062_));
  AOI21_X1   g14986(.A1(new_n3989_), .A2(new_n12809_), .B(new_n17370_), .ZN(new_n18063_));
  NAND2_X1   g14987(.A1(new_n18063_), .A2(pi0215), .ZN(new_n18064_));
  NAND2_X1   g14988(.A1(new_n18064_), .A2(new_n5741_), .ZN(new_n18065_));
  AOI22_X1   g14989(.A1(new_n18055_), .A2(pi0299), .B1(new_n12784_), .B2(new_n18065_), .ZN(new_n18066_));
  NOR3_X1    g14990(.A1(new_n17368_), .A2(new_n18062_), .A3(new_n18066_), .ZN(new_n18067_));
  NOR3_X1    g14991(.A1(new_n17263_), .A2(new_n3259_), .A3(new_n18051_), .ZN(new_n18068_));
  OAI21_X1   g14992(.A1(new_n18067_), .A2(pi0171), .B(new_n18068_), .ZN(new_n18069_));
  AOI21_X1   g14993(.A1(new_n3183_), .A2(new_n18061_), .B(new_n18069_), .ZN(new_n18070_));
  OAI21_X1   g14994(.A1(new_n18070_), .A2(new_n18053_), .B(new_n16970_), .ZN(new_n18071_));
  NOR2_X1    g14995(.A1(new_n13081_), .A2(new_n18051_), .ZN(new_n18072_));
  OAI21_X1   g14996(.A1(new_n17380_), .A2(pi0171), .B(new_n18072_), .ZN(new_n18073_));
  NAND2_X1   g14997(.A1(new_n18073_), .A2(new_n17070_), .ZN(new_n18074_));
  NOR3_X1    g14998(.A1(new_n18062_), .A2(new_n17384_), .A3(new_n18063_), .ZN(new_n18075_));
  AOI21_X1   g14999(.A1(new_n18074_), .A2(new_n18075_), .B(pi0171), .ZN(new_n18076_));
  NAND2_X1   g15000(.A1(new_n3183_), .A2(new_n3989_), .ZN(new_n18077_));
  OAI22_X1   g15001(.A1(new_n18053_), .A2(pi0038), .B1(pi0764), .B2(new_n18077_), .ZN(new_n18078_));
  OR3_X2     g15002(.A1(new_n18078_), .A2(new_n17127_), .A3(new_n17003_), .Z(new_n18079_));
  NOR2_X1    g15003(.A1(new_n17123_), .A2(pi0691), .ZN(new_n18080_));
  OAI21_X1   g15004(.A1(new_n18076_), .A2(new_n18079_), .B(new_n18080_), .ZN(new_n18081_));
  INV_X1     g15005(.I(pi0691), .ZN(new_n18082_));
  AOI21_X1   g15006(.A1(pi0764), .A2(pi0947), .B(new_n2723_), .ZN(new_n18083_));
  AOI21_X1   g15007(.A1(new_n5503_), .A2(new_n18083_), .B(pi0038), .ZN(new_n18084_));
  NOR4_X1    g15008(.A1(new_n13625_), .A2(new_n3989_), .A3(new_n18082_), .A4(new_n18084_), .ZN(new_n18085_));
  NAND2_X1   g15009(.A1(new_n18081_), .A2(new_n18085_), .ZN(new_n18086_));
  NOR3_X1    g15010(.A1(new_n17176_), .A2(new_n18051_), .A3(new_n5800_), .ZN(new_n18087_));
  NAND2_X1   g15011(.A1(new_n5371_), .A2(pi0171), .ZN(new_n18091_));
  NOR2_X1    g15012(.A1(new_n13109_), .A2(new_n18091_), .ZN(new_n18092_));
  OAI21_X1   g15013(.A1(new_n18087_), .A2(pi0038), .B(new_n18092_), .ZN(new_n18093_));
  AOI21_X1   g15014(.A1(new_n18071_), .A2(new_n18086_), .B(new_n18093_), .ZN(po0328));
  INV_X1     g15015(.I(pi0739), .ZN(new_n18095_));
  NOR2_X1    g15016(.A1(new_n18095_), .A2(new_n5800_), .ZN(new_n18096_));
  NAND3_X1   g15017(.A1(new_n14874_), .A2(pi0039), .A3(new_n18096_), .ZN(new_n18097_));
  INV_X1     g15018(.I(new_n18096_), .ZN(new_n18098_));
  NAND3_X1   g15019(.A1(new_n14874_), .A2(new_n3183_), .A3(new_n18098_), .ZN(new_n18099_));
  AOI21_X1   g15020(.A1(new_n18097_), .A2(new_n18099_), .B(new_n3827_), .ZN(new_n18100_));
  NOR2_X1    g15021(.A1(new_n17358_), .A2(pi0172), .ZN(new_n18101_));
  AOI21_X1   g15022(.A1(pi0172), .A2(new_n13081_), .B(new_n17073_), .ZN(new_n18102_));
  NOR2_X1    g15023(.A1(new_n18102_), .A2(new_n17034_), .ZN(new_n18103_));
  OAI22_X1   g15024(.A1(new_n18101_), .A2(new_n12809_), .B1(new_n18103_), .B2(new_n17362_), .ZN(new_n18104_));
  NOR2_X1    g15025(.A1(new_n16971_), .A2(pi0172), .ZN(new_n18105_));
  OAI21_X1   g15026(.A1(new_n16973_), .A2(new_n18105_), .B(new_n18095_), .ZN(new_n18106_));
  AOI21_X1   g15027(.A1(new_n17238_), .A2(new_n3827_), .B(new_n12831_), .ZN(new_n18107_));
  NAND4_X1   g15028(.A1(new_n18104_), .A2(pi0299), .A3(new_n18106_), .A4(new_n18107_), .ZN(new_n18108_));
  INV_X1     g15029(.I(new_n18107_), .ZN(new_n18109_));
  AOI21_X1   g15030(.A1(new_n3827_), .A2(new_n12809_), .B(new_n17370_), .ZN(new_n18110_));
  NAND2_X1   g15031(.A1(new_n18110_), .A2(pi0215), .ZN(new_n18111_));
  NAND2_X1   g15032(.A1(new_n18111_), .A2(new_n5741_), .ZN(new_n18112_));
  AOI22_X1   g15033(.A1(new_n18102_), .A2(pi0299), .B1(new_n12784_), .B2(new_n18112_), .ZN(new_n18113_));
  NOR3_X1    g15034(.A1(new_n17368_), .A2(new_n18109_), .A3(new_n18113_), .ZN(new_n18114_));
  NOR3_X1    g15035(.A1(new_n17263_), .A2(new_n3259_), .A3(new_n18095_), .ZN(new_n18115_));
  OAI21_X1   g15036(.A1(new_n18114_), .A2(pi0172), .B(new_n18115_), .ZN(new_n18116_));
  AOI21_X1   g15037(.A1(new_n3183_), .A2(new_n18108_), .B(new_n18116_), .ZN(new_n18117_));
  OAI21_X1   g15038(.A1(new_n18117_), .A2(new_n18100_), .B(new_n16970_), .ZN(new_n18118_));
  NOR2_X1    g15039(.A1(new_n13081_), .A2(new_n18095_), .ZN(new_n18119_));
  OAI21_X1   g15040(.A1(new_n17380_), .A2(pi0172), .B(new_n18119_), .ZN(new_n18120_));
  NAND2_X1   g15041(.A1(new_n18120_), .A2(new_n17070_), .ZN(new_n18121_));
  NOR3_X1    g15042(.A1(new_n18109_), .A2(new_n17384_), .A3(new_n18110_), .ZN(new_n18122_));
  AOI21_X1   g15043(.A1(new_n18121_), .A2(new_n18122_), .B(pi0172), .ZN(new_n18123_));
  NAND2_X1   g15044(.A1(new_n3183_), .A2(new_n3827_), .ZN(new_n18124_));
  OAI22_X1   g15045(.A1(new_n18100_), .A2(pi0038), .B1(pi0739), .B2(new_n18124_), .ZN(new_n18125_));
  OR3_X2     g15046(.A1(new_n17127_), .A2(new_n18125_), .A3(new_n17003_), .Z(new_n18126_));
  NOR2_X1    g15047(.A1(new_n17123_), .A2(pi0690), .ZN(new_n18127_));
  OAI21_X1   g15048(.A1(new_n18123_), .A2(new_n18126_), .B(new_n18127_), .ZN(new_n18128_));
  INV_X1     g15049(.I(pi0690), .ZN(new_n18129_));
  NOR2_X1    g15050(.A1(new_n18096_), .A2(new_n2723_), .ZN(new_n18130_));
  AOI21_X1   g15051(.A1(new_n5503_), .A2(new_n18130_), .B(pi0038), .ZN(new_n18131_));
  NOR4_X1    g15052(.A1(new_n13625_), .A2(new_n3827_), .A3(new_n18129_), .A4(new_n18131_), .ZN(new_n18132_));
  NAND2_X1   g15053(.A1(new_n18128_), .A2(new_n18132_), .ZN(new_n18133_));
  OAI21_X1   g15054(.A1(new_n17176_), .A2(new_n18098_), .B(new_n3259_), .ZN(new_n18134_));
  NOR2_X1    g15055(.A1(new_n3827_), .A2(pi0057), .ZN(new_n18139_));
  NAND3_X1   g15056(.A1(new_n18134_), .A2(new_n13108_), .A3(new_n18139_), .ZN(new_n18140_));
  AOI21_X1   g15057(.A1(new_n18118_), .A2(new_n18133_), .B(new_n18140_), .ZN(po0329));
  INV_X1     g15058(.I(new_n14051_), .ZN(new_n18142_));
  NOR3_X1    g15059(.A1(new_n13219_), .A2(pi0625), .A3(pi0723), .ZN(new_n18143_));
  INV_X1     g15060(.I(new_n18143_), .ZN(new_n18144_));
  NOR2_X1    g15061(.A1(new_n9992_), .A2(pi0173), .ZN(new_n18145_));
  NOR2_X1    g15062(.A1(new_n18145_), .A2(pi1153), .ZN(new_n18146_));
  NAND2_X1   g15063(.A1(new_n18144_), .A2(new_n18146_), .ZN(new_n18147_));
  INV_X1     g15064(.I(new_n18147_), .ZN(new_n18148_));
  NOR2_X1    g15065(.A1(new_n18148_), .A2(new_n13748_), .ZN(new_n18149_));
  AOI21_X1   g15066(.A1(new_n13218_), .A2(new_n17227_), .B(new_n18145_), .ZN(new_n18150_));
  INV_X1     g15067(.I(new_n18150_), .ZN(new_n18151_));
  AOI21_X1   g15068(.A1(new_n18144_), .A2(new_n18151_), .B(new_n13614_), .ZN(new_n18152_));
  INV_X1     g15069(.I(new_n18152_), .ZN(new_n18153_));
  NOR3_X1    g15070(.A1(new_n18153_), .A2(new_n13748_), .A3(new_n18151_), .ZN(new_n18154_));
  INV_X1     g15071(.I(new_n18154_), .ZN(new_n18155_));
  NOR2_X1    g15072(.A1(new_n18155_), .A2(new_n18149_), .ZN(new_n18156_));
  NAND2_X1   g15073(.A1(new_n18155_), .A2(new_n18149_), .ZN(new_n18157_));
  INV_X1     g15074(.I(new_n18157_), .ZN(new_n18158_));
  NOR2_X1    g15075(.A1(new_n18158_), .A2(new_n18156_), .ZN(new_n18159_));
  INV_X1     g15076(.I(new_n18159_), .ZN(new_n18160_));
  NOR2_X1    g15077(.A1(new_n18160_), .A2(new_n14048_), .ZN(new_n18161_));
  NAND2_X1   g15078(.A1(new_n18161_), .A2(new_n18142_), .ZN(new_n18162_));
  INV_X1     g15079(.I(new_n18162_), .ZN(new_n18163_));
  NOR2_X1    g15080(.A1(new_n18150_), .A2(new_n13203_), .ZN(new_n18164_));
  NAND2_X1   g15081(.A1(new_n18164_), .A2(pi0625), .ZN(new_n18165_));
  NOR2_X1    g15082(.A1(new_n13105_), .A2(pi0745), .ZN(new_n18166_));
  NOR2_X1    g15083(.A1(new_n18166_), .A2(new_n18145_), .ZN(new_n18167_));
  NAND3_X1   g15084(.A1(new_n18165_), .A2(pi1153), .A3(new_n18167_), .ZN(new_n18168_));
  NOR2_X1    g15085(.A1(new_n18148_), .A2(new_n14081_), .ZN(new_n18169_));
  AOI21_X1   g15086(.A1(new_n18169_), .A2(new_n18168_), .B(new_n13748_), .ZN(new_n18170_));
  INV_X1     g15087(.I(new_n18167_), .ZN(new_n18171_));
  NOR2_X1    g15088(.A1(new_n18171_), .A2(new_n18164_), .ZN(new_n18172_));
  INV_X1     g15089(.I(new_n18165_), .ZN(new_n18173_));
  OAI21_X1   g15090(.A1(new_n18172_), .A2(new_n18173_), .B(new_n18146_), .ZN(new_n18174_));
  NAND4_X1   g15091(.A1(new_n18174_), .A2(new_n13749_), .A3(new_n18153_), .A4(new_n18172_), .ZN(new_n18175_));
  XOR2_X1    g15092(.A1(new_n18175_), .A2(new_n18170_), .Z(new_n18176_));
  NAND2_X1   g15093(.A1(new_n18176_), .A2(pi1155), .ZN(new_n18177_));
  XOR2_X1    g15094(.A1(new_n18177_), .A2(new_n14090_), .Z(new_n18178_));
  NOR2_X1    g15095(.A1(new_n18178_), .A2(new_n18159_), .ZN(new_n18179_));
  INV_X1     g15096(.I(new_n18166_), .ZN(new_n18180_));
  NOR2_X1    g15097(.A1(new_n18145_), .A2(pi1155), .ZN(new_n18181_));
  NOR3_X1    g15098(.A1(new_n18180_), .A2(new_n16444_), .A3(new_n18181_), .ZN(new_n18182_));
  NOR3_X1    g15099(.A1(new_n18179_), .A2(new_n13783_), .A3(new_n18182_), .ZN(new_n18183_));
  INV_X1     g15100(.I(new_n14096_), .ZN(new_n18184_));
  NAND3_X1   g15101(.A1(new_n18171_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n18185_));
  AOI21_X1   g15102(.A1(new_n18185_), .A2(new_n16444_), .B(new_n18180_), .ZN(new_n18186_));
  NOR3_X1    g15103(.A1(new_n18183_), .A2(pi0660), .A3(new_n18186_), .ZN(new_n18187_));
  NAND2_X1   g15104(.A1(new_n18176_), .A2(pi0609), .ZN(new_n18188_));
  XOR2_X1    g15105(.A1(new_n18188_), .A2(new_n14694_), .Z(new_n18189_));
  NAND3_X1   g15106(.A1(new_n18189_), .A2(pi0785), .A3(new_n18160_), .ZN(new_n18190_));
  OAI22_X1   g15107(.A1(new_n18187_), .A2(new_n18190_), .B1(pi0785), .B2(new_n18176_), .ZN(new_n18191_));
  AND2_X2    g15108(.A1(new_n18191_), .A2(new_n13855_), .Z(new_n18192_));
  NOR2_X1    g15109(.A1(new_n18191_), .A2(new_n13816_), .ZN(new_n18193_));
  XOR2_X1    g15110(.A1(new_n18193_), .A2(new_n13818_), .Z(new_n18194_));
  NAND2_X1   g15111(.A1(new_n18194_), .A2(new_n18161_), .ZN(new_n18195_));
  NOR2_X1    g15112(.A1(new_n18186_), .A2(new_n13801_), .ZN(new_n18196_));
  NAND4_X1   g15113(.A1(new_n18182_), .A2(new_n18171_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n18197_));
  XOR2_X1    g15114(.A1(new_n18196_), .A2(new_n18197_), .Z(new_n18198_));
  NOR2_X1    g15115(.A1(new_n18198_), .A2(new_n13817_), .ZN(new_n18199_));
  OAI21_X1   g15116(.A1(new_n18199_), .A2(new_n9992_), .B(pi0618), .ZN(new_n18200_));
  NAND3_X1   g15117(.A1(new_n18195_), .A2(new_n13823_), .A3(new_n18200_), .ZN(new_n18201_));
  OAI21_X1   g15118(.A1(new_n18199_), .A2(pi0618), .B(new_n9992_), .ZN(new_n18202_));
  AND2_X2    g15119(.A1(new_n18202_), .A2(new_n13823_), .Z(new_n18203_));
  NOR2_X1    g15120(.A1(new_n18191_), .A2(new_n13817_), .ZN(new_n18204_));
  XOR2_X1    g15121(.A1(new_n18204_), .A2(new_n13818_), .Z(new_n18205_));
  NAND3_X1   g15122(.A1(new_n18205_), .A2(pi0781), .A3(new_n18161_), .ZN(new_n18206_));
  AOI21_X1   g15123(.A1(new_n18201_), .A2(new_n18203_), .B(new_n18206_), .ZN(new_n18207_));
  NOR2_X1    g15124(.A1(new_n18207_), .A2(new_n18192_), .ZN(new_n18208_));
  NAND2_X1   g15125(.A1(new_n18208_), .A2(pi0619), .ZN(new_n18209_));
  XOR2_X1    g15126(.A1(new_n18209_), .A2(new_n13904_), .Z(new_n18210_));
  NAND2_X1   g15127(.A1(new_n18210_), .A2(new_n18163_), .ZN(new_n18211_));
  NAND2_X1   g15128(.A1(new_n18202_), .A2(pi0781), .ZN(new_n18212_));
  NOR3_X1    g15129(.A1(new_n18200_), .A2(new_n13855_), .A3(new_n18198_), .ZN(new_n18213_));
  XOR2_X1    g15130(.A1(new_n18213_), .A2(new_n18212_), .Z(new_n18214_));
  NOR2_X1    g15131(.A1(new_n18214_), .A2(new_n13868_), .ZN(new_n18215_));
  NOR2_X1    g15132(.A1(new_n18215_), .A2(new_n9992_), .ZN(new_n18216_));
  NOR2_X1    g15133(.A1(new_n18216_), .A2(new_n13860_), .ZN(new_n18217_));
  NOR2_X1    g15134(.A1(new_n18217_), .A2(pi0648), .ZN(new_n18218_));
  INV_X1     g15135(.I(new_n18208_), .ZN(new_n18219_));
  OAI21_X1   g15136(.A1(new_n18219_), .A2(new_n15479_), .B(new_n13896_), .ZN(new_n18220_));
  AOI21_X1   g15137(.A1(new_n18211_), .A2(new_n18218_), .B(new_n18220_), .ZN(new_n18221_));
  NAND2_X1   g15138(.A1(new_n18208_), .A2(pi1159), .ZN(new_n18222_));
  XOR2_X1    g15139(.A1(new_n18222_), .A2(new_n13904_), .Z(new_n18223_));
  NAND2_X1   g15140(.A1(new_n18223_), .A2(new_n18163_), .ZN(new_n18224_));
  OAI21_X1   g15141(.A1(new_n18215_), .A2(pi0619), .B(new_n9992_), .ZN(new_n18225_));
  NAND4_X1   g15142(.A1(new_n18224_), .A2(pi0648), .A3(new_n16423_), .A4(new_n18225_), .ZN(new_n18226_));
  OAI21_X1   g15143(.A1(new_n18226_), .A2(new_n18221_), .B(new_n13937_), .ZN(new_n18227_));
  NAND2_X1   g15144(.A1(new_n18225_), .A2(pi0789), .ZN(new_n18228_));
  NOR4_X1    g15145(.A1(new_n18216_), .A2(new_n13860_), .A3(new_n13896_), .A4(new_n18214_), .ZN(new_n18229_));
  XOR2_X1    g15146(.A1(new_n18229_), .A2(new_n18228_), .Z(new_n18230_));
  NOR2_X1    g15147(.A1(new_n18230_), .A2(pi0788), .ZN(new_n18231_));
  NAND2_X1   g15148(.A1(new_n18230_), .A2(new_n14153_), .ZN(new_n18232_));
  NAND2_X1   g15149(.A1(new_n14153_), .A2(new_n18145_), .ZN(new_n18233_));
  XOR2_X1    g15150(.A1(new_n18232_), .A2(new_n18233_), .Z(new_n18234_));
  AOI21_X1   g15151(.A1(new_n18234_), .A2(pi0788), .B(new_n18231_), .ZN(new_n18235_));
  NAND2_X1   g15152(.A1(new_n18163_), .A2(new_n9992_), .ZN(new_n18236_));
  AOI21_X1   g15153(.A1(new_n18236_), .A2(new_n13966_), .B(new_n13919_), .ZN(new_n18237_));
  INV_X1     g15154(.I(new_n18237_), .ZN(new_n18238_));
  NOR2_X1    g15155(.A1(new_n18235_), .A2(new_n18238_), .ZN(new_n18239_));
  NOR2_X1    g15156(.A1(new_n18239_), .A2(new_n16570_), .ZN(new_n18240_));
  XOR2_X1    g15157(.A1(new_n18240_), .A2(new_n16572_), .Z(new_n18241_));
  OAI21_X1   g15158(.A1(new_n16547_), .A2(new_n18239_), .B(new_n18241_), .ZN(new_n18242_));
  INV_X1     g15159(.I(new_n18145_), .ZN(new_n18243_));
  NAND2_X1   g15160(.A1(new_n13993_), .A2(new_n18243_), .ZN(new_n18244_));
  NAND2_X1   g15161(.A1(new_n18235_), .A2(new_n13994_), .ZN(new_n18245_));
  NAND2_X1   g15162(.A1(new_n18245_), .A2(new_n18244_), .ZN(new_n18246_));
  INV_X1     g15163(.I(new_n18246_), .ZN(new_n18247_));
  NOR2_X1    g15164(.A1(new_n18243_), .A2(pi0647), .ZN(new_n18248_));
  NOR2_X1    g15165(.A1(new_n18238_), .A2(new_n14060_), .ZN(new_n18249_));
  AOI21_X1   g15166(.A1(new_n18249_), .A2(pi0647), .B(new_n18248_), .ZN(new_n18250_));
  NAND2_X1   g15167(.A1(new_n18250_), .A2(pi0630), .ZN(new_n18251_));
  NOR2_X1    g15168(.A1(new_n18249_), .A2(new_n14005_), .ZN(new_n18252_));
  XOR2_X1    g15169(.A1(new_n18252_), .A2(new_n14007_), .Z(new_n18253_));
  NAND2_X1   g15170(.A1(new_n18253_), .A2(new_n18145_), .ZN(new_n18254_));
  NOR2_X1    g15171(.A1(new_n18254_), .A2(new_n14012_), .ZN(new_n18255_));
  XOR2_X1    g15172(.A1(new_n18255_), .A2(new_n18251_), .Z(new_n18256_));
  OAI21_X1   g15173(.A1(new_n12776_), .A2(new_n18256_), .B(new_n18247_), .ZN(new_n18257_));
  AOI21_X1   g15174(.A1(new_n18257_), .A2(new_n16576_), .B(new_n16574_), .ZN(new_n18258_));
  AOI21_X1   g15175(.A1(new_n18162_), .A2(new_n14162_), .B(new_n14164_), .ZN(new_n18259_));
  NOR2_X1    g15176(.A1(new_n18259_), .A2(new_n13929_), .ZN(new_n18260_));
  NAND2_X1   g15177(.A1(new_n18259_), .A2(new_n13929_), .ZN(new_n18261_));
  NAND2_X1   g15178(.A1(new_n18261_), .A2(new_n13922_), .ZN(new_n18262_));
  OAI21_X1   g15179(.A1(new_n18260_), .A2(new_n18262_), .B(new_n18234_), .ZN(new_n18263_));
  AOI21_X1   g15180(.A1(new_n18242_), .A2(new_n18258_), .B(new_n18263_), .ZN(new_n18264_));
  NAND2_X1   g15181(.A1(new_n18264_), .A2(new_n18227_), .ZN(new_n18265_));
  AOI21_X1   g15182(.A1(new_n18250_), .A2(pi1157), .B(new_n12776_), .ZN(new_n18266_));
  AOI22_X1   g15183(.A1(new_n18254_), .A2(new_n18266_), .B1(new_n12776_), .B2(new_n18249_), .ZN(new_n18267_));
  NAND2_X1   g15184(.A1(new_n18265_), .A2(pi0644), .ZN(new_n18268_));
  XOR2_X1    g15185(.A1(new_n18268_), .A2(new_n14205_), .Z(new_n18269_));
  NOR2_X1    g15186(.A1(new_n18269_), .A2(new_n18267_), .ZN(new_n18270_));
  NOR2_X1    g15187(.A1(new_n14211_), .A2(new_n18145_), .ZN(new_n18271_));
  AOI21_X1   g15188(.A1(new_n18246_), .A2(new_n14211_), .B(new_n18271_), .ZN(new_n18272_));
  NAND2_X1   g15189(.A1(new_n18272_), .A2(pi0715), .ZN(new_n18273_));
  XOR2_X1    g15190(.A1(new_n18273_), .A2(new_n14205_), .Z(new_n18274_));
  OAI21_X1   g15191(.A1(new_n18274_), .A2(new_n18243_), .B(new_n14203_), .ZN(new_n18275_));
  NAND2_X1   g15192(.A1(new_n18272_), .A2(pi0644), .ZN(new_n18276_));
  XOR2_X1    g15193(.A1(new_n18276_), .A2(new_n14217_), .Z(new_n18277_));
  AOI21_X1   g15194(.A1(new_n18277_), .A2(new_n18145_), .B(pi1160), .ZN(new_n18278_));
  OAI21_X1   g15195(.A1(new_n18270_), .A2(new_n18275_), .B(new_n18278_), .ZN(new_n18279_));
  NAND2_X1   g15196(.A1(new_n18265_), .A2(pi0715), .ZN(new_n18280_));
  XOR2_X1    g15197(.A1(new_n18280_), .A2(new_n14205_), .Z(new_n18281_));
  NOR2_X1    g15198(.A1(new_n18281_), .A2(new_n18267_), .ZN(new_n18282_));
  AOI21_X1   g15199(.A1(new_n18279_), .A2(new_n18282_), .B(new_n14799_), .ZN(new_n18283_));
  XOR2_X1    g15200(.A1(new_n18283_), .A2(new_n14801_), .Z(new_n18284_));
  NOR2_X1    g15201(.A1(new_n18284_), .A2(new_n18265_), .ZN(new_n18285_));
  NOR2_X1    g15202(.A1(new_n14428_), .A2(pi0173), .ZN(new_n18286_));
  NOR2_X1    g15203(.A1(new_n18286_), .A2(new_n13994_), .ZN(new_n18287_));
  NAND2_X1   g15204(.A1(new_n13109_), .A2(new_n10664_), .ZN(new_n18288_));
  NAND2_X1   g15205(.A1(new_n18288_), .A2(pi0038), .ZN(new_n18289_));
  INV_X1     g15206(.I(pi0745), .ZN(new_n18290_));
  NOR4_X1    g15207(.A1(new_n15562_), .A2(new_n10664_), .A3(new_n18290_), .A4(new_n14362_), .ZN(new_n18291_));
  NOR4_X1    g15208(.A1(new_n13107_), .A2(new_n3259_), .A3(new_n10664_), .A4(pi0745), .ZN(new_n18292_));
  OAI21_X1   g15209(.A1(new_n18291_), .A2(new_n13097_), .B(new_n18292_), .ZN(new_n18293_));
  XOR2_X1    g15210(.A1(new_n18293_), .A2(new_n18289_), .Z(new_n18294_));
  NOR2_X1    g15211(.A1(new_n3289_), .A2(pi0173), .ZN(new_n18295_));
  AOI21_X1   g15212(.A1(new_n18294_), .A2(new_n3289_), .B(new_n18295_), .ZN(new_n18296_));
  NAND2_X1   g15213(.A1(new_n18296_), .A2(new_n13776_), .ZN(new_n18297_));
  OAI21_X1   g15214(.A1(new_n15147_), .A2(new_n18286_), .B(new_n18297_), .ZN(new_n18298_));
  NAND2_X1   g15215(.A1(new_n18298_), .A2(pi0609), .ZN(new_n18299_));
  NAND2_X1   g15216(.A1(new_n18299_), .A2(pi0785), .ZN(new_n18300_));
  INV_X1     g15217(.I(new_n18296_), .ZN(new_n18301_));
  INV_X1     g15218(.I(new_n18286_), .ZN(new_n18302_));
  NOR2_X1    g15219(.A1(new_n18302_), .A2(new_n13776_), .ZN(new_n18303_));
  AOI21_X1   g15220(.A1(new_n18301_), .A2(new_n13776_), .B(new_n18303_), .ZN(new_n18304_));
  AOI21_X1   g15221(.A1(new_n18302_), .A2(new_n14467_), .B(pi0609), .ZN(new_n18305_));
  NOR2_X1    g15222(.A1(new_n18297_), .A2(new_n18305_), .ZN(new_n18306_));
  INV_X1     g15223(.I(new_n18306_), .ZN(new_n18307_));
  NOR3_X1    g15224(.A1(new_n18307_), .A2(new_n13801_), .A3(new_n18304_), .ZN(new_n18308_));
  XOR2_X1    g15225(.A1(new_n18300_), .A2(new_n18308_), .Z(new_n18309_));
  NOR2_X1    g15226(.A1(new_n18309_), .A2(pi0781), .ZN(new_n18310_));
  XNOR2_X1   g15227(.A1(new_n18300_), .A2(new_n18308_), .ZN(new_n18311_));
  NAND3_X1   g15228(.A1(new_n18311_), .A2(new_n16689_), .A3(new_n18286_), .ZN(new_n18312_));
  NAND3_X1   g15229(.A1(new_n18309_), .A2(new_n16689_), .A3(new_n18302_), .ZN(new_n18313_));
  NAND2_X1   g15230(.A1(new_n18312_), .A2(new_n18313_), .ZN(new_n18314_));
  AOI21_X1   g15231(.A1(new_n18314_), .A2(pi0781), .B(new_n18310_), .ZN(new_n18315_));
  NOR2_X1    g15232(.A1(new_n18315_), .A2(pi0789), .ZN(new_n18316_));
  NAND2_X1   g15233(.A1(new_n18315_), .A2(new_n16697_), .ZN(new_n18317_));
  NAND2_X1   g15234(.A1(new_n18286_), .A2(new_n16697_), .ZN(new_n18318_));
  XOR2_X1    g15235(.A1(new_n18317_), .A2(new_n18318_), .Z(new_n18319_));
  AOI21_X1   g15236(.A1(new_n18319_), .A2(pi0789), .B(new_n18316_), .ZN(new_n18320_));
  NOR2_X1    g15237(.A1(new_n18320_), .A2(pi0788), .ZN(new_n18321_));
  OR3_X2     g15238(.A1(new_n18320_), .A2(new_n14141_), .A3(new_n18302_), .Z(new_n18322_));
  NAND3_X1   g15239(.A1(new_n18320_), .A2(new_n14153_), .A3(new_n18302_), .ZN(new_n18323_));
  AOI21_X1   g15240(.A1(new_n18322_), .A2(new_n18323_), .B(new_n13937_), .ZN(new_n18324_));
  NOR3_X1    g15241(.A1(new_n18324_), .A2(new_n18321_), .A3(new_n13993_), .ZN(new_n18325_));
  OAI21_X1   g15242(.A1(new_n18325_), .A2(new_n18287_), .B(new_n14211_), .ZN(new_n18326_));
  NOR2_X1    g15243(.A1(new_n18286_), .A2(new_n14211_), .ZN(new_n18327_));
  INV_X1     g15244(.I(new_n18327_), .ZN(new_n18328_));
  AOI21_X1   g15245(.A1(new_n18302_), .A2(new_n14254_), .B(pi0644), .ZN(new_n18329_));
  AOI21_X1   g15246(.A1(new_n18326_), .A2(new_n18328_), .B(new_n18329_), .ZN(new_n18330_));
  INV_X1     g15247(.I(new_n18330_), .ZN(new_n18331_));
  NAND2_X1   g15248(.A1(new_n18288_), .A2(new_n13720_), .ZN(new_n18332_));
  NAND2_X1   g15249(.A1(new_n16715_), .A2(new_n10664_), .ZN(new_n18333_));
  NAND4_X1   g15250(.A1(new_n15655_), .A2(new_n17227_), .A3(new_n18332_), .A4(new_n18333_), .ZN(new_n18334_));
  AOI21_X1   g15251(.A1(new_n18334_), .A2(new_n14424_), .B(new_n10664_), .ZN(new_n18335_));
  NAND2_X1   g15252(.A1(new_n18286_), .A2(new_n18335_), .ZN(new_n18336_));
  NAND2_X1   g15253(.A1(new_n18336_), .A2(new_n3290_), .ZN(new_n18337_));
  NAND2_X1   g15254(.A1(new_n18337_), .A2(pi0723), .ZN(new_n18338_));
  NAND2_X1   g15255(.A1(new_n18338_), .A2(pi0625), .ZN(new_n18339_));
  XOR2_X1    g15256(.A1(new_n18339_), .A2(new_n13620_), .Z(new_n18340_));
  NAND2_X1   g15257(.A1(new_n18340_), .A2(new_n18286_), .ZN(new_n18341_));
  NAND2_X1   g15258(.A1(new_n18341_), .A2(pi0778), .ZN(new_n18342_));
  NAND2_X1   g15259(.A1(new_n18338_), .A2(pi1153), .ZN(new_n18343_));
  XOR2_X1    g15260(.A1(new_n18343_), .A2(new_n13620_), .Z(new_n18344_));
  NAND2_X1   g15261(.A1(new_n18344_), .A2(new_n18286_), .ZN(new_n18345_));
  NOR3_X1    g15262(.A1(new_n18345_), .A2(new_n13748_), .A3(new_n18338_), .ZN(new_n18346_));
  XNOR2_X1   g15263(.A1(new_n18346_), .A2(new_n18342_), .ZN(new_n18347_));
  INV_X1     g15264(.I(new_n18347_), .ZN(new_n18348_));
  INV_X1     g15265(.I(new_n18294_), .ZN(new_n18349_));
  NOR2_X1    g15266(.A1(new_n10664_), .A2(new_n18290_), .ZN(new_n18350_));
  NOR2_X1    g15267(.A1(new_n13453_), .A2(new_n10664_), .ZN(new_n18351_));
  XOR2_X1    g15268(.A1(new_n18351_), .A2(new_n18350_), .Z(new_n18352_));
  NAND2_X1   g15269(.A1(new_n18352_), .A2(new_n13521_), .ZN(new_n18353_));
  NAND3_X1   g15270(.A1(new_n14270_), .A2(pi0173), .A3(pi0745), .ZN(new_n18354_));
  NAND3_X1   g15271(.A1(new_n14272_), .A2(new_n10664_), .A3(pi0745), .ZN(new_n18355_));
  AOI21_X1   g15272(.A1(new_n18354_), .A2(new_n18355_), .B(new_n13152_), .ZN(new_n18356_));
  NAND3_X1   g15273(.A1(new_n13198_), .A2(pi0173), .A3(pi0745), .ZN(new_n18357_));
  NAND3_X1   g15274(.A1(new_n13200_), .A2(pi0173), .A3(new_n18290_), .ZN(new_n18358_));
  AOI21_X1   g15275(.A1(new_n18358_), .A2(new_n18357_), .B(new_n13191_), .ZN(new_n18359_));
  OAI21_X1   g15276(.A1(new_n18356_), .A2(new_n3262_), .B(new_n18359_), .ZN(new_n18360_));
  NAND3_X1   g15277(.A1(new_n18353_), .A2(new_n3183_), .A3(new_n18360_), .ZN(new_n18361_));
  NOR2_X1    g15278(.A1(new_n14284_), .A2(new_n18290_), .ZN(new_n18362_));
  XOR2_X1    g15279(.A1(new_n18362_), .A2(new_n18350_), .Z(new_n18363_));
  NAND3_X1   g15280(.A1(new_n18361_), .A2(new_n18363_), .A3(new_n13359_), .ZN(new_n18364_));
  NAND3_X1   g15281(.A1(new_n18364_), .A2(new_n17227_), .A3(new_n3290_), .ZN(new_n18365_));
  OAI21_X1   g15282(.A1(new_n15587_), .A2(new_n10664_), .B(new_n18290_), .ZN(new_n18366_));
  NAND2_X1   g15283(.A1(new_n18366_), .A2(new_n13209_), .ZN(new_n18367_));
  NAND2_X1   g15284(.A1(new_n18180_), .A2(new_n16751_), .ZN(new_n18368_));
  NAND4_X1   g15285(.A1(new_n5503_), .A2(new_n18368_), .A3(pi0173), .A4(new_n3290_), .ZN(new_n18369_));
  AOI21_X1   g15286(.A1(new_n18367_), .A2(new_n3259_), .B(new_n18369_), .ZN(new_n18370_));
  NAND2_X1   g15287(.A1(new_n18365_), .A2(new_n18370_), .ZN(new_n18371_));
  AOI21_X1   g15288(.A1(new_n18371_), .A2(new_n17227_), .B(new_n18349_), .ZN(new_n18372_));
  NAND3_X1   g15289(.A1(new_n18372_), .A2(pi0625), .A3(pi1153), .ZN(new_n18373_));
  NOR2_X1    g15290(.A1(new_n18372_), .A2(new_n13613_), .ZN(new_n18374_));
  NAND2_X1   g15291(.A1(new_n18374_), .A2(new_n13620_), .ZN(new_n18375_));
  NAND2_X1   g15292(.A1(new_n18375_), .A2(new_n18373_), .ZN(new_n18376_));
  NAND2_X1   g15293(.A1(new_n18345_), .A2(new_n14081_), .ZN(new_n18377_));
  AOI21_X1   g15294(.A1(new_n18376_), .A2(new_n18301_), .B(new_n18377_), .ZN(new_n18378_));
  NOR2_X1    g15295(.A1(new_n18372_), .A2(new_n13614_), .ZN(new_n18379_));
  NOR2_X1    g15296(.A1(new_n18379_), .A2(new_n13620_), .ZN(new_n18380_));
  NOR3_X1    g15297(.A1(new_n18372_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n18381_));
  OAI21_X1   g15298(.A1(new_n18380_), .A2(new_n18381_), .B(new_n18301_), .ZN(new_n18382_));
  NAND2_X1   g15299(.A1(new_n18382_), .A2(new_n14081_), .ZN(new_n18383_));
  NOR2_X1    g15300(.A1(new_n18341_), .A2(new_n13748_), .ZN(new_n18384_));
  OAI21_X1   g15301(.A1(new_n18383_), .A2(new_n18378_), .B(new_n18384_), .ZN(new_n18385_));
  NOR2_X1    g15302(.A1(new_n18372_), .A2(pi0778), .ZN(new_n18386_));
  INV_X1     g15303(.I(new_n18386_), .ZN(new_n18387_));
  NAND2_X1   g15304(.A1(new_n18385_), .A2(new_n18387_), .ZN(new_n18388_));
  NAND3_X1   g15305(.A1(new_n18388_), .A2(pi0609), .A3(pi1155), .ZN(new_n18389_));
  NAND4_X1   g15306(.A1(new_n18385_), .A2(new_n13766_), .A3(pi1155), .A4(new_n18387_), .ZN(new_n18390_));
  AOI21_X1   g15307(.A1(new_n18389_), .A2(new_n18390_), .B(new_n18348_), .ZN(new_n18391_));
  NAND2_X1   g15308(.A1(new_n18299_), .A2(pi0660), .ZN(new_n18392_));
  OAI21_X1   g15309(.A1(new_n18391_), .A2(new_n18392_), .B(pi0785), .ZN(new_n18393_));
  NAND3_X1   g15310(.A1(new_n18385_), .A2(pi0609), .A3(new_n18387_), .ZN(new_n18394_));
  XOR2_X1    g15311(.A1(new_n18394_), .A2(new_n14694_), .Z(new_n18395_));
  NAND3_X1   g15312(.A1(new_n18388_), .A2(new_n16780_), .A3(new_n18307_), .ZN(new_n18396_));
  AOI21_X1   g15313(.A1(new_n18395_), .A2(new_n18347_), .B(new_n18396_), .ZN(new_n18397_));
  NAND2_X1   g15314(.A1(new_n18397_), .A2(new_n18393_), .ZN(new_n18398_));
  INV_X1     g15315(.I(new_n18398_), .ZN(new_n18399_));
  NOR2_X1    g15316(.A1(new_n18397_), .A2(new_n18393_), .ZN(new_n18400_));
  NOR2_X1    g15317(.A1(new_n18302_), .A2(new_n13805_), .ZN(new_n18401_));
  AOI21_X1   g15318(.A1(new_n18347_), .A2(new_n13805_), .B(new_n18401_), .ZN(new_n18402_));
  OAI21_X1   g15319(.A1(new_n18302_), .A2(new_n13816_), .B(new_n13877_), .ZN(new_n18403_));
  AOI21_X1   g15320(.A1(new_n18309_), .A2(new_n18403_), .B(new_n13819_), .ZN(new_n18404_));
  AOI21_X1   g15321(.A1(new_n18402_), .A2(new_n18404_), .B(pi0618), .ZN(new_n18405_));
  INV_X1     g15322(.I(new_n18405_), .ZN(new_n18406_));
  OAI21_X1   g15323(.A1(new_n18399_), .A2(new_n18400_), .B(new_n18406_), .ZN(new_n18407_));
  AOI21_X1   g15324(.A1(new_n18302_), .A2(new_n13824_), .B(pi0618), .ZN(new_n18408_));
  NOR3_X1    g15325(.A1(new_n18309_), .A2(pi1154), .A3(new_n18408_), .ZN(new_n18409_));
  OAI21_X1   g15326(.A1(new_n18402_), .A2(new_n13816_), .B(new_n18409_), .ZN(new_n18410_));
  INV_X1     g15327(.I(new_n18410_), .ZN(new_n18411_));
  NOR2_X1    g15328(.A1(new_n18411_), .A2(pi0618), .ZN(new_n18412_));
  NOR2_X1    g15329(.A1(new_n18412_), .A2(new_n13855_), .ZN(new_n18413_));
  OAI21_X1   g15330(.A1(new_n18399_), .A2(new_n18400_), .B(new_n18413_), .ZN(new_n18414_));
  AOI21_X1   g15331(.A1(pi0781), .A2(new_n18407_), .B(new_n18414_), .ZN(new_n18415_));
  INV_X1     g15332(.I(new_n18400_), .ZN(new_n18416_));
  AOI21_X1   g15333(.A1(new_n18416_), .A2(new_n18398_), .B(new_n18405_), .ZN(new_n18417_));
  INV_X1     g15334(.I(new_n18413_), .ZN(new_n18418_));
  AOI21_X1   g15335(.A1(new_n18416_), .A2(new_n18398_), .B(new_n18418_), .ZN(new_n18419_));
  NOR3_X1    g15336(.A1(new_n18417_), .A2(new_n18419_), .A3(new_n13855_), .ZN(new_n18420_));
  OAI21_X1   g15337(.A1(new_n18415_), .A2(new_n18420_), .B(new_n13896_), .ZN(new_n18421_));
  NAND2_X1   g15338(.A1(new_n18421_), .A2(new_n14143_), .ZN(new_n18422_));
  OAI21_X1   g15339(.A1(new_n13855_), .A2(new_n18417_), .B(new_n18419_), .ZN(new_n18423_));
  NAND3_X1   g15340(.A1(new_n18407_), .A2(new_n18414_), .A3(pi0781), .ZN(new_n18424_));
  NAND2_X1   g15341(.A1(new_n18423_), .A2(new_n18424_), .ZN(new_n18425_));
  INV_X1     g15342(.I(new_n18402_), .ZN(new_n18426_));
  NOR2_X1    g15343(.A1(new_n18426_), .A2(new_n13879_), .ZN(new_n18427_));
  AOI21_X1   g15344(.A1(new_n13879_), .A2(new_n18302_), .B(new_n18427_), .ZN(new_n18428_));
  INV_X1     g15345(.I(new_n18428_), .ZN(new_n18429_));
  NOR2_X1    g15346(.A1(new_n18429_), .A2(new_n13860_), .ZN(new_n18430_));
  AOI21_X1   g15347(.A1(new_n18302_), .A2(new_n13885_), .B(pi0619), .ZN(new_n18431_));
  OR3_X2     g15348(.A1(new_n18315_), .A2(pi1159), .A3(new_n18431_), .Z(new_n18432_));
  OAI21_X1   g15349(.A1(new_n18430_), .A2(new_n18432_), .B(new_n13860_), .ZN(new_n18433_));
  AOI21_X1   g15350(.A1(new_n18425_), .A2(new_n18433_), .B(pi0789), .ZN(new_n18434_));
  OAI21_X1   g15351(.A1(new_n18302_), .A2(new_n13860_), .B(new_n13916_), .ZN(new_n18435_));
  AOI21_X1   g15352(.A1(new_n18315_), .A2(new_n18435_), .B(new_n13904_), .ZN(new_n18436_));
  AOI21_X1   g15353(.A1(new_n18429_), .A2(new_n18436_), .B(pi0619), .ZN(new_n18437_));
  AOI21_X1   g15354(.A1(new_n18423_), .A2(new_n18424_), .B(new_n18437_), .ZN(new_n18438_));
  INV_X1     g15355(.I(new_n18438_), .ZN(new_n18439_));
  AOI21_X1   g15356(.A1(new_n18422_), .A2(new_n18434_), .B(new_n18439_), .ZN(new_n18440_));
  INV_X1     g15357(.I(new_n18324_), .ZN(new_n18441_));
  NAND2_X1   g15358(.A1(new_n18428_), .A2(new_n16639_), .ZN(new_n18442_));
  XOR2_X1    g15359(.A1(new_n18442_), .A2(new_n16829_), .Z(new_n18443_));
  NAND2_X1   g15360(.A1(new_n18443_), .A2(new_n18286_), .ZN(new_n18444_));
  OAI21_X1   g15361(.A1(new_n18444_), .A2(pi1158), .B(new_n13922_), .ZN(new_n18445_));
  AOI21_X1   g15362(.A1(pi1158), .A2(new_n18444_), .B(new_n18445_), .ZN(new_n18446_));
  NOR2_X1    g15363(.A1(new_n18446_), .A2(new_n18441_), .ZN(new_n18447_));
  OAI21_X1   g15364(.A1(new_n18440_), .A2(new_n16423_), .B(new_n18447_), .ZN(new_n18448_));
  NOR2_X1    g15365(.A1(new_n18325_), .A2(new_n18287_), .ZN(new_n18449_));
  INV_X1     g15366(.I(new_n18449_), .ZN(new_n18450_));
  NAND4_X1   g15367(.A1(new_n18402_), .A2(new_n13880_), .A3(new_n15395_), .A4(new_n18286_), .ZN(new_n18451_));
  NOR4_X1    g15368(.A1(new_n18402_), .A2(new_n13879_), .A3(new_n16839_), .A4(new_n18286_), .ZN(new_n18452_));
  INV_X1     g15369(.I(new_n18452_), .ZN(new_n18453_));
  NAND2_X1   g15370(.A1(new_n18453_), .A2(new_n18451_), .ZN(new_n18454_));
  NAND3_X1   g15371(.A1(new_n18454_), .A2(pi0628), .A3(pi1156), .ZN(new_n18455_));
  NOR3_X1    g15372(.A1(new_n18454_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n18456_));
  INV_X1     g15373(.I(new_n18456_), .ZN(new_n18457_));
  AOI21_X1   g15374(.A1(new_n18457_), .A2(new_n18455_), .B(new_n18302_), .ZN(new_n18458_));
  NAND3_X1   g15375(.A1(new_n18454_), .A2(pi0628), .A3(pi1156), .ZN(new_n18459_));
  NAND4_X1   g15376(.A1(new_n18453_), .A2(new_n13942_), .A3(pi1156), .A4(new_n18451_), .ZN(new_n18460_));
  AOI21_X1   g15377(.A1(new_n18459_), .A2(new_n18460_), .B(new_n18302_), .ZN(new_n18461_));
  NAND4_X1   g15378(.A1(new_n18458_), .A2(pi0792), .A3(new_n18454_), .A4(new_n18461_), .ZN(new_n18462_));
  INV_X1     g15379(.I(new_n18455_), .ZN(new_n18463_));
  OAI21_X1   g15380(.A1(new_n18463_), .A2(new_n18456_), .B(new_n18286_), .ZN(new_n18464_));
  NAND3_X1   g15381(.A1(new_n18461_), .A2(pi0792), .A3(new_n18454_), .ZN(new_n18465_));
  NAND3_X1   g15382(.A1(new_n18465_), .A2(pi0792), .A3(new_n18464_), .ZN(new_n18466_));
  AOI21_X1   g15383(.A1(new_n18466_), .A2(new_n18462_), .B(pi0647), .ZN(new_n18467_));
  NOR2_X1    g15384(.A1(new_n18302_), .A2(new_n14005_), .ZN(new_n18468_));
  OAI21_X1   g15385(.A1(new_n18467_), .A2(new_n18468_), .B(new_n14011_), .ZN(new_n18469_));
  NAND2_X1   g15386(.A1(new_n18466_), .A2(new_n18462_), .ZN(new_n18470_));
  AOI21_X1   g15387(.A1(new_n18286_), .A2(new_n14005_), .B(new_n14006_), .ZN(new_n18471_));
  INV_X1     g15388(.I(new_n18471_), .ZN(new_n18472_));
  AOI21_X1   g15389(.A1(new_n18470_), .A2(pi0647), .B(new_n18472_), .ZN(new_n18473_));
  NAND3_X1   g15390(.A1(new_n18469_), .A2(new_n18473_), .A3(new_n14010_), .ZN(new_n18474_));
  NOR2_X1    g15391(.A1(new_n18467_), .A2(new_n18468_), .ZN(new_n18475_));
  NOR3_X1    g15392(.A1(new_n18475_), .A2(new_n14010_), .A3(new_n14006_), .ZN(new_n18476_));
  INV_X1     g15393(.I(new_n18476_), .ZN(new_n18477_));
  AOI21_X1   g15394(.A1(new_n18477_), .A2(new_n18474_), .B(new_n12776_), .ZN(new_n18478_));
  OAI21_X1   g15395(.A1(new_n18478_), .A2(new_n18450_), .B(new_n16868_), .ZN(new_n18479_));
  NAND2_X1   g15396(.A1(new_n18479_), .A2(new_n18448_), .ZN(new_n18480_));
  INV_X1     g15397(.I(new_n18321_), .ZN(new_n18481_));
  NOR2_X1    g15398(.A1(new_n18458_), .A2(new_n13976_), .ZN(new_n18482_));
  NOR2_X1    g15399(.A1(new_n18461_), .A2(pi0629), .ZN(new_n18483_));
  OAI21_X1   g15400(.A1(new_n18482_), .A2(new_n18483_), .B(pi0792), .ZN(new_n18484_));
  AOI22_X1   g15401(.A1(new_n18441_), .A2(new_n18481_), .B1(new_n16875_), .B2(new_n18484_), .ZN(new_n18485_));
  NAND3_X1   g15402(.A1(new_n18480_), .A2(pi0790), .A3(new_n18485_), .ZN(new_n18486_));
  AOI21_X1   g15403(.A1(new_n18486_), .A2(new_n14204_), .B(new_n18331_), .ZN(new_n18487_));
  NAND4_X1   g15404(.A1(new_n18480_), .A2(pi0644), .A3(pi0715), .A4(new_n18485_), .ZN(new_n18488_));
  AOI21_X1   g15405(.A1(new_n18425_), .A2(new_n13896_), .B(new_n15479_), .ZN(new_n18489_));
  OAI21_X1   g15406(.A1(new_n18415_), .A2(new_n18420_), .B(new_n18433_), .ZN(new_n18490_));
  NAND2_X1   g15407(.A1(new_n18490_), .A2(new_n13896_), .ZN(new_n18491_));
  OAI21_X1   g15408(.A1(new_n18491_), .A2(new_n18489_), .B(new_n18438_), .ZN(new_n18492_));
  INV_X1     g15409(.I(new_n18447_), .ZN(new_n18493_));
  AOI21_X1   g15410(.A1(new_n18492_), .A2(new_n16424_), .B(new_n18493_), .ZN(new_n18494_));
  INV_X1     g15411(.I(new_n18474_), .ZN(new_n18495_));
  OAI21_X1   g15412(.A1(new_n18495_), .A2(new_n18476_), .B(pi0787), .ZN(new_n18496_));
  AOI21_X1   g15413(.A1(new_n18496_), .A2(new_n18449_), .B(new_n16891_), .ZN(new_n18497_));
  OAI21_X1   g15414(.A1(new_n18497_), .A2(new_n18494_), .B(new_n18485_), .ZN(new_n18498_));
  NAND3_X1   g15415(.A1(new_n18498_), .A2(pi0644), .A3(new_n14200_), .ZN(new_n18499_));
  AOI21_X1   g15416(.A1(new_n14006_), .A2(new_n18475_), .B(new_n18473_), .ZN(new_n18500_));
  NOR2_X1    g15417(.A1(new_n18500_), .A2(new_n12776_), .ZN(new_n18501_));
  NOR2_X1    g15418(.A1(new_n18470_), .A2(pi0787), .ZN(new_n18502_));
  AOI21_X1   g15419(.A1(new_n18450_), .A2(new_n14211_), .B(new_n18327_), .ZN(new_n18503_));
  NOR2_X1    g15420(.A1(new_n14243_), .A2(pi0644), .ZN(new_n18504_));
  AOI21_X1   g15421(.A1(new_n18330_), .A2(pi0715), .B(pi0644), .ZN(new_n18505_));
  OAI21_X1   g15422(.A1(new_n18501_), .A2(new_n18502_), .B(pi0790), .ZN(new_n18506_));
  OAI22_X1   g15423(.A1(new_n18506_), .A2(new_n18505_), .B1(new_n18503_), .B2(new_n18504_), .ZN(new_n18507_));
  OAI21_X1   g15424(.A1(new_n18501_), .A2(new_n18502_), .B(new_n18507_), .ZN(new_n18508_));
  AOI21_X1   g15425(.A1(new_n18499_), .A2(new_n18488_), .B(new_n18508_), .ZN(new_n18509_));
  OAI21_X1   g15426(.A1(new_n18509_), .A2(new_n18487_), .B(new_n7240_), .ZN(new_n18510_));
  AOI21_X1   g15427(.A1(po1038), .A2(new_n10664_), .B(pi0832), .ZN(new_n18511_));
  AOI21_X1   g15428(.A1(new_n18510_), .A2(new_n18511_), .B(new_n18285_), .ZN(po0330));
  NOR3_X1    g15429(.A1(new_n13085_), .A2(new_n16088_), .A3(new_n17309_), .ZN(new_n18513_));
  NOR3_X1    g15430(.A1(new_n12977_), .A2(new_n16086_), .A3(new_n17309_), .ZN(new_n18514_));
  NAND3_X1   g15431(.A1(new_n14356_), .A2(pi0039), .A3(pi0759), .ZN(new_n18515_));
  NAND3_X1   g15432(.A1(new_n14338_), .A2(new_n3183_), .A3(pi0759), .ZN(new_n18516_));
  NAND2_X1   g15433(.A1(new_n14874_), .A2(pi0174), .ZN(new_n18517_));
  AOI21_X1   g15434(.A1(new_n18515_), .A2(new_n18516_), .B(new_n18517_), .ZN(new_n18518_));
  OAI22_X1   g15435(.A1(new_n18514_), .A2(new_n18513_), .B1(pi0039), .B2(new_n18518_), .ZN(new_n18519_));
  AOI21_X1   g15436(.A1(new_n13203_), .A2(pi0759), .B(new_n3259_), .ZN(new_n18520_));
  XOR2_X1    g15437(.A1(new_n13723_), .A2(new_n18520_), .Z(new_n18521_));
  NAND2_X1   g15438(.A1(new_n18521_), .A2(pi0174), .ZN(new_n18522_));
  OAI21_X1   g15439(.A1(new_n3259_), .A2(new_n18522_), .B(new_n18519_), .ZN(new_n18523_));
  NAND4_X1   g15440(.A1(new_n18523_), .A2(new_n7378_), .A3(pi0759), .A4(new_n16114_), .ZN(new_n18524_));
  NOR2_X1    g15441(.A1(new_n18524_), .A2(new_n3290_), .ZN(new_n18525_));
  NOR2_X1    g15442(.A1(new_n3289_), .A2(pi0174), .ZN(new_n18526_));
  OR2_X2     g15443(.A1(new_n18525_), .A2(new_n18526_), .Z(new_n18527_));
  NAND3_X1   g15444(.A1(new_n14270_), .A2(pi0174), .A3(pi0759), .ZN(new_n18528_));
  NAND3_X1   g15445(.A1(new_n14272_), .A2(pi0174), .A3(new_n17309_), .ZN(new_n18529_));
  NAND2_X1   g15446(.A1(new_n18529_), .A2(new_n18528_), .ZN(new_n18530_));
  AOI21_X1   g15447(.A1(new_n14269_), .A2(new_n18530_), .B(new_n3212_), .ZN(new_n18531_));
  NOR3_X1    g15448(.A1(new_n13200_), .A2(new_n7378_), .A3(new_n17309_), .ZN(new_n18532_));
  NOR3_X1    g15449(.A1(new_n13198_), .A2(pi0174), .A3(new_n17309_), .ZN(new_n18533_));
  OAI21_X1   g15450(.A1(new_n18532_), .A2(new_n18533_), .B(new_n13190_), .ZN(new_n18534_));
  NOR2_X1    g15451(.A1(new_n3290_), .A2(new_n17327_), .ZN(new_n18535_));
  NAND3_X1   g15452(.A1(new_n18522_), .A2(new_n15630_), .A3(new_n18535_), .ZN(new_n18536_));
  OAI21_X1   g15453(.A1(new_n18531_), .A2(new_n18534_), .B(new_n18536_), .ZN(new_n18537_));
  INV_X1     g15454(.I(new_n13359_), .ZN(new_n18538_));
  NAND4_X1   g15455(.A1(new_n18537_), .A2(pi0174), .A3(new_n3290_), .A4(new_n14284_), .ZN(new_n18544_));
  AOI21_X1   g15456(.A1(new_n18544_), .A2(new_n18524_), .B(new_n17327_), .ZN(new_n18545_));
  NAND3_X1   g15457(.A1(new_n18545_), .A2(pi0625), .A3(pi1153), .ZN(new_n18546_));
  INV_X1     g15458(.I(new_n18545_), .ZN(new_n18547_));
  NAND3_X1   g15459(.A1(new_n18547_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n18548_));
  NAND2_X1   g15460(.A1(new_n18548_), .A2(new_n18546_), .ZN(new_n18549_));
  NAND3_X1   g15461(.A1(new_n14422_), .A2(pi0038), .A3(pi0174), .ZN(new_n18550_));
  NAND3_X1   g15462(.A1(new_n14424_), .A2(new_n3259_), .A3(pi0174), .ZN(new_n18551_));
  AOI21_X1   g15463(.A1(new_n18551_), .A2(new_n18550_), .B(new_n14404_), .ZN(new_n18552_));
  OAI21_X1   g15464(.A1(new_n16149_), .A2(new_n7378_), .B(new_n18535_), .ZN(new_n18553_));
  NOR2_X1    g15465(.A1(new_n18552_), .A2(new_n18553_), .ZN(new_n18554_));
  NOR2_X1    g15466(.A1(new_n18554_), .A2(pi0174), .ZN(new_n18555_));
  NOR2_X1    g15467(.A1(new_n18555_), .A2(new_n13627_), .ZN(new_n18556_));
  NOR2_X1    g15468(.A1(new_n14428_), .A2(new_n7378_), .ZN(new_n18557_));
  NOR2_X1    g15469(.A1(new_n18557_), .A2(new_n13613_), .ZN(new_n18558_));
  XOR2_X1    g15470(.A1(new_n18558_), .A2(new_n13615_), .Z(new_n18559_));
  NAND2_X1   g15471(.A1(new_n18559_), .A2(new_n18556_), .ZN(new_n18560_));
  NAND2_X1   g15472(.A1(new_n18560_), .A2(pi0608), .ZN(new_n18561_));
  AOI21_X1   g15473(.A1(new_n18549_), .A2(new_n18527_), .B(new_n18561_), .ZN(new_n18562_));
  NOR2_X1    g15474(.A1(new_n18562_), .A2(new_n13748_), .ZN(new_n18563_));
  INV_X1     g15475(.I(new_n18527_), .ZN(new_n18564_));
  NAND3_X1   g15476(.A1(new_n18545_), .A2(pi0625), .A3(pi1153), .ZN(new_n18565_));
  NAND3_X1   g15477(.A1(new_n18547_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n18566_));
  AOI21_X1   g15478(.A1(new_n18566_), .A2(new_n18565_), .B(new_n18564_), .ZN(new_n18567_));
  NOR2_X1    g15479(.A1(new_n18557_), .A2(new_n13614_), .ZN(new_n18568_));
  XOR2_X1    g15480(.A1(new_n18568_), .A2(new_n13615_), .Z(new_n18569_));
  AND2_X2    g15481(.A1(new_n18569_), .A2(new_n18556_), .Z(new_n18570_));
  NOR4_X1    g15482(.A1(new_n18567_), .A2(new_n13750_), .A3(new_n18547_), .A4(new_n18570_), .ZN(new_n18571_));
  XOR2_X1    g15483(.A1(new_n18563_), .A2(new_n18571_), .Z(new_n18572_));
  INV_X1     g15484(.I(new_n18572_), .ZN(new_n18573_));
  NAND2_X1   g15485(.A1(new_n18560_), .A2(pi0778), .ZN(new_n18574_));
  NAND3_X1   g15486(.A1(new_n18569_), .A2(pi0778), .A3(new_n18556_), .ZN(new_n18575_));
  XNOR2_X1   g15487(.A1(new_n18574_), .A2(new_n18575_), .ZN(new_n18576_));
  INV_X1     g15488(.I(new_n18557_), .ZN(new_n18577_));
  NAND2_X1   g15489(.A1(new_n18557_), .A2(new_n13775_), .ZN(new_n18578_));
  OAI21_X1   g15490(.A1(new_n18527_), .A2(new_n13775_), .B(new_n18578_), .ZN(new_n18579_));
  NAND3_X1   g15491(.A1(new_n18579_), .A2(pi0609), .A3(pi1155), .ZN(new_n18580_));
  INV_X1     g15492(.I(new_n18579_), .ZN(new_n18581_));
  NAND3_X1   g15493(.A1(new_n18581_), .A2(pi0609), .A3(new_n14694_), .ZN(new_n18582_));
  AOI21_X1   g15494(.A1(new_n18582_), .A2(new_n18580_), .B(new_n18577_), .ZN(new_n18583_));
  NOR2_X1    g15495(.A1(new_n18583_), .A2(new_n13785_), .ZN(new_n18584_));
  AOI21_X1   g15496(.A1(new_n18584_), .A2(new_n18576_), .B(pi0609), .ZN(new_n18585_));
  OAI21_X1   g15497(.A1(new_n18573_), .A2(new_n18585_), .B(pi0785), .ZN(new_n18586_));
  NOR2_X1    g15498(.A1(new_n18576_), .A2(new_n13766_), .ZN(new_n18587_));
  NAND3_X1   g15499(.A1(new_n18579_), .A2(pi0609), .A3(pi1155), .ZN(new_n18588_));
  INV_X1     g15500(.I(new_n18588_), .ZN(new_n18589_));
  NOR3_X1    g15501(.A1(new_n18579_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n18590_));
  OAI21_X1   g15502(.A1(new_n18589_), .A2(new_n18590_), .B(new_n18557_), .ZN(new_n18591_));
  NAND2_X1   g15503(.A1(new_n18591_), .A2(new_n13793_), .ZN(new_n18592_));
  OAI21_X1   g15504(.A1(new_n18587_), .A2(new_n18592_), .B(new_n13766_), .ZN(new_n18593_));
  NAND3_X1   g15505(.A1(new_n18572_), .A2(new_n18593_), .A3(pi0785), .ZN(new_n18594_));
  XNOR2_X1   g15506(.A1(new_n18586_), .A2(new_n18594_), .ZN(new_n18595_));
  INV_X1     g15507(.I(new_n18590_), .ZN(new_n18596_));
  AOI21_X1   g15508(.A1(new_n18596_), .A2(new_n18588_), .B(new_n18577_), .ZN(new_n18597_));
  NAND4_X1   g15509(.A1(new_n18597_), .A2(new_n18583_), .A3(pi0785), .A4(new_n18579_), .ZN(new_n18598_));
  INV_X1     g15510(.I(new_n18598_), .ZN(new_n18599_));
  NOR3_X1    g15511(.A1(new_n18591_), .A2(new_n13801_), .A3(new_n18581_), .ZN(new_n18600_));
  NOR3_X1    g15512(.A1(new_n18600_), .A2(new_n13801_), .A3(new_n18583_), .ZN(new_n18601_));
  NOR2_X1    g15513(.A1(new_n18601_), .A2(new_n18599_), .ZN(new_n18602_));
  AOI21_X1   g15514(.A1(new_n18602_), .A2(pi0618), .B(new_n13819_), .ZN(new_n18603_));
  NOR2_X1    g15515(.A1(new_n18583_), .A2(new_n13801_), .ZN(new_n18604_));
  NOR2_X1    g15516(.A1(new_n18581_), .A2(new_n13801_), .ZN(new_n18605_));
  NAND2_X1   g15517(.A1(new_n18597_), .A2(new_n18605_), .ZN(new_n18606_));
  NAND2_X1   g15518(.A1(new_n18606_), .A2(new_n18604_), .ZN(new_n18607_));
  NAND2_X1   g15519(.A1(new_n18607_), .A2(new_n18598_), .ZN(new_n18608_));
  NOR3_X1    g15520(.A1(new_n18608_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n18609_));
  OAI21_X1   g15521(.A1(new_n18603_), .A2(new_n18609_), .B(new_n18557_), .ZN(new_n18610_));
  NOR2_X1    g15522(.A1(new_n18577_), .A2(new_n13805_), .ZN(new_n18611_));
  AOI21_X1   g15523(.A1(new_n18576_), .A2(new_n13805_), .B(new_n18611_), .ZN(new_n18612_));
  AOI21_X1   g15524(.A1(new_n18612_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n18613_));
  AOI21_X1   g15525(.A1(new_n18610_), .A2(new_n18613_), .B(pi0618), .ZN(new_n18614_));
  OAI21_X1   g15526(.A1(new_n18595_), .A2(new_n18614_), .B(pi0781), .ZN(new_n18615_));
  XOR2_X1    g15527(.A1(new_n18586_), .A2(new_n18594_), .Z(new_n18616_));
  NAND3_X1   g15528(.A1(new_n18608_), .A2(pi0618), .A3(pi1154), .ZN(new_n18617_));
  NAND4_X1   g15529(.A1(new_n18607_), .A2(new_n13816_), .A3(pi1154), .A4(new_n18598_), .ZN(new_n18618_));
  AOI21_X1   g15530(.A1(new_n18617_), .A2(new_n18618_), .B(new_n18577_), .ZN(new_n18619_));
  NAND2_X1   g15531(.A1(new_n18612_), .A2(pi0618), .ZN(new_n18620_));
  NAND2_X1   g15532(.A1(new_n18620_), .A2(new_n13836_), .ZN(new_n18621_));
  OAI21_X1   g15533(.A1(new_n18619_), .A2(new_n18621_), .B(new_n13816_), .ZN(new_n18622_));
  NAND3_X1   g15534(.A1(new_n18616_), .A2(new_n18622_), .A3(pi0781), .ZN(new_n18623_));
  XOR2_X1    g15535(.A1(new_n18615_), .A2(new_n18623_), .Z(new_n18624_));
  NAND3_X1   g15536(.A1(new_n18608_), .A2(pi0618), .A3(pi1154), .ZN(new_n18625_));
  NAND3_X1   g15537(.A1(new_n18602_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n18626_));
  AOI21_X1   g15538(.A1(new_n18626_), .A2(new_n18625_), .B(new_n18577_), .ZN(new_n18627_));
  NAND4_X1   g15539(.A1(new_n18627_), .A2(new_n18619_), .A3(pi0781), .A4(new_n18608_), .ZN(new_n18628_));
  NOR2_X1    g15540(.A1(new_n18602_), .A2(new_n13855_), .ZN(new_n18629_));
  NAND2_X1   g15541(.A1(new_n18619_), .A2(new_n18629_), .ZN(new_n18630_));
  NAND3_X1   g15542(.A1(new_n18630_), .A2(pi0781), .A3(new_n18610_), .ZN(new_n18631_));
  NAND2_X1   g15543(.A1(new_n18631_), .A2(new_n18628_), .ZN(new_n18632_));
  NAND3_X1   g15544(.A1(new_n18632_), .A2(pi0619), .A3(pi1159), .ZN(new_n18633_));
  NAND4_X1   g15545(.A1(new_n18631_), .A2(pi0619), .A3(new_n13868_), .A4(new_n18628_), .ZN(new_n18634_));
  AOI21_X1   g15546(.A1(new_n18633_), .A2(new_n18634_), .B(new_n18577_), .ZN(new_n18635_));
  NOR2_X1    g15547(.A1(new_n18557_), .A2(new_n13880_), .ZN(new_n18636_));
  AOI21_X1   g15548(.A1(new_n18612_), .A2(new_n13880_), .B(new_n18636_), .ZN(new_n18637_));
  INV_X1     g15549(.I(new_n18637_), .ZN(new_n18638_));
  AOI21_X1   g15550(.A1(new_n18638_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n18639_));
  INV_X1     g15551(.I(new_n18639_), .ZN(new_n18640_));
  OAI21_X1   g15552(.A1(new_n18635_), .A2(new_n18640_), .B(new_n13860_), .ZN(new_n18641_));
  NAND3_X1   g15553(.A1(new_n18632_), .A2(pi0619), .A3(pi1159), .ZN(new_n18642_));
  NAND4_X1   g15554(.A1(new_n18631_), .A2(new_n13860_), .A3(pi1159), .A4(new_n18628_), .ZN(new_n18643_));
  AOI21_X1   g15555(.A1(new_n18642_), .A2(new_n18643_), .B(new_n18577_), .ZN(new_n18644_));
  AOI21_X1   g15556(.A1(new_n18638_), .A2(pi0619), .B(new_n15217_), .ZN(new_n18645_));
  INV_X1     g15557(.I(new_n18645_), .ZN(new_n18646_));
  OAI21_X1   g15558(.A1(new_n18644_), .A2(new_n18646_), .B(new_n13860_), .ZN(new_n18647_));
  NAND4_X1   g15559(.A1(new_n18641_), .A2(new_n18647_), .A3(pi0789), .A4(new_n18624_), .ZN(new_n18648_));
  NAND2_X1   g15560(.A1(new_n18641_), .A2(new_n18624_), .ZN(new_n18649_));
  NAND3_X1   g15561(.A1(new_n18647_), .A2(pi0789), .A3(new_n18624_), .ZN(new_n18650_));
  NAND3_X1   g15562(.A1(new_n18650_), .A2(new_n18649_), .A3(pi0789), .ZN(new_n18651_));
  NAND2_X1   g15563(.A1(new_n18651_), .A2(new_n18648_), .ZN(new_n18652_));
  NAND4_X1   g15564(.A1(new_n18635_), .A2(new_n18644_), .A3(pi0789), .A4(new_n18632_), .ZN(new_n18653_));
  AOI21_X1   g15565(.A1(new_n18602_), .A2(pi1154), .B(new_n13819_), .ZN(new_n18654_));
  INV_X1     g15566(.I(new_n18618_), .ZN(new_n18655_));
  OAI21_X1   g15567(.A1(new_n18654_), .A2(new_n18655_), .B(new_n18557_), .ZN(new_n18656_));
  NOR4_X1    g15568(.A1(new_n18610_), .A2(new_n18656_), .A3(new_n13855_), .A4(new_n18602_), .ZN(new_n18657_));
  NAND2_X1   g15569(.A1(new_n18610_), .A2(pi0781), .ZN(new_n18658_));
  NOR3_X1    g15570(.A1(new_n18656_), .A2(new_n13855_), .A3(new_n18602_), .ZN(new_n18659_));
  NOR2_X1    g15571(.A1(new_n18659_), .A2(new_n18658_), .ZN(new_n18660_));
  NOR2_X1    g15572(.A1(new_n18660_), .A2(new_n18657_), .ZN(new_n18661_));
  AOI21_X1   g15573(.A1(new_n18661_), .A2(pi0619), .B(new_n13904_), .ZN(new_n18662_));
  INV_X1     g15574(.I(new_n18634_), .ZN(new_n18663_));
  OAI21_X1   g15575(.A1(new_n18662_), .A2(new_n18663_), .B(new_n18557_), .ZN(new_n18664_));
  NOR2_X1    g15576(.A1(new_n18661_), .A2(new_n13896_), .ZN(new_n18665_));
  NAND2_X1   g15577(.A1(new_n18644_), .A2(new_n18665_), .ZN(new_n18666_));
  NAND3_X1   g15578(.A1(new_n18666_), .A2(pi0789), .A3(new_n18664_), .ZN(new_n18667_));
  NOR2_X1    g15579(.A1(new_n18577_), .A2(new_n13919_), .ZN(new_n18668_));
  AOI21_X1   g15580(.A1(new_n18637_), .A2(new_n13919_), .B(new_n18668_), .ZN(new_n18669_));
  NOR2_X1    g15581(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n18670_));
  INV_X1     g15582(.I(new_n18670_), .ZN(new_n18671_));
  AOI21_X1   g15583(.A1(new_n18667_), .A2(new_n18653_), .B(new_n18671_), .ZN(new_n18672_));
  AND3_X2    g15584(.A1(new_n18652_), .A2(pi0626), .A3(pi0788), .Z(new_n18676_));
  INV_X1     g15585(.I(new_n18653_), .ZN(new_n18677_));
  NAND2_X1   g15586(.A1(new_n18664_), .A2(pi0789), .ZN(new_n18678_));
  AOI21_X1   g15587(.A1(new_n18661_), .A2(pi1159), .B(new_n13904_), .ZN(new_n18679_));
  INV_X1     g15588(.I(new_n18643_), .ZN(new_n18680_));
  OAI21_X1   g15589(.A1(new_n18679_), .A2(new_n18680_), .B(new_n18557_), .ZN(new_n18681_));
  NOR3_X1    g15590(.A1(new_n18681_), .A2(new_n13896_), .A3(new_n18661_), .ZN(new_n18682_));
  NOR2_X1    g15591(.A1(new_n18682_), .A2(new_n18678_), .ZN(new_n18683_));
  OAI21_X1   g15592(.A1(new_n18683_), .A2(new_n18677_), .B(new_n18670_), .ZN(new_n18684_));
  AOI22_X1   g15593(.A1(new_n18684_), .A2(new_n13901_), .B1(new_n18648_), .B2(new_n18651_), .ZN(new_n18685_));
  AOI21_X1   g15594(.A1(new_n18651_), .A2(new_n18648_), .B(new_n15258_), .ZN(new_n18686_));
  NOR3_X1    g15595(.A1(new_n18685_), .A2(new_n13937_), .A3(new_n18686_), .ZN(new_n18687_));
  NOR2_X1    g15596(.A1(new_n18687_), .A2(new_n18676_), .ZN(new_n18688_));
  NAND2_X1   g15597(.A1(new_n18667_), .A2(new_n18653_), .ZN(new_n18689_));
  NOR2_X1    g15598(.A1(new_n18557_), .A2(new_n16372_), .ZN(new_n18690_));
  AOI21_X1   g15599(.A1(new_n18689_), .A2(new_n16372_), .B(new_n18690_), .ZN(new_n18691_));
  NOR2_X1    g15600(.A1(new_n18557_), .A2(new_n13966_), .ZN(new_n18693_));
  AOI21_X1   g15601(.A1(new_n18669_), .A2(new_n13966_), .B(new_n18693_), .ZN(new_n18694_));
  AOI21_X1   g15602(.A1(new_n18694_), .A2(pi0628), .B(new_n13971_), .ZN(new_n18695_));
  INV_X1     g15603(.I(new_n18694_), .ZN(new_n18696_));
  NOR3_X1    g15604(.A1(new_n18696_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n18697_));
  OAI21_X1   g15605(.A1(new_n18697_), .A2(new_n18695_), .B(new_n18557_), .ZN(new_n18698_));
  INV_X1     g15606(.I(new_n18698_), .ZN(new_n18699_));
  NOR2_X1    g15607(.A1(new_n18699_), .A2(new_n15270_), .ZN(new_n18700_));
  AOI21_X1   g15608(.A1(new_n18694_), .A2(pi1156), .B(new_n13971_), .ZN(new_n18703_));
  NOR3_X1    g15609(.A1(new_n18696_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n18704_));
  OAI21_X1   g15610(.A1(new_n18704_), .A2(new_n18703_), .B(new_n18557_), .ZN(new_n18705_));
  NOR3_X1    g15611(.A1(new_n18688_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n18708_));
  NAND3_X1   g15612(.A1(new_n18652_), .A2(pi0626), .A3(pi0788), .ZN(new_n18709_));
  INV_X1     g15613(.I(new_n18648_), .ZN(new_n18710_));
  INV_X1     g15614(.I(new_n18624_), .ZN(new_n18711_));
  AOI21_X1   g15615(.A1(new_n18664_), .A2(new_n18639_), .B(pi0619), .ZN(new_n18712_));
  OAI21_X1   g15616(.A1(new_n18712_), .A2(new_n18711_), .B(pi0789), .ZN(new_n18713_));
  AOI21_X1   g15617(.A1(new_n18681_), .A2(new_n18645_), .B(pi0619), .ZN(new_n18714_));
  INV_X1     g15618(.I(new_n18614_), .ZN(new_n18715_));
  AOI21_X1   g15619(.A1(new_n18616_), .A2(new_n18715_), .B(new_n13855_), .ZN(new_n18716_));
  NOR2_X1    g15620(.A1(new_n18716_), .A2(new_n18623_), .ZN(new_n18717_));
  NAND2_X1   g15621(.A1(new_n18716_), .A2(new_n18623_), .ZN(new_n18718_));
  INV_X1     g15622(.I(new_n18718_), .ZN(new_n18719_));
  OAI21_X1   g15623(.A1(new_n18719_), .A2(new_n18717_), .B(pi0789), .ZN(new_n18720_));
  NOR2_X1    g15624(.A1(new_n18714_), .A2(new_n18720_), .ZN(new_n18721_));
  NOR2_X1    g15625(.A1(new_n18713_), .A2(new_n18721_), .ZN(new_n18722_));
  OAI22_X1   g15626(.A1(new_n18722_), .A2(new_n18710_), .B1(pi0626), .B2(new_n18672_), .ZN(new_n18723_));
  OAI21_X1   g15627(.A1(new_n18722_), .A2(new_n18710_), .B(new_n14577_), .ZN(new_n18724_));
  NAND3_X1   g15628(.A1(new_n18723_), .A2(new_n18724_), .A3(pi0788), .ZN(new_n18725_));
  AOI21_X1   g15629(.A1(new_n18691_), .A2(new_n18700_), .B(pi0628), .ZN(new_n18726_));
  AOI21_X1   g15630(.A1(new_n18725_), .A2(new_n18709_), .B(new_n18726_), .ZN(new_n18727_));
  AOI21_X1   g15631(.A1(new_n18725_), .A2(new_n18709_), .B(new_n15296_), .ZN(new_n18728_));
  NOR3_X1    g15632(.A1(new_n18727_), .A2(new_n18728_), .A3(new_n12777_), .ZN(new_n18729_));
  NOR2_X1    g15633(.A1(new_n18729_), .A2(new_n18708_), .ZN(new_n18730_));
  NOR2_X1    g15634(.A1(new_n18557_), .A2(new_n13994_), .ZN(new_n18731_));
  INV_X1     g15635(.I(new_n18731_), .ZN(new_n18732_));
  OAI21_X1   g15636(.A1(new_n18691_), .A2(new_n13993_), .B(new_n18732_), .ZN(new_n18733_));
  NOR2_X1    g15637(.A1(new_n18699_), .A2(new_n12777_), .ZN(new_n18734_));
  NOR3_X1    g15638(.A1(new_n18705_), .A2(new_n12777_), .A3(new_n18694_), .ZN(new_n18735_));
  INV_X1     g15639(.I(new_n18735_), .ZN(new_n18736_));
  NOR2_X1    g15640(.A1(new_n18736_), .A2(new_n18734_), .ZN(new_n18737_));
  NAND2_X1   g15641(.A1(new_n18736_), .A2(new_n18734_), .ZN(new_n18738_));
  INV_X1     g15642(.I(new_n18738_), .ZN(new_n18739_));
  NOR2_X1    g15643(.A1(new_n18739_), .A2(new_n18737_), .ZN(new_n18740_));
  AOI21_X1   g15644(.A1(new_n18740_), .A2(pi0647), .B(new_n14008_), .ZN(new_n18741_));
  INV_X1     g15645(.I(new_n18737_), .ZN(new_n18742_));
  NAND2_X1   g15646(.A1(new_n18742_), .A2(new_n18738_), .ZN(new_n18743_));
  NOR3_X1    g15647(.A1(new_n18743_), .A2(new_n14005_), .A3(new_n14007_), .ZN(new_n18744_));
  OAI21_X1   g15648(.A1(new_n18744_), .A2(new_n18741_), .B(new_n18557_), .ZN(new_n18745_));
  NAND2_X1   g15649(.A1(new_n18745_), .A2(new_n14011_), .ZN(new_n18746_));
  OAI21_X1   g15650(.A1(new_n18746_), .A2(new_n18733_), .B(new_n14005_), .ZN(new_n18747_));
  INV_X1     g15651(.I(new_n18747_), .ZN(new_n18748_));
  AOI21_X1   g15652(.A1(new_n18740_), .A2(pi1157), .B(new_n14008_), .ZN(new_n18749_));
  NAND4_X1   g15653(.A1(new_n18742_), .A2(new_n18738_), .A3(new_n14005_), .A4(pi1157), .ZN(new_n18750_));
  INV_X1     g15654(.I(new_n18750_), .ZN(new_n18751_));
  OAI21_X1   g15655(.A1(new_n18749_), .A2(new_n18751_), .B(new_n18557_), .ZN(new_n18752_));
  NAND2_X1   g15656(.A1(new_n18752_), .A2(new_n14027_), .ZN(new_n18753_));
  AOI21_X1   g15657(.A1(pi0647), .A2(new_n18733_), .B(new_n18753_), .ZN(new_n18754_));
  NOR2_X1    g15658(.A1(new_n18754_), .A2(pi0647), .ZN(new_n18755_));
  NOR4_X1    g15659(.A1(new_n18730_), .A2(new_n12776_), .A3(new_n18748_), .A4(new_n18755_), .ZN(new_n18756_));
  NAND2_X1   g15660(.A1(new_n18725_), .A2(new_n18709_), .ZN(new_n18757_));
  NAND3_X1   g15661(.A1(new_n18757_), .A2(pi0628), .A3(pi0792), .ZN(new_n18758_));
  INV_X1     g15662(.I(new_n18726_), .ZN(new_n18759_));
  OAI21_X1   g15663(.A1(new_n18687_), .A2(new_n18676_), .B(new_n18759_), .ZN(new_n18760_));
  OAI21_X1   g15664(.A1(new_n18687_), .A2(new_n18676_), .B(new_n14606_), .ZN(new_n18761_));
  NAND3_X1   g15665(.A1(new_n18760_), .A2(new_n18761_), .A3(pi0792), .ZN(new_n18762_));
  AOI21_X1   g15666(.A1(new_n18762_), .A2(new_n18758_), .B(new_n18748_), .ZN(new_n18763_));
  OAI21_X1   g15667(.A1(new_n18754_), .A2(pi0647), .B(pi0787), .ZN(new_n18764_));
  AOI21_X1   g15668(.A1(new_n18762_), .A2(new_n18758_), .B(new_n18764_), .ZN(new_n18765_));
  NOR3_X1    g15669(.A1(new_n18765_), .A2(new_n18763_), .A3(new_n12776_), .ZN(new_n18766_));
  OAI21_X1   g15670(.A1(new_n18766_), .A2(new_n18756_), .B(new_n12775_), .ZN(new_n18767_));
  NAND2_X1   g15671(.A1(new_n18767_), .A2(new_n5787_), .ZN(new_n18768_));
  NAND2_X1   g15672(.A1(new_n18762_), .A2(new_n18758_), .ZN(new_n18769_));
  INV_X1     g15673(.I(new_n18755_), .ZN(new_n18770_));
  NAND4_X1   g15674(.A1(new_n18769_), .A2(pi0787), .A3(new_n18747_), .A4(new_n18770_), .ZN(new_n18771_));
  OAI21_X1   g15675(.A1(new_n18729_), .A2(new_n18708_), .B(new_n18747_), .ZN(new_n18772_));
  NAND2_X1   g15676(.A1(new_n18733_), .A2(pi0647), .ZN(new_n18773_));
  NAND3_X1   g15677(.A1(new_n18743_), .A2(pi0647), .A3(pi1157), .ZN(new_n18774_));
  NAND2_X1   g15678(.A1(new_n18774_), .A2(new_n18750_), .ZN(new_n18775_));
  AOI21_X1   g15679(.A1(new_n18775_), .A2(new_n18557_), .B(new_n16329_), .ZN(new_n18776_));
  NAND2_X1   g15680(.A1(new_n18773_), .A2(new_n18776_), .ZN(new_n18777_));
  AOI21_X1   g15681(.A1(new_n18777_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n18778_));
  OAI21_X1   g15682(.A1(new_n18729_), .A2(new_n18708_), .B(new_n18778_), .ZN(new_n18779_));
  NAND3_X1   g15683(.A1(new_n18772_), .A2(new_n18779_), .A3(pi0787), .ZN(new_n18780_));
  NAND2_X1   g15684(.A1(new_n18780_), .A2(new_n18771_), .ZN(new_n18781_));
  NOR4_X1    g15685(.A1(new_n18745_), .A2(new_n18752_), .A3(new_n12776_), .A4(new_n18740_), .ZN(new_n18782_));
  NAND2_X1   g15686(.A1(new_n18745_), .A2(pi0787), .ZN(new_n18783_));
  NOR3_X1    g15687(.A1(new_n18752_), .A2(new_n12776_), .A3(new_n18740_), .ZN(new_n18784_));
  NOR2_X1    g15688(.A1(new_n18784_), .A2(new_n18783_), .ZN(new_n18785_));
  OR2_X2     g15689(.A1(new_n18785_), .A2(new_n18782_), .Z(new_n18786_));
  NAND2_X1   g15690(.A1(new_n18557_), .A2(new_n14210_), .ZN(new_n18787_));
  OAI21_X1   g15691(.A1(new_n18733_), .A2(new_n14210_), .B(new_n18787_), .ZN(new_n18788_));
  NOR2_X1    g15692(.A1(new_n14204_), .A2(new_n14200_), .ZN(new_n18789_));
  NAND2_X1   g15693(.A1(new_n18788_), .A2(new_n18789_), .ZN(new_n18790_));
  OAI21_X1   g15694(.A1(new_n18786_), .A2(new_n18790_), .B(new_n14204_), .ZN(new_n18791_));
  AOI21_X1   g15695(.A1(new_n18781_), .A2(new_n18791_), .B(pi0790), .ZN(new_n18792_));
  OAI21_X1   g15696(.A1(new_n18785_), .A2(new_n18782_), .B(pi0644), .ZN(new_n18793_));
  NOR2_X1    g15697(.A1(new_n14204_), .A2(pi0715), .ZN(new_n18794_));
  NAND3_X1   g15698(.A1(new_n18793_), .A2(new_n18788_), .A3(new_n18794_), .ZN(new_n18795_));
  NAND2_X1   g15699(.A1(new_n5788_), .A2(new_n7378_), .ZN(new_n18796_));
  NOR2_X1    g15700(.A1(new_n13105_), .A2(new_n17309_), .ZN(new_n18797_));
  INV_X1     g15701(.I(new_n18797_), .ZN(new_n18798_));
  NOR2_X1    g15702(.A1(new_n18798_), .A2(new_n16376_), .ZN(new_n18799_));
  INV_X1     g15703(.I(new_n18799_), .ZN(new_n18800_));
  NOR2_X1    g15704(.A1(new_n16388_), .A2(new_n18800_), .ZN(new_n18801_));
  INV_X1     g15705(.I(new_n18801_), .ZN(new_n18802_));
  NOR2_X1    g15706(.A1(new_n18802_), .A2(new_n14142_), .ZN(new_n18803_));
  NOR2_X1    g15707(.A1(new_n13993_), .A2(new_n14210_), .ZN(new_n18804_));
  NOR2_X1    g15708(.A1(new_n9992_), .A2(new_n7378_), .ZN(new_n18805_));
  INV_X1     g15709(.I(new_n18805_), .ZN(new_n18806_));
  NAND2_X1   g15710(.A1(new_n18806_), .A2(new_n14200_), .ZN(new_n18807_));
  NAND4_X1   g15711(.A1(new_n18803_), .A2(pi0644), .A3(new_n18804_), .A4(new_n18807_), .ZN(new_n18808_));
  NOR2_X1    g15712(.A1(new_n13219_), .A2(new_n17327_), .ZN(new_n18809_));
  AOI21_X1   g15713(.A1(new_n18806_), .A2(new_n13614_), .B(new_n13613_), .ZN(new_n18810_));
  AOI21_X1   g15714(.A1(new_n18810_), .A2(new_n18809_), .B(new_n13748_), .ZN(new_n18811_));
  NOR4_X1    g15715(.A1(new_n13219_), .A2(new_n13613_), .A3(new_n17327_), .A4(new_n13614_), .ZN(new_n18812_));
  NOR4_X1    g15716(.A1(new_n13219_), .A2(pi0625), .A3(new_n17327_), .A4(pi1153), .ZN(new_n18813_));
  OAI21_X1   g15717(.A1(new_n18812_), .A2(new_n18813_), .B(new_n18805_), .ZN(new_n18814_));
  NOR4_X1    g15718(.A1(new_n18814_), .A2(new_n13748_), .A3(new_n18805_), .A4(new_n18809_), .ZN(new_n18815_));
  XNOR2_X1   g15719(.A1(new_n18815_), .A2(new_n18811_), .ZN(new_n18816_));
  NOR2_X1    g15720(.A1(new_n18816_), .A2(new_n15396_), .ZN(new_n18817_));
  INV_X1     g15721(.I(new_n18817_), .ZN(new_n18818_));
  NOR2_X1    g15722(.A1(new_n18818_), .A2(new_n14058_), .ZN(new_n18819_));
  AOI21_X1   g15723(.A1(new_n18819_), .A2(new_n15402_), .B(new_n18805_), .ZN(new_n18820_));
  NOR2_X1    g15724(.A1(new_n16435_), .A2(new_n17327_), .ZN(new_n18821_));
  NAND4_X1   g15725(.A1(new_n18821_), .A2(pi1153), .A3(new_n18797_), .A4(new_n18805_), .ZN(new_n18822_));
  NAND3_X1   g15726(.A1(new_n18822_), .A2(pi0608), .A3(new_n18814_), .ZN(new_n18823_));
  NAND2_X1   g15727(.A1(new_n18823_), .A2(pi0778), .ZN(new_n18824_));
  NOR2_X1    g15728(.A1(new_n18824_), .A2(pi0785), .ZN(new_n18825_));
  NAND2_X1   g15729(.A1(new_n18824_), .A2(pi1155), .ZN(new_n18826_));
  XOR2_X1    g15730(.A1(new_n18826_), .A2(new_n14090_), .Z(new_n18827_));
  NOR2_X1    g15731(.A1(new_n18805_), .A2(pi1155), .ZN(new_n18828_));
  NOR2_X1    g15732(.A1(new_n16444_), .A2(new_n18828_), .ZN(new_n18829_));
  AOI21_X1   g15733(.A1(new_n18829_), .A2(new_n18797_), .B(new_n13783_), .ZN(new_n18830_));
  OAI21_X1   g15734(.A1(new_n18827_), .A2(new_n18816_), .B(new_n18830_), .ZN(new_n18831_));
  NOR2_X1    g15735(.A1(new_n14102_), .A2(new_n18828_), .ZN(new_n18832_));
  AOI21_X1   g15736(.A1(new_n18832_), .A2(new_n18797_), .B(pi0660), .ZN(new_n18833_));
  INV_X1     g15737(.I(new_n18816_), .ZN(new_n18834_));
  NAND2_X1   g15738(.A1(new_n18824_), .A2(pi0609), .ZN(new_n18835_));
  XOR2_X1    g15739(.A1(new_n18835_), .A2(new_n14694_), .Z(new_n18836_));
  NAND3_X1   g15740(.A1(new_n18836_), .A2(pi0785), .A3(new_n18834_), .ZN(new_n18837_));
  AOI21_X1   g15741(.A1(new_n18831_), .A2(new_n18833_), .B(new_n18837_), .ZN(new_n18838_));
  NOR2_X1    g15742(.A1(new_n18838_), .A2(new_n18825_), .ZN(new_n18839_));
  AOI21_X1   g15743(.A1(new_n18834_), .A2(new_n13805_), .B(new_n18805_), .ZN(new_n18840_));
  INV_X1     g15744(.I(new_n18840_), .ZN(new_n18841_));
  NAND2_X1   g15745(.A1(new_n18839_), .A2(pi1154), .ZN(new_n18842_));
  XOR2_X1    g15746(.A1(new_n18842_), .A2(new_n13818_), .Z(new_n18843_));
  NOR2_X1    g15747(.A1(new_n18805_), .A2(pi1154), .ZN(new_n18844_));
  NOR2_X1    g15748(.A1(new_n16460_), .A2(new_n18844_), .ZN(new_n18845_));
  AOI21_X1   g15749(.A1(new_n18799_), .A2(new_n18845_), .B(new_n13823_), .ZN(new_n18846_));
  OAI21_X1   g15750(.A1(new_n18843_), .A2(new_n18841_), .B(new_n18846_), .ZN(new_n18847_));
  NOR2_X1    g15751(.A1(new_n16464_), .A2(new_n18844_), .ZN(new_n18848_));
  AOI21_X1   g15752(.A1(new_n18799_), .A2(new_n18848_), .B(pi0627), .ZN(new_n18849_));
  NAND2_X1   g15753(.A1(new_n18847_), .A2(new_n18849_), .ZN(new_n18850_));
  NAND2_X1   g15754(.A1(new_n18839_), .A2(pi0618), .ZN(new_n18851_));
  XOR2_X1    g15755(.A1(new_n18851_), .A2(new_n13818_), .Z(new_n18852_));
  NOR2_X1    g15756(.A1(new_n18852_), .A2(new_n18841_), .ZN(new_n18853_));
  AOI21_X1   g15757(.A1(new_n18850_), .A2(new_n18853_), .B(new_n13855_), .ZN(new_n18854_));
  XNOR2_X1   g15758(.A1(pi0619), .A2(pi0648), .ZN(new_n18855_));
  AOI21_X1   g15759(.A1(new_n13917_), .A2(new_n18855_), .B(new_n13896_), .ZN(new_n18856_));
  NAND2_X1   g15760(.A1(new_n18856_), .A2(pi0781), .ZN(new_n18857_));
  XOR2_X1    g15761(.A1(new_n18854_), .A2(new_n18857_), .Z(new_n18858_));
  NAND2_X1   g15762(.A1(new_n18834_), .A2(new_n15437_), .ZN(new_n18859_));
  OAI21_X1   g15763(.A1(new_n18859_), .A2(new_n13918_), .B(new_n18806_), .ZN(new_n18860_));
  NAND3_X1   g15764(.A1(new_n13901_), .A2(pi0641), .A3(pi1158), .ZN(new_n18861_));
  NOR2_X1    g15765(.A1(new_n16423_), .A2(pi0788), .ZN(new_n18862_));
  OAI21_X1   g15766(.A1(new_n18860_), .A2(new_n18861_), .B(new_n18862_), .ZN(new_n18863_));
  AOI21_X1   g15767(.A1(new_n18805_), .A2(pi1158), .B(pi0626), .ZN(new_n18864_));
  OAI21_X1   g15768(.A1(new_n18802_), .A2(new_n18864_), .B(new_n13922_), .ZN(new_n18865_));
  NAND2_X1   g15769(.A1(new_n18865_), .A2(new_n14140_), .ZN(new_n18866_));
  NOR2_X1    g15770(.A1(new_n18866_), .A2(new_n18860_), .ZN(new_n18867_));
  INV_X1     g15771(.I(new_n18855_), .ZN(new_n18868_));
  NAND4_X1   g15772(.A1(new_n13775_), .A2(new_n16382_), .A3(pi0619), .A4(new_n13885_), .ZN(new_n18869_));
  NOR2_X1    g15773(.A1(new_n18800_), .A2(new_n18869_), .ZN(new_n18870_));
  OAI21_X1   g15774(.A1(new_n18800_), .A2(new_n16476_), .B(new_n13915_), .ZN(new_n18871_));
  XNOR2_X1   g15775(.A1(new_n18871_), .A2(new_n18870_), .ZN(new_n18872_));
  NAND2_X1   g15776(.A1(new_n18806_), .A2(new_n13896_), .ZN(new_n18873_));
  NAND4_X1   g15777(.A1(new_n18872_), .A2(new_n16697_), .A3(new_n18868_), .A4(new_n18873_), .ZN(new_n18874_));
  OAI21_X1   g15778(.A1(new_n18874_), .A2(new_n18859_), .B(new_n15479_), .ZN(new_n18875_));
  AOI21_X1   g15779(.A1(new_n18867_), .A2(new_n18863_), .B(new_n18875_), .ZN(new_n18876_));
  NOR3_X1    g15780(.A1(new_n18858_), .A2(new_n18839_), .A3(new_n18876_), .ZN(new_n18877_));
  NOR3_X1    g15781(.A1(new_n18803_), .A2(pi0630), .A3(pi0647), .ZN(new_n18878_));
  NAND2_X1   g15782(.A1(new_n13993_), .A2(pi1157), .ZN(new_n18879_));
  OAI21_X1   g15783(.A1(new_n18878_), .A2(new_n18879_), .B(new_n14010_), .ZN(new_n18880_));
  NOR3_X1    g15784(.A1(new_n18803_), .A2(pi0630), .A3(pi1157), .ZN(new_n18881_));
  NAND2_X1   g15785(.A1(new_n13993_), .A2(pi0647), .ZN(new_n18882_));
  OAI22_X1   g15786(.A1(new_n18881_), .A2(new_n18882_), .B1(new_n14058_), .B2(new_n18818_), .ZN(new_n18883_));
  AND3_X2    g15787(.A1(new_n16418_), .A2(pi0630), .A3(pi0787), .Z(new_n18884_));
  AND4_X2    g15788(.A1(new_n18819_), .A2(new_n18883_), .A3(new_n18880_), .A4(new_n18884_), .Z(new_n18885_));
  NOR2_X1    g15789(.A1(new_n18818_), .A2(new_n13942_), .ZN(new_n18886_));
  NOR2_X1    g15790(.A1(new_n18886_), .A2(new_n13969_), .ZN(new_n18887_));
  INV_X1     g15791(.I(new_n18803_), .ZN(new_n18888_));
  AOI21_X1   g15792(.A1(new_n18818_), .A2(new_n13976_), .B(new_n18888_), .ZN(new_n18889_));
  AOI21_X1   g15793(.A1(new_n18888_), .A2(new_n13942_), .B(new_n15270_), .ZN(new_n18890_));
  OAI21_X1   g15794(.A1(new_n18889_), .A2(new_n18886_), .B(new_n18890_), .ZN(new_n18891_));
  NOR2_X1    g15795(.A1(new_n18805_), .A2(new_n12777_), .ZN(new_n18892_));
  OAI21_X1   g15796(.A1(new_n18891_), .A2(new_n18887_), .B(new_n18892_), .ZN(new_n18893_));
  AOI21_X1   g15797(.A1(new_n18887_), .A2(new_n18891_), .B(new_n18893_), .ZN(new_n18894_));
  OAI21_X1   g15798(.A1(new_n18877_), .A2(new_n18885_), .B(new_n18894_), .ZN(new_n18895_));
  NAND2_X1   g15799(.A1(new_n18895_), .A2(pi0644), .ZN(new_n18896_));
  XOR2_X1    g15800(.A1(new_n18896_), .A2(new_n14217_), .Z(new_n18897_));
  NAND4_X1   g15801(.A1(new_n18897_), .A2(new_n14203_), .A3(new_n18808_), .A4(new_n18820_), .ZN(new_n18898_));
  INV_X1     g15802(.I(new_n18820_), .ZN(new_n18899_));
  NAND2_X1   g15803(.A1(new_n18895_), .A2(pi0715), .ZN(new_n18900_));
  XOR2_X1    g15804(.A1(new_n18900_), .A2(new_n14205_), .Z(new_n18901_));
  NOR2_X1    g15805(.A1(new_n18901_), .A2(new_n18899_), .ZN(new_n18902_));
  AOI21_X1   g15806(.A1(new_n18898_), .A2(new_n18902_), .B(new_n14799_), .ZN(new_n18903_));
  XOR2_X1    g15807(.A1(new_n18903_), .A2(new_n14800_), .Z(new_n18904_));
  OAI21_X1   g15808(.A1(new_n5371_), .A2(new_n7378_), .B(new_n14799_), .ZN(new_n18905_));
  NOR2_X1    g15809(.A1(new_n18895_), .A2(new_n18905_), .ZN(new_n18906_));
  AOI22_X1   g15810(.A1(new_n18904_), .A2(new_n18906_), .B1(new_n5371_), .B2(new_n18796_), .ZN(new_n18907_));
  AOI21_X1   g15811(.A1(new_n18795_), .A2(new_n14204_), .B(new_n18907_), .ZN(new_n18908_));
  NAND2_X1   g15812(.A1(new_n18781_), .A2(new_n18908_), .ZN(new_n18909_));
  AOI21_X1   g15813(.A1(new_n18768_), .A2(new_n18792_), .B(new_n18909_), .ZN(po0331));
  NOR2_X1    g15814(.A1(new_n14652_), .A2(new_n17392_), .ZN(new_n18911_));
  INV_X1     g15815(.I(new_n18911_), .ZN(new_n18912_));
  NOR2_X1    g15816(.A1(new_n9992_), .A2(pi0175), .ZN(new_n18913_));
  NOR2_X1    g15817(.A1(new_n18913_), .A2(pi1153), .ZN(new_n18914_));
  NAND2_X1   g15818(.A1(new_n18912_), .A2(new_n18914_), .ZN(new_n18915_));
  INV_X1     g15819(.I(new_n18915_), .ZN(new_n18916_));
  NOR2_X1    g15820(.A1(new_n18916_), .A2(new_n13748_), .ZN(new_n18917_));
  AOI21_X1   g15821(.A1(new_n13218_), .A2(pi0700), .B(new_n18913_), .ZN(new_n18918_));
  INV_X1     g15822(.I(new_n18918_), .ZN(new_n18919_));
  AOI21_X1   g15823(.A1(new_n18912_), .A2(new_n18919_), .B(new_n13614_), .ZN(new_n18920_));
  INV_X1     g15824(.I(new_n18920_), .ZN(new_n18921_));
  NOR3_X1    g15825(.A1(new_n18921_), .A2(new_n13748_), .A3(new_n18919_), .ZN(new_n18922_));
  XNOR2_X1   g15826(.A1(new_n18922_), .A2(new_n18917_), .ZN(new_n18923_));
  NAND2_X1   g15827(.A1(new_n18923_), .A2(new_n14049_), .ZN(new_n18924_));
  NOR2_X1    g15828(.A1(new_n18924_), .A2(new_n14051_), .ZN(new_n18925_));
  INV_X1     g15829(.I(new_n18925_), .ZN(new_n18926_));
  NOR2_X1    g15830(.A1(new_n18926_), .A2(new_n14163_), .ZN(new_n18927_));
  NOR2_X1    g15831(.A1(new_n13966_), .A2(new_n2723_), .ZN(new_n18928_));
  INV_X1     g15832(.I(new_n18928_), .ZN(new_n18929_));
  NAND2_X1   g15833(.A1(new_n18927_), .A2(new_n18929_), .ZN(new_n18930_));
  NOR2_X1    g15834(.A1(new_n18930_), .A2(new_n14060_), .ZN(new_n18931_));
  INV_X1     g15835(.I(new_n18913_), .ZN(new_n18932_));
  NAND3_X1   g15836(.A1(new_n18931_), .A2(pi0647), .A3(pi1157), .ZN(new_n18933_));
  OR3_X2     g15837(.A1(new_n18931_), .A2(new_n14005_), .A3(pi1157), .Z(new_n18934_));
  AOI21_X1   g15838(.A1(new_n18934_), .A2(new_n18933_), .B(new_n18932_), .ZN(new_n18935_));
  INV_X1     g15839(.I(new_n18935_), .ZN(new_n18936_));
  NOR2_X1    g15840(.A1(new_n18932_), .A2(pi0647), .ZN(new_n18937_));
  AOI21_X1   g15841(.A1(new_n18931_), .A2(pi0647), .B(new_n18937_), .ZN(new_n18938_));
  AOI21_X1   g15842(.A1(new_n18938_), .A2(pi1157), .B(new_n12776_), .ZN(new_n18939_));
  AOI22_X1   g15843(.A1(new_n18936_), .A2(new_n18939_), .B1(new_n12776_), .B2(new_n18931_), .ZN(new_n18940_));
  INV_X1     g15844(.I(new_n18940_), .ZN(new_n18941_));
  NOR2_X1    g15845(.A1(new_n13105_), .A2(new_n17355_), .ZN(new_n18942_));
  INV_X1     g15846(.I(new_n18942_), .ZN(new_n18943_));
  NOR2_X1    g15847(.A1(new_n18942_), .A2(new_n18913_), .ZN(new_n18944_));
  INV_X1     g15848(.I(new_n18944_), .ZN(new_n18945_));
  NAND3_X1   g15849(.A1(new_n18945_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n18946_));
  AOI21_X1   g15850(.A1(new_n18946_), .A2(new_n16444_), .B(new_n18943_), .ZN(new_n18947_));
  NOR2_X1    g15851(.A1(new_n18947_), .A2(new_n13801_), .ZN(new_n18948_));
  NOR2_X1    g15852(.A1(new_n18913_), .A2(pi1155), .ZN(new_n18949_));
  NOR3_X1    g15853(.A1(new_n18943_), .A2(new_n16444_), .A3(new_n18949_), .ZN(new_n18950_));
  NAND4_X1   g15854(.A1(new_n18950_), .A2(new_n18945_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n18951_));
  XOR2_X1    g15855(.A1(new_n18948_), .A2(new_n18951_), .Z(new_n18952_));
  NOR2_X1    g15856(.A1(new_n18952_), .A2(new_n13817_), .ZN(new_n18953_));
  OAI21_X1   g15857(.A1(new_n18953_), .A2(pi0618), .B(new_n9992_), .ZN(new_n18954_));
  NAND2_X1   g15858(.A1(new_n18954_), .A2(pi0781), .ZN(new_n18955_));
  OAI21_X1   g15859(.A1(new_n18953_), .A2(new_n9992_), .B(pi0618), .ZN(new_n18956_));
  NOR3_X1    g15860(.A1(new_n18956_), .A2(new_n13855_), .A3(new_n18952_), .ZN(new_n18957_));
  XOR2_X1    g15861(.A1(new_n18957_), .A2(new_n18955_), .Z(new_n18958_));
  NOR2_X1    g15862(.A1(new_n18958_), .A2(new_n13868_), .ZN(new_n18959_));
  OAI21_X1   g15863(.A1(new_n18959_), .A2(pi0619), .B(new_n9992_), .ZN(new_n18960_));
  NAND2_X1   g15864(.A1(new_n18960_), .A2(pi0789), .ZN(new_n18961_));
  OAI21_X1   g15865(.A1(new_n18959_), .A2(new_n9992_), .B(pi0619), .ZN(new_n18962_));
  NOR3_X1    g15866(.A1(new_n18962_), .A2(new_n13896_), .A3(new_n18958_), .ZN(new_n18963_));
  XOR2_X1    g15867(.A1(new_n18963_), .A2(new_n18961_), .Z(new_n18964_));
  NAND2_X1   g15868(.A1(new_n18964_), .A2(new_n16372_), .ZN(new_n18965_));
  OAI21_X1   g15869(.A1(new_n16372_), .A2(new_n18913_), .B(new_n18965_), .ZN(new_n18966_));
  NOR2_X1    g15870(.A1(new_n13994_), .A2(new_n14211_), .ZN(new_n18967_));
  INV_X1     g15871(.I(new_n18967_), .ZN(new_n18968_));
  NOR2_X1    g15872(.A1(new_n18966_), .A2(new_n18968_), .ZN(new_n18969_));
  NAND2_X1   g15873(.A1(new_n18967_), .A2(new_n18913_), .ZN(new_n18970_));
  XOR2_X1    g15874(.A1(new_n18969_), .A2(new_n18970_), .Z(new_n18971_));
  AOI21_X1   g15875(.A1(new_n18932_), .A2(new_n14254_), .B(pi0644), .ZN(new_n18972_));
  NAND2_X1   g15876(.A1(new_n18964_), .A2(new_n13962_), .ZN(new_n18973_));
  INV_X1     g15877(.I(new_n13962_), .ZN(new_n18974_));
  NOR2_X1    g15878(.A1(new_n18974_), .A2(new_n13901_), .ZN(new_n18975_));
  INV_X1     g15879(.I(new_n18975_), .ZN(new_n18976_));
  XOR2_X1    g15880(.A1(new_n18973_), .A2(new_n18976_), .Z(new_n18977_));
  AOI22_X1   g15881(.A1(new_n18977_), .A2(new_n18913_), .B1(new_n16639_), .B2(new_n18927_), .ZN(new_n18978_));
  NOR2_X1    g15882(.A1(new_n18918_), .A2(new_n13203_), .ZN(new_n18979_));
  NAND2_X1   g15883(.A1(new_n18979_), .A2(pi0625), .ZN(new_n18980_));
  NAND3_X1   g15884(.A1(new_n18980_), .A2(pi1153), .A3(new_n18944_), .ZN(new_n18981_));
  NOR2_X1    g15885(.A1(new_n18916_), .A2(new_n14081_), .ZN(new_n18982_));
  AOI21_X1   g15886(.A1(new_n18982_), .A2(new_n18981_), .B(new_n13748_), .ZN(new_n18983_));
  NOR2_X1    g15887(.A1(new_n18945_), .A2(new_n18979_), .ZN(new_n18984_));
  INV_X1     g15888(.I(new_n18980_), .ZN(new_n18985_));
  OAI21_X1   g15889(.A1(new_n18984_), .A2(new_n18985_), .B(new_n18914_), .ZN(new_n18986_));
  NAND4_X1   g15890(.A1(new_n18986_), .A2(new_n13749_), .A3(new_n18921_), .A4(new_n18984_), .ZN(new_n18987_));
  XNOR2_X1   g15891(.A1(new_n18987_), .A2(new_n18983_), .ZN(new_n18988_));
  NAND2_X1   g15892(.A1(new_n18988_), .A2(new_n13801_), .ZN(new_n18989_));
  NOR2_X1    g15893(.A1(new_n18947_), .A2(pi0660), .ZN(new_n18992_));
  NOR2_X1    g15894(.A1(new_n18988_), .A2(new_n13766_), .ZN(new_n18993_));
  XOR2_X1    g15895(.A1(new_n18993_), .A2(new_n14090_), .Z(new_n18994_));
  NOR2_X1    g15896(.A1(new_n18923_), .A2(new_n13801_), .ZN(new_n18995_));
  NAND2_X1   g15897(.A1(new_n18994_), .A2(new_n18995_), .ZN(new_n18996_));
  OAI21_X1   g15898(.A1(new_n18996_), .A2(new_n18992_), .B(new_n18989_), .ZN(new_n18997_));
  NAND2_X1   g15899(.A1(new_n18997_), .A2(new_n13855_), .ZN(new_n18998_));
  INV_X1     g15900(.I(new_n18924_), .ZN(new_n18999_));
  NOR2_X1    g15901(.A1(new_n18997_), .A2(new_n13816_), .ZN(new_n19000_));
  XOR2_X1    g15902(.A1(new_n19000_), .A2(new_n13818_), .Z(new_n19001_));
  NAND2_X1   g15903(.A1(new_n19001_), .A2(new_n18999_), .ZN(new_n19002_));
  NAND3_X1   g15904(.A1(new_n19002_), .A2(new_n13823_), .A3(new_n18956_), .ZN(new_n19003_));
  NAND3_X1   g15905(.A1(new_n19003_), .A2(new_n13823_), .A3(new_n18954_), .ZN(new_n19004_));
  NOR2_X1    g15906(.A1(new_n18997_), .A2(new_n13817_), .ZN(new_n19005_));
  XOR2_X1    g15907(.A1(new_n19005_), .A2(new_n13818_), .Z(new_n19006_));
  NAND4_X1   g15908(.A1(new_n19004_), .A2(pi0781), .A3(new_n18999_), .A4(new_n19006_), .ZN(new_n19007_));
  NAND2_X1   g15909(.A1(new_n19007_), .A2(new_n18998_), .ZN(new_n19008_));
  NOR2_X1    g15910(.A1(new_n19008_), .A2(new_n13860_), .ZN(new_n19009_));
  XOR2_X1    g15911(.A1(new_n19009_), .A2(new_n13904_), .Z(new_n19010_));
  NOR2_X1    g15912(.A1(new_n19010_), .A2(new_n18926_), .ZN(new_n19011_));
  NAND2_X1   g15913(.A1(new_n18962_), .A2(new_n13884_), .ZN(new_n19012_));
  INV_X1     g15914(.I(new_n19008_), .ZN(new_n19013_));
  AOI21_X1   g15915(.A1(new_n19013_), .A2(new_n14143_), .B(pi0789), .ZN(new_n19014_));
  OAI21_X1   g15916(.A1(new_n19011_), .A2(new_n19012_), .B(new_n19014_), .ZN(new_n19015_));
  NOR2_X1    g15917(.A1(new_n19008_), .A2(new_n13868_), .ZN(new_n19016_));
  XOR2_X1    g15918(.A1(new_n19016_), .A2(new_n13903_), .Z(new_n19017_));
  NOR2_X1    g15919(.A1(new_n13884_), .A2(new_n13937_), .ZN(new_n19018_));
  NAND2_X1   g15920(.A1(new_n18960_), .A2(new_n19018_), .ZN(new_n19019_));
  AOI21_X1   g15921(.A1(new_n19017_), .A2(new_n18925_), .B(new_n19019_), .ZN(new_n19020_));
  AOI21_X1   g15922(.A1(new_n19015_), .A2(new_n19020_), .B(new_n18978_), .ZN(new_n19021_));
  INV_X1     g15923(.I(new_n16547_), .ZN(new_n19022_));
  NAND3_X1   g15924(.A1(new_n18966_), .A2(new_n18927_), .A3(new_n18929_), .ZN(new_n19023_));
  NAND2_X1   g15925(.A1(new_n19023_), .A2(new_n16569_), .ZN(new_n19024_));
  XOR2_X1    g15926(.A1(new_n19024_), .A2(new_n16572_), .Z(new_n19025_));
  AOI21_X1   g15927(.A1(new_n19022_), .A2(new_n19023_), .B(new_n19025_), .ZN(new_n19026_));
  NAND2_X1   g15928(.A1(new_n18964_), .A2(new_n13963_), .ZN(new_n19027_));
  NAND2_X1   g15929(.A1(new_n13963_), .A2(pi0626), .ZN(new_n19028_));
  XNOR2_X1   g15930(.A1(new_n19027_), .A2(new_n19028_), .ZN(new_n19029_));
  NOR3_X1    g15931(.A1(new_n19029_), .A2(new_n16424_), .A3(new_n18932_), .ZN(new_n19030_));
  OAI21_X1   g15932(.A1(new_n19026_), .A2(new_n16574_), .B(new_n19030_), .ZN(new_n19031_));
  NOR2_X1    g15933(.A1(new_n18966_), .A2(new_n13994_), .ZN(new_n19032_));
  NAND2_X1   g15934(.A1(new_n13993_), .A2(new_n16576_), .ZN(new_n19033_));
  XNOR2_X1   g15935(.A1(new_n19032_), .A2(new_n19033_), .ZN(new_n19034_));
  AOI22_X1   g15936(.A1(new_n19034_), .A2(new_n18913_), .B1(new_n14206_), .B2(new_n18938_), .ZN(new_n19035_));
  NOR3_X1    g15937(.A1(new_n19035_), .A2(new_n14010_), .A3(new_n18936_), .ZN(new_n19036_));
  OAI22_X1   g15938(.A1(new_n19021_), .A2(new_n19031_), .B1(new_n12776_), .B2(new_n19036_), .ZN(new_n19037_));
  NAND2_X1   g15939(.A1(new_n19037_), .A2(pi0644), .ZN(new_n19038_));
  XOR2_X1    g15940(.A1(new_n19038_), .A2(new_n14205_), .Z(new_n19039_));
  NOR2_X1    g15941(.A1(new_n19039_), .A2(new_n18940_), .ZN(new_n19040_));
  NAND2_X1   g15942(.A1(new_n18971_), .A2(pi0715), .ZN(new_n19041_));
  XOR2_X1    g15943(.A1(new_n19041_), .A2(new_n14205_), .Z(new_n19042_));
  NOR2_X1    g15944(.A1(new_n12775_), .A2(pi1160), .ZN(new_n19043_));
  OAI21_X1   g15945(.A1(new_n19042_), .A2(new_n18932_), .B(new_n19043_), .ZN(new_n19044_));
  OAI22_X1   g15946(.A1(new_n19040_), .A2(new_n19044_), .B1(new_n18971_), .B2(new_n18972_), .ZN(new_n19045_));
  NAND2_X1   g15947(.A1(new_n19037_), .A2(pi0715), .ZN(new_n19046_));
  XOR2_X1    g15948(.A1(new_n19046_), .A2(new_n14217_), .Z(new_n19047_));
  AOI21_X1   g15949(.A1(po1038), .A2(new_n9486_), .B(pi0832), .ZN(new_n19048_));
  NAND4_X1   g15950(.A1(new_n19045_), .A2(new_n18941_), .A3(new_n19047_), .A4(new_n19048_), .ZN(new_n19049_));
  NOR2_X1    g15951(.A1(new_n14428_), .A2(pi0175), .ZN(new_n19050_));
  INV_X1     g15952(.I(new_n19050_), .ZN(new_n19051_));
  INV_X1     g15953(.I(new_n14389_), .ZN(new_n19052_));
  OAI22_X1   g15954(.A1(new_n17127_), .A2(new_n9486_), .B1(new_n17355_), .B2(new_n19052_), .ZN(new_n19053_));
  OAI21_X1   g15955(.A1(pi0175), .A2(new_n14299_), .B(new_n14301_), .ZN(new_n19054_));
  NAND2_X1   g15956(.A1(new_n14299_), .A2(pi0766), .ZN(new_n19055_));
  NAND4_X1   g15957(.A1(new_n19054_), .A2(new_n17355_), .A3(new_n14362_), .A4(new_n19055_), .ZN(new_n19056_));
  NAND3_X1   g15958(.A1(new_n19056_), .A2(pi0038), .A3(pi0175), .ZN(new_n19057_));
  NAND2_X1   g15959(.A1(new_n19057_), .A2(new_n3183_), .ZN(new_n19058_));
  NAND2_X1   g15960(.A1(new_n13109_), .A2(new_n9486_), .ZN(new_n19059_));
  NAND4_X1   g15961(.A1(new_n19058_), .A2(pi0038), .A3(new_n19053_), .A4(new_n19059_), .ZN(new_n19060_));
  AOI21_X1   g15962(.A1(new_n19060_), .A2(new_n17355_), .B(new_n13107_), .ZN(new_n19061_));
  NAND2_X1   g15963(.A1(new_n19061_), .A2(new_n3289_), .ZN(new_n19062_));
  NAND2_X1   g15964(.A1(new_n3290_), .A2(new_n9486_), .ZN(new_n19063_));
  NAND3_X1   g15965(.A1(new_n19062_), .A2(new_n13776_), .A3(new_n19063_), .ZN(new_n19064_));
  NAND2_X1   g15966(.A1(new_n19051_), .A2(new_n13780_), .ZN(new_n19065_));
  NAND2_X1   g15967(.A1(new_n19064_), .A2(new_n19065_), .ZN(new_n19066_));
  NAND2_X1   g15968(.A1(new_n19066_), .A2(pi0609), .ZN(new_n19067_));
  NAND2_X1   g15969(.A1(new_n19067_), .A2(pi0785), .ZN(new_n19068_));
  NAND2_X1   g15970(.A1(new_n19062_), .A2(new_n19063_), .ZN(new_n19069_));
  NOR2_X1    g15971(.A1(new_n19051_), .A2(new_n13776_), .ZN(new_n19070_));
  AOI21_X1   g15972(.A1(new_n19069_), .A2(new_n13776_), .B(new_n19070_), .ZN(new_n19071_));
  AOI21_X1   g15973(.A1(new_n19051_), .A2(new_n14467_), .B(pi0609), .ZN(new_n19072_));
  OR2_X2     g15974(.A1(new_n19064_), .A2(new_n19072_), .Z(new_n19073_));
  NOR3_X1    g15975(.A1(new_n19073_), .A2(new_n13801_), .A3(new_n19071_), .ZN(new_n19074_));
  XNOR2_X1   g15976(.A1(new_n19074_), .A2(new_n19068_), .ZN(new_n19075_));
  NAND3_X1   g15977(.A1(new_n19075_), .A2(pi0618), .A3(pi1154), .ZN(new_n19076_));
  XOR2_X1    g15978(.A1(new_n19074_), .A2(new_n19068_), .Z(new_n19077_));
  NAND3_X1   g15979(.A1(new_n19077_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n19078_));
  NAND2_X1   g15980(.A1(new_n19076_), .A2(new_n19078_), .ZN(new_n19079_));
  NAND2_X1   g15981(.A1(new_n19079_), .A2(new_n19050_), .ZN(new_n19080_));
  NAND2_X1   g15982(.A1(new_n19080_), .A2(pi0781), .ZN(new_n19081_));
  NAND3_X1   g15983(.A1(new_n19075_), .A2(pi0618), .A3(pi1154), .ZN(new_n19082_));
  NAND3_X1   g15984(.A1(new_n19077_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n19083_));
  NAND2_X1   g15985(.A1(new_n19082_), .A2(new_n19083_), .ZN(new_n19084_));
  NAND2_X1   g15986(.A1(new_n19084_), .A2(new_n19050_), .ZN(new_n19085_));
  NOR3_X1    g15987(.A1(new_n19085_), .A2(new_n13855_), .A3(new_n19077_), .ZN(new_n19086_));
  NAND2_X1   g15988(.A1(new_n19086_), .A2(new_n19081_), .ZN(new_n19087_));
  OR2_X2     g15989(.A1(new_n19086_), .A2(new_n19081_), .Z(new_n19088_));
  NAND2_X1   g15990(.A1(new_n19088_), .A2(new_n19087_), .ZN(new_n19089_));
  NAND3_X1   g15991(.A1(new_n19089_), .A2(pi0619), .A3(pi1159), .ZN(new_n19090_));
  NOR3_X1    g15992(.A1(new_n19089_), .A2(new_n13860_), .A3(pi1159), .ZN(new_n19091_));
  INV_X1     g15993(.I(new_n19091_), .ZN(new_n19092_));
  AOI21_X1   g15994(.A1(new_n19092_), .A2(new_n19090_), .B(new_n19051_), .ZN(new_n19093_));
  NAND2_X1   g15995(.A1(new_n19051_), .A2(new_n13879_), .ZN(new_n19094_));
  OAI21_X1   g15996(.A1(new_n13721_), .A2(new_n17392_), .B(new_n9486_), .ZN(new_n19095_));
  NAND2_X1   g15997(.A1(new_n19095_), .A2(new_n13108_), .ZN(new_n19096_));
  NAND2_X1   g15998(.A1(new_n9486_), .A2(new_n17392_), .ZN(new_n19097_));
  NAND4_X1   g15999(.A1(new_n13634_), .A2(pi0175), .A3(new_n3290_), .A4(new_n19097_), .ZN(new_n19098_));
  NOR3_X1    g16000(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n9486_), .ZN(new_n19099_));
  NOR3_X1    g16001(.A1(new_n14422_), .A2(pi0038), .A3(new_n9486_), .ZN(new_n19100_));
  OAI21_X1   g16002(.A1(new_n19099_), .A2(new_n19100_), .B(new_n15655_), .ZN(new_n19101_));
  AOI21_X1   g16003(.A1(new_n19096_), .A2(new_n19098_), .B(new_n19101_), .ZN(new_n19102_));
  NOR2_X1    g16004(.A1(new_n19050_), .A2(new_n13613_), .ZN(new_n19103_));
  XOR2_X1    g16005(.A1(new_n19103_), .A2(new_n13615_), .Z(new_n19104_));
  NAND2_X1   g16006(.A1(new_n19104_), .A2(new_n19102_), .ZN(new_n19105_));
  NAND2_X1   g16007(.A1(new_n19105_), .A2(pi0778), .ZN(new_n19106_));
  NOR2_X1    g16008(.A1(new_n19050_), .A2(new_n13614_), .ZN(new_n19107_));
  XOR2_X1    g16009(.A1(new_n19107_), .A2(new_n13615_), .Z(new_n19108_));
  NAND3_X1   g16010(.A1(new_n19108_), .A2(pi0778), .A3(new_n19102_), .ZN(new_n19109_));
  XOR2_X1    g16011(.A1(new_n19106_), .A2(new_n19109_), .Z(new_n19110_));
  INV_X1     g16012(.I(new_n19110_), .ZN(new_n19111_));
  NAND2_X1   g16013(.A1(new_n19050_), .A2(new_n13803_), .ZN(new_n19112_));
  OAI21_X1   g16014(.A1(new_n19111_), .A2(new_n13803_), .B(new_n19112_), .ZN(new_n19113_));
  OAI21_X1   g16015(.A1(new_n19113_), .A2(new_n13879_), .B(new_n19094_), .ZN(new_n19114_));
  INV_X1     g16016(.I(new_n19061_), .ZN(new_n19115_));
  NOR2_X1    g16017(.A1(new_n9486_), .A2(new_n17355_), .ZN(new_n19116_));
  INV_X1     g16018(.I(new_n19116_), .ZN(new_n19117_));
  NAND2_X1   g16019(.A1(new_n13461_), .A2(pi0766), .ZN(new_n19118_));
  XOR2_X1    g16020(.A1(new_n19118_), .A2(new_n19117_), .Z(new_n19119_));
  NAND2_X1   g16021(.A1(new_n19119_), .A2(new_n13521_), .ZN(new_n19120_));
  NAND3_X1   g16022(.A1(new_n14270_), .A2(pi0175), .A3(pi0766), .ZN(new_n19121_));
  NAND3_X1   g16023(.A1(new_n14272_), .A2(pi0175), .A3(new_n17355_), .ZN(new_n19122_));
  AOI21_X1   g16024(.A1(new_n19121_), .A2(new_n19122_), .B(new_n13152_), .ZN(new_n19123_));
  NAND3_X1   g16025(.A1(new_n13198_), .A2(pi0175), .A3(pi0766), .ZN(new_n19124_));
  NAND3_X1   g16026(.A1(new_n13200_), .A2(new_n9486_), .A3(pi0766), .ZN(new_n19125_));
  AOI21_X1   g16027(.A1(new_n19125_), .A2(new_n19124_), .B(new_n13191_), .ZN(new_n19126_));
  OAI21_X1   g16028(.A1(new_n19123_), .A2(new_n3212_), .B(new_n19126_), .ZN(new_n19127_));
  NAND3_X1   g16029(.A1(new_n19120_), .A2(new_n3183_), .A3(new_n19127_), .ZN(new_n19128_));
  NOR2_X1    g16030(.A1(new_n14284_), .A2(new_n9486_), .ZN(new_n19129_));
  XOR2_X1    g16031(.A1(new_n19129_), .A2(new_n19116_), .Z(new_n19130_));
  NAND3_X1   g16032(.A1(new_n19128_), .A2(new_n19130_), .A3(new_n13359_), .ZN(new_n19131_));
  NAND3_X1   g16033(.A1(new_n19131_), .A2(new_n17392_), .A3(new_n3290_), .ZN(new_n19132_));
  NAND2_X1   g16034(.A1(new_n3290_), .A2(pi0175), .ZN(new_n19133_));
  NOR2_X1    g16035(.A1(new_n14291_), .A2(new_n13211_), .ZN(new_n19134_));
  AOI21_X1   g16036(.A1(new_n13209_), .A2(pi0039), .B(new_n19134_), .ZN(new_n19135_));
  NAND2_X1   g16037(.A1(new_n5504_), .A2(new_n9486_), .ZN(new_n19136_));
  NOR2_X1    g16038(.A1(new_n18943_), .A2(new_n16751_), .ZN(new_n19137_));
  AOI21_X1   g16039(.A1(new_n19136_), .A2(new_n19137_), .B(pi0038), .ZN(new_n19138_));
  NOR4_X1    g16040(.A1(new_n19135_), .A2(new_n19138_), .A3(new_n19133_), .A4(new_n19117_), .ZN(new_n19139_));
  NAND2_X1   g16041(.A1(new_n19132_), .A2(new_n19139_), .ZN(new_n19140_));
  AOI21_X1   g16042(.A1(new_n19140_), .A2(new_n19115_), .B(new_n17392_), .ZN(new_n19141_));
  NOR2_X1    g16043(.A1(new_n19069_), .A2(new_n13613_), .ZN(new_n19142_));
  XOR2_X1    g16044(.A1(new_n19142_), .A2(new_n13615_), .Z(new_n19143_));
  NAND2_X1   g16045(.A1(new_n19143_), .A2(new_n19141_), .ZN(new_n19144_));
  AOI21_X1   g16046(.A1(new_n19108_), .A2(new_n19102_), .B(pi0608), .ZN(new_n19145_));
  NAND2_X1   g16047(.A1(new_n19105_), .A2(new_n14081_), .ZN(new_n19146_));
  AOI21_X1   g16048(.A1(new_n19144_), .A2(new_n19145_), .B(new_n19146_), .ZN(new_n19147_));
  NOR2_X1    g16049(.A1(new_n19069_), .A2(new_n13614_), .ZN(new_n19148_));
  XOR2_X1    g16050(.A1(new_n19148_), .A2(new_n13615_), .Z(new_n19149_));
  NAND3_X1   g16051(.A1(new_n19149_), .A2(new_n19141_), .A3(pi0778), .ZN(new_n19150_));
  OAI22_X1   g16052(.A1(new_n19147_), .A2(new_n19150_), .B1(pi0778), .B2(new_n19141_), .ZN(new_n19151_));
  NAND3_X1   g16053(.A1(new_n19151_), .A2(pi0609), .A3(pi1155), .ZN(new_n19152_));
  INV_X1     g16054(.I(new_n19151_), .ZN(new_n19153_));
  NAND3_X1   g16055(.A1(new_n19153_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n19154_));
  AOI21_X1   g16056(.A1(new_n19154_), .A2(new_n19152_), .B(new_n19111_), .ZN(new_n19155_));
  NAND2_X1   g16057(.A1(new_n19067_), .A2(pi0660), .ZN(new_n19156_));
  NAND2_X1   g16058(.A1(new_n19073_), .A2(new_n13783_), .ZN(new_n19157_));
  INV_X1     g16059(.I(new_n19157_), .ZN(new_n19158_));
  OAI21_X1   g16060(.A1(new_n19155_), .A2(new_n19156_), .B(new_n19158_), .ZN(new_n19159_));
  AOI21_X1   g16061(.A1(new_n19153_), .A2(pi0609), .B(new_n14694_), .ZN(new_n19160_));
  NOR3_X1    g16062(.A1(new_n19151_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n19161_));
  NOR2_X1    g16063(.A1(new_n19111_), .A2(new_n13801_), .ZN(new_n19162_));
  OAI21_X1   g16064(.A1(new_n19160_), .A2(new_n19161_), .B(new_n19162_), .ZN(new_n19163_));
  INV_X1     g16065(.I(new_n19163_), .ZN(new_n19164_));
  AOI22_X1   g16066(.A1(new_n19159_), .A2(new_n19164_), .B1(new_n13801_), .B2(new_n19151_), .ZN(new_n19165_));
  AOI21_X1   g16067(.A1(new_n19165_), .A2(pi1154), .B(new_n13819_), .ZN(new_n19166_));
  INV_X1     g16068(.I(new_n19165_), .ZN(new_n19167_));
  NOR3_X1    g16069(.A1(new_n19167_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n19168_));
  OAI21_X1   g16070(.A1(new_n19168_), .A2(new_n19166_), .B(new_n19113_), .ZN(new_n19169_));
  NAND2_X1   g16071(.A1(new_n19080_), .A2(pi0627), .ZN(new_n19170_));
  INV_X1     g16072(.I(new_n19170_), .ZN(new_n19171_));
  AOI21_X1   g16073(.A1(new_n19169_), .A2(new_n19171_), .B(new_n13855_), .ZN(new_n19172_));
  NAND3_X1   g16074(.A1(new_n19167_), .A2(pi0618), .A3(pi1154), .ZN(new_n19173_));
  NAND3_X1   g16075(.A1(new_n19165_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n19174_));
  NAND2_X1   g16076(.A1(new_n19173_), .A2(new_n19174_), .ZN(new_n19175_));
  AND2_X2    g16077(.A1(new_n19175_), .A2(new_n19113_), .Z(new_n19176_));
  NOR2_X1    g16078(.A1(new_n13855_), .A2(pi0627), .ZN(new_n19177_));
  NAND3_X1   g16079(.A1(new_n19167_), .A2(new_n19085_), .A3(new_n19177_), .ZN(new_n19178_));
  NOR3_X1    g16080(.A1(new_n19176_), .A2(new_n19172_), .A3(new_n19178_), .ZN(new_n19179_));
  INV_X1     g16081(.I(new_n19172_), .ZN(new_n19180_));
  NOR2_X1    g16082(.A1(new_n19176_), .A2(new_n19178_), .ZN(new_n19181_));
  NOR2_X1    g16083(.A1(new_n19181_), .A2(new_n19180_), .ZN(new_n19182_));
  NOR2_X1    g16084(.A1(new_n19182_), .A2(new_n19179_), .ZN(new_n19183_));
  AOI21_X1   g16085(.A1(new_n19183_), .A2(pi1159), .B(new_n13904_), .ZN(new_n19184_));
  NOR4_X1    g16086(.A1(new_n19182_), .A2(pi0619), .A3(new_n13868_), .A4(new_n19179_), .ZN(new_n19185_));
  OAI21_X1   g16087(.A1(new_n19184_), .A2(new_n19185_), .B(new_n19114_), .ZN(new_n19186_));
  NAND2_X1   g16088(.A1(new_n19186_), .A2(new_n16474_), .ZN(new_n19187_));
  NAND3_X1   g16089(.A1(new_n19089_), .A2(pi0619), .A3(pi1159), .ZN(new_n19188_));
  NAND4_X1   g16090(.A1(new_n19088_), .A2(new_n13860_), .A3(pi1159), .A4(new_n19087_), .ZN(new_n19189_));
  AOI21_X1   g16091(.A1(new_n19188_), .A2(new_n19189_), .B(new_n19051_), .ZN(new_n19190_));
  NAND4_X1   g16092(.A1(new_n19093_), .A2(pi0789), .A3(new_n19190_), .A4(new_n19089_), .ZN(new_n19191_));
  NOR2_X1    g16093(.A1(new_n19093_), .A2(new_n13896_), .ZN(new_n19192_));
  NAND3_X1   g16094(.A1(new_n19190_), .A2(pi0789), .A3(new_n19089_), .ZN(new_n19193_));
  NAND2_X1   g16095(.A1(new_n19192_), .A2(new_n19193_), .ZN(new_n19194_));
  NAND2_X1   g16096(.A1(new_n19194_), .A2(new_n19191_), .ZN(new_n19195_));
  NAND3_X1   g16097(.A1(new_n19195_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n19196_));
  INV_X1     g16098(.I(new_n19195_), .ZN(new_n19197_));
  NAND3_X1   g16099(.A1(new_n19197_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n19198_));
  AOI21_X1   g16100(.A1(new_n19198_), .A2(new_n19196_), .B(new_n19051_), .ZN(new_n19199_));
  NOR2_X1    g16101(.A1(new_n19114_), .A2(new_n13918_), .ZN(new_n19200_));
  AOI21_X1   g16102(.A1(new_n13918_), .A2(new_n19050_), .B(new_n19200_), .ZN(new_n19201_));
  NOR2_X1    g16103(.A1(new_n19201_), .A2(new_n14162_), .ZN(new_n19202_));
  NOR2_X1    g16104(.A1(new_n16424_), .A2(new_n13937_), .ZN(new_n19203_));
  INV_X1     g16105(.I(new_n19203_), .ZN(new_n19204_));
  OAI21_X1   g16106(.A1(new_n19199_), .A2(new_n19202_), .B(new_n19204_), .ZN(new_n19205_));
  NOR2_X1    g16107(.A1(new_n19183_), .A2(pi0789), .ZN(new_n19206_));
  AOI21_X1   g16108(.A1(new_n19197_), .A2(new_n13963_), .B(new_n19028_), .ZN(new_n19207_));
  INV_X1     g16109(.I(new_n13963_), .ZN(new_n19208_));
  NOR3_X1    g16110(.A1(new_n19195_), .A2(pi0626), .A3(new_n19208_), .ZN(new_n19209_));
  NOR2_X1    g16111(.A1(new_n19207_), .A2(new_n19209_), .ZN(new_n19210_));
  NOR4_X1    g16112(.A1(new_n19210_), .A2(new_n15479_), .A3(new_n19051_), .A4(new_n19206_), .ZN(new_n19211_));
  AOI22_X1   g16113(.A1(new_n19187_), .A2(new_n19093_), .B1(new_n19211_), .B2(new_n19205_), .ZN(new_n19212_));
  AOI21_X1   g16114(.A1(new_n19183_), .A2(pi0619), .B(new_n13904_), .ZN(new_n19213_));
  NOR4_X1    g16115(.A1(new_n19182_), .A2(new_n13860_), .A3(pi1159), .A4(new_n19179_), .ZN(new_n19214_));
  OAI21_X1   g16116(.A1(new_n19213_), .A2(new_n19214_), .B(new_n19114_), .ZN(new_n19215_));
  NOR2_X1    g16117(.A1(new_n19190_), .A2(pi0648), .ZN(new_n19216_));
  NAND2_X1   g16118(.A1(new_n19215_), .A2(new_n19216_), .ZN(new_n19217_));
  NOR2_X1    g16119(.A1(new_n19050_), .A2(new_n16372_), .ZN(new_n19218_));
  INV_X1     g16120(.I(new_n19218_), .ZN(new_n19219_));
  NAND3_X1   g16121(.A1(new_n19194_), .A2(new_n19191_), .A3(new_n16372_), .ZN(new_n19220_));
  AOI21_X1   g16122(.A1(new_n19220_), .A2(new_n19219_), .B(new_n13993_), .ZN(new_n19221_));
  NOR2_X1    g16123(.A1(new_n19050_), .A2(new_n13994_), .ZN(new_n19222_));
  OR2_X2     g16124(.A1(new_n19221_), .A2(new_n19222_), .Z(new_n19223_));
  NAND2_X1   g16125(.A1(new_n19201_), .A2(new_n13966_), .ZN(new_n19224_));
  OAI21_X1   g16126(.A1(new_n13966_), .A2(new_n19050_), .B(new_n19224_), .ZN(new_n19225_));
  NAND2_X1   g16127(.A1(new_n19225_), .A2(new_n12777_), .ZN(new_n19226_));
  NOR2_X1    g16128(.A1(new_n19050_), .A2(new_n13942_), .ZN(new_n19227_));
  AOI21_X1   g16129(.A1(new_n19225_), .A2(new_n13942_), .B(new_n19227_), .ZN(new_n19228_));
  NOR2_X1    g16130(.A1(new_n19228_), .A2(pi1156), .ZN(new_n19229_));
  NOR2_X1    g16131(.A1(new_n19050_), .A2(pi0628), .ZN(new_n19230_));
  AOI21_X1   g16132(.A1(new_n19225_), .A2(pi0628), .B(new_n19230_), .ZN(new_n19231_));
  NOR2_X1    g16133(.A1(new_n19231_), .A2(new_n13969_), .ZN(new_n19232_));
  OAI21_X1   g16134(.A1(new_n19229_), .A2(new_n19232_), .B(pi0792), .ZN(new_n19233_));
  NAND2_X1   g16135(.A1(new_n19233_), .A2(new_n19226_), .ZN(new_n19234_));
  NAND2_X1   g16136(.A1(new_n19234_), .A2(new_n14005_), .ZN(new_n19235_));
  NAND2_X1   g16137(.A1(new_n19051_), .A2(pi0647), .ZN(new_n19236_));
  AOI21_X1   g16138(.A1(new_n19235_), .A2(new_n19236_), .B(new_n14012_), .ZN(new_n19237_));
  NOR2_X1    g16139(.A1(new_n19050_), .A2(pi0647), .ZN(new_n19238_));
  AOI21_X1   g16140(.A1(new_n19234_), .A2(pi0647), .B(new_n19238_), .ZN(new_n19239_));
  NAND2_X1   g16141(.A1(new_n19239_), .A2(new_n14206_), .ZN(new_n19240_));
  OR2_X2     g16142(.A1(new_n19237_), .A2(new_n19240_), .Z(new_n19241_));
  NAND2_X1   g16143(.A1(new_n19237_), .A2(new_n19240_), .ZN(new_n19242_));
  AOI21_X1   g16144(.A1(new_n19241_), .A2(new_n19242_), .B(new_n12776_), .ZN(new_n19243_));
  NOR2_X1    g16145(.A1(new_n19223_), .A2(new_n19243_), .ZN(new_n19244_));
  OAI22_X1   g16146(.A1(new_n19212_), .A2(new_n19217_), .B1(new_n16891_), .B2(new_n19244_), .ZN(new_n19245_));
  AOI21_X1   g16147(.A1(new_n19197_), .A2(new_n16372_), .B(new_n19218_), .ZN(new_n19246_));
  NOR2_X1    g16148(.A1(new_n19228_), .A2(new_n15270_), .ZN(new_n19247_));
  NAND2_X1   g16149(.A1(new_n19231_), .A2(new_n13990_), .ZN(new_n19248_));
  XNOR2_X1   g16150(.A1(new_n19247_), .A2(new_n19248_), .ZN(new_n19249_));
  NAND2_X1   g16151(.A1(new_n19249_), .A2(pi0792), .ZN(new_n19250_));
  AOI21_X1   g16152(.A1(new_n19246_), .A2(new_n19250_), .B(new_n16875_), .ZN(new_n19251_));
  NAND2_X1   g16153(.A1(new_n19234_), .A2(new_n12776_), .ZN(new_n19252_));
  AOI21_X1   g16154(.A1(new_n19235_), .A2(new_n19236_), .B(pi1157), .ZN(new_n19253_));
  NOR2_X1    g16155(.A1(new_n19239_), .A2(new_n14006_), .ZN(new_n19254_));
  OAI21_X1   g16156(.A1(new_n19254_), .A2(new_n19253_), .B(pi0787), .ZN(new_n19255_));
  NAND2_X1   g16157(.A1(new_n19255_), .A2(new_n19252_), .ZN(new_n19256_));
  INV_X1     g16158(.I(new_n19256_), .ZN(new_n19257_));
  OAI21_X1   g16159(.A1(new_n19221_), .A2(new_n19222_), .B(new_n14211_), .ZN(new_n19258_));
  NOR2_X1    g16160(.A1(new_n19050_), .A2(new_n14211_), .ZN(new_n19259_));
  INV_X1     g16161(.I(new_n19259_), .ZN(new_n19260_));
  NOR2_X1    g16162(.A1(new_n14243_), .A2(pi0644), .ZN(new_n19261_));
  AOI21_X1   g16163(.A1(new_n19258_), .A2(new_n19260_), .B(new_n19261_), .ZN(new_n19262_));
  AOI21_X1   g16164(.A1(new_n19262_), .A2(pi0715), .B(pi0644), .ZN(new_n19263_));
  AOI21_X1   g16165(.A1(new_n19050_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n19264_));
  NOR2_X1    g16166(.A1(new_n19264_), .A2(pi0644), .ZN(new_n19265_));
  AOI21_X1   g16167(.A1(new_n19258_), .A2(new_n19260_), .B(new_n19265_), .ZN(new_n19266_));
  AOI21_X1   g16168(.A1(new_n19266_), .A2(pi0715), .B(new_n19256_), .ZN(new_n19267_));
  OAI22_X1   g16169(.A1(new_n14204_), .A2(new_n19267_), .B1(new_n19263_), .B2(new_n19257_), .ZN(new_n19268_));
  NOR2_X1    g16170(.A1(new_n7240_), .A2(new_n12775_), .ZN(new_n19269_));
  AOI22_X1   g16171(.A1(new_n19245_), .A2(new_n19251_), .B1(new_n19268_), .B2(new_n19269_), .ZN(new_n19270_));
  AOI21_X1   g16172(.A1(new_n19223_), .A2(new_n14211_), .B(new_n19259_), .ZN(new_n19271_));
  NOR3_X1    g16173(.A1(new_n19271_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n19272_));
  NOR3_X1    g16174(.A1(new_n19266_), .A2(pi0644), .A3(new_n12775_), .ZN(new_n19273_));
  NOR2_X1    g16175(.A1(new_n19037_), .A2(pi0790), .ZN(new_n19274_));
  NOR4_X1    g16176(.A1(new_n19271_), .A2(new_n14799_), .A3(new_n19261_), .A4(new_n19274_), .ZN(new_n19275_));
  OAI21_X1   g16177(.A1(new_n19272_), .A2(new_n19273_), .B(new_n19275_), .ZN(new_n19276_));
  OAI21_X1   g16178(.A1(new_n19270_), .A2(new_n19276_), .B(new_n19049_), .ZN(po0332));
  NOR2_X1    g16179(.A1(new_n14428_), .A2(pi0176), .ZN(new_n19278_));
  NOR2_X1    g16180(.A1(new_n19278_), .A2(new_n13880_), .ZN(new_n19279_));
  NAND2_X1   g16181(.A1(new_n14422_), .A2(new_n13723_), .ZN(new_n19280_));
  XNOR2_X1   g16182(.A1(new_n19280_), .A2(new_n16146_), .ZN(new_n19281_));
  NOR3_X1    g16183(.A1(new_n3289_), .A2(pi0176), .A3(pi0704), .ZN(new_n19282_));
  NOR3_X1    g16184(.A1(new_n14396_), .A2(new_n17414_), .A3(new_n19282_), .ZN(new_n19283_));
  NOR2_X1    g16185(.A1(new_n19281_), .A2(new_n19283_), .ZN(new_n19284_));
  AOI21_X1   g16186(.A1(new_n14404_), .A2(new_n3289_), .B(new_n16715_), .ZN(new_n19285_));
  NOR3_X1    g16187(.A1(new_n15655_), .A2(pi0038), .A3(new_n3290_), .ZN(new_n19286_));
  OAI21_X1   g16188(.A1(new_n19285_), .A2(new_n19286_), .B(new_n13719_), .ZN(new_n19287_));
  INV_X1     g16189(.I(new_n19287_), .ZN(new_n19288_));
  AOI21_X1   g16190(.A1(new_n19284_), .A2(new_n19288_), .B(new_n7459_), .ZN(new_n19289_));
  NAND2_X1   g16191(.A1(new_n19289_), .A2(pi0625), .ZN(new_n19290_));
  XOR2_X1    g16192(.A1(new_n19290_), .A2(new_n13620_), .Z(new_n19291_));
  NAND2_X1   g16193(.A1(new_n19291_), .A2(new_n19278_), .ZN(new_n19292_));
  NAND2_X1   g16194(.A1(new_n19292_), .A2(pi0778), .ZN(new_n19293_));
  NAND2_X1   g16195(.A1(new_n19289_), .A2(pi1153), .ZN(new_n19294_));
  XOR2_X1    g16196(.A1(new_n19294_), .A2(new_n13620_), .Z(new_n19295_));
  NAND2_X1   g16197(.A1(new_n19295_), .A2(new_n19278_), .ZN(new_n19296_));
  NOR3_X1    g16198(.A1(new_n19296_), .A2(new_n13748_), .A3(new_n19289_), .ZN(new_n19297_));
  XNOR2_X1   g16199(.A1(new_n19297_), .A2(new_n19293_), .ZN(new_n19298_));
  INV_X1     g16200(.I(new_n19278_), .ZN(new_n19299_));
  NOR2_X1    g16201(.A1(new_n19299_), .A2(new_n13805_), .ZN(new_n19300_));
  AOI21_X1   g16202(.A1(new_n19298_), .A2(new_n13805_), .B(new_n19300_), .ZN(new_n19301_));
  AOI21_X1   g16203(.A1(new_n19301_), .A2(new_n13880_), .B(new_n19279_), .ZN(new_n19302_));
  NAND2_X1   g16204(.A1(new_n19302_), .A2(new_n15395_), .ZN(new_n19303_));
  NAND2_X1   g16205(.A1(new_n19278_), .A2(new_n15395_), .ZN(new_n19304_));
  XOR2_X1    g16206(.A1(new_n19303_), .A2(new_n19304_), .Z(new_n19305_));
  NAND2_X1   g16207(.A1(new_n19305_), .A2(new_n12777_), .ZN(new_n19306_));
  NOR2_X1    g16208(.A1(new_n19305_), .A2(new_n14057_), .ZN(new_n19307_));
  NOR2_X1    g16209(.A1(new_n19299_), .A2(new_n14057_), .ZN(new_n19308_));
  XNOR2_X1   g16210(.A1(new_n19307_), .A2(new_n19308_), .ZN(new_n19309_));
  OAI21_X1   g16211(.A1(new_n19309_), .A2(new_n12777_), .B(new_n19306_), .ZN(new_n19310_));
  AND2_X2    g16212(.A1(new_n19310_), .A2(new_n12776_), .Z(new_n19311_));
  NOR2_X1    g16213(.A1(new_n19278_), .A2(new_n14005_), .ZN(new_n19312_));
  AOI21_X1   g16214(.A1(new_n19310_), .A2(new_n14005_), .B(new_n19312_), .ZN(new_n19313_));
  OR2_X2     g16215(.A1(new_n19313_), .A2(pi1157), .Z(new_n19314_));
  NOR2_X1    g16216(.A1(new_n19278_), .A2(pi0647), .ZN(new_n19315_));
  AOI21_X1   g16217(.A1(new_n19310_), .A2(pi0647), .B(new_n19315_), .ZN(new_n19316_));
  OAI21_X1   g16218(.A1(new_n14006_), .A2(new_n19316_), .B(new_n19314_), .ZN(new_n19317_));
  AOI21_X1   g16219(.A1(new_n19317_), .A2(pi0787), .B(new_n19311_), .ZN(new_n19318_));
  NOR2_X1    g16220(.A1(new_n19278_), .A2(new_n16372_), .ZN(new_n19319_));
  NOR2_X1    g16221(.A1(new_n13634_), .A2(new_n17409_), .ZN(new_n19320_));
  NOR2_X1    g16222(.A1(new_n7499_), .A2(new_n13105_), .ZN(new_n19321_));
  NOR2_X1    g16223(.A1(new_n19321_), .A2(new_n3259_), .ZN(new_n19322_));
  AOI21_X1   g16224(.A1(new_n15562_), .A2(new_n3259_), .B(new_n19322_), .ZN(new_n19323_));
  NAND2_X1   g16225(.A1(new_n19323_), .A2(pi0176), .ZN(new_n19324_));
  NAND3_X1   g16226(.A1(new_n14355_), .A2(new_n14356_), .A3(new_n14360_), .ZN(new_n19325_));
  OAI21_X1   g16227(.A1(new_n14348_), .A2(new_n14338_), .B(new_n14330_), .ZN(new_n19326_));
  NAND2_X1   g16228(.A1(new_n19325_), .A2(new_n19326_), .ZN(new_n19327_));
  INV_X1     g16229(.I(new_n15555_), .ZN(new_n19328_));
  OAI21_X1   g16230(.A1(new_n19327_), .A2(pi0038), .B(new_n19328_), .ZN(new_n19329_));
  NAND2_X1   g16231(.A1(new_n19329_), .A2(new_n7459_), .ZN(new_n19330_));
  NAND2_X1   g16232(.A1(pi0176), .A2(pi0742), .ZN(new_n19331_));
  AOI21_X1   g16233(.A1(new_n19324_), .A2(new_n19330_), .B(new_n19331_), .ZN(new_n19332_));
  XOR2_X1    g16234(.A1(new_n19332_), .A2(new_n19320_), .Z(new_n19333_));
  NAND2_X1   g16235(.A1(new_n19333_), .A2(new_n3289_), .ZN(new_n19334_));
  OAI21_X1   g16236(.A1(pi0176), .A2(new_n3289_), .B(new_n19334_), .ZN(new_n19335_));
  NOR2_X1    g16237(.A1(new_n19335_), .A2(new_n13775_), .ZN(new_n19336_));
  NOR2_X1    g16238(.A1(new_n19278_), .A2(new_n15147_), .ZN(new_n19337_));
  OAI21_X1   g16239(.A1(new_n19336_), .A2(new_n19337_), .B(pi0609), .ZN(new_n19338_));
  NAND2_X1   g16240(.A1(new_n19338_), .A2(pi0785), .ZN(new_n19339_));
  NOR2_X1    g16241(.A1(new_n19299_), .A2(new_n13776_), .ZN(new_n19340_));
  AOI21_X1   g16242(.A1(new_n19335_), .A2(new_n13776_), .B(new_n19340_), .ZN(new_n19341_));
  AOI21_X1   g16243(.A1(new_n19299_), .A2(new_n14467_), .B(pi0609), .ZN(new_n19342_));
  INV_X1     g16244(.I(new_n19342_), .ZN(new_n19343_));
  NAND2_X1   g16245(.A1(new_n19336_), .A2(new_n19343_), .ZN(new_n19344_));
  NOR3_X1    g16246(.A1(new_n19344_), .A2(new_n13801_), .A3(new_n19341_), .ZN(new_n19345_));
  XOR2_X1    g16247(.A1(new_n19345_), .A2(new_n19339_), .Z(new_n19346_));
  NAND2_X1   g16248(.A1(new_n19346_), .A2(pi0618), .ZN(new_n19347_));
  XOR2_X1    g16249(.A1(new_n19347_), .A2(new_n13819_), .Z(new_n19348_));
  NAND2_X1   g16250(.A1(new_n19348_), .A2(new_n19278_), .ZN(new_n19349_));
  NAND2_X1   g16251(.A1(new_n19349_), .A2(pi0781), .ZN(new_n19350_));
  AND2_X2    g16252(.A1(new_n19346_), .A2(pi1154), .Z(new_n19351_));
  XOR2_X1    g16253(.A1(new_n19351_), .A2(new_n13819_), .Z(new_n19352_));
  NOR2_X1    g16254(.A1(new_n19352_), .A2(new_n19299_), .ZN(new_n19353_));
  NOR2_X1    g16255(.A1(new_n19346_), .A2(new_n13855_), .ZN(new_n19354_));
  NAND2_X1   g16256(.A1(new_n19353_), .A2(new_n19354_), .ZN(new_n19355_));
  XOR2_X1    g16257(.A1(new_n19355_), .A2(new_n19350_), .Z(new_n19356_));
  INV_X1     g16258(.I(new_n19356_), .ZN(new_n19357_));
  NOR2_X1    g16259(.A1(new_n19357_), .A2(pi0789), .ZN(new_n19358_));
  NAND3_X1   g16260(.A1(new_n19356_), .A2(new_n16697_), .A3(new_n19278_), .ZN(new_n19359_));
  NAND3_X1   g16261(.A1(new_n19350_), .A2(new_n16697_), .A3(new_n19299_), .ZN(new_n19360_));
  AOI21_X1   g16262(.A1(new_n19359_), .A2(new_n19360_), .B(new_n13896_), .ZN(new_n19361_));
  NOR3_X1    g16263(.A1(new_n19361_), .A2(new_n14142_), .A3(new_n19358_), .ZN(new_n19362_));
  NOR2_X1    g16264(.A1(new_n19362_), .A2(new_n19319_), .ZN(new_n19363_));
  NOR2_X1    g16265(.A1(new_n19363_), .A2(new_n13993_), .ZN(new_n19364_));
  NOR2_X1    g16266(.A1(new_n19278_), .A2(new_n13994_), .ZN(new_n19365_));
  NOR2_X1    g16267(.A1(new_n19364_), .A2(new_n19365_), .ZN(new_n19366_));
  NOR2_X1    g16268(.A1(new_n19278_), .A2(new_n14211_), .ZN(new_n19367_));
  INV_X1     g16269(.I(new_n19367_), .ZN(new_n19368_));
  OAI21_X1   g16270(.A1(new_n19366_), .A2(new_n14210_), .B(new_n19368_), .ZN(new_n19369_));
  INV_X1     g16271(.I(new_n14243_), .ZN(new_n19370_));
  NAND2_X1   g16272(.A1(new_n19370_), .A2(new_n14204_), .ZN(new_n19371_));
  AND2_X2    g16273(.A1(new_n19369_), .A2(new_n19371_), .Z(new_n19372_));
  NAND2_X1   g16274(.A1(new_n19372_), .A2(pi0715), .ZN(new_n19373_));
  AOI21_X1   g16275(.A1(new_n19373_), .A2(new_n14204_), .B(new_n19318_), .ZN(new_n19374_));
  OAI21_X1   g16276(.A1(new_n19278_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n19375_));
  NAND3_X1   g16277(.A1(new_n19369_), .A2(pi0715), .A3(new_n19375_), .ZN(new_n19376_));
  AOI21_X1   g16278(.A1(new_n19376_), .A2(new_n19318_), .B(new_n14204_), .ZN(new_n19377_));
  OAI21_X1   g16279(.A1(new_n19374_), .A2(new_n19377_), .B(pi0790), .ZN(new_n19378_));
  NOR2_X1    g16280(.A1(new_n14204_), .A2(new_n12775_), .ZN(new_n19379_));
  AOI21_X1   g16281(.A1(new_n19369_), .A2(new_n19375_), .B(new_n12775_), .ZN(new_n19380_));
  XOR2_X1    g16282(.A1(new_n19380_), .A2(new_n19379_), .Z(new_n19381_));
  NOR2_X1    g16283(.A1(new_n19313_), .A2(new_n14012_), .ZN(new_n19382_));
  NAND2_X1   g16284(.A1(new_n19316_), .A2(new_n14206_), .ZN(new_n19383_));
  XNOR2_X1   g16285(.A1(new_n19382_), .A2(new_n19383_), .ZN(new_n19384_));
  NAND2_X1   g16286(.A1(new_n19384_), .A2(pi0787), .ZN(new_n19385_));
  AOI21_X1   g16287(.A1(new_n19385_), .A2(new_n19366_), .B(new_n16867_), .ZN(new_n19386_));
  AOI21_X1   g16288(.A1(new_n19381_), .A2(new_n19372_), .B(new_n19386_), .ZN(new_n19387_));
  AOI21_X1   g16289(.A1(new_n19333_), .A2(pi0704), .B(new_n3290_), .ZN(new_n19388_));
  INV_X1     g16290(.I(new_n19388_), .ZN(new_n19389_));
  NOR2_X1    g16291(.A1(new_n15615_), .A2(new_n15629_), .ZN(new_n19390_));
  NAND2_X1   g16292(.A1(new_n15595_), .A2(pi0742), .ZN(new_n19391_));
  XOR2_X1    g16293(.A1(new_n19391_), .A2(new_n19331_), .Z(new_n19392_));
  NOR3_X1    g16294(.A1(new_n15625_), .A2(new_n15616_), .A3(new_n15626_), .ZN(new_n19393_));
  AOI21_X1   g16295(.A1(new_n15619_), .A2(new_n15622_), .B(new_n15617_), .ZN(new_n19394_));
  NOR2_X1    g16296(.A1(new_n19394_), .A2(new_n19393_), .ZN(new_n19395_));
  NAND2_X1   g16297(.A1(new_n19395_), .A2(pi0176), .ZN(new_n19396_));
  XOR2_X1    g16298(.A1(new_n19396_), .A2(new_n19331_), .Z(new_n19397_));
  NAND2_X1   g16299(.A1(new_n19397_), .A2(new_n15607_), .ZN(new_n19398_));
  NAND4_X1   g16300(.A1(new_n19398_), .A2(pi0176), .A3(new_n17414_), .A4(new_n3289_), .ZN(new_n19399_));
  AOI21_X1   g16301(.A1(new_n19390_), .A2(new_n19392_), .B(new_n19399_), .ZN(new_n19400_));
  NAND2_X1   g16302(.A1(new_n19400_), .A2(new_n19389_), .ZN(new_n19401_));
  AND2_X2    g16303(.A1(new_n19392_), .A2(new_n19390_), .Z(new_n19402_));
  OAI21_X1   g16304(.A1(new_n19402_), .A2(new_n19399_), .B(new_n19388_), .ZN(new_n19403_));
  NAND2_X1   g16305(.A1(new_n19403_), .A2(new_n19401_), .ZN(new_n19404_));
  NOR2_X1    g16306(.A1(new_n19404_), .A2(new_n13613_), .ZN(new_n19405_));
  XOR2_X1    g16307(.A1(new_n19405_), .A2(new_n13615_), .Z(new_n19406_));
  NAND2_X1   g16308(.A1(new_n19406_), .A2(new_n19335_), .ZN(new_n19407_));
  NAND3_X1   g16309(.A1(new_n19407_), .A2(new_n14081_), .A3(new_n19296_), .ZN(new_n19408_));
  NOR2_X1    g16310(.A1(new_n19404_), .A2(new_n13614_), .ZN(new_n19409_));
  XOR2_X1    g16311(.A1(new_n19409_), .A2(new_n13615_), .Z(new_n19410_));
  AOI21_X1   g16312(.A1(new_n19410_), .A2(new_n19335_), .B(pi0608), .ZN(new_n19411_));
  NAND2_X1   g16313(.A1(new_n19408_), .A2(new_n19411_), .ZN(new_n19412_));
  NAND4_X1   g16314(.A1(new_n19412_), .A2(pi0778), .A3(new_n19278_), .A4(new_n19291_), .ZN(new_n19413_));
  NAND3_X1   g16315(.A1(new_n19403_), .A2(new_n19401_), .A3(new_n13748_), .ZN(new_n19414_));
  NAND2_X1   g16316(.A1(new_n19413_), .A2(new_n19414_), .ZN(new_n19415_));
  NAND2_X1   g16317(.A1(new_n19415_), .A2(new_n13801_), .ZN(new_n19416_));
  NAND3_X1   g16318(.A1(new_n19415_), .A2(pi0609), .A3(pi1155), .ZN(new_n19417_));
  INV_X1     g16319(.I(new_n19417_), .ZN(new_n19418_));
  NOR3_X1    g16320(.A1(new_n19415_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n19419_));
  OAI21_X1   g16321(.A1(new_n19418_), .A2(new_n19419_), .B(new_n19298_), .ZN(new_n19420_));
  NAND2_X1   g16322(.A1(new_n19338_), .A2(pi0660), .ZN(new_n19421_));
  INV_X1     g16323(.I(new_n19421_), .ZN(new_n19422_));
  NAND2_X1   g16324(.A1(new_n19344_), .A2(new_n13783_), .ZN(new_n19423_));
  AOI21_X1   g16325(.A1(new_n19420_), .A2(new_n19422_), .B(new_n19423_), .ZN(new_n19424_));
  NOR2_X1    g16326(.A1(new_n19415_), .A2(new_n13766_), .ZN(new_n19425_));
  NOR2_X1    g16327(.A1(new_n19425_), .A2(new_n14694_), .ZN(new_n19426_));
  NAND2_X1   g16328(.A1(new_n19425_), .A2(new_n14694_), .ZN(new_n19427_));
  INV_X1     g16329(.I(new_n19427_), .ZN(new_n19428_));
  INV_X1     g16330(.I(new_n19298_), .ZN(new_n19429_));
  NOR2_X1    g16331(.A1(new_n19429_), .A2(new_n13801_), .ZN(new_n19430_));
  OAI21_X1   g16332(.A1(new_n19428_), .A2(new_n19426_), .B(new_n19430_), .ZN(new_n19431_));
  OAI21_X1   g16333(.A1(new_n19424_), .A2(new_n19431_), .B(new_n19416_), .ZN(new_n19432_));
  NAND3_X1   g16334(.A1(new_n19432_), .A2(pi0618), .A3(pi1154), .ZN(new_n19433_));
  INV_X1     g16335(.I(new_n19415_), .ZN(new_n19434_));
  NAND3_X1   g16336(.A1(new_n19434_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n19435_));
  AOI21_X1   g16337(.A1(new_n19435_), .A2(new_n19417_), .B(new_n19429_), .ZN(new_n19436_));
  INV_X1     g16338(.I(new_n19423_), .ZN(new_n19437_));
  OAI21_X1   g16339(.A1(new_n19436_), .A2(new_n19421_), .B(new_n19437_), .ZN(new_n19438_));
  INV_X1     g16340(.I(new_n19426_), .ZN(new_n19439_));
  INV_X1     g16341(.I(new_n19430_), .ZN(new_n19440_));
  AOI21_X1   g16342(.A1(new_n19439_), .A2(new_n19427_), .B(new_n19440_), .ZN(new_n19441_));
  AOI22_X1   g16343(.A1(new_n19438_), .A2(new_n19441_), .B1(new_n13801_), .B2(new_n19415_), .ZN(new_n19442_));
  NAND3_X1   g16344(.A1(new_n19442_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n19443_));
  AOI21_X1   g16345(.A1(new_n19443_), .A2(new_n19433_), .B(new_n19301_), .ZN(new_n19444_));
  NAND2_X1   g16346(.A1(new_n19349_), .A2(pi0627), .ZN(new_n19445_));
  OAI21_X1   g16347(.A1(new_n19444_), .A2(new_n19445_), .B(pi0781), .ZN(new_n19446_));
  INV_X1     g16348(.I(new_n19301_), .ZN(new_n19447_));
  NAND3_X1   g16349(.A1(new_n19432_), .A2(pi0618), .A3(pi1154), .ZN(new_n19448_));
  NAND3_X1   g16350(.A1(new_n19442_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n19449_));
  NAND2_X1   g16351(.A1(new_n19449_), .A2(new_n19448_), .ZN(new_n19450_));
  INV_X1     g16352(.I(new_n19353_), .ZN(new_n19451_));
  NAND3_X1   g16353(.A1(new_n19432_), .A2(new_n19177_), .A3(new_n19451_), .ZN(new_n19452_));
  AOI21_X1   g16354(.A1(new_n19450_), .A2(new_n19447_), .B(new_n19452_), .ZN(new_n19453_));
  NAND2_X1   g16355(.A1(new_n19446_), .A2(new_n19453_), .ZN(new_n19454_));
  AOI21_X1   g16356(.A1(new_n19442_), .A2(pi1154), .B(new_n13819_), .ZN(new_n19455_));
  NOR3_X1    g16357(.A1(new_n19432_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n19456_));
  OAI21_X1   g16358(.A1(new_n19455_), .A2(new_n19456_), .B(new_n19447_), .ZN(new_n19457_));
  INV_X1     g16359(.I(new_n19445_), .ZN(new_n19458_));
  AOI21_X1   g16360(.A1(new_n19457_), .A2(new_n19458_), .B(new_n13855_), .ZN(new_n19459_));
  AOI21_X1   g16361(.A1(new_n19442_), .A2(pi0618), .B(new_n13819_), .ZN(new_n19460_));
  NOR3_X1    g16362(.A1(new_n19432_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n19461_));
  OAI21_X1   g16363(.A1(new_n19460_), .A2(new_n19461_), .B(new_n19447_), .ZN(new_n19462_));
  NAND4_X1   g16364(.A1(new_n19462_), .A2(new_n19177_), .A3(new_n19451_), .A4(new_n19432_), .ZN(new_n19463_));
  NAND2_X1   g16365(.A1(new_n19463_), .A2(new_n19459_), .ZN(new_n19464_));
  NAND2_X1   g16366(.A1(new_n19464_), .A2(new_n19454_), .ZN(new_n19465_));
  AOI21_X1   g16367(.A1(new_n19465_), .A2(new_n13896_), .B(new_n15479_), .ZN(new_n19466_));
  XOR2_X1    g16368(.A1(new_n19446_), .A2(new_n19453_), .Z(new_n19467_));
  OAI21_X1   g16369(.A1(new_n19278_), .A2(new_n14538_), .B(new_n13860_), .ZN(new_n19468_));
  NAND2_X1   g16370(.A1(new_n19468_), .A2(new_n13868_), .ZN(new_n19469_));
  AOI21_X1   g16371(.A1(new_n19302_), .A2(pi0619), .B(new_n19469_), .ZN(new_n19470_));
  AOI21_X1   g16372(.A1(new_n19356_), .A2(new_n19470_), .B(pi0619), .ZN(new_n19471_));
  OAI21_X1   g16373(.A1(new_n19467_), .A2(new_n19471_), .B(new_n13896_), .ZN(new_n19472_));
  NOR2_X1    g16374(.A1(new_n19361_), .A2(new_n19358_), .ZN(new_n19473_));
  AOI21_X1   g16375(.A1(new_n19473_), .A2(new_n13963_), .B(new_n19028_), .ZN(new_n19474_));
  NOR4_X1    g16376(.A1(new_n19361_), .A2(pi0626), .A3(new_n19208_), .A4(new_n19358_), .ZN(new_n19475_));
  OAI21_X1   g16377(.A1(new_n19474_), .A2(new_n19475_), .B(new_n19278_), .ZN(new_n19476_));
  NAND2_X1   g16378(.A1(new_n19302_), .A2(new_n16639_), .ZN(new_n19477_));
  XOR2_X1    g16379(.A1(new_n19477_), .A2(new_n16829_), .Z(new_n19478_));
  AOI21_X1   g16380(.A1(new_n19478_), .A2(new_n19278_), .B(pi0788), .ZN(new_n19479_));
  AOI21_X1   g16381(.A1(new_n19473_), .A2(new_n13962_), .B(new_n18976_), .ZN(new_n19480_));
  NOR4_X1    g16382(.A1(new_n19361_), .A2(pi0626), .A3(new_n18974_), .A4(new_n19358_), .ZN(new_n19481_));
  OAI21_X1   g16383(.A1(new_n19480_), .A2(new_n19481_), .B(new_n19278_), .ZN(new_n19482_));
  AOI21_X1   g16384(.A1(new_n19476_), .A2(new_n19479_), .B(new_n19482_), .ZN(new_n19483_));
  INV_X1     g16385(.I(new_n13991_), .ZN(new_n19484_));
  NOR2_X1    g16386(.A1(new_n19305_), .A2(new_n19484_), .ZN(new_n19485_));
  NAND2_X1   g16387(.A1(new_n13991_), .A2(pi0628), .ZN(new_n19486_));
  XOR2_X1    g16388(.A1(new_n19485_), .A2(new_n19486_), .Z(new_n19487_));
  NOR2_X1    g16389(.A1(new_n19487_), .A2(new_n19299_), .ZN(new_n19488_));
  INV_X1     g16390(.I(new_n13990_), .ZN(new_n19489_));
  NAND2_X1   g16391(.A1(new_n19305_), .A2(pi0628), .ZN(new_n19490_));
  NAND2_X1   g16392(.A1(new_n19299_), .A2(new_n13942_), .ZN(new_n19491_));
  AOI21_X1   g16393(.A1(new_n19490_), .A2(new_n19491_), .B(new_n19489_), .ZN(new_n19492_));
  OAI21_X1   g16394(.A1(new_n19488_), .A2(new_n19492_), .B(new_n16874_), .ZN(new_n19493_));
  NOR2_X1    g16395(.A1(new_n19363_), .A2(new_n19493_), .ZN(new_n19494_));
  NOR3_X1    g16396(.A1(new_n19363_), .A2(new_n16424_), .A3(new_n19493_), .ZN(new_n19495_));
  NOR4_X1    g16397(.A1(new_n19495_), .A2(new_n19494_), .A3(new_n12777_), .A4(new_n16574_), .ZN(new_n19496_));
  OAI21_X1   g16398(.A1(new_n19299_), .A2(new_n13860_), .B(new_n13916_), .ZN(new_n19497_));
  NAND2_X1   g16399(.A1(new_n19357_), .A2(new_n19497_), .ZN(new_n19498_));
  NOR2_X1    g16400(.A1(new_n13860_), .A2(new_n13868_), .ZN(new_n19499_));
  NAND2_X1   g16401(.A1(new_n19498_), .A2(new_n19499_), .ZN(new_n19500_));
  NOR2_X1    g16402(.A1(new_n9992_), .A2(pi0176), .ZN(new_n19501_));
  AOI21_X1   g16403(.A1(new_n13218_), .A2(new_n17414_), .B(new_n19501_), .ZN(new_n19502_));
  INV_X1     g16404(.I(new_n19502_), .ZN(new_n19503_));
  NOR3_X1    g16405(.A1(new_n13219_), .A2(pi0625), .A3(pi0704), .ZN(new_n19504_));
  NAND3_X1   g16406(.A1(new_n19503_), .A2(new_n19504_), .A3(new_n19501_), .ZN(new_n19505_));
  NOR3_X1    g16407(.A1(new_n19504_), .A2(new_n13614_), .A3(new_n19502_), .ZN(new_n19506_));
  XOR2_X1    g16408(.A1(new_n19505_), .A2(new_n19506_), .Z(new_n19507_));
  NAND2_X1   g16409(.A1(new_n19503_), .A2(new_n13748_), .ZN(new_n19508_));
  OAI21_X1   g16410(.A1(new_n19507_), .A2(new_n13748_), .B(new_n19508_), .ZN(new_n19509_));
  NAND2_X1   g16411(.A1(new_n19509_), .A2(new_n14049_), .ZN(new_n19510_));
  NOR2_X1    g16412(.A1(new_n19510_), .A2(new_n14051_), .ZN(new_n19511_));
  INV_X1     g16413(.I(new_n19511_), .ZN(new_n19512_));
  NOR2_X1    g16414(.A1(new_n19512_), .A2(new_n14163_), .ZN(new_n19513_));
  AOI21_X1   g16415(.A1(new_n13104_), .A2(new_n17409_), .B(new_n19501_), .ZN(new_n19514_));
  NOR2_X1    g16416(.A1(new_n14096_), .A2(new_n19514_), .ZN(new_n19515_));
  AOI21_X1   g16417(.A1(new_n19515_), .A2(new_n14094_), .B(pi1155), .ZN(new_n19516_));
  NOR2_X1    g16418(.A1(new_n19516_), .A2(new_n13801_), .ZN(new_n19517_));
  NAND2_X1   g16419(.A1(new_n19514_), .A2(pi1155), .ZN(new_n19518_));
  AOI21_X1   g16420(.A1(new_n19518_), .A2(new_n2723_), .B(new_n14102_), .ZN(new_n19519_));
  NAND3_X1   g16421(.A1(new_n19519_), .A2(pi0785), .A3(new_n19515_), .ZN(new_n19520_));
  XOR2_X1    g16422(.A1(new_n19517_), .A2(new_n19520_), .Z(new_n19521_));
  NOR2_X1    g16423(.A1(new_n19521_), .A2(new_n13817_), .ZN(new_n19522_));
  OAI21_X1   g16424(.A1(new_n19522_), .A2(pi0618), .B(new_n9992_), .ZN(new_n19523_));
  NAND2_X1   g16425(.A1(new_n19523_), .A2(pi0781), .ZN(new_n19524_));
  OAI21_X1   g16426(.A1(new_n19522_), .A2(new_n9992_), .B(pi0618), .ZN(new_n19525_));
  NOR3_X1    g16427(.A1(new_n19525_), .A2(new_n13855_), .A3(new_n19521_), .ZN(new_n19526_));
  XOR2_X1    g16428(.A1(new_n19526_), .A2(new_n19524_), .Z(new_n19527_));
  NAND2_X1   g16429(.A1(new_n19527_), .A2(pi0619), .ZN(new_n19528_));
  XOR2_X1    g16430(.A1(new_n19528_), .A2(new_n13904_), .Z(new_n19529_));
  NAND2_X1   g16431(.A1(new_n19529_), .A2(new_n19501_), .ZN(new_n19530_));
  NAND2_X1   g16432(.A1(new_n19530_), .A2(pi0789), .ZN(new_n19531_));
  NAND2_X1   g16433(.A1(new_n19527_), .A2(pi1159), .ZN(new_n19532_));
  XOR2_X1    g16434(.A1(new_n19532_), .A2(new_n13904_), .Z(new_n19533_));
  NAND2_X1   g16435(.A1(new_n19533_), .A2(new_n19501_), .ZN(new_n19534_));
  NOR3_X1    g16436(.A1(new_n19534_), .A2(new_n13896_), .A3(new_n19527_), .ZN(new_n19535_));
  XOR2_X1    g16437(.A1(new_n19535_), .A2(new_n19531_), .Z(new_n19536_));
  NAND2_X1   g16438(.A1(new_n19536_), .A2(new_n13962_), .ZN(new_n19537_));
  XOR2_X1    g16439(.A1(new_n19537_), .A2(new_n18976_), .Z(new_n19538_));
  AOI22_X1   g16440(.A1(new_n19538_), .A2(new_n19501_), .B1(new_n16639_), .B2(new_n19513_), .ZN(new_n19539_));
  NOR3_X1    g16441(.A1(new_n19502_), .A2(new_n13613_), .A3(new_n13203_), .ZN(new_n19540_));
  INV_X1     g16442(.I(new_n19514_), .ZN(new_n19541_));
  NOR2_X1    g16443(.A1(new_n19501_), .A2(pi1153), .ZN(new_n19542_));
  INV_X1     g16444(.I(new_n19542_), .ZN(new_n19543_));
  OAI21_X1   g16445(.A1(new_n19504_), .A2(new_n19543_), .B(pi0608), .ZN(new_n19544_));
  NAND3_X1   g16446(.A1(new_n19544_), .A2(new_n13614_), .A3(new_n19541_), .ZN(new_n19545_));
  AOI21_X1   g16447(.A1(new_n19545_), .A2(new_n19540_), .B(new_n13748_), .ZN(new_n19546_));
  NOR2_X1    g16448(.A1(new_n19502_), .A2(new_n13203_), .ZN(new_n19547_));
  NAND2_X1   g16449(.A1(new_n19504_), .A2(new_n19542_), .ZN(new_n19548_));
  AOI21_X1   g16450(.A1(new_n14083_), .A2(new_n19503_), .B(new_n19548_), .ZN(new_n19549_));
  NOR2_X1    g16451(.A1(new_n19549_), .A2(new_n19540_), .ZN(new_n19550_));
  NOR4_X1    g16452(.A1(new_n19550_), .A2(new_n13748_), .A3(new_n19541_), .A4(new_n19547_), .ZN(new_n19551_));
  XOR2_X1    g16453(.A1(new_n19551_), .A2(new_n19546_), .Z(new_n19552_));
  NAND2_X1   g16454(.A1(new_n19552_), .A2(new_n13801_), .ZN(new_n19553_));
  NOR2_X1    g16455(.A1(new_n19552_), .A2(new_n13778_), .ZN(new_n19554_));
  XOR2_X1    g16456(.A1(new_n19554_), .A2(new_n14090_), .Z(new_n19555_));
  NAND2_X1   g16457(.A1(new_n19555_), .A2(new_n19509_), .ZN(new_n19556_));
  NOR2_X1    g16458(.A1(new_n19516_), .A2(new_n13783_), .ZN(new_n19557_));
  NAND2_X1   g16459(.A1(new_n19556_), .A2(new_n19557_), .ZN(new_n19558_));
  NOR2_X1    g16460(.A1(new_n19519_), .A2(pi0660), .ZN(new_n19559_));
  NAND2_X1   g16461(.A1(new_n19558_), .A2(new_n19559_), .ZN(new_n19560_));
  NOR2_X1    g16462(.A1(new_n19552_), .A2(new_n13766_), .ZN(new_n19561_));
  XOR2_X1    g16463(.A1(new_n19561_), .A2(new_n14090_), .Z(new_n19562_));
  NAND4_X1   g16464(.A1(new_n19560_), .A2(pi0785), .A3(new_n19509_), .A4(new_n19562_), .ZN(new_n19563_));
  NAND2_X1   g16465(.A1(new_n19563_), .A2(new_n19553_), .ZN(new_n19564_));
  NAND2_X1   g16466(.A1(new_n19564_), .A2(new_n13855_), .ZN(new_n19565_));
  NOR2_X1    g16467(.A1(new_n19564_), .A2(new_n13816_), .ZN(new_n19566_));
  XOR2_X1    g16468(.A1(new_n19566_), .A2(new_n13818_), .Z(new_n19567_));
  NAND3_X1   g16469(.A1(new_n19567_), .A2(new_n14049_), .A3(new_n19509_), .ZN(new_n19568_));
  NAND3_X1   g16470(.A1(new_n19568_), .A2(new_n13823_), .A3(new_n19525_), .ZN(new_n19569_));
  AND3_X2    g16471(.A1(new_n19569_), .A2(new_n13823_), .A3(new_n19523_), .Z(new_n19570_));
  NOR2_X1    g16472(.A1(new_n19564_), .A2(new_n13817_), .ZN(new_n19571_));
  XOR2_X1    g16473(.A1(new_n19571_), .A2(new_n13819_), .Z(new_n19572_));
  NOR3_X1    g16474(.A1(new_n19572_), .A2(new_n13855_), .A3(new_n19510_), .ZN(new_n19573_));
  INV_X1     g16475(.I(new_n19573_), .ZN(new_n19574_));
  OAI21_X1   g16476(.A1(new_n19570_), .A2(new_n19574_), .B(new_n19565_), .ZN(new_n19575_));
  NOR2_X1    g16477(.A1(new_n19575_), .A2(new_n13860_), .ZN(new_n19576_));
  XOR2_X1    g16478(.A1(new_n19576_), .A2(new_n13904_), .Z(new_n19577_));
  NOR2_X1    g16479(.A1(new_n19577_), .A2(new_n19512_), .ZN(new_n19578_));
  NAND2_X1   g16480(.A1(new_n19534_), .A2(new_n13884_), .ZN(new_n19579_));
  INV_X1     g16481(.I(new_n19575_), .ZN(new_n19580_));
  AOI21_X1   g16482(.A1(new_n19580_), .A2(new_n14143_), .B(pi0789), .ZN(new_n19581_));
  OAI21_X1   g16483(.A1(new_n19578_), .A2(new_n19579_), .B(new_n19581_), .ZN(new_n19582_));
  NOR2_X1    g16484(.A1(new_n19575_), .A2(new_n13868_), .ZN(new_n19583_));
  XOR2_X1    g16485(.A1(new_n19583_), .A2(new_n13903_), .Z(new_n19584_));
  NAND2_X1   g16486(.A1(new_n19530_), .A2(new_n19018_), .ZN(new_n19585_));
  AOI21_X1   g16487(.A1(new_n19584_), .A2(new_n19511_), .B(new_n19585_), .ZN(new_n19586_));
  AOI21_X1   g16488(.A1(new_n19582_), .A2(new_n19586_), .B(new_n19539_), .ZN(new_n19587_));
  NAND2_X1   g16489(.A1(new_n19536_), .A2(new_n16372_), .ZN(new_n19588_));
  OAI21_X1   g16490(.A1(new_n16372_), .A2(new_n19501_), .B(new_n19588_), .ZN(new_n19589_));
  NAND3_X1   g16491(.A1(new_n19589_), .A2(new_n18929_), .A3(new_n19513_), .ZN(new_n19590_));
  NAND2_X1   g16492(.A1(new_n19590_), .A2(new_n16569_), .ZN(new_n19591_));
  XOR2_X1    g16493(.A1(new_n19591_), .A2(new_n16572_), .Z(new_n19592_));
  AOI21_X1   g16494(.A1(new_n19022_), .A2(new_n19590_), .B(new_n19592_), .ZN(new_n19593_));
  INV_X1     g16495(.I(new_n19501_), .ZN(new_n19594_));
  NAND2_X1   g16496(.A1(new_n19536_), .A2(new_n13963_), .ZN(new_n19595_));
  XNOR2_X1   g16497(.A1(new_n19595_), .A2(new_n19028_), .ZN(new_n19596_));
  NOR3_X1    g16498(.A1(new_n19596_), .A2(new_n16424_), .A3(new_n19594_), .ZN(new_n19597_));
  OAI21_X1   g16499(.A1(new_n19593_), .A2(new_n16574_), .B(new_n19597_), .ZN(new_n19598_));
  NOR4_X1    g16500(.A1(new_n19512_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n19599_));
  NOR2_X1    g16501(.A1(new_n19599_), .A2(new_n14005_), .ZN(new_n19600_));
  XOR2_X1    g16502(.A1(new_n19600_), .A2(new_n14007_), .Z(new_n19601_));
  NAND2_X1   g16503(.A1(new_n19601_), .A2(new_n19501_), .ZN(new_n19602_));
  NOR2_X1    g16504(.A1(new_n19594_), .A2(pi0647), .ZN(new_n19603_));
  AOI21_X1   g16505(.A1(new_n19599_), .A2(pi0647), .B(new_n19603_), .ZN(new_n19604_));
  NOR2_X1    g16506(.A1(new_n19589_), .A2(new_n13994_), .ZN(new_n19605_));
  XNOR2_X1   g16507(.A1(new_n19605_), .A2(new_n19033_), .ZN(new_n19606_));
  AOI22_X1   g16508(.A1(new_n19606_), .A2(new_n19501_), .B1(new_n14206_), .B2(new_n19604_), .ZN(new_n19607_));
  NOR3_X1    g16509(.A1(new_n19607_), .A2(new_n14010_), .A3(new_n19602_), .ZN(new_n19608_));
  OAI22_X1   g16510(.A1(new_n19587_), .A2(new_n19598_), .B1(new_n12776_), .B2(new_n19608_), .ZN(new_n19609_));
  AOI21_X1   g16511(.A1(new_n19604_), .A2(pi1157), .B(new_n12776_), .ZN(new_n19610_));
  AOI22_X1   g16512(.A1(new_n19602_), .A2(new_n19610_), .B1(new_n12776_), .B2(new_n19599_), .ZN(new_n19611_));
  NAND2_X1   g16513(.A1(new_n19609_), .A2(pi0644), .ZN(new_n19612_));
  XOR2_X1    g16514(.A1(new_n19612_), .A2(new_n14205_), .Z(new_n19613_));
  NOR2_X1    g16515(.A1(new_n19613_), .A2(new_n19611_), .ZN(new_n19614_));
  NOR2_X1    g16516(.A1(new_n19589_), .A2(new_n18968_), .ZN(new_n19615_));
  NAND2_X1   g16517(.A1(new_n18967_), .A2(new_n19501_), .ZN(new_n19616_));
  XOR2_X1    g16518(.A1(new_n19615_), .A2(new_n19616_), .Z(new_n19617_));
  NAND2_X1   g16519(.A1(new_n19617_), .A2(pi0715), .ZN(new_n19618_));
  XOR2_X1    g16520(.A1(new_n19618_), .A2(new_n14205_), .Z(new_n19619_));
  OAI21_X1   g16521(.A1(new_n19619_), .A2(new_n19594_), .B(new_n14203_), .ZN(new_n19620_));
  NAND2_X1   g16522(.A1(new_n19617_), .A2(pi0644), .ZN(new_n19621_));
  XOR2_X1    g16523(.A1(new_n19621_), .A2(new_n14217_), .Z(new_n19622_));
  AOI21_X1   g16524(.A1(new_n19622_), .A2(new_n19501_), .B(pi1160), .ZN(new_n19623_));
  OAI21_X1   g16525(.A1(new_n19614_), .A2(new_n19620_), .B(new_n19623_), .ZN(new_n19624_));
  NAND2_X1   g16526(.A1(new_n19609_), .A2(pi0715), .ZN(new_n19625_));
  XOR2_X1    g16527(.A1(new_n19625_), .A2(new_n14205_), .Z(new_n19626_));
  NOR2_X1    g16528(.A1(new_n19626_), .A2(new_n19611_), .ZN(new_n19627_));
  AOI21_X1   g16529(.A1(new_n19624_), .A2(new_n19627_), .B(new_n14799_), .ZN(new_n19628_));
  XOR2_X1    g16530(.A1(new_n19628_), .A2(new_n14801_), .Z(new_n19629_));
  OAI21_X1   g16531(.A1(new_n7240_), .A2(pi0176), .B(new_n14799_), .ZN(new_n19630_));
  OR3_X2     g16532(.A1(new_n19629_), .A2(new_n19609_), .A3(new_n19630_), .Z(new_n19631_));
  AOI22_X1   g16533(.A1(new_n19500_), .A2(new_n13860_), .B1(new_n7240_), .B2(new_n19631_), .ZN(new_n19632_));
  OAI21_X1   g16534(.A1(new_n19483_), .A2(new_n19496_), .B(new_n19632_), .ZN(new_n19633_));
  NOR2_X1    g16535(.A1(new_n19467_), .A2(new_n19633_), .ZN(new_n19634_));
  OAI21_X1   g16536(.A1(new_n19472_), .A2(new_n19466_), .B(new_n19634_), .ZN(new_n19635_));
  AOI21_X1   g16537(.A1(new_n19378_), .A2(new_n19387_), .B(new_n19635_), .ZN(po0333));
  NOR2_X1    g16538(.A1(new_n15562_), .A2(pi0038), .ZN(new_n19637_));
  NAND3_X1   g16539(.A1(new_n13097_), .A2(pi0038), .A3(pi0757), .ZN(new_n19638_));
  NAND3_X1   g16540(.A1(new_n13632_), .A2(new_n3259_), .A3(pi0757), .ZN(new_n19639_));
  NAND2_X1   g16541(.A1(new_n19639_), .A2(new_n19638_), .ZN(new_n19640_));
  INV_X1     g16542(.I(new_n19321_), .ZN(new_n19641_));
  NOR2_X1    g16543(.A1(new_n19641_), .A2(new_n3259_), .ZN(new_n19642_));
  AOI22_X1   g16544(.A1(new_n19640_), .A2(new_n13624_), .B1(pi0177), .B2(new_n19637_), .ZN(new_n19645_));
  NOR2_X1    g16545(.A1(new_n15556_), .A2(pi0757), .ZN(new_n19646_));
  INV_X1     g16546(.I(new_n19646_), .ZN(new_n19647_));
  NOR2_X1    g16547(.A1(new_n19645_), .A2(new_n19647_), .ZN(new_n19648_));
  INV_X1     g16548(.I(new_n19648_), .ZN(new_n19649_));
  NAND2_X1   g16549(.A1(new_n13359_), .A2(pi0039), .ZN(new_n19650_));
  OAI21_X1   g16550(.A1(pi0039), .A2(new_n13152_), .B(new_n19650_), .ZN(new_n19651_));
  NAND2_X1   g16551(.A1(new_n19651_), .A2(pi0177), .ZN(new_n19652_));
  AOI21_X1   g16552(.A1(new_n14293_), .A2(pi0757), .B(pi0177), .ZN(new_n19653_));
  NOR3_X1    g16553(.A1(new_n19653_), .A2(pi0038), .A3(new_n13109_), .ZN(new_n19654_));
  AOI22_X1   g16554(.A1(new_n19652_), .A2(new_n19654_), .B1(new_n15578_), .B2(new_n15585_), .ZN(new_n19655_));
  OAI22_X1   g16555(.A1(new_n19655_), .A2(new_n8010_), .B1(new_n17440_), .B2(new_n3290_), .ZN(new_n19656_));
  OAI21_X1   g16556(.A1(pi0039), .A2(new_n13191_), .B(new_n13522_), .ZN(new_n19657_));
  NAND2_X1   g16557(.A1(new_n13198_), .A2(new_n3183_), .ZN(new_n19658_));
  AOI21_X1   g16558(.A1(new_n15625_), .A2(new_n19658_), .B(new_n8010_), .ZN(new_n19659_));
  NAND2_X1   g16559(.A1(pi0038), .A2(pi0177), .ZN(new_n19660_));
  XNOR2_X1   g16560(.A1(new_n19659_), .A2(new_n19660_), .ZN(new_n19661_));
  NAND2_X1   g16561(.A1(new_n13209_), .A2(new_n3183_), .ZN(new_n19662_));
  NAND2_X1   g16562(.A1(new_n19662_), .A2(pi0038), .ZN(new_n19663_));
  XOR2_X1    g16563(.A1(new_n19663_), .A2(new_n19660_), .Z(new_n19664_));
  NAND2_X1   g16564(.A1(new_n19664_), .A2(new_n15620_), .ZN(new_n19665_));
  NAND4_X1   g16565(.A1(new_n19665_), .A2(pi0177), .A3(new_n17446_), .A4(new_n3290_), .ZN(new_n19666_));
  AOI21_X1   g16566(.A1(new_n19661_), .A2(new_n19657_), .B(new_n19666_), .ZN(new_n19667_));
  NAND2_X1   g16567(.A1(new_n19656_), .A2(new_n19667_), .ZN(new_n19668_));
  AOI21_X1   g16568(.A1(new_n19668_), .A2(new_n17440_), .B(new_n19649_), .ZN(new_n19669_));
  NOR2_X1    g16569(.A1(new_n3289_), .A2(pi0177), .ZN(new_n19670_));
  INV_X1     g16570(.I(new_n19670_), .ZN(new_n19671_));
  OAI21_X1   g16571(.A1(new_n19648_), .A2(new_n3290_), .B(new_n19671_), .ZN(new_n19672_));
  OAI21_X1   g16572(.A1(new_n13721_), .A2(new_n17440_), .B(new_n8010_), .ZN(new_n19673_));
  NAND2_X1   g16573(.A1(new_n19673_), .A2(new_n13108_), .ZN(new_n19674_));
  NAND2_X1   g16574(.A1(new_n8010_), .A2(new_n17440_), .ZN(new_n19675_));
  NAND4_X1   g16575(.A1(new_n13634_), .A2(pi0177), .A3(new_n3290_), .A4(new_n19675_), .ZN(new_n19676_));
  AOI21_X1   g16576(.A1(new_n14424_), .A2(pi0177), .B(new_n19660_), .ZN(new_n19677_));
  NOR3_X1    g16577(.A1(new_n14422_), .A2(pi0038), .A3(new_n8010_), .ZN(new_n19678_));
  OAI21_X1   g16578(.A1(new_n19677_), .A2(new_n19678_), .B(new_n15655_), .ZN(new_n19679_));
  AOI21_X1   g16579(.A1(new_n19674_), .A2(new_n19676_), .B(new_n19679_), .ZN(new_n19680_));
  NOR3_X1    g16580(.A1(new_n14431_), .A2(new_n8010_), .A3(new_n14081_), .ZN(new_n19681_));
  OAI21_X1   g16581(.A1(new_n19680_), .A2(new_n19681_), .B(new_n13615_), .ZN(new_n19682_));
  OAI21_X1   g16582(.A1(new_n19672_), .A2(new_n19682_), .B(new_n13613_), .ZN(new_n19683_));
  AOI21_X1   g16583(.A1(new_n19669_), .A2(new_n19683_), .B(new_n13748_), .ZN(new_n19684_));
  NAND3_X1   g16584(.A1(new_n19669_), .A2(pi0625), .A3(pi0778), .ZN(new_n19689_));
  XOR2_X1    g16585(.A1(new_n19684_), .A2(new_n19689_), .Z(new_n19690_));
  NOR2_X1    g16586(.A1(new_n19672_), .A2(new_n13775_), .ZN(new_n19691_));
  NOR2_X1    g16587(.A1(new_n14428_), .A2(pi0177), .ZN(new_n19692_));
  NOR2_X1    g16588(.A1(new_n19692_), .A2(new_n15147_), .ZN(new_n19693_));
  OAI21_X1   g16589(.A1(new_n19691_), .A2(new_n19693_), .B(pi0609), .ZN(new_n19694_));
  NAND2_X1   g16590(.A1(new_n19680_), .A2(new_n13748_), .ZN(new_n19695_));
  NOR2_X1    g16591(.A1(new_n19680_), .A2(new_n14452_), .ZN(new_n19696_));
  INV_X1     g16592(.I(new_n19692_), .ZN(new_n19697_));
  NOR2_X1    g16593(.A1(new_n19697_), .A2(new_n14452_), .ZN(new_n19698_));
  XNOR2_X1   g16594(.A1(new_n19696_), .A2(new_n19698_), .ZN(new_n19699_));
  OAI21_X1   g16595(.A1(new_n19699_), .A2(new_n13748_), .B(new_n19695_), .ZN(new_n19700_));
  AOI21_X1   g16596(.A1(new_n19700_), .A2(new_n13766_), .B(new_n13785_), .ZN(new_n19701_));
  AOI21_X1   g16597(.A1(new_n19701_), .A2(new_n19694_), .B(pi0609), .ZN(new_n19702_));
  OAI21_X1   g16598(.A1(new_n19690_), .A2(new_n19702_), .B(pi0785), .ZN(new_n19703_));
  NAND2_X1   g16599(.A1(new_n19700_), .A2(pi0609), .ZN(new_n19704_));
  AOI21_X1   g16600(.A1(new_n19697_), .A2(new_n14467_), .B(pi0609), .ZN(new_n19705_));
  INV_X1     g16601(.I(new_n19705_), .ZN(new_n19706_));
  AOI21_X1   g16602(.A1(new_n19691_), .A2(new_n19706_), .B(new_n14465_), .ZN(new_n19707_));
  AOI21_X1   g16603(.A1(new_n19704_), .A2(new_n19707_), .B(pi0609), .ZN(new_n19708_));
  NOR3_X1    g16604(.A1(new_n19690_), .A2(new_n13801_), .A3(new_n19708_), .ZN(new_n19709_));
  XOR2_X1    g16605(.A1(new_n19709_), .A2(new_n19703_), .Z(new_n19710_));
  NAND2_X1   g16606(.A1(new_n19694_), .A2(pi0785), .ZN(new_n19711_));
  NOR2_X1    g16607(.A1(new_n19697_), .A2(new_n13776_), .ZN(new_n19712_));
  AOI21_X1   g16608(.A1(new_n19672_), .A2(new_n13776_), .B(new_n19712_), .ZN(new_n19713_));
  NAND3_X1   g16609(.A1(new_n19691_), .A2(pi0785), .A3(new_n19706_), .ZN(new_n19714_));
  NOR2_X1    g16610(.A1(new_n19714_), .A2(new_n19713_), .ZN(new_n19715_));
  NAND2_X1   g16611(.A1(new_n19711_), .A2(new_n19715_), .ZN(new_n19716_));
  NOR2_X1    g16612(.A1(new_n19711_), .A2(new_n19715_), .ZN(new_n19717_));
  INV_X1     g16613(.I(new_n19717_), .ZN(new_n19718_));
  NAND2_X1   g16614(.A1(new_n19718_), .A2(new_n19716_), .ZN(new_n19719_));
  NAND3_X1   g16615(.A1(new_n19719_), .A2(pi0618), .A3(pi1154), .ZN(new_n19720_));
  INV_X1     g16616(.I(new_n19720_), .ZN(new_n19721_));
  NOR3_X1    g16617(.A1(new_n19719_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n19722_));
  OAI21_X1   g16618(.A1(new_n19721_), .A2(new_n19722_), .B(new_n19692_), .ZN(new_n19723_));
  NOR2_X1    g16619(.A1(new_n19697_), .A2(new_n13805_), .ZN(new_n19724_));
  AOI21_X1   g16620(.A1(new_n19700_), .A2(new_n13805_), .B(new_n19724_), .ZN(new_n19725_));
  INV_X1     g16621(.I(new_n19725_), .ZN(new_n19726_));
  AOI21_X1   g16622(.A1(new_n19726_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n19727_));
  AOI21_X1   g16623(.A1(new_n19723_), .A2(new_n19727_), .B(pi0618), .ZN(new_n19728_));
  NAND3_X1   g16624(.A1(new_n19719_), .A2(pi0618), .A3(pi1154), .ZN(new_n19729_));
  NAND4_X1   g16625(.A1(new_n19718_), .A2(new_n19716_), .A3(new_n13816_), .A4(pi1154), .ZN(new_n19730_));
  AOI21_X1   g16626(.A1(new_n19729_), .A2(new_n19730_), .B(new_n19697_), .ZN(new_n19731_));
  INV_X1     g16627(.I(new_n19731_), .ZN(new_n19732_));
  AOI21_X1   g16628(.A1(new_n19726_), .A2(pi0618), .B(new_n13837_), .ZN(new_n19733_));
  AOI21_X1   g16629(.A1(new_n19732_), .A2(new_n19733_), .B(pi0618), .ZN(new_n19734_));
  NOR4_X1    g16630(.A1(new_n19710_), .A2(new_n19734_), .A3(new_n19728_), .A4(new_n13855_), .ZN(new_n19735_));
  OAI21_X1   g16631(.A1(new_n19710_), .A2(new_n19728_), .B(pi0781), .ZN(new_n19736_));
  NOR3_X1    g16632(.A1(new_n19710_), .A2(new_n19734_), .A3(new_n13855_), .ZN(new_n19737_));
  NOR2_X1    g16633(.A1(new_n19737_), .A2(new_n19736_), .ZN(new_n19738_));
  NOR2_X1    g16634(.A1(new_n19738_), .A2(new_n19735_), .ZN(new_n19739_));
  INV_X1     g16635(.I(new_n19739_), .ZN(new_n19740_));
  INV_X1     g16636(.I(new_n19722_), .ZN(new_n19741_));
  AOI21_X1   g16637(.A1(new_n19741_), .A2(new_n19720_), .B(new_n19697_), .ZN(new_n19742_));
  NAND4_X1   g16638(.A1(new_n19742_), .A2(new_n19731_), .A3(pi0781), .A4(new_n19719_), .ZN(new_n19743_));
  NAND3_X1   g16639(.A1(new_n19731_), .A2(pi0781), .A3(new_n19719_), .ZN(new_n19744_));
  NAND3_X1   g16640(.A1(new_n19744_), .A2(pi0781), .A3(new_n19723_), .ZN(new_n19745_));
  NAND2_X1   g16641(.A1(new_n19745_), .A2(new_n19743_), .ZN(new_n19746_));
  NAND3_X1   g16642(.A1(new_n19746_), .A2(pi0619), .A3(pi1159), .ZN(new_n19747_));
  NAND4_X1   g16643(.A1(new_n19745_), .A2(new_n19743_), .A3(pi0619), .A4(new_n13868_), .ZN(new_n19748_));
  AOI21_X1   g16644(.A1(new_n19747_), .A2(new_n19748_), .B(new_n19697_), .ZN(new_n19749_));
  NOR2_X1    g16645(.A1(new_n19692_), .A2(new_n13880_), .ZN(new_n19750_));
  AOI21_X1   g16646(.A1(new_n19725_), .A2(new_n13880_), .B(new_n19750_), .ZN(new_n19751_));
  AOI21_X1   g16647(.A1(new_n19751_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n19752_));
  INV_X1     g16648(.I(new_n19752_), .ZN(new_n19753_));
  OAI21_X1   g16649(.A1(new_n19749_), .A2(new_n19753_), .B(new_n13860_), .ZN(new_n19754_));
  NAND3_X1   g16650(.A1(new_n19746_), .A2(pi0619), .A3(pi1159), .ZN(new_n19755_));
  NAND4_X1   g16651(.A1(new_n19745_), .A2(new_n19743_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n19756_));
  AOI21_X1   g16652(.A1(new_n19755_), .A2(new_n19756_), .B(new_n19697_), .ZN(new_n19757_));
  AOI21_X1   g16653(.A1(new_n19751_), .A2(pi0619), .B(new_n15217_), .ZN(new_n19758_));
  INV_X1     g16654(.I(new_n19758_), .ZN(new_n19759_));
  OAI21_X1   g16655(.A1(new_n19757_), .A2(new_n19759_), .B(new_n13860_), .ZN(new_n19760_));
  NAND4_X1   g16656(.A1(new_n19754_), .A2(new_n19760_), .A3(pi0789), .A4(new_n19740_), .ZN(new_n19761_));
  AOI21_X1   g16657(.A1(new_n19754_), .A2(new_n19740_), .B(new_n13896_), .ZN(new_n19762_));
  NAND3_X1   g16658(.A1(new_n19760_), .A2(pi0789), .A3(new_n19740_), .ZN(new_n19763_));
  NAND2_X1   g16659(.A1(new_n19762_), .A2(new_n19763_), .ZN(new_n19764_));
  NAND2_X1   g16660(.A1(new_n19764_), .A2(new_n19761_), .ZN(new_n19765_));
  NAND4_X1   g16661(.A1(new_n19749_), .A2(new_n19757_), .A3(pi0789), .A4(new_n19746_), .ZN(new_n19766_));
  INV_X1     g16662(.I(new_n19749_), .ZN(new_n19767_));
  NAND3_X1   g16663(.A1(new_n19757_), .A2(pi0789), .A3(new_n19746_), .ZN(new_n19768_));
  NAND3_X1   g16664(.A1(new_n19768_), .A2(pi0789), .A3(new_n19767_), .ZN(new_n19769_));
  NOR2_X1    g16665(.A1(new_n19697_), .A2(new_n13919_), .ZN(new_n19770_));
  AOI21_X1   g16666(.A1(new_n19751_), .A2(new_n13919_), .B(new_n19770_), .ZN(new_n19771_));
  NOR2_X1    g16667(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n19772_));
  INV_X1     g16668(.I(new_n19772_), .ZN(new_n19773_));
  AOI21_X1   g16669(.A1(new_n19769_), .A2(new_n19766_), .B(new_n19773_), .ZN(new_n19774_));
  INV_X1     g16670(.I(new_n19766_), .ZN(new_n19775_));
  AND3_X2    g16671(.A1(new_n19768_), .A2(pi0789), .A3(new_n19767_), .Z(new_n19776_));
  NOR2_X1    g16672(.A1(new_n19776_), .A2(new_n19775_), .ZN(new_n19777_));
  NAND3_X1   g16673(.A1(new_n19765_), .A2(pi0626), .A3(pi0788), .ZN(new_n19782_));
  INV_X1     g16674(.I(new_n19782_), .ZN(new_n19783_));
  OAI21_X1   g16675(.A1(new_n19776_), .A2(new_n19775_), .B(new_n19772_), .ZN(new_n19784_));
  AOI22_X1   g16676(.A1(new_n19784_), .A2(new_n13901_), .B1(new_n19764_), .B2(new_n19761_), .ZN(new_n19785_));
  AOI21_X1   g16677(.A1(new_n19764_), .A2(new_n19761_), .B(new_n15258_), .ZN(new_n19786_));
  NOR3_X1    g16678(.A1(new_n19785_), .A2(new_n13937_), .A3(new_n19786_), .ZN(new_n19787_));
  NOR2_X1    g16679(.A1(new_n19787_), .A2(new_n19783_), .ZN(new_n19788_));
  NOR2_X1    g16680(.A1(new_n19692_), .A2(new_n16372_), .ZN(new_n19789_));
  AOI21_X1   g16681(.A1(new_n19777_), .A2(new_n16372_), .B(new_n19789_), .ZN(new_n19790_));
  NOR2_X1    g16682(.A1(new_n19692_), .A2(new_n13966_), .ZN(new_n19791_));
  AOI21_X1   g16683(.A1(new_n19771_), .A2(new_n13966_), .B(new_n19791_), .ZN(new_n19792_));
  NAND2_X1   g16684(.A1(new_n19792_), .A2(pi0628), .ZN(new_n19793_));
  NAND2_X1   g16685(.A1(new_n19793_), .A2(new_n13970_), .ZN(new_n19794_));
  NAND3_X1   g16686(.A1(new_n19792_), .A2(pi0628), .A3(new_n13971_), .ZN(new_n19795_));
  AOI21_X1   g16687(.A1(new_n19794_), .A2(new_n19795_), .B(new_n19697_), .ZN(new_n19796_));
  NOR2_X1    g16688(.A1(new_n19796_), .A2(new_n15270_), .ZN(new_n19797_));
  INV_X1     g16689(.I(new_n19797_), .ZN(new_n19798_));
  NAND2_X1   g16690(.A1(new_n19792_), .A2(pi1156), .ZN(new_n19800_));
  XOR2_X1    g16691(.A1(new_n19800_), .A2(new_n13971_), .Z(new_n19801_));
  NAND2_X1   g16692(.A1(new_n19801_), .A2(new_n19692_), .ZN(new_n19802_));
  NOR3_X1    g16693(.A1(new_n19788_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n19805_));
  INV_X1     g16694(.I(new_n19761_), .ZN(new_n19806_));
  AND2_X2    g16695(.A1(new_n19762_), .A2(new_n19763_), .Z(new_n19807_));
  OAI22_X1   g16696(.A1(new_n19807_), .A2(new_n19806_), .B1(new_n19774_), .B2(pi0626), .ZN(new_n19808_));
  NAND2_X1   g16697(.A1(new_n19765_), .A2(new_n14577_), .ZN(new_n19809_));
  NAND3_X1   g16698(.A1(new_n19808_), .A2(new_n19809_), .A3(pi0788), .ZN(new_n19810_));
  NAND3_X1   g16699(.A1(new_n19769_), .A2(new_n16372_), .A3(new_n19766_), .ZN(new_n19811_));
  OAI21_X1   g16700(.A1(new_n16372_), .A2(new_n19692_), .B(new_n19811_), .ZN(new_n19812_));
  AOI21_X1   g16701(.A1(new_n19812_), .A2(new_n19797_), .B(pi0628), .ZN(new_n19813_));
  AOI21_X1   g16702(.A1(new_n19810_), .A2(new_n19782_), .B(new_n19813_), .ZN(new_n19814_));
  AOI21_X1   g16703(.A1(new_n19810_), .A2(new_n19782_), .B(new_n15296_), .ZN(new_n19815_));
  NOR3_X1    g16704(.A1(new_n19814_), .A2(new_n19815_), .A3(new_n12777_), .ZN(new_n19816_));
  NOR2_X1    g16705(.A1(new_n19816_), .A2(new_n19805_), .ZN(new_n19817_));
  NOR2_X1    g16706(.A1(new_n19692_), .A2(new_n13994_), .ZN(new_n19818_));
  AOI21_X1   g16707(.A1(new_n19812_), .A2(new_n13994_), .B(new_n19818_), .ZN(new_n19819_));
  INV_X1     g16708(.I(new_n19819_), .ZN(new_n19820_));
  NOR2_X1    g16709(.A1(new_n19796_), .A2(new_n12777_), .ZN(new_n19821_));
  NOR4_X1    g16710(.A1(new_n19802_), .A2(new_n12777_), .A3(new_n19821_), .A4(new_n19792_), .ZN(new_n19822_));
  NOR3_X1    g16711(.A1(new_n19802_), .A2(new_n12777_), .A3(new_n19792_), .ZN(new_n19823_));
  NOR3_X1    g16712(.A1(new_n19823_), .A2(new_n12777_), .A3(new_n19796_), .ZN(new_n19824_));
  NOR2_X1    g16713(.A1(new_n19824_), .A2(new_n19822_), .ZN(new_n19825_));
  NAND2_X1   g16714(.A1(new_n19825_), .A2(pi0647), .ZN(new_n19826_));
  XOR2_X1    g16715(.A1(new_n19826_), .A2(new_n14008_), .Z(new_n19827_));
  AOI21_X1   g16716(.A1(new_n19827_), .A2(new_n19692_), .B(new_n14012_), .ZN(new_n19828_));
  AOI21_X1   g16717(.A1(new_n19820_), .A2(new_n19828_), .B(pi0647), .ZN(new_n19829_));
  AOI21_X1   g16718(.A1(new_n19825_), .A2(pi1157), .B(new_n14008_), .ZN(new_n19830_));
  NOR4_X1    g16719(.A1(new_n19824_), .A2(new_n19822_), .A3(pi0647), .A4(new_n14006_), .ZN(new_n19831_));
  OAI21_X1   g16720(.A1(new_n19830_), .A2(new_n19831_), .B(new_n19692_), .ZN(new_n19832_));
  NAND2_X1   g16721(.A1(new_n19832_), .A2(new_n14027_), .ZN(new_n19833_));
  AOI21_X1   g16722(.A1(new_n19819_), .A2(pi0647), .B(new_n19833_), .ZN(new_n19834_));
  NOR2_X1    g16723(.A1(new_n19834_), .A2(pi0647), .ZN(new_n19835_));
  NOR4_X1    g16724(.A1(new_n19817_), .A2(new_n12776_), .A3(new_n19829_), .A4(new_n19835_), .ZN(new_n19836_));
  NAND2_X1   g16725(.A1(new_n19810_), .A2(new_n19782_), .ZN(new_n19837_));
  NAND3_X1   g16726(.A1(new_n19837_), .A2(pi0628), .A3(pi0792), .ZN(new_n19838_));
  OAI21_X1   g16727(.A1(new_n19790_), .A2(new_n19798_), .B(new_n13942_), .ZN(new_n19839_));
  OAI21_X1   g16728(.A1(new_n19787_), .A2(new_n19783_), .B(new_n19839_), .ZN(new_n19840_));
  OAI21_X1   g16729(.A1(new_n19787_), .A2(new_n19783_), .B(new_n14606_), .ZN(new_n19841_));
  NAND3_X1   g16730(.A1(new_n19840_), .A2(new_n19841_), .A3(pi0792), .ZN(new_n19842_));
  AOI21_X1   g16731(.A1(new_n19842_), .A2(new_n19838_), .B(new_n19829_), .ZN(new_n19843_));
  OAI21_X1   g16732(.A1(new_n19834_), .A2(pi0647), .B(pi0787), .ZN(new_n19844_));
  AOI21_X1   g16733(.A1(new_n19842_), .A2(new_n19838_), .B(new_n19844_), .ZN(new_n19845_));
  NOR3_X1    g16734(.A1(new_n19843_), .A2(new_n19845_), .A3(new_n12776_), .ZN(new_n19846_));
  OAI21_X1   g16735(.A1(new_n19846_), .A2(new_n19836_), .B(new_n12775_), .ZN(new_n19847_));
  NOR2_X1    g16736(.A1(new_n9992_), .A2(pi0177), .ZN(new_n19848_));
  AOI21_X1   g16737(.A1(new_n13218_), .A2(new_n17440_), .B(new_n19848_), .ZN(new_n19849_));
  INV_X1     g16738(.I(new_n19849_), .ZN(new_n19850_));
  NOR3_X1    g16739(.A1(new_n13219_), .A2(pi0625), .A3(pi0686), .ZN(new_n19851_));
  NAND3_X1   g16740(.A1(new_n19850_), .A2(new_n19851_), .A3(new_n19848_), .ZN(new_n19852_));
  NOR3_X1    g16741(.A1(new_n19851_), .A2(new_n13614_), .A3(new_n19849_), .ZN(new_n19853_));
  XOR2_X1    g16742(.A1(new_n19852_), .A2(new_n19853_), .Z(new_n19854_));
  NAND2_X1   g16743(.A1(new_n19850_), .A2(new_n13748_), .ZN(new_n19855_));
  OAI21_X1   g16744(.A1(new_n19854_), .A2(new_n13748_), .B(new_n19855_), .ZN(new_n19856_));
  NAND2_X1   g16745(.A1(new_n19856_), .A2(new_n14049_), .ZN(new_n19857_));
  NOR2_X1    g16746(.A1(new_n19857_), .A2(new_n14051_), .ZN(new_n19858_));
  INV_X1     g16747(.I(new_n19858_), .ZN(new_n19859_));
  NOR2_X1    g16748(.A1(new_n19859_), .A2(new_n14163_), .ZN(new_n19860_));
  AOI21_X1   g16749(.A1(new_n13104_), .A2(new_n17446_), .B(new_n19848_), .ZN(new_n19861_));
  NOR2_X1    g16750(.A1(new_n14096_), .A2(new_n19861_), .ZN(new_n19862_));
  AOI21_X1   g16751(.A1(new_n19862_), .A2(new_n14094_), .B(pi1155), .ZN(new_n19863_));
  NOR2_X1    g16752(.A1(new_n19863_), .A2(new_n13801_), .ZN(new_n19864_));
  NAND2_X1   g16753(.A1(new_n19861_), .A2(pi1155), .ZN(new_n19865_));
  AOI21_X1   g16754(.A1(new_n19865_), .A2(new_n2723_), .B(new_n14102_), .ZN(new_n19866_));
  NAND3_X1   g16755(.A1(new_n19866_), .A2(pi0785), .A3(new_n19862_), .ZN(new_n19867_));
  XOR2_X1    g16756(.A1(new_n19864_), .A2(new_n19867_), .Z(new_n19868_));
  NOR2_X1    g16757(.A1(new_n19868_), .A2(new_n13817_), .ZN(new_n19869_));
  OAI21_X1   g16758(.A1(new_n19869_), .A2(pi0618), .B(new_n9992_), .ZN(new_n19870_));
  NAND2_X1   g16759(.A1(new_n19870_), .A2(pi0781), .ZN(new_n19871_));
  OAI21_X1   g16760(.A1(new_n19869_), .A2(new_n9992_), .B(pi0618), .ZN(new_n19872_));
  NOR3_X1    g16761(.A1(new_n19872_), .A2(new_n13855_), .A3(new_n19868_), .ZN(new_n19873_));
  XOR2_X1    g16762(.A1(new_n19873_), .A2(new_n19871_), .Z(new_n19874_));
  NAND2_X1   g16763(.A1(new_n19874_), .A2(pi0619), .ZN(new_n19875_));
  XOR2_X1    g16764(.A1(new_n19875_), .A2(new_n13904_), .Z(new_n19876_));
  NAND2_X1   g16765(.A1(new_n19876_), .A2(new_n19848_), .ZN(new_n19877_));
  NAND2_X1   g16766(.A1(new_n19877_), .A2(pi0789), .ZN(new_n19878_));
  NAND2_X1   g16767(.A1(new_n19874_), .A2(pi1159), .ZN(new_n19879_));
  XOR2_X1    g16768(.A1(new_n19879_), .A2(new_n13904_), .Z(new_n19880_));
  NAND2_X1   g16769(.A1(new_n19880_), .A2(new_n19848_), .ZN(new_n19881_));
  NOR3_X1    g16770(.A1(new_n19881_), .A2(new_n13896_), .A3(new_n19874_), .ZN(new_n19882_));
  XOR2_X1    g16771(.A1(new_n19882_), .A2(new_n19878_), .Z(new_n19883_));
  NAND2_X1   g16772(.A1(new_n19883_), .A2(new_n13962_), .ZN(new_n19884_));
  XOR2_X1    g16773(.A1(new_n19884_), .A2(new_n18976_), .Z(new_n19885_));
  AOI22_X1   g16774(.A1(new_n19885_), .A2(new_n19848_), .B1(new_n16639_), .B2(new_n19860_), .ZN(new_n19886_));
  NOR3_X1    g16775(.A1(new_n19849_), .A2(new_n13613_), .A3(new_n13203_), .ZN(new_n19887_));
  INV_X1     g16776(.I(new_n19861_), .ZN(new_n19888_));
  NOR2_X1    g16777(.A1(new_n19848_), .A2(pi1153), .ZN(new_n19889_));
  INV_X1     g16778(.I(new_n19889_), .ZN(new_n19890_));
  OAI21_X1   g16779(.A1(new_n19851_), .A2(new_n19890_), .B(pi0608), .ZN(new_n19891_));
  NAND3_X1   g16780(.A1(new_n19891_), .A2(new_n13614_), .A3(new_n19888_), .ZN(new_n19892_));
  AOI21_X1   g16781(.A1(new_n19892_), .A2(new_n19887_), .B(new_n13748_), .ZN(new_n19893_));
  NOR2_X1    g16782(.A1(new_n19849_), .A2(new_n13203_), .ZN(new_n19894_));
  NAND2_X1   g16783(.A1(new_n19851_), .A2(new_n19889_), .ZN(new_n19895_));
  AOI21_X1   g16784(.A1(new_n14083_), .A2(new_n19850_), .B(new_n19895_), .ZN(new_n19896_));
  NOR2_X1    g16785(.A1(new_n19896_), .A2(new_n19887_), .ZN(new_n19897_));
  NOR4_X1    g16786(.A1(new_n19897_), .A2(new_n13748_), .A3(new_n19888_), .A4(new_n19894_), .ZN(new_n19898_));
  XOR2_X1    g16787(.A1(new_n19898_), .A2(new_n19893_), .Z(new_n19899_));
  NAND2_X1   g16788(.A1(new_n19899_), .A2(new_n13801_), .ZN(new_n19900_));
  NOR2_X1    g16789(.A1(new_n19899_), .A2(new_n13778_), .ZN(new_n19901_));
  XOR2_X1    g16790(.A1(new_n19901_), .A2(new_n14090_), .Z(new_n19902_));
  NAND2_X1   g16791(.A1(new_n19902_), .A2(new_n19856_), .ZN(new_n19903_));
  NOR2_X1    g16792(.A1(new_n19863_), .A2(new_n13783_), .ZN(new_n19904_));
  NAND2_X1   g16793(.A1(new_n19903_), .A2(new_n19904_), .ZN(new_n19905_));
  NOR2_X1    g16794(.A1(new_n19866_), .A2(pi0660), .ZN(new_n19906_));
  NAND2_X1   g16795(.A1(new_n19905_), .A2(new_n19906_), .ZN(new_n19907_));
  NOR2_X1    g16796(.A1(new_n19899_), .A2(new_n13766_), .ZN(new_n19908_));
  XOR2_X1    g16797(.A1(new_n19908_), .A2(new_n14090_), .Z(new_n19909_));
  NAND4_X1   g16798(.A1(new_n19907_), .A2(pi0785), .A3(new_n19856_), .A4(new_n19909_), .ZN(new_n19910_));
  NAND2_X1   g16799(.A1(new_n19910_), .A2(new_n19900_), .ZN(new_n19911_));
  NAND2_X1   g16800(.A1(new_n19911_), .A2(new_n13855_), .ZN(new_n19912_));
  NOR2_X1    g16801(.A1(new_n19911_), .A2(new_n13816_), .ZN(new_n19913_));
  XOR2_X1    g16802(.A1(new_n19913_), .A2(new_n13818_), .Z(new_n19914_));
  NAND3_X1   g16803(.A1(new_n19914_), .A2(new_n14049_), .A3(new_n19856_), .ZN(new_n19915_));
  NAND3_X1   g16804(.A1(new_n19915_), .A2(new_n13823_), .A3(new_n19872_), .ZN(new_n19916_));
  AND3_X2    g16805(.A1(new_n19916_), .A2(new_n13823_), .A3(new_n19870_), .Z(new_n19917_));
  NOR2_X1    g16806(.A1(new_n19911_), .A2(new_n13817_), .ZN(new_n19918_));
  XOR2_X1    g16807(.A1(new_n19918_), .A2(new_n13819_), .Z(new_n19919_));
  NOR3_X1    g16808(.A1(new_n19919_), .A2(new_n13855_), .A3(new_n19857_), .ZN(new_n19920_));
  INV_X1     g16809(.I(new_n19920_), .ZN(new_n19921_));
  OAI21_X1   g16810(.A1(new_n19917_), .A2(new_n19921_), .B(new_n19912_), .ZN(new_n19922_));
  NOR2_X1    g16811(.A1(new_n19922_), .A2(new_n13860_), .ZN(new_n19923_));
  XOR2_X1    g16812(.A1(new_n19923_), .A2(new_n13904_), .Z(new_n19924_));
  NOR2_X1    g16813(.A1(new_n19924_), .A2(new_n19859_), .ZN(new_n19925_));
  NAND2_X1   g16814(.A1(new_n19881_), .A2(new_n13884_), .ZN(new_n19926_));
  INV_X1     g16815(.I(new_n19922_), .ZN(new_n19927_));
  AOI21_X1   g16816(.A1(new_n19927_), .A2(new_n14143_), .B(pi0789), .ZN(new_n19928_));
  OAI21_X1   g16817(.A1(new_n19925_), .A2(new_n19926_), .B(new_n19928_), .ZN(new_n19929_));
  NOR2_X1    g16818(.A1(new_n19922_), .A2(new_n13868_), .ZN(new_n19930_));
  XOR2_X1    g16819(.A1(new_n19930_), .A2(new_n13903_), .Z(new_n19931_));
  NAND2_X1   g16820(.A1(new_n19877_), .A2(new_n19018_), .ZN(new_n19932_));
  AOI21_X1   g16821(.A1(new_n19931_), .A2(new_n19858_), .B(new_n19932_), .ZN(new_n19933_));
  AOI21_X1   g16822(.A1(new_n19929_), .A2(new_n19933_), .B(new_n19886_), .ZN(new_n19934_));
  NAND2_X1   g16823(.A1(new_n19883_), .A2(new_n16372_), .ZN(new_n19935_));
  OAI21_X1   g16824(.A1(new_n16372_), .A2(new_n19848_), .B(new_n19935_), .ZN(new_n19936_));
  NAND3_X1   g16825(.A1(new_n19936_), .A2(new_n18929_), .A3(new_n19860_), .ZN(new_n19937_));
  NAND2_X1   g16826(.A1(new_n19937_), .A2(new_n16569_), .ZN(new_n19938_));
  XOR2_X1    g16827(.A1(new_n19938_), .A2(new_n16572_), .Z(new_n19939_));
  AOI21_X1   g16828(.A1(new_n19022_), .A2(new_n19937_), .B(new_n19939_), .ZN(new_n19940_));
  INV_X1     g16829(.I(new_n19848_), .ZN(new_n19941_));
  NAND2_X1   g16830(.A1(new_n19883_), .A2(new_n13963_), .ZN(new_n19942_));
  XNOR2_X1   g16831(.A1(new_n19942_), .A2(new_n19028_), .ZN(new_n19943_));
  NOR3_X1    g16832(.A1(new_n19943_), .A2(new_n16424_), .A3(new_n19941_), .ZN(new_n19944_));
  OAI21_X1   g16833(.A1(new_n19940_), .A2(new_n16574_), .B(new_n19944_), .ZN(new_n19945_));
  NOR4_X1    g16834(.A1(new_n19859_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n19946_));
  NOR2_X1    g16835(.A1(new_n19946_), .A2(new_n14005_), .ZN(new_n19947_));
  XOR2_X1    g16836(.A1(new_n19947_), .A2(new_n14007_), .Z(new_n19948_));
  NAND2_X1   g16837(.A1(new_n19948_), .A2(new_n19848_), .ZN(new_n19949_));
  NOR2_X1    g16838(.A1(new_n19941_), .A2(pi0647), .ZN(new_n19950_));
  AOI21_X1   g16839(.A1(new_n19946_), .A2(pi0647), .B(new_n19950_), .ZN(new_n19951_));
  NOR2_X1    g16840(.A1(new_n19936_), .A2(new_n13994_), .ZN(new_n19952_));
  XNOR2_X1   g16841(.A1(new_n19952_), .A2(new_n19033_), .ZN(new_n19953_));
  AOI22_X1   g16842(.A1(new_n19953_), .A2(new_n19848_), .B1(new_n14206_), .B2(new_n19951_), .ZN(new_n19954_));
  NOR3_X1    g16843(.A1(new_n19954_), .A2(new_n14010_), .A3(new_n19949_), .ZN(new_n19955_));
  OAI22_X1   g16844(.A1(new_n19934_), .A2(new_n19945_), .B1(new_n12776_), .B2(new_n19955_), .ZN(new_n19956_));
  AOI21_X1   g16845(.A1(new_n19951_), .A2(pi1157), .B(new_n12776_), .ZN(new_n19957_));
  AOI22_X1   g16846(.A1(new_n19949_), .A2(new_n19957_), .B1(new_n12776_), .B2(new_n19946_), .ZN(new_n19958_));
  NAND2_X1   g16847(.A1(new_n19956_), .A2(pi0644), .ZN(new_n19959_));
  XOR2_X1    g16848(.A1(new_n19959_), .A2(new_n14205_), .Z(new_n19960_));
  NOR2_X1    g16849(.A1(new_n19960_), .A2(new_n19958_), .ZN(new_n19961_));
  NOR2_X1    g16850(.A1(new_n19936_), .A2(new_n18968_), .ZN(new_n19962_));
  NAND2_X1   g16851(.A1(new_n18967_), .A2(new_n19848_), .ZN(new_n19963_));
  XOR2_X1    g16852(.A1(new_n19962_), .A2(new_n19963_), .Z(new_n19964_));
  NAND2_X1   g16853(.A1(new_n19964_), .A2(pi0715), .ZN(new_n19965_));
  XOR2_X1    g16854(.A1(new_n19965_), .A2(new_n14205_), .Z(new_n19966_));
  OAI21_X1   g16855(.A1(new_n19966_), .A2(new_n19941_), .B(new_n14203_), .ZN(new_n19967_));
  NAND2_X1   g16856(.A1(new_n19964_), .A2(pi0644), .ZN(new_n19968_));
  XOR2_X1    g16857(.A1(new_n19968_), .A2(new_n14217_), .Z(new_n19969_));
  AOI21_X1   g16858(.A1(new_n19969_), .A2(new_n19848_), .B(pi1160), .ZN(new_n19970_));
  OAI21_X1   g16859(.A1(new_n19961_), .A2(new_n19967_), .B(new_n19970_), .ZN(new_n19971_));
  NAND2_X1   g16860(.A1(new_n19956_), .A2(pi0715), .ZN(new_n19972_));
  XOR2_X1    g16861(.A1(new_n19972_), .A2(new_n14205_), .Z(new_n19973_));
  NOR2_X1    g16862(.A1(new_n19973_), .A2(new_n19958_), .ZN(new_n19974_));
  AOI21_X1   g16863(.A1(new_n19971_), .A2(new_n19974_), .B(new_n14799_), .ZN(new_n19975_));
  XOR2_X1    g16864(.A1(new_n19975_), .A2(new_n14801_), .Z(new_n19976_));
  NOR2_X1    g16865(.A1(new_n7240_), .A2(pi0177), .ZN(new_n19977_));
  NOR4_X1    g16866(.A1(new_n19976_), .A2(pi0832), .A3(new_n19956_), .A4(new_n19977_), .ZN(new_n19978_));
  AOI21_X1   g16867(.A1(new_n19847_), .A2(new_n7240_), .B(new_n19978_), .ZN(new_n19979_));
  NOR2_X1    g16868(.A1(new_n19846_), .A2(new_n19836_), .ZN(new_n19980_));
  AOI21_X1   g16869(.A1(new_n19980_), .A2(pi0715), .B(new_n14217_), .ZN(new_n19981_));
  NOR4_X1    g16870(.A1(new_n19846_), .A2(new_n19836_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n19982_));
  NOR2_X1    g16871(.A1(new_n19981_), .A2(new_n19982_), .ZN(new_n19983_));
  OAI21_X1   g16872(.A1(new_n12776_), .A2(new_n19843_), .B(new_n19845_), .ZN(new_n19984_));
  INV_X1     g16873(.I(new_n19829_), .ZN(new_n19985_));
  OAI21_X1   g16874(.A1(new_n19816_), .A2(new_n19805_), .B(new_n19985_), .ZN(new_n19986_));
  INV_X1     g16875(.I(new_n19844_), .ZN(new_n19987_));
  OAI21_X1   g16876(.A1(new_n19805_), .A2(new_n19816_), .B(new_n19987_), .ZN(new_n19988_));
  NAND3_X1   g16877(.A1(new_n19988_), .A2(new_n19986_), .A3(pi0787), .ZN(new_n19989_));
  NOR2_X1    g16878(.A1(new_n19697_), .A2(new_n14211_), .ZN(new_n19990_));
  AOI21_X1   g16879(.A1(new_n19819_), .A2(new_n14211_), .B(new_n19990_), .ZN(new_n19991_));
  OAI21_X1   g16880(.A1(new_n19697_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n19992_));
  NAND2_X1   g16881(.A1(new_n19991_), .A2(new_n19992_), .ZN(new_n19993_));
  AOI21_X1   g16882(.A1(new_n19827_), .A2(new_n19692_), .B(new_n12776_), .ZN(new_n19994_));
  NOR3_X1    g16883(.A1(new_n19832_), .A2(new_n12776_), .A3(new_n19825_), .ZN(new_n19995_));
  XNOR2_X1   g16884(.A1(new_n19994_), .A2(new_n19995_), .ZN(new_n19996_));
  AOI21_X1   g16885(.A1(new_n19993_), .A2(new_n14815_), .B(pi0644), .ZN(new_n19997_));
  AOI21_X1   g16886(.A1(new_n19984_), .A2(new_n19989_), .B(new_n19997_), .ZN(new_n19998_));
  AOI21_X1   g16887(.A1(new_n19697_), .A2(new_n14254_), .B(pi0644), .ZN(new_n19999_));
  NOR3_X1    g16888(.A1(new_n19996_), .A2(new_n19991_), .A3(new_n19999_), .ZN(new_n20000_));
  OAI21_X1   g16889(.A1(new_n19998_), .A2(pi0790), .B(new_n20000_), .ZN(new_n20001_));
  NOR3_X1    g16890(.A1(new_n19983_), .A2(new_n19979_), .A3(new_n20001_), .ZN(po0334));
  INV_X1     g16891(.I(new_n16474_), .ZN(new_n20003_));
  NAND2_X1   g16892(.A1(new_n13627_), .A2(new_n7510_), .ZN(new_n20004_));
  INV_X1     g16893(.I(new_n20004_), .ZN(new_n20005_));
  AOI21_X1   g16894(.A1(new_n7510_), .A2(new_n17500_), .B(pi0038), .ZN(new_n20006_));
  NOR2_X1    g16895(.A1(new_n13107_), .A2(new_n13109_), .ZN(new_n20007_));
  NOR2_X1    g16896(.A1(new_n7510_), .A2(new_n17500_), .ZN(new_n20008_));
  OAI21_X1   g16897(.A1(new_n20007_), .A2(new_n20008_), .B(pi0038), .ZN(new_n20009_));
  INV_X1     g16898(.I(new_n20009_), .ZN(new_n20010_));
  AOI21_X1   g16899(.A1(new_n13097_), .A2(new_n20006_), .B(new_n20010_), .ZN(new_n20011_));
  NOR2_X1    g16900(.A1(new_n3289_), .A2(pi0178), .ZN(new_n20012_));
  AOI21_X1   g16901(.A1(new_n20011_), .A2(new_n3289_), .B(new_n20012_), .ZN(new_n20013_));
  NAND2_X1   g16902(.A1(new_n20013_), .A2(new_n13776_), .ZN(new_n20014_));
  OAI21_X1   g16903(.A1(new_n15147_), .A2(new_n20005_), .B(new_n20014_), .ZN(new_n20015_));
  NAND2_X1   g16904(.A1(new_n20015_), .A2(pi0609), .ZN(new_n20016_));
  NAND2_X1   g16905(.A1(new_n20016_), .A2(pi0785), .ZN(new_n20017_));
  AOI21_X1   g16906(.A1(new_n20004_), .A2(new_n14467_), .B(pi0609), .ZN(new_n20018_));
  NOR2_X1    g16907(.A1(new_n20018_), .A2(new_n20014_), .ZN(new_n20019_));
  NAND2_X1   g16908(.A1(new_n20005_), .A2(new_n13775_), .ZN(new_n20020_));
  OAI21_X1   g16909(.A1(new_n13775_), .A2(new_n20013_), .B(new_n20020_), .ZN(new_n20021_));
  NAND3_X1   g16910(.A1(new_n20021_), .A2(pi0785), .A3(new_n20019_), .ZN(new_n20022_));
  XNOR2_X1   g16911(.A1(new_n20017_), .A2(new_n20022_), .ZN(new_n20023_));
  NAND2_X1   g16912(.A1(new_n20023_), .A2(pi0618), .ZN(new_n20024_));
  XOR2_X1    g16913(.A1(new_n20024_), .A2(new_n13819_), .Z(new_n20025_));
  NAND2_X1   g16914(.A1(new_n20025_), .A2(new_n20005_), .ZN(new_n20026_));
  NAND2_X1   g16915(.A1(new_n20026_), .A2(pi0781), .ZN(new_n20027_));
  NAND2_X1   g16916(.A1(new_n20023_), .A2(pi1154), .ZN(new_n20028_));
  XOR2_X1    g16917(.A1(new_n20028_), .A2(new_n13819_), .Z(new_n20029_));
  NAND2_X1   g16918(.A1(new_n20029_), .A2(new_n20005_), .ZN(new_n20030_));
  NOR3_X1    g16919(.A1(new_n20030_), .A2(new_n13855_), .A3(new_n20023_), .ZN(new_n20031_));
  XNOR2_X1   g16920(.A1(new_n20031_), .A2(new_n20027_), .ZN(new_n20032_));
  NAND3_X1   g16921(.A1(new_n20032_), .A2(pi0619), .A3(pi1159), .ZN(new_n20033_));
  XOR2_X1    g16922(.A1(new_n20031_), .A2(new_n20027_), .Z(new_n20034_));
  NAND3_X1   g16923(.A1(new_n20034_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n20035_));
  AOI21_X1   g16924(.A1(new_n20033_), .A2(new_n20035_), .B(new_n20004_), .ZN(new_n20036_));
  NOR2_X1    g16925(.A1(new_n20005_), .A2(new_n13880_), .ZN(new_n20037_));
  OAI21_X1   g16926(.A1(new_n13721_), .A2(new_n17495_), .B(new_n7510_), .ZN(new_n20038_));
  NAND2_X1   g16927(.A1(new_n16715_), .A2(new_n7510_), .ZN(new_n20039_));
  NAND4_X1   g16928(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n20038_), .A4(new_n20039_), .ZN(new_n20040_));
  NAND2_X1   g16929(.A1(new_n20040_), .A2(new_n14424_), .ZN(new_n20041_));
  NAND2_X1   g16930(.A1(new_n20041_), .A2(pi0178), .ZN(new_n20042_));
  OAI21_X1   g16931(.A1(new_n20042_), .A2(new_n20004_), .B(new_n3290_), .ZN(new_n20043_));
  NAND2_X1   g16932(.A1(new_n20043_), .A2(pi0688), .ZN(new_n20044_));
  NAND2_X1   g16933(.A1(new_n20044_), .A2(pi0625), .ZN(new_n20045_));
  XOR2_X1    g16934(.A1(new_n20045_), .A2(new_n13620_), .Z(new_n20046_));
  NAND2_X1   g16935(.A1(new_n20046_), .A2(new_n20005_), .ZN(new_n20047_));
  NAND2_X1   g16936(.A1(new_n20047_), .A2(pi0778), .ZN(new_n20048_));
  NAND2_X1   g16937(.A1(new_n20044_), .A2(pi1153), .ZN(new_n20049_));
  XOR2_X1    g16938(.A1(new_n20049_), .A2(new_n13620_), .Z(new_n20050_));
  NAND2_X1   g16939(.A1(new_n20050_), .A2(new_n20005_), .ZN(new_n20051_));
  NOR3_X1    g16940(.A1(new_n20051_), .A2(new_n13748_), .A3(new_n20044_), .ZN(new_n20052_));
  XNOR2_X1   g16941(.A1(new_n20052_), .A2(new_n20048_), .ZN(new_n20053_));
  NOR2_X1    g16942(.A1(new_n20004_), .A2(new_n13805_), .ZN(new_n20054_));
  AOI21_X1   g16943(.A1(new_n20053_), .A2(new_n13805_), .B(new_n20054_), .ZN(new_n20055_));
  AOI21_X1   g16944(.A1(new_n20055_), .A2(new_n13880_), .B(new_n20037_), .ZN(new_n20056_));
  NOR2_X1    g16945(.A1(new_n13453_), .A2(new_n7510_), .ZN(new_n20057_));
  XOR2_X1    g16946(.A1(new_n20057_), .A2(new_n20008_), .Z(new_n20058_));
  NAND2_X1   g16947(.A1(new_n20058_), .A2(new_n13521_), .ZN(new_n20059_));
  NAND3_X1   g16948(.A1(new_n14270_), .A2(pi0178), .A3(pi0760), .ZN(new_n20060_));
  NAND3_X1   g16949(.A1(new_n14272_), .A2(new_n7510_), .A3(pi0760), .ZN(new_n20061_));
  AOI21_X1   g16950(.A1(new_n20060_), .A2(new_n20061_), .B(new_n13152_), .ZN(new_n20062_));
  NAND3_X1   g16951(.A1(new_n13198_), .A2(pi0178), .A3(pi0760), .ZN(new_n20063_));
  NAND3_X1   g16952(.A1(new_n13200_), .A2(pi0178), .A3(new_n17500_), .ZN(new_n20064_));
  AOI21_X1   g16953(.A1(new_n20064_), .A2(new_n20063_), .B(new_n13191_), .ZN(new_n20065_));
  OAI21_X1   g16954(.A1(new_n20062_), .A2(new_n3262_), .B(new_n20065_), .ZN(new_n20066_));
  NAND3_X1   g16955(.A1(new_n20059_), .A2(new_n3183_), .A3(new_n20066_), .ZN(new_n20067_));
  NOR2_X1    g16956(.A1(new_n14284_), .A2(new_n17500_), .ZN(new_n20068_));
  XOR2_X1    g16957(.A1(new_n20068_), .A2(new_n20008_), .Z(new_n20069_));
  NAND3_X1   g16958(.A1(new_n20067_), .A2(new_n20069_), .A3(new_n13359_), .ZN(new_n20070_));
  NAND3_X1   g16959(.A1(new_n20070_), .A2(new_n17495_), .A3(new_n3290_), .ZN(new_n20071_));
  OAI21_X1   g16960(.A1(new_n15587_), .A2(new_n7510_), .B(new_n17500_), .ZN(new_n20072_));
  NAND2_X1   g16961(.A1(new_n20072_), .A2(new_n13209_), .ZN(new_n20073_));
  NOR2_X1    g16962(.A1(new_n13105_), .A2(pi0760), .ZN(new_n20074_));
  INV_X1     g16963(.I(new_n20074_), .ZN(new_n20075_));
  NAND2_X1   g16964(.A1(new_n20075_), .A2(new_n16751_), .ZN(new_n20076_));
  NAND4_X1   g16965(.A1(new_n5503_), .A2(new_n20076_), .A3(pi0178), .A4(new_n3290_), .ZN(new_n20077_));
  AOI21_X1   g16966(.A1(new_n20073_), .A2(new_n3259_), .B(new_n20077_), .ZN(new_n20078_));
  AOI21_X1   g16967(.A1(new_n20071_), .A2(new_n20078_), .B(pi0688), .ZN(new_n20079_));
  NOR2_X1    g16968(.A1(new_n20079_), .A2(new_n20011_), .ZN(new_n20080_));
  INV_X1     g16969(.I(new_n20080_), .ZN(new_n20081_));
  INV_X1     g16970(.I(new_n20013_), .ZN(new_n20082_));
  NOR2_X1    g16971(.A1(new_n20080_), .A2(new_n13613_), .ZN(new_n20083_));
  XOR2_X1    g16972(.A1(new_n20083_), .A2(new_n13615_), .Z(new_n20084_));
  NAND2_X1   g16973(.A1(new_n20051_), .A2(new_n14081_), .ZN(new_n20085_));
  AOI21_X1   g16974(.A1(new_n20084_), .A2(new_n20082_), .B(new_n20085_), .ZN(new_n20086_));
  INV_X1     g16975(.I(new_n20086_), .ZN(new_n20087_));
  NOR2_X1    g16976(.A1(new_n20080_), .A2(new_n13614_), .ZN(new_n20088_));
  XOR2_X1    g16977(.A1(new_n20088_), .A2(new_n13615_), .Z(new_n20089_));
  AOI21_X1   g16978(.A1(new_n20089_), .A2(new_n20082_), .B(pi0608), .ZN(new_n20090_));
  NAND2_X1   g16979(.A1(new_n20087_), .A2(new_n20090_), .ZN(new_n20091_));
  NOR2_X1    g16980(.A1(new_n20047_), .A2(new_n13748_), .ZN(new_n20092_));
  AOI22_X1   g16981(.A1(new_n20091_), .A2(new_n20092_), .B1(new_n13748_), .B2(new_n20081_), .ZN(new_n20093_));
  AOI21_X1   g16982(.A1(new_n20093_), .A2(pi1155), .B(new_n14694_), .ZN(new_n20094_));
  INV_X1     g16983(.I(new_n20090_), .ZN(new_n20095_));
  NOR2_X1    g16984(.A1(new_n20095_), .A2(new_n20086_), .ZN(new_n20096_));
  INV_X1     g16985(.I(new_n20092_), .ZN(new_n20097_));
  OAI22_X1   g16986(.A1(new_n20096_), .A2(new_n20097_), .B1(pi0778), .B2(new_n20080_), .ZN(new_n20098_));
  NOR3_X1    g16987(.A1(new_n20098_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n20099_));
  OAI21_X1   g16988(.A1(new_n20099_), .A2(new_n20094_), .B(new_n20053_), .ZN(new_n20100_));
  NAND2_X1   g16989(.A1(new_n20016_), .A2(pi0660), .ZN(new_n20101_));
  INV_X1     g16990(.I(new_n20101_), .ZN(new_n20102_));
  NOR2_X1    g16991(.A1(new_n20019_), .A2(pi0660), .ZN(new_n20103_));
  INV_X1     g16992(.I(new_n20103_), .ZN(new_n20104_));
  AOI21_X1   g16993(.A1(new_n20100_), .A2(new_n20102_), .B(new_n20104_), .ZN(new_n20105_));
  NOR2_X1    g16994(.A1(new_n20098_), .A2(new_n13766_), .ZN(new_n20106_));
  NOR2_X1    g16995(.A1(new_n20106_), .A2(new_n14694_), .ZN(new_n20107_));
  NAND2_X1   g16996(.A1(new_n20106_), .A2(new_n14694_), .ZN(new_n20108_));
  INV_X1     g16997(.I(new_n20108_), .ZN(new_n20109_));
  INV_X1     g16998(.I(new_n20053_), .ZN(new_n20110_));
  NOR2_X1    g16999(.A1(new_n20110_), .A2(new_n13801_), .ZN(new_n20111_));
  OAI21_X1   g17000(.A1(new_n20109_), .A2(new_n20107_), .B(new_n20111_), .ZN(new_n20112_));
  OAI22_X1   g17001(.A1(new_n20112_), .A2(new_n20105_), .B1(pi0785), .B2(new_n20093_), .ZN(new_n20113_));
  NAND3_X1   g17002(.A1(new_n20113_), .A2(pi0618), .A3(pi1154), .ZN(new_n20114_));
  NAND3_X1   g17003(.A1(new_n20098_), .A2(pi0609), .A3(pi1155), .ZN(new_n20115_));
  NAND3_X1   g17004(.A1(new_n20093_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n20116_));
  AOI21_X1   g17005(.A1(new_n20115_), .A2(new_n20116_), .B(new_n20110_), .ZN(new_n20117_));
  OAI21_X1   g17006(.A1(new_n20117_), .A2(new_n20101_), .B(new_n20103_), .ZN(new_n20118_));
  NAND2_X1   g17007(.A1(new_n20093_), .A2(pi0609), .ZN(new_n20119_));
  NAND2_X1   g17008(.A1(new_n20119_), .A2(new_n14090_), .ZN(new_n20120_));
  INV_X1     g17009(.I(new_n20111_), .ZN(new_n20121_));
  AOI21_X1   g17010(.A1(new_n20108_), .A2(new_n20120_), .B(new_n20121_), .ZN(new_n20122_));
  AOI22_X1   g17011(.A1(new_n20118_), .A2(new_n20122_), .B1(new_n13801_), .B2(new_n20098_), .ZN(new_n20123_));
  NAND3_X1   g17012(.A1(new_n20123_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n20124_));
  AOI21_X1   g17013(.A1(new_n20114_), .A2(new_n20124_), .B(new_n20055_), .ZN(new_n20125_));
  NAND2_X1   g17014(.A1(new_n20026_), .A2(pi0627), .ZN(new_n20126_));
  OAI21_X1   g17015(.A1(new_n20125_), .A2(new_n20126_), .B(pi0781), .ZN(new_n20127_));
  INV_X1     g17016(.I(new_n20055_), .ZN(new_n20128_));
  AOI21_X1   g17017(.A1(new_n20123_), .A2(pi0618), .B(new_n13819_), .ZN(new_n20129_));
  NOR3_X1    g17018(.A1(new_n20113_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n20130_));
  OAI21_X1   g17019(.A1(new_n20130_), .A2(new_n20129_), .B(new_n20128_), .ZN(new_n20131_));
  AND3_X2    g17020(.A1(new_n20113_), .A2(new_n19177_), .A3(new_n20030_), .Z(new_n20132_));
  NAND3_X1   g17021(.A1(new_n20127_), .A2(new_n20131_), .A3(new_n20132_), .ZN(new_n20133_));
  AOI21_X1   g17022(.A1(new_n20123_), .A2(pi1154), .B(new_n13819_), .ZN(new_n20134_));
  NOR3_X1    g17023(.A1(new_n20113_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n20135_));
  OAI21_X1   g17024(.A1(new_n20135_), .A2(new_n20134_), .B(new_n20128_), .ZN(new_n20136_));
  INV_X1     g17025(.I(new_n20126_), .ZN(new_n20137_));
  AOI21_X1   g17026(.A1(new_n20136_), .A2(new_n20137_), .B(new_n13855_), .ZN(new_n20138_));
  NAND4_X1   g17027(.A1(new_n20131_), .A2(new_n19177_), .A3(new_n20030_), .A4(new_n20113_), .ZN(new_n20139_));
  NAND2_X1   g17028(.A1(new_n20139_), .A2(new_n20138_), .ZN(new_n20140_));
  NAND2_X1   g17029(.A1(new_n20140_), .A2(new_n20133_), .ZN(new_n20141_));
  NAND3_X1   g17030(.A1(new_n20141_), .A2(pi0619), .A3(pi1159), .ZN(new_n20142_));
  NAND4_X1   g17031(.A1(new_n20140_), .A2(new_n20133_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n20143_));
  AOI21_X1   g17032(.A1(new_n20142_), .A2(new_n20143_), .B(new_n20056_), .ZN(new_n20144_));
  OAI21_X1   g17033(.A1(new_n20144_), .A2(new_n20003_), .B(new_n20036_), .ZN(new_n20145_));
  NAND2_X1   g17034(.A1(new_n20141_), .A2(new_n13896_), .ZN(new_n20146_));
  NOR2_X1    g17035(.A1(new_n20036_), .A2(new_n13896_), .ZN(new_n20147_));
  NAND3_X1   g17036(.A1(new_n20032_), .A2(pi0619), .A3(pi1159), .ZN(new_n20148_));
  NAND3_X1   g17037(.A1(new_n20034_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n20149_));
  NAND2_X1   g17038(.A1(new_n20148_), .A2(new_n20149_), .ZN(new_n20150_));
  NAND4_X1   g17039(.A1(new_n20150_), .A2(pi0789), .A3(new_n20005_), .A4(new_n20032_), .ZN(new_n20151_));
  OR2_X2     g17040(.A1(new_n20151_), .A2(new_n20147_), .Z(new_n20152_));
  NAND2_X1   g17041(.A1(new_n20151_), .A2(new_n20147_), .ZN(new_n20153_));
  NAND2_X1   g17042(.A1(new_n20152_), .A2(new_n20153_), .ZN(new_n20154_));
  NAND3_X1   g17043(.A1(new_n20154_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n20155_));
  NAND4_X1   g17044(.A1(new_n20152_), .A2(new_n13901_), .A3(new_n13962_), .A4(new_n20153_), .ZN(new_n20156_));
  AOI21_X1   g17045(.A1(new_n20155_), .A2(new_n20156_), .B(new_n20004_), .ZN(new_n20157_));
  NOR2_X1    g17046(.A1(new_n20004_), .A2(new_n13919_), .ZN(new_n20158_));
  NAND2_X1   g17047(.A1(new_n20056_), .A2(new_n13919_), .ZN(new_n20159_));
  INV_X1     g17048(.I(new_n20159_), .ZN(new_n20160_));
  NOR2_X1    g17049(.A1(new_n20160_), .A2(new_n20158_), .ZN(new_n20161_));
  NOR2_X1    g17050(.A1(new_n20161_), .A2(new_n14162_), .ZN(new_n20162_));
  OAI21_X1   g17051(.A1(new_n20157_), .A2(new_n20162_), .B(new_n19204_), .ZN(new_n20163_));
  NOR2_X1    g17052(.A1(new_n20154_), .A2(new_n19208_), .ZN(new_n20164_));
  XNOR2_X1   g17053(.A1(new_n20164_), .A2(new_n19028_), .ZN(new_n20165_));
  NOR2_X1    g17054(.A1(new_n20004_), .A2(new_n15479_), .ZN(new_n20166_));
  NAND4_X1   g17055(.A1(new_n20146_), .A2(new_n20163_), .A3(new_n20165_), .A4(new_n20166_), .ZN(new_n20167_));
  NAND2_X1   g17056(.A1(new_n20145_), .A2(new_n20167_), .ZN(new_n20168_));
  INV_X1     g17057(.I(new_n20056_), .ZN(new_n20169_));
  NAND3_X1   g17058(.A1(new_n20140_), .A2(new_n20133_), .A3(pi0619), .ZN(new_n20170_));
  XOR2_X1    g17059(.A1(new_n20170_), .A2(new_n13904_), .Z(new_n20171_));
  NAND2_X1   g17060(.A1(new_n20150_), .A2(new_n20005_), .ZN(new_n20172_));
  NOR2_X1    g17061(.A1(new_n16419_), .A2(pi0648), .ZN(new_n20173_));
  NAND2_X1   g17062(.A1(new_n20172_), .A2(new_n20173_), .ZN(new_n20174_));
  AOI21_X1   g17063(.A1(new_n20171_), .A2(new_n20169_), .B(new_n20174_), .ZN(new_n20175_));
  AOI21_X1   g17064(.A1(new_n20168_), .A2(new_n20175_), .B(pi0792), .ZN(new_n20176_));
  NOR2_X1    g17065(.A1(new_n20005_), .A2(new_n13966_), .ZN(new_n20177_));
  NOR3_X1    g17066(.A1(new_n20160_), .A2(new_n13965_), .A3(new_n20158_), .ZN(new_n20178_));
  NOR2_X1    g17067(.A1(new_n20178_), .A2(new_n20177_), .ZN(new_n20179_));
  INV_X1     g17068(.I(new_n20179_), .ZN(new_n20180_));
  NAND3_X1   g17069(.A1(new_n20180_), .A2(pi0628), .A3(pi1156), .ZN(new_n20181_));
  NAND3_X1   g17070(.A1(new_n20179_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n20182_));
  AOI21_X1   g17071(.A1(new_n20181_), .A2(new_n20182_), .B(new_n20004_), .ZN(new_n20183_));
  NOR2_X1    g17072(.A1(new_n20183_), .A2(new_n12777_), .ZN(new_n20184_));
  NAND3_X1   g17073(.A1(new_n20180_), .A2(pi0628), .A3(pi1156), .ZN(new_n20185_));
  NAND3_X1   g17074(.A1(new_n20179_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n20186_));
  AOI21_X1   g17075(.A1(new_n20185_), .A2(new_n20186_), .B(new_n20004_), .ZN(new_n20187_));
  NAND3_X1   g17076(.A1(new_n20187_), .A2(pi0792), .A3(new_n20180_), .ZN(new_n20188_));
  NOR2_X1    g17077(.A1(new_n20188_), .A2(new_n20184_), .ZN(new_n20189_));
  INV_X1     g17078(.I(new_n20189_), .ZN(new_n20190_));
  NAND2_X1   g17079(.A1(new_n20188_), .A2(new_n20184_), .ZN(new_n20191_));
  NAND2_X1   g17080(.A1(new_n20190_), .A2(new_n20191_), .ZN(new_n20192_));
  NAND2_X1   g17081(.A1(new_n20005_), .A2(new_n14005_), .ZN(new_n20193_));
  NAND2_X1   g17082(.A1(new_n20193_), .A2(pi1157), .ZN(new_n20194_));
  AOI21_X1   g17083(.A1(new_n20192_), .A2(pi0647), .B(new_n20194_), .ZN(new_n20195_));
  AOI21_X1   g17084(.A1(new_n20190_), .A2(new_n20191_), .B(pi0647), .ZN(new_n20196_));
  NOR2_X1    g17085(.A1(new_n20004_), .A2(new_n14005_), .ZN(new_n20197_));
  NOR3_X1    g17086(.A1(new_n20196_), .A2(pi1157), .A3(new_n20197_), .ZN(new_n20198_));
  OAI21_X1   g17087(.A1(new_n20198_), .A2(new_n20195_), .B(pi0787), .ZN(new_n20199_));
  OAI21_X1   g17088(.A1(pi0787), .A2(new_n20192_), .B(new_n20199_), .ZN(new_n20200_));
  NOR2_X1    g17089(.A1(new_n20005_), .A2(new_n16372_), .ZN(new_n20201_));
  NOR2_X1    g17090(.A1(new_n20154_), .A2(new_n14142_), .ZN(new_n20202_));
  OAI21_X1   g17091(.A1(new_n20202_), .A2(new_n20201_), .B(new_n13994_), .ZN(new_n20203_));
  NOR2_X1    g17092(.A1(new_n20005_), .A2(new_n13994_), .ZN(new_n20204_));
  INV_X1     g17093(.I(new_n20204_), .ZN(new_n20205_));
  AOI21_X1   g17094(.A1(new_n20203_), .A2(new_n20205_), .B(new_n14210_), .ZN(new_n20206_));
  NOR2_X1    g17095(.A1(new_n20005_), .A2(new_n14211_), .ZN(new_n20207_));
  NOR2_X1    g17096(.A1(new_n20206_), .A2(new_n20207_), .ZN(new_n20208_));
  NOR2_X1    g17097(.A1(new_n14243_), .A2(pi0644), .ZN(new_n20209_));
  NOR2_X1    g17098(.A1(new_n20208_), .A2(new_n20209_), .ZN(new_n20210_));
  NAND2_X1   g17099(.A1(new_n20210_), .A2(pi0715), .ZN(new_n20211_));
  NAND2_X1   g17100(.A1(new_n20211_), .A2(new_n14204_), .ZN(new_n20212_));
  NAND2_X1   g17101(.A1(new_n20200_), .A2(new_n20212_), .ZN(new_n20213_));
  AOI21_X1   g17102(.A1(new_n20005_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n20214_));
  NOR2_X1    g17103(.A1(new_n20214_), .A2(pi0644), .ZN(new_n20215_));
  NOR3_X1    g17104(.A1(new_n20208_), .A2(new_n14200_), .A3(new_n20215_), .ZN(new_n20216_));
  OAI21_X1   g17105(.A1(new_n20200_), .A2(new_n20216_), .B(pi0644), .ZN(new_n20217_));
  AOI21_X1   g17106(.A1(new_n20217_), .A2(new_n20213_), .B(new_n12775_), .ZN(new_n20218_));
  NOR3_X1    g17107(.A1(new_n20208_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n20219_));
  OAI21_X1   g17108(.A1(new_n20208_), .A2(new_n20215_), .B(pi0790), .ZN(new_n20220_));
  NOR2_X1    g17109(.A1(new_n20220_), .A2(new_n19379_), .ZN(new_n20221_));
  OAI21_X1   g17110(.A1(new_n20221_), .A2(new_n20219_), .B(new_n20210_), .ZN(new_n20222_));
  NAND2_X1   g17111(.A1(new_n20203_), .A2(new_n20205_), .ZN(new_n20223_));
  INV_X1     g17112(.I(new_n20191_), .ZN(new_n20224_));
  OAI21_X1   g17113(.A1(new_n20224_), .A2(new_n20189_), .B(pi0647), .ZN(new_n20225_));
  NOR2_X1    g17114(.A1(new_n20224_), .A2(new_n20189_), .ZN(new_n20226_));
  INV_X1     g17115(.I(new_n20197_), .ZN(new_n20227_));
  OAI21_X1   g17116(.A1(new_n20226_), .A2(pi0647), .B(new_n20227_), .ZN(new_n20228_));
  NAND4_X1   g17117(.A1(new_n20225_), .A2(new_n14010_), .A3(pi1157), .A4(new_n20193_), .ZN(new_n20230_));
  NAND4_X1   g17118(.A1(new_n20225_), .A2(new_n14010_), .A3(pi1157), .A4(new_n20193_), .ZN(new_n20231_));
  NAND3_X1   g17119(.A1(new_n20231_), .A2(new_n20228_), .A3(new_n14011_), .ZN(new_n20232_));
  AOI21_X1   g17120(.A1(new_n20232_), .A2(new_n20230_), .B(new_n12776_), .ZN(new_n20233_));
  OAI21_X1   g17121(.A1(new_n20233_), .A2(new_n20223_), .B(new_n16576_), .ZN(new_n20234_));
  NAND2_X1   g17122(.A1(new_n20234_), .A2(new_n20222_), .ZN(new_n20235_));
  NOR2_X1    g17123(.A1(new_n20183_), .A2(new_n13976_), .ZN(new_n20236_));
  NOR2_X1    g17124(.A1(new_n20187_), .A2(pi0629), .ZN(new_n20237_));
  NOR2_X1    g17125(.A1(new_n20236_), .A2(new_n20237_), .ZN(new_n20238_));
  NOR2_X1    g17126(.A1(new_n20202_), .A2(new_n20201_), .ZN(new_n20239_));
  NOR2_X1    g17127(.A1(new_n20239_), .A2(new_n16874_), .ZN(new_n20240_));
  NOR3_X1    g17128(.A1(new_n13219_), .A2(pi0625), .A3(pi0688), .ZN(new_n20241_));
  INV_X1     g17129(.I(new_n20241_), .ZN(new_n20242_));
  NOR2_X1    g17130(.A1(new_n9992_), .A2(pi0178), .ZN(new_n20243_));
  NOR2_X1    g17131(.A1(new_n20243_), .A2(pi1153), .ZN(new_n20244_));
  NAND2_X1   g17132(.A1(new_n20242_), .A2(new_n20244_), .ZN(new_n20245_));
  INV_X1     g17133(.I(new_n20245_), .ZN(new_n20246_));
  NOR2_X1    g17134(.A1(new_n20246_), .A2(new_n13748_), .ZN(new_n20247_));
  AOI21_X1   g17135(.A1(new_n13218_), .A2(new_n17495_), .B(new_n20243_), .ZN(new_n20248_));
  INV_X1     g17136(.I(new_n20248_), .ZN(new_n20249_));
  AOI21_X1   g17137(.A1(new_n20242_), .A2(new_n20249_), .B(new_n13614_), .ZN(new_n20250_));
  INV_X1     g17138(.I(new_n20250_), .ZN(new_n20251_));
  NOR3_X1    g17139(.A1(new_n20251_), .A2(new_n13748_), .A3(new_n20249_), .ZN(new_n20252_));
  XNOR2_X1   g17140(.A1(new_n20252_), .A2(new_n20247_), .ZN(new_n20253_));
  NAND2_X1   g17141(.A1(new_n20253_), .A2(new_n14049_), .ZN(new_n20254_));
  NOR2_X1    g17142(.A1(new_n20254_), .A2(new_n14051_), .ZN(new_n20255_));
  INV_X1     g17143(.I(new_n20255_), .ZN(new_n20256_));
  NOR4_X1    g17144(.A1(new_n20256_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n20257_));
  NOR2_X1    g17145(.A1(new_n20257_), .A2(new_n14005_), .ZN(new_n20258_));
  XOR2_X1    g17146(.A1(new_n20258_), .A2(new_n14007_), .Z(new_n20259_));
  NAND2_X1   g17147(.A1(new_n20259_), .A2(new_n20243_), .ZN(new_n20260_));
  INV_X1     g17148(.I(new_n20243_), .ZN(new_n20261_));
  NOR2_X1    g17149(.A1(new_n20261_), .A2(pi0647), .ZN(new_n20262_));
  AOI21_X1   g17150(.A1(new_n20257_), .A2(pi0647), .B(new_n20262_), .ZN(new_n20263_));
  AOI21_X1   g17151(.A1(new_n20263_), .A2(pi1157), .B(new_n12776_), .ZN(new_n20264_));
  AOI22_X1   g17152(.A1(new_n20260_), .A2(new_n20264_), .B1(new_n12776_), .B2(new_n20257_), .ZN(new_n20265_));
  NOR2_X1    g17153(.A1(new_n20256_), .A2(new_n14163_), .ZN(new_n20266_));
  NOR2_X1    g17154(.A1(new_n20074_), .A2(new_n20243_), .ZN(new_n20267_));
  INV_X1     g17155(.I(new_n20267_), .ZN(new_n20268_));
  NAND3_X1   g17156(.A1(new_n20268_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n20269_));
  AOI21_X1   g17157(.A1(new_n20269_), .A2(new_n16444_), .B(new_n20075_), .ZN(new_n20270_));
  NOR2_X1    g17158(.A1(new_n20270_), .A2(new_n13801_), .ZN(new_n20271_));
  NOR2_X1    g17159(.A1(new_n20243_), .A2(pi1155), .ZN(new_n20272_));
  NOR3_X1    g17160(.A1(new_n20075_), .A2(new_n16444_), .A3(new_n20272_), .ZN(new_n20273_));
  NAND4_X1   g17161(.A1(new_n20273_), .A2(new_n20268_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n20274_));
  XOR2_X1    g17162(.A1(new_n20271_), .A2(new_n20274_), .Z(new_n20275_));
  NOR2_X1    g17163(.A1(new_n20275_), .A2(new_n13817_), .ZN(new_n20276_));
  OAI21_X1   g17164(.A1(new_n20276_), .A2(pi0618), .B(new_n9992_), .ZN(new_n20277_));
  NAND2_X1   g17165(.A1(new_n20277_), .A2(pi0781), .ZN(new_n20278_));
  OAI21_X1   g17166(.A1(new_n20276_), .A2(new_n9992_), .B(pi0618), .ZN(new_n20279_));
  NOR3_X1    g17167(.A1(new_n20279_), .A2(new_n13855_), .A3(new_n20275_), .ZN(new_n20280_));
  XOR2_X1    g17168(.A1(new_n20280_), .A2(new_n20278_), .Z(new_n20281_));
  NOR2_X1    g17169(.A1(new_n20281_), .A2(new_n13868_), .ZN(new_n20282_));
  OAI21_X1   g17170(.A1(new_n20282_), .A2(pi0619), .B(new_n9992_), .ZN(new_n20283_));
  NAND2_X1   g17171(.A1(new_n20283_), .A2(pi0789), .ZN(new_n20284_));
  OAI21_X1   g17172(.A1(new_n20282_), .A2(new_n9992_), .B(pi0619), .ZN(new_n20285_));
  NOR3_X1    g17173(.A1(new_n20285_), .A2(new_n13896_), .A3(new_n20281_), .ZN(new_n20286_));
  XOR2_X1    g17174(.A1(new_n20286_), .A2(new_n20284_), .Z(new_n20287_));
  NAND2_X1   g17175(.A1(new_n20287_), .A2(new_n13962_), .ZN(new_n20288_));
  XOR2_X1    g17176(.A1(new_n20288_), .A2(new_n18976_), .Z(new_n20289_));
  AOI22_X1   g17177(.A1(new_n20289_), .A2(new_n20243_), .B1(new_n16639_), .B2(new_n20266_), .ZN(new_n20290_));
  NOR2_X1    g17178(.A1(new_n20248_), .A2(new_n13203_), .ZN(new_n20291_));
  NAND2_X1   g17179(.A1(new_n20291_), .A2(pi0625), .ZN(new_n20292_));
  NAND3_X1   g17180(.A1(new_n20292_), .A2(pi1153), .A3(new_n20267_), .ZN(new_n20293_));
  NOR2_X1    g17181(.A1(new_n20246_), .A2(new_n14081_), .ZN(new_n20294_));
  AOI21_X1   g17182(.A1(new_n20294_), .A2(new_n20293_), .B(new_n13748_), .ZN(new_n20295_));
  NOR2_X1    g17183(.A1(new_n20268_), .A2(new_n20291_), .ZN(new_n20296_));
  INV_X1     g17184(.I(new_n20292_), .ZN(new_n20297_));
  OAI21_X1   g17185(.A1(new_n20296_), .A2(new_n20297_), .B(new_n20244_), .ZN(new_n20298_));
  NAND4_X1   g17186(.A1(new_n20298_), .A2(new_n13749_), .A3(new_n20251_), .A4(new_n20296_), .ZN(new_n20299_));
  XNOR2_X1   g17187(.A1(new_n20299_), .A2(new_n20295_), .ZN(new_n20300_));
  NAND2_X1   g17188(.A1(new_n20300_), .A2(new_n13801_), .ZN(new_n20301_));
  NOR2_X1    g17189(.A1(new_n20270_), .A2(pi0660), .ZN(new_n20305_));
  NOR2_X1    g17190(.A1(new_n20300_), .A2(new_n13766_), .ZN(new_n20306_));
  XOR2_X1    g17191(.A1(new_n20306_), .A2(new_n14090_), .Z(new_n20307_));
  NOR2_X1    g17192(.A1(new_n20253_), .A2(new_n13801_), .ZN(new_n20308_));
  NAND2_X1   g17193(.A1(new_n20307_), .A2(new_n20308_), .ZN(new_n20309_));
  OAI21_X1   g17194(.A1(new_n20309_), .A2(new_n20305_), .B(new_n20301_), .ZN(new_n20310_));
  NAND2_X1   g17195(.A1(new_n20310_), .A2(new_n13855_), .ZN(new_n20311_));
  INV_X1     g17196(.I(new_n20254_), .ZN(new_n20312_));
  NOR2_X1    g17197(.A1(new_n20310_), .A2(new_n13816_), .ZN(new_n20313_));
  XOR2_X1    g17198(.A1(new_n20313_), .A2(new_n13818_), .Z(new_n20314_));
  NAND2_X1   g17199(.A1(new_n20314_), .A2(new_n20312_), .ZN(new_n20315_));
  NAND3_X1   g17200(.A1(new_n20315_), .A2(new_n13823_), .A3(new_n20279_), .ZN(new_n20316_));
  NAND3_X1   g17201(.A1(new_n20316_), .A2(new_n13823_), .A3(new_n20277_), .ZN(new_n20317_));
  NOR2_X1    g17202(.A1(new_n20310_), .A2(new_n13817_), .ZN(new_n20318_));
  XOR2_X1    g17203(.A1(new_n20318_), .A2(new_n13818_), .Z(new_n20319_));
  NAND4_X1   g17204(.A1(new_n20317_), .A2(pi0781), .A3(new_n20312_), .A4(new_n20319_), .ZN(new_n20320_));
  NAND2_X1   g17205(.A1(new_n20320_), .A2(new_n20311_), .ZN(new_n20321_));
  NOR2_X1    g17206(.A1(new_n20321_), .A2(new_n13860_), .ZN(new_n20322_));
  XOR2_X1    g17207(.A1(new_n20322_), .A2(new_n13904_), .Z(new_n20323_));
  NOR2_X1    g17208(.A1(new_n20323_), .A2(new_n20256_), .ZN(new_n20324_));
  NAND2_X1   g17209(.A1(new_n20285_), .A2(new_n13884_), .ZN(new_n20325_));
  INV_X1     g17210(.I(new_n20321_), .ZN(new_n20326_));
  AOI21_X1   g17211(.A1(new_n20326_), .A2(new_n14143_), .B(pi0789), .ZN(new_n20327_));
  OAI21_X1   g17212(.A1(new_n20324_), .A2(new_n20325_), .B(new_n20327_), .ZN(new_n20328_));
  NOR2_X1    g17213(.A1(new_n20321_), .A2(new_n13868_), .ZN(new_n20329_));
  XOR2_X1    g17214(.A1(new_n20329_), .A2(new_n13903_), .Z(new_n20330_));
  NAND2_X1   g17215(.A1(new_n20283_), .A2(new_n19018_), .ZN(new_n20331_));
  AOI21_X1   g17216(.A1(new_n20330_), .A2(new_n20255_), .B(new_n20331_), .ZN(new_n20332_));
  AOI21_X1   g17217(.A1(new_n20328_), .A2(new_n20332_), .B(new_n20290_), .ZN(new_n20333_));
  NAND2_X1   g17218(.A1(new_n20287_), .A2(new_n16372_), .ZN(new_n20334_));
  OAI21_X1   g17219(.A1(new_n16372_), .A2(new_n20243_), .B(new_n20334_), .ZN(new_n20335_));
  NAND3_X1   g17220(.A1(new_n20335_), .A2(new_n18929_), .A3(new_n20266_), .ZN(new_n20336_));
  NAND2_X1   g17221(.A1(new_n20336_), .A2(new_n16569_), .ZN(new_n20337_));
  XOR2_X1    g17222(.A1(new_n20337_), .A2(new_n16572_), .Z(new_n20338_));
  AOI21_X1   g17223(.A1(new_n19022_), .A2(new_n20336_), .B(new_n20338_), .ZN(new_n20339_));
  NAND2_X1   g17224(.A1(new_n20287_), .A2(new_n13963_), .ZN(new_n20340_));
  XNOR2_X1   g17225(.A1(new_n20340_), .A2(new_n19028_), .ZN(new_n20341_));
  NOR3_X1    g17226(.A1(new_n20341_), .A2(new_n16424_), .A3(new_n20261_), .ZN(new_n20342_));
  OAI21_X1   g17227(.A1(new_n20339_), .A2(new_n16574_), .B(new_n20342_), .ZN(new_n20343_));
  NOR2_X1    g17228(.A1(new_n20335_), .A2(new_n13994_), .ZN(new_n20344_));
  XNOR2_X1   g17229(.A1(new_n20344_), .A2(new_n19033_), .ZN(new_n20345_));
  AOI22_X1   g17230(.A1(new_n20345_), .A2(new_n20243_), .B1(new_n14206_), .B2(new_n20263_), .ZN(new_n20346_));
  NOR3_X1    g17231(.A1(new_n20346_), .A2(new_n14010_), .A3(new_n20260_), .ZN(new_n20347_));
  OAI22_X1   g17232(.A1(new_n20333_), .A2(new_n20343_), .B1(new_n12776_), .B2(new_n20347_), .ZN(new_n20348_));
  NAND2_X1   g17233(.A1(new_n20348_), .A2(pi0644), .ZN(new_n20349_));
  XOR2_X1    g17234(.A1(new_n20349_), .A2(new_n14205_), .Z(new_n20350_));
  NOR2_X1    g17235(.A1(new_n20350_), .A2(new_n20265_), .ZN(new_n20351_));
  NOR2_X1    g17236(.A1(new_n20335_), .A2(new_n18968_), .ZN(new_n20352_));
  NAND2_X1   g17237(.A1(new_n18967_), .A2(new_n20243_), .ZN(new_n20353_));
  XOR2_X1    g17238(.A1(new_n20352_), .A2(new_n20353_), .Z(new_n20354_));
  NAND2_X1   g17239(.A1(new_n20354_), .A2(pi0715), .ZN(new_n20355_));
  XOR2_X1    g17240(.A1(new_n20355_), .A2(new_n14205_), .Z(new_n20356_));
  OAI21_X1   g17241(.A1(new_n20356_), .A2(new_n20261_), .B(new_n14203_), .ZN(new_n20357_));
  NAND2_X1   g17242(.A1(new_n20354_), .A2(pi0644), .ZN(new_n20358_));
  XOR2_X1    g17243(.A1(new_n20358_), .A2(new_n14217_), .Z(new_n20359_));
  AOI21_X1   g17244(.A1(new_n20359_), .A2(new_n20243_), .B(pi1160), .ZN(new_n20360_));
  OAI21_X1   g17245(.A1(new_n20351_), .A2(new_n20357_), .B(new_n20360_), .ZN(new_n20361_));
  NAND2_X1   g17246(.A1(new_n20348_), .A2(pi0715), .ZN(new_n20362_));
  XOR2_X1    g17247(.A1(new_n20362_), .A2(new_n14205_), .Z(new_n20363_));
  NOR2_X1    g17248(.A1(new_n20363_), .A2(new_n20265_), .ZN(new_n20364_));
  AOI21_X1   g17249(.A1(new_n20361_), .A2(new_n20364_), .B(new_n14799_), .ZN(new_n20365_));
  XOR2_X1    g17250(.A1(new_n20365_), .A2(new_n14800_), .Z(new_n20366_));
  OAI21_X1   g17251(.A1(new_n7240_), .A2(pi0178), .B(new_n14799_), .ZN(new_n20367_));
  NOR2_X1    g17252(.A1(new_n20348_), .A2(new_n20367_), .ZN(new_n20368_));
  AOI21_X1   g17253(.A1(new_n20366_), .A2(new_n20368_), .B(po1038), .ZN(new_n20369_));
  NOR3_X1    g17254(.A1(new_n20240_), .A2(new_n20238_), .A3(new_n20369_), .ZN(new_n20370_));
  OAI21_X1   g17255(.A1(new_n20218_), .A2(new_n20235_), .B(new_n20370_), .ZN(new_n20371_));
  NOR2_X1    g17256(.A1(new_n20371_), .A2(new_n20176_), .ZN(po0335));
  NOR2_X1    g17257(.A1(new_n15628_), .A2(new_n9545_), .ZN(new_n20373_));
  NOR2_X1    g17258(.A1(new_n9545_), .A2(new_n17475_), .ZN(new_n20374_));
  XOR2_X1    g17259(.A1(new_n20373_), .A2(new_n20374_), .Z(new_n20375_));
  NAND2_X1   g17260(.A1(new_n20375_), .A2(new_n15607_), .ZN(new_n20376_));
  NOR2_X1    g17261(.A1(new_n14396_), .A2(new_n17475_), .ZN(new_n20377_));
  NAND3_X1   g17262(.A1(new_n15556_), .A2(new_n19642_), .A3(new_n20374_), .ZN(new_n20378_));
  AOI21_X1   g17263(.A1(new_n20378_), .A2(new_n17475_), .B(new_n19323_), .ZN(new_n20379_));
  NOR3_X1    g17264(.A1(new_n20379_), .A2(pi0724), .A3(new_n3289_), .ZN(new_n20380_));
  NOR3_X1    g17265(.A1(new_n20380_), .A2(new_n9545_), .A3(new_n3289_), .ZN(new_n20381_));
  AOI22_X1   g17266(.A1(new_n20376_), .A2(new_n17474_), .B1(new_n20377_), .B2(new_n20381_), .ZN(new_n20382_));
  NAND3_X1   g17267(.A1(new_n14284_), .A2(pi0039), .A3(pi0179), .ZN(new_n20383_));
  NAND3_X1   g17268(.A1(new_n14285_), .A2(pi0039), .A3(new_n9545_), .ZN(new_n20384_));
  AOI21_X1   g17269(.A1(new_n20384_), .A2(new_n20383_), .B(new_n18538_), .ZN(new_n20385_));
  NAND2_X1   g17270(.A1(pi0038), .A2(pi0039), .ZN(new_n20386_));
  AOI21_X1   g17271(.A1(new_n13109_), .A2(new_n9545_), .B(new_n20386_), .ZN(new_n20387_));
  NAND3_X1   g17272(.A1(new_n14270_), .A2(pi0039), .A3(pi0179), .ZN(new_n20388_));
  NAND3_X1   g17273(.A1(new_n14272_), .A2(new_n3183_), .A3(pi0179), .ZN(new_n20389_));
  AOI21_X1   g17274(.A1(new_n20388_), .A2(new_n20389_), .B(new_n13152_), .ZN(new_n20390_));
  OAI21_X1   g17275(.A1(new_n20385_), .A2(new_n20387_), .B(new_n20390_), .ZN(new_n20391_));
  NAND2_X1   g17276(.A1(new_n20391_), .A2(pi0741), .ZN(new_n20392_));
  NOR2_X1    g17277(.A1(new_n20382_), .A2(new_n20392_), .ZN(new_n20393_));
  AOI21_X1   g17278(.A1(new_n3289_), .A2(new_n17474_), .B(pi0179), .ZN(new_n20397_));
  OR2_X2     g17279(.A1(new_n13627_), .A2(new_n20397_), .Z(new_n20398_));
  INV_X1     g17280(.I(new_n20398_), .ZN(new_n20399_));
  NOR3_X1    g17281(.A1(new_n14431_), .A2(new_n9545_), .A3(new_n14081_), .ZN(new_n20400_));
  OAI21_X1   g17282(.A1(new_n20400_), .A2(pi0625), .B(new_n20399_), .ZN(new_n20401_));
  NOR2_X1    g17283(.A1(new_n20377_), .A2(new_n3290_), .ZN(new_n20402_));
  NAND3_X1   g17284(.A1(new_n20379_), .A2(pi0179), .A3(new_n3289_), .ZN(new_n20403_));
  XNOR2_X1   g17285(.A1(new_n20403_), .A2(new_n20402_), .ZN(new_n20404_));
  INV_X1     g17286(.I(new_n20404_), .ZN(new_n20405_));
  OAI21_X1   g17287(.A1(new_n20405_), .A2(pi0625), .B(pi1153), .ZN(new_n20406_));
  OAI21_X1   g17288(.A1(new_n20406_), .A2(new_n20401_), .B(new_n13613_), .ZN(new_n20407_));
  AOI21_X1   g17289(.A1(new_n20407_), .A2(new_n20393_), .B(new_n13748_), .ZN(new_n20408_));
  NOR2_X1    g17290(.A1(new_n13613_), .A2(new_n13748_), .ZN(new_n20409_));
  NAND2_X1   g17291(.A1(new_n20393_), .A2(new_n20409_), .ZN(new_n20412_));
  INV_X1     g17292(.I(new_n20412_), .ZN(new_n20413_));
  XOR2_X1    g17293(.A1(new_n20408_), .A2(new_n20413_), .Z(new_n20414_));
  NOR2_X1    g17294(.A1(new_n14428_), .A2(pi0179), .ZN(new_n20415_));
  INV_X1     g17295(.I(new_n20415_), .ZN(new_n20416_));
  NOR3_X1    g17296(.A1(new_n20416_), .A2(new_n14452_), .A3(new_n20398_), .ZN(new_n20417_));
  NOR3_X1    g17297(.A1(new_n20399_), .A2(new_n14452_), .A3(new_n20415_), .ZN(new_n20418_));
  OAI21_X1   g17298(.A1(new_n20417_), .A2(new_n20418_), .B(pi0778), .ZN(new_n20419_));
  OAI21_X1   g17299(.A1(pi0778), .A2(new_n20399_), .B(new_n20419_), .ZN(new_n20420_));
  NOR2_X1    g17300(.A1(new_n20404_), .A2(new_n13775_), .ZN(new_n20421_));
  NOR2_X1    g17301(.A1(new_n20415_), .A2(new_n15147_), .ZN(new_n20422_));
  OAI21_X1   g17302(.A1(new_n20420_), .A2(new_n13785_), .B(new_n13766_), .ZN(new_n20423_));
  AOI21_X1   g17303(.A1(new_n20414_), .A2(new_n20423_), .B(new_n13801_), .ZN(new_n20424_));
  OAI21_X1   g17304(.A1(new_n20415_), .A2(new_n15707_), .B(new_n13766_), .ZN(new_n20425_));
  NAND2_X1   g17305(.A1(new_n20421_), .A2(new_n20425_), .ZN(new_n20426_));
  NAND2_X1   g17306(.A1(new_n20426_), .A2(new_n13793_), .ZN(new_n20427_));
  AOI21_X1   g17307(.A1(pi0609), .A2(new_n20420_), .B(new_n20427_), .ZN(new_n20428_));
  NOR2_X1    g17308(.A1(new_n20428_), .A2(pi0609), .ZN(new_n20429_));
  NOR2_X1    g17309(.A1(new_n20429_), .A2(new_n13801_), .ZN(new_n20430_));
  NAND2_X1   g17310(.A1(new_n20414_), .A2(new_n20430_), .ZN(new_n20431_));
  XOR2_X1    g17311(.A1(new_n20424_), .A2(new_n20431_), .Z(new_n20432_));
  OAI21_X1   g17312(.A1(new_n20421_), .A2(new_n20422_), .B(pi0609), .ZN(new_n20433_));
  NAND2_X1   g17313(.A1(new_n20433_), .A2(pi0785), .ZN(new_n20434_));
  NOR2_X1    g17314(.A1(new_n20416_), .A2(new_n13776_), .ZN(new_n20435_));
  AOI21_X1   g17315(.A1(new_n20404_), .A2(new_n13776_), .B(new_n20435_), .ZN(new_n20436_));
  NOR3_X1    g17316(.A1(new_n20426_), .A2(new_n13801_), .A3(new_n20436_), .ZN(new_n20437_));
  NAND2_X1   g17317(.A1(new_n20437_), .A2(new_n20434_), .ZN(new_n20438_));
  OR2_X2     g17318(.A1(new_n20437_), .A2(new_n20434_), .Z(new_n20439_));
  NAND2_X1   g17319(.A1(new_n20439_), .A2(new_n20438_), .ZN(new_n20440_));
  NAND3_X1   g17320(.A1(new_n20440_), .A2(pi0618), .A3(pi1154), .ZN(new_n20441_));
  INV_X1     g17321(.I(new_n20441_), .ZN(new_n20442_));
  NOR3_X1    g17322(.A1(new_n20440_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n20443_));
  OAI21_X1   g17323(.A1(new_n20442_), .A2(new_n20443_), .B(new_n20415_), .ZN(new_n20444_));
  NOR2_X1    g17324(.A1(new_n20416_), .A2(new_n13805_), .ZN(new_n20445_));
  AOI21_X1   g17325(.A1(new_n20420_), .A2(new_n13805_), .B(new_n20445_), .ZN(new_n20446_));
  INV_X1     g17326(.I(new_n20446_), .ZN(new_n20447_));
  AOI21_X1   g17327(.A1(new_n20447_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n20448_));
  AOI21_X1   g17328(.A1(new_n20444_), .A2(new_n20448_), .B(pi0618), .ZN(new_n20449_));
  OAI21_X1   g17329(.A1(new_n20432_), .A2(new_n20449_), .B(pi0781), .ZN(new_n20450_));
  XNOR2_X1   g17330(.A1(new_n20424_), .A2(new_n20431_), .ZN(new_n20451_));
  NAND3_X1   g17331(.A1(new_n20440_), .A2(pi0618), .A3(pi1154), .ZN(new_n20452_));
  NAND4_X1   g17332(.A1(new_n20439_), .A2(new_n13816_), .A3(new_n20438_), .A4(pi1154), .ZN(new_n20453_));
  AOI21_X1   g17333(.A1(new_n20452_), .A2(new_n20453_), .B(new_n20416_), .ZN(new_n20454_));
  INV_X1     g17334(.I(new_n20454_), .ZN(new_n20455_));
  AOI21_X1   g17335(.A1(new_n20447_), .A2(pi0618), .B(new_n13837_), .ZN(new_n20456_));
  AOI21_X1   g17336(.A1(new_n20455_), .A2(new_n20456_), .B(pi0618), .ZN(new_n20457_));
  INV_X1     g17337(.I(new_n20457_), .ZN(new_n20458_));
  NAND3_X1   g17338(.A1(new_n20451_), .A2(pi0781), .A3(new_n20458_), .ZN(new_n20459_));
  XOR2_X1    g17339(.A1(new_n20459_), .A2(new_n20450_), .Z(new_n20460_));
  INV_X1     g17340(.I(new_n20443_), .ZN(new_n20461_));
  AOI21_X1   g17341(.A1(new_n20461_), .A2(new_n20441_), .B(new_n20416_), .ZN(new_n20462_));
  NAND4_X1   g17342(.A1(new_n20462_), .A2(new_n20454_), .A3(pi0781), .A4(new_n20440_), .ZN(new_n20463_));
  NAND3_X1   g17343(.A1(new_n20454_), .A2(pi0781), .A3(new_n20440_), .ZN(new_n20464_));
  NAND3_X1   g17344(.A1(new_n20464_), .A2(pi0781), .A3(new_n20444_), .ZN(new_n20465_));
  NAND2_X1   g17345(.A1(new_n20465_), .A2(new_n20463_), .ZN(new_n20466_));
  NAND3_X1   g17346(.A1(new_n20466_), .A2(pi0619), .A3(pi1159), .ZN(new_n20467_));
  NAND4_X1   g17347(.A1(new_n20465_), .A2(new_n20463_), .A3(pi0619), .A4(new_n13868_), .ZN(new_n20468_));
  AOI21_X1   g17348(.A1(new_n20467_), .A2(new_n20468_), .B(new_n20416_), .ZN(new_n20469_));
  NOR2_X1    g17349(.A1(new_n20415_), .A2(new_n13880_), .ZN(new_n20470_));
  AOI21_X1   g17350(.A1(new_n20446_), .A2(new_n13880_), .B(new_n20470_), .ZN(new_n20471_));
  AOI21_X1   g17351(.A1(new_n20471_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n20472_));
  INV_X1     g17352(.I(new_n20472_), .ZN(new_n20473_));
  OAI21_X1   g17353(.A1(new_n20469_), .A2(new_n20473_), .B(new_n13860_), .ZN(new_n20474_));
  NAND3_X1   g17354(.A1(new_n20466_), .A2(pi0619), .A3(pi1159), .ZN(new_n20475_));
  NAND4_X1   g17355(.A1(new_n20465_), .A2(new_n20463_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n20476_));
  AOI21_X1   g17356(.A1(new_n20475_), .A2(new_n20476_), .B(new_n20416_), .ZN(new_n20477_));
  AOI21_X1   g17357(.A1(new_n20471_), .A2(pi0619), .B(new_n15217_), .ZN(new_n20478_));
  INV_X1     g17358(.I(new_n20478_), .ZN(new_n20479_));
  OAI21_X1   g17359(.A1(new_n20477_), .A2(new_n20479_), .B(new_n13860_), .ZN(new_n20480_));
  NAND4_X1   g17360(.A1(new_n20460_), .A2(new_n20474_), .A3(new_n20480_), .A4(pi0789), .ZN(new_n20481_));
  AOI21_X1   g17361(.A1(new_n20460_), .A2(new_n20474_), .B(new_n13896_), .ZN(new_n20482_));
  NAND3_X1   g17362(.A1(new_n20460_), .A2(new_n20480_), .A3(pi0789), .ZN(new_n20483_));
  NAND2_X1   g17363(.A1(new_n20482_), .A2(new_n20483_), .ZN(new_n20484_));
  NAND2_X1   g17364(.A1(new_n20484_), .A2(new_n20481_), .ZN(new_n20485_));
  NAND4_X1   g17365(.A1(new_n20469_), .A2(new_n20477_), .A3(pi0789), .A4(new_n20466_), .ZN(new_n20486_));
  INV_X1     g17366(.I(new_n20469_), .ZN(new_n20487_));
  NAND3_X1   g17367(.A1(new_n20477_), .A2(pi0789), .A3(new_n20466_), .ZN(new_n20488_));
  NAND3_X1   g17368(.A1(new_n20488_), .A2(pi0789), .A3(new_n20487_), .ZN(new_n20489_));
  NOR2_X1    g17369(.A1(new_n20416_), .A2(new_n13919_), .ZN(new_n20490_));
  AOI21_X1   g17370(.A1(new_n20471_), .A2(new_n13919_), .B(new_n20490_), .ZN(new_n20491_));
  NOR2_X1    g17371(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n20492_));
  INV_X1     g17372(.I(new_n20492_), .ZN(new_n20493_));
  AOI21_X1   g17373(.A1(new_n20489_), .A2(new_n20486_), .B(new_n20493_), .ZN(new_n20494_));
  INV_X1     g17374(.I(new_n20486_), .ZN(new_n20495_));
  INV_X1     g17375(.I(new_n20489_), .ZN(new_n20496_));
  NOR2_X1    g17376(.A1(new_n20496_), .A2(new_n20495_), .ZN(new_n20497_));
  NAND3_X1   g17377(.A1(new_n20485_), .A2(pi0626), .A3(pi0788), .ZN(new_n20502_));
  INV_X1     g17378(.I(new_n20502_), .ZN(new_n20503_));
  INV_X1     g17379(.I(new_n20494_), .ZN(new_n20504_));
  AOI22_X1   g17380(.A1(new_n20504_), .A2(new_n13901_), .B1(new_n20484_), .B2(new_n20481_), .ZN(new_n20505_));
  AOI21_X1   g17381(.A1(new_n20484_), .A2(new_n20481_), .B(new_n15258_), .ZN(new_n20506_));
  NOR3_X1    g17382(.A1(new_n20505_), .A2(new_n13937_), .A3(new_n20506_), .ZN(new_n20507_));
  NOR2_X1    g17383(.A1(new_n20507_), .A2(new_n20503_), .ZN(new_n20508_));
  NOR2_X1    g17384(.A1(new_n20415_), .A2(new_n16372_), .ZN(new_n20509_));
  AOI21_X1   g17385(.A1(new_n20497_), .A2(new_n16372_), .B(new_n20509_), .ZN(new_n20510_));
  NAND2_X1   g17386(.A1(new_n20491_), .A2(new_n13966_), .ZN(new_n20511_));
  OAI21_X1   g17387(.A1(new_n13966_), .A2(new_n20415_), .B(new_n20511_), .ZN(new_n20512_));
  NOR2_X1    g17388(.A1(new_n20512_), .A2(new_n13942_), .ZN(new_n20513_));
  XOR2_X1    g17389(.A1(new_n20513_), .A2(new_n13970_), .Z(new_n20514_));
  NAND2_X1   g17390(.A1(new_n20514_), .A2(new_n20415_), .ZN(new_n20515_));
  NAND2_X1   g17391(.A1(new_n20515_), .A2(new_n13977_), .ZN(new_n20516_));
  AOI21_X1   g17392(.A1(new_n20510_), .A2(new_n13942_), .B(new_n20516_), .ZN(new_n20517_));
  NOR2_X1    g17393(.A1(new_n20512_), .A2(new_n13969_), .ZN(new_n20518_));
  XOR2_X1    g17394(.A1(new_n20518_), .A2(new_n13970_), .Z(new_n20519_));
  NAND2_X1   g17395(.A1(new_n20519_), .A2(new_n20415_), .ZN(new_n20520_));
  NOR3_X1    g17396(.A1(new_n20508_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n20523_));
  INV_X1     g17397(.I(new_n20481_), .ZN(new_n20524_));
  AND2_X2    g17398(.A1(new_n20482_), .A2(new_n20483_), .Z(new_n20525_));
  OAI22_X1   g17399(.A1(new_n20525_), .A2(new_n20524_), .B1(pi0626), .B2(new_n20494_), .ZN(new_n20526_));
  NAND2_X1   g17400(.A1(new_n20485_), .A2(new_n14577_), .ZN(new_n20527_));
  NAND3_X1   g17401(.A1(new_n20526_), .A2(new_n20527_), .A3(pi0788), .ZN(new_n20528_));
  NAND3_X1   g17402(.A1(new_n20489_), .A2(new_n16372_), .A3(new_n20486_), .ZN(new_n20529_));
  OAI21_X1   g17403(.A1(new_n16372_), .A2(new_n20415_), .B(new_n20529_), .ZN(new_n20530_));
  INV_X1     g17404(.I(new_n20516_), .ZN(new_n20531_));
  AOI21_X1   g17405(.A1(new_n20530_), .A2(new_n20531_), .B(pi0628), .ZN(new_n20532_));
  AOI21_X1   g17406(.A1(new_n20528_), .A2(new_n20502_), .B(new_n20532_), .ZN(new_n20533_));
  AOI21_X1   g17407(.A1(new_n20528_), .A2(new_n20502_), .B(new_n15296_), .ZN(new_n20534_));
  NOR3_X1    g17408(.A1(new_n20533_), .A2(new_n20534_), .A3(new_n12777_), .ZN(new_n20535_));
  NOR2_X1    g17409(.A1(new_n20535_), .A2(new_n20523_), .ZN(new_n20536_));
  NOR2_X1    g17410(.A1(new_n20415_), .A2(new_n13994_), .ZN(new_n20537_));
  AOI21_X1   g17411(.A1(new_n20530_), .A2(new_n13994_), .B(new_n20537_), .ZN(new_n20538_));
  INV_X1     g17412(.I(new_n20538_), .ZN(new_n20539_));
  NAND2_X1   g17413(.A1(new_n20515_), .A2(pi0792), .ZN(new_n20540_));
  INV_X1     g17414(.I(new_n20512_), .ZN(new_n20541_));
  NOR3_X1    g17415(.A1(new_n20520_), .A2(new_n12777_), .A3(new_n20541_), .ZN(new_n20542_));
  XOR2_X1    g17416(.A1(new_n20542_), .A2(new_n20540_), .Z(new_n20543_));
  NAND2_X1   g17417(.A1(new_n20543_), .A2(pi0647), .ZN(new_n20544_));
  XOR2_X1    g17418(.A1(new_n20544_), .A2(new_n14008_), .Z(new_n20545_));
  AOI21_X1   g17419(.A1(new_n20545_), .A2(new_n20415_), .B(new_n14012_), .ZN(new_n20546_));
  AOI21_X1   g17420(.A1(new_n20539_), .A2(new_n20546_), .B(pi0647), .ZN(new_n20547_));
  AOI21_X1   g17421(.A1(new_n20543_), .A2(pi1157), .B(new_n14008_), .ZN(new_n20548_));
  NAND2_X1   g17422(.A1(new_n20543_), .A2(pi1157), .ZN(new_n20549_));
  NOR2_X1    g17423(.A1(new_n20549_), .A2(new_n14007_), .ZN(new_n20550_));
  OAI21_X1   g17424(.A1(new_n20550_), .A2(new_n20548_), .B(new_n20415_), .ZN(new_n20551_));
  NAND2_X1   g17425(.A1(new_n20551_), .A2(new_n14027_), .ZN(new_n20552_));
  AOI21_X1   g17426(.A1(new_n20538_), .A2(pi0647), .B(new_n20552_), .ZN(new_n20553_));
  NOR2_X1    g17427(.A1(new_n20553_), .A2(pi0647), .ZN(new_n20554_));
  NOR4_X1    g17428(.A1(new_n20536_), .A2(new_n12776_), .A3(new_n20547_), .A4(new_n20554_), .ZN(new_n20555_));
  NAND2_X1   g17429(.A1(new_n20528_), .A2(new_n20502_), .ZN(new_n20556_));
  NAND3_X1   g17430(.A1(new_n20556_), .A2(pi0628), .A3(pi0792), .ZN(new_n20557_));
  OAI22_X1   g17431(.A1(new_n20507_), .A2(new_n20503_), .B1(pi0628), .B2(new_n20517_), .ZN(new_n20558_));
  OAI21_X1   g17432(.A1(new_n20507_), .A2(new_n20503_), .B(new_n14606_), .ZN(new_n20559_));
  NAND3_X1   g17433(.A1(new_n20558_), .A2(new_n20559_), .A3(pi0792), .ZN(new_n20560_));
  AOI21_X1   g17434(.A1(new_n20560_), .A2(new_n20557_), .B(new_n20547_), .ZN(new_n20561_));
  OAI21_X1   g17435(.A1(new_n20553_), .A2(pi0647), .B(pi0787), .ZN(new_n20562_));
  AOI21_X1   g17436(.A1(new_n20560_), .A2(new_n20557_), .B(new_n20562_), .ZN(new_n20563_));
  NOR3_X1    g17437(.A1(new_n20561_), .A2(new_n20563_), .A3(new_n12776_), .ZN(new_n20564_));
  OAI21_X1   g17438(.A1(new_n20564_), .A2(new_n20555_), .B(new_n12775_), .ZN(new_n20565_));
  NOR2_X1    g17439(.A1(new_n9992_), .A2(pi0179), .ZN(new_n20566_));
  AOI21_X1   g17440(.A1(new_n13218_), .A2(new_n17474_), .B(new_n20566_), .ZN(new_n20567_));
  INV_X1     g17441(.I(new_n20567_), .ZN(new_n20568_));
  NOR3_X1    g17442(.A1(new_n13219_), .A2(pi0625), .A3(pi0724), .ZN(new_n20569_));
  NAND3_X1   g17443(.A1(new_n20568_), .A2(new_n20569_), .A3(new_n20566_), .ZN(new_n20570_));
  NOR3_X1    g17444(.A1(new_n20569_), .A2(new_n13614_), .A3(new_n20567_), .ZN(new_n20571_));
  XOR2_X1    g17445(.A1(new_n20570_), .A2(new_n20571_), .Z(new_n20572_));
  NAND2_X1   g17446(.A1(new_n20568_), .A2(new_n13748_), .ZN(new_n20573_));
  OAI21_X1   g17447(.A1(new_n20572_), .A2(new_n13748_), .B(new_n20573_), .ZN(new_n20574_));
  NAND2_X1   g17448(.A1(new_n20574_), .A2(new_n14049_), .ZN(new_n20575_));
  NOR2_X1    g17449(.A1(new_n20575_), .A2(new_n14051_), .ZN(new_n20576_));
  INV_X1     g17450(.I(new_n20576_), .ZN(new_n20577_));
  NOR2_X1    g17451(.A1(new_n20577_), .A2(new_n14163_), .ZN(new_n20578_));
  AOI21_X1   g17452(.A1(new_n13104_), .A2(new_n17475_), .B(new_n20566_), .ZN(new_n20579_));
  NOR2_X1    g17453(.A1(new_n14096_), .A2(new_n20579_), .ZN(new_n20580_));
  AOI21_X1   g17454(.A1(new_n20580_), .A2(new_n14094_), .B(pi1155), .ZN(new_n20581_));
  NOR2_X1    g17455(.A1(new_n20581_), .A2(new_n13801_), .ZN(new_n20582_));
  NAND2_X1   g17456(.A1(new_n20579_), .A2(pi1155), .ZN(new_n20583_));
  AOI21_X1   g17457(.A1(new_n20583_), .A2(new_n2723_), .B(new_n14102_), .ZN(new_n20584_));
  NAND3_X1   g17458(.A1(new_n20584_), .A2(pi0785), .A3(new_n20580_), .ZN(new_n20585_));
  XOR2_X1    g17459(.A1(new_n20582_), .A2(new_n20585_), .Z(new_n20586_));
  NOR2_X1    g17460(.A1(new_n20586_), .A2(new_n13817_), .ZN(new_n20587_));
  OAI21_X1   g17461(.A1(new_n20587_), .A2(pi0618), .B(new_n9992_), .ZN(new_n20588_));
  NAND2_X1   g17462(.A1(new_n20588_), .A2(pi0781), .ZN(new_n20589_));
  OAI21_X1   g17463(.A1(new_n20587_), .A2(new_n9992_), .B(pi0618), .ZN(new_n20590_));
  NOR3_X1    g17464(.A1(new_n20590_), .A2(new_n13855_), .A3(new_n20586_), .ZN(new_n20591_));
  XOR2_X1    g17465(.A1(new_n20591_), .A2(new_n20589_), .Z(new_n20592_));
  NAND2_X1   g17466(.A1(new_n20592_), .A2(pi0619), .ZN(new_n20593_));
  XOR2_X1    g17467(.A1(new_n20593_), .A2(new_n13904_), .Z(new_n20594_));
  NAND2_X1   g17468(.A1(new_n20594_), .A2(new_n20566_), .ZN(new_n20595_));
  NAND2_X1   g17469(.A1(new_n20595_), .A2(pi0789), .ZN(new_n20596_));
  NAND2_X1   g17470(.A1(new_n20592_), .A2(pi1159), .ZN(new_n20597_));
  XOR2_X1    g17471(.A1(new_n20597_), .A2(new_n13904_), .Z(new_n20598_));
  NAND2_X1   g17472(.A1(new_n20598_), .A2(new_n20566_), .ZN(new_n20599_));
  NOR3_X1    g17473(.A1(new_n20599_), .A2(new_n13896_), .A3(new_n20592_), .ZN(new_n20600_));
  XOR2_X1    g17474(.A1(new_n20600_), .A2(new_n20596_), .Z(new_n20601_));
  NAND2_X1   g17475(.A1(new_n20601_), .A2(new_n13962_), .ZN(new_n20602_));
  XOR2_X1    g17476(.A1(new_n20602_), .A2(new_n18976_), .Z(new_n20603_));
  AOI22_X1   g17477(.A1(new_n20603_), .A2(new_n20566_), .B1(new_n16639_), .B2(new_n20578_), .ZN(new_n20604_));
  NOR3_X1    g17478(.A1(new_n20567_), .A2(new_n13613_), .A3(new_n13203_), .ZN(new_n20605_));
  INV_X1     g17479(.I(new_n20579_), .ZN(new_n20606_));
  NOR2_X1    g17480(.A1(new_n20566_), .A2(pi1153), .ZN(new_n20607_));
  INV_X1     g17481(.I(new_n20607_), .ZN(new_n20608_));
  OAI21_X1   g17482(.A1(new_n20569_), .A2(new_n20608_), .B(pi0608), .ZN(new_n20609_));
  NAND3_X1   g17483(.A1(new_n20609_), .A2(new_n13614_), .A3(new_n20606_), .ZN(new_n20610_));
  AOI21_X1   g17484(.A1(new_n20610_), .A2(new_n20605_), .B(new_n13748_), .ZN(new_n20611_));
  NOR2_X1    g17485(.A1(new_n20567_), .A2(new_n13203_), .ZN(new_n20612_));
  NAND2_X1   g17486(.A1(new_n20569_), .A2(new_n20607_), .ZN(new_n20613_));
  AOI21_X1   g17487(.A1(new_n14083_), .A2(new_n20568_), .B(new_n20613_), .ZN(new_n20614_));
  NOR2_X1    g17488(.A1(new_n20614_), .A2(new_n20605_), .ZN(new_n20615_));
  NOR4_X1    g17489(.A1(new_n20615_), .A2(new_n13748_), .A3(new_n20606_), .A4(new_n20612_), .ZN(new_n20616_));
  XOR2_X1    g17490(.A1(new_n20616_), .A2(new_n20611_), .Z(new_n20617_));
  NAND2_X1   g17491(.A1(new_n20617_), .A2(new_n13801_), .ZN(new_n20618_));
  NOR2_X1    g17492(.A1(new_n20617_), .A2(new_n13778_), .ZN(new_n20619_));
  XOR2_X1    g17493(.A1(new_n20619_), .A2(new_n14090_), .Z(new_n20620_));
  NAND2_X1   g17494(.A1(new_n20620_), .A2(new_n20574_), .ZN(new_n20621_));
  NOR2_X1    g17495(.A1(new_n20581_), .A2(new_n13783_), .ZN(new_n20622_));
  NAND2_X1   g17496(.A1(new_n20621_), .A2(new_n20622_), .ZN(new_n20623_));
  NOR2_X1    g17497(.A1(new_n20584_), .A2(pi0660), .ZN(new_n20624_));
  NAND2_X1   g17498(.A1(new_n20623_), .A2(new_n20624_), .ZN(new_n20625_));
  NOR2_X1    g17499(.A1(new_n20617_), .A2(new_n13766_), .ZN(new_n20626_));
  XOR2_X1    g17500(.A1(new_n20626_), .A2(new_n14090_), .Z(new_n20627_));
  NAND4_X1   g17501(.A1(new_n20625_), .A2(pi0785), .A3(new_n20574_), .A4(new_n20627_), .ZN(new_n20628_));
  NAND2_X1   g17502(.A1(new_n20628_), .A2(new_n20618_), .ZN(new_n20629_));
  NAND2_X1   g17503(.A1(new_n20629_), .A2(new_n13855_), .ZN(new_n20630_));
  NOR2_X1    g17504(.A1(new_n20629_), .A2(new_n13816_), .ZN(new_n20631_));
  XOR2_X1    g17505(.A1(new_n20631_), .A2(new_n13818_), .Z(new_n20632_));
  NAND3_X1   g17506(.A1(new_n20632_), .A2(new_n14049_), .A3(new_n20574_), .ZN(new_n20633_));
  NAND3_X1   g17507(.A1(new_n20633_), .A2(new_n13823_), .A3(new_n20590_), .ZN(new_n20634_));
  AND3_X2    g17508(.A1(new_n20634_), .A2(new_n13823_), .A3(new_n20588_), .Z(new_n20635_));
  NOR2_X1    g17509(.A1(new_n20629_), .A2(new_n13817_), .ZN(new_n20636_));
  XOR2_X1    g17510(.A1(new_n20636_), .A2(new_n13819_), .Z(new_n20637_));
  NOR3_X1    g17511(.A1(new_n20637_), .A2(new_n13855_), .A3(new_n20575_), .ZN(new_n20638_));
  INV_X1     g17512(.I(new_n20638_), .ZN(new_n20639_));
  OAI21_X1   g17513(.A1(new_n20635_), .A2(new_n20639_), .B(new_n20630_), .ZN(new_n20640_));
  NOR2_X1    g17514(.A1(new_n20640_), .A2(new_n13860_), .ZN(new_n20641_));
  XOR2_X1    g17515(.A1(new_n20641_), .A2(new_n13904_), .Z(new_n20642_));
  NOR2_X1    g17516(.A1(new_n20642_), .A2(new_n20577_), .ZN(new_n20643_));
  NAND2_X1   g17517(.A1(new_n20599_), .A2(new_n13884_), .ZN(new_n20644_));
  INV_X1     g17518(.I(new_n20640_), .ZN(new_n20645_));
  AOI21_X1   g17519(.A1(new_n20645_), .A2(new_n14143_), .B(pi0789), .ZN(new_n20646_));
  OAI21_X1   g17520(.A1(new_n20643_), .A2(new_n20644_), .B(new_n20646_), .ZN(new_n20647_));
  NOR2_X1    g17521(.A1(new_n20640_), .A2(new_n13868_), .ZN(new_n20648_));
  XOR2_X1    g17522(.A1(new_n20648_), .A2(new_n13903_), .Z(new_n20649_));
  NAND2_X1   g17523(.A1(new_n20595_), .A2(new_n19018_), .ZN(new_n20650_));
  AOI21_X1   g17524(.A1(new_n20649_), .A2(new_n20576_), .B(new_n20650_), .ZN(new_n20651_));
  AOI21_X1   g17525(.A1(new_n20647_), .A2(new_n20651_), .B(new_n20604_), .ZN(new_n20652_));
  NAND2_X1   g17526(.A1(new_n20601_), .A2(new_n16372_), .ZN(new_n20653_));
  OAI21_X1   g17527(.A1(new_n16372_), .A2(new_n20566_), .B(new_n20653_), .ZN(new_n20654_));
  NAND3_X1   g17528(.A1(new_n20654_), .A2(new_n18929_), .A3(new_n20578_), .ZN(new_n20655_));
  NAND2_X1   g17529(.A1(new_n20655_), .A2(new_n16569_), .ZN(new_n20656_));
  XOR2_X1    g17530(.A1(new_n20656_), .A2(new_n16572_), .Z(new_n20657_));
  AOI21_X1   g17531(.A1(new_n19022_), .A2(new_n20655_), .B(new_n20657_), .ZN(new_n20658_));
  INV_X1     g17532(.I(new_n20566_), .ZN(new_n20659_));
  NAND2_X1   g17533(.A1(new_n20601_), .A2(new_n13963_), .ZN(new_n20660_));
  XNOR2_X1   g17534(.A1(new_n20660_), .A2(new_n19028_), .ZN(new_n20661_));
  NOR3_X1    g17535(.A1(new_n20661_), .A2(new_n16424_), .A3(new_n20659_), .ZN(new_n20662_));
  OAI21_X1   g17536(.A1(new_n20658_), .A2(new_n16574_), .B(new_n20662_), .ZN(new_n20663_));
  NOR4_X1    g17537(.A1(new_n20577_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n20664_));
  NOR2_X1    g17538(.A1(new_n20664_), .A2(new_n14005_), .ZN(new_n20665_));
  XOR2_X1    g17539(.A1(new_n20665_), .A2(new_n14007_), .Z(new_n20666_));
  NAND2_X1   g17540(.A1(new_n20666_), .A2(new_n20566_), .ZN(new_n20667_));
  NOR2_X1    g17541(.A1(new_n20659_), .A2(pi0647), .ZN(new_n20668_));
  AOI21_X1   g17542(.A1(new_n20664_), .A2(pi0647), .B(new_n20668_), .ZN(new_n20669_));
  NOR2_X1    g17543(.A1(new_n20654_), .A2(new_n13994_), .ZN(new_n20670_));
  XNOR2_X1   g17544(.A1(new_n20670_), .A2(new_n19033_), .ZN(new_n20671_));
  AOI22_X1   g17545(.A1(new_n20671_), .A2(new_n20566_), .B1(new_n14206_), .B2(new_n20669_), .ZN(new_n20672_));
  NOR3_X1    g17546(.A1(new_n20672_), .A2(new_n14010_), .A3(new_n20667_), .ZN(new_n20673_));
  OAI22_X1   g17547(.A1(new_n20652_), .A2(new_n20663_), .B1(new_n12776_), .B2(new_n20673_), .ZN(new_n20674_));
  AOI21_X1   g17548(.A1(new_n20669_), .A2(pi1157), .B(new_n12776_), .ZN(new_n20675_));
  AOI22_X1   g17549(.A1(new_n20667_), .A2(new_n20675_), .B1(new_n12776_), .B2(new_n20664_), .ZN(new_n20676_));
  NAND2_X1   g17550(.A1(new_n20674_), .A2(pi0644), .ZN(new_n20677_));
  XOR2_X1    g17551(.A1(new_n20677_), .A2(new_n14205_), .Z(new_n20678_));
  NOR2_X1    g17552(.A1(new_n20678_), .A2(new_n20676_), .ZN(new_n20679_));
  NOR2_X1    g17553(.A1(new_n20654_), .A2(new_n18968_), .ZN(new_n20680_));
  NAND2_X1   g17554(.A1(new_n18967_), .A2(new_n20566_), .ZN(new_n20681_));
  XOR2_X1    g17555(.A1(new_n20680_), .A2(new_n20681_), .Z(new_n20682_));
  NAND2_X1   g17556(.A1(new_n20682_), .A2(pi0715), .ZN(new_n20683_));
  XOR2_X1    g17557(.A1(new_n20683_), .A2(new_n14205_), .Z(new_n20684_));
  OAI21_X1   g17558(.A1(new_n20684_), .A2(new_n20659_), .B(new_n14203_), .ZN(new_n20685_));
  NAND2_X1   g17559(.A1(new_n20682_), .A2(pi0644), .ZN(new_n20686_));
  XOR2_X1    g17560(.A1(new_n20686_), .A2(new_n14217_), .Z(new_n20687_));
  AOI21_X1   g17561(.A1(new_n20687_), .A2(new_n20566_), .B(pi1160), .ZN(new_n20688_));
  OAI21_X1   g17562(.A1(new_n20679_), .A2(new_n20685_), .B(new_n20688_), .ZN(new_n20689_));
  NAND2_X1   g17563(.A1(new_n20674_), .A2(pi0715), .ZN(new_n20690_));
  XOR2_X1    g17564(.A1(new_n20690_), .A2(new_n14205_), .Z(new_n20691_));
  NOR2_X1    g17565(.A1(new_n20691_), .A2(new_n20676_), .ZN(new_n20692_));
  AOI21_X1   g17566(.A1(new_n20689_), .A2(new_n20692_), .B(new_n14799_), .ZN(new_n20693_));
  XOR2_X1    g17567(.A1(new_n20693_), .A2(new_n14801_), .Z(new_n20694_));
  NOR2_X1    g17568(.A1(new_n7240_), .A2(pi0179), .ZN(new_n20695_));
  NOR4_X1    g17569(.A1(new_n20694_), .A2(pi0832), .A3(new_n20674_), .A4(new_n20695_), .ZN(new_n20696_));
  AOI21_X1   g17570(.A1(new_n20565_), .A2(new_n7240_), .B(new_n20696_), .ZN(new_n20697_));
  NOR3_X1    g17571(.A1(new_n20564_), .A2(new_n20555_), .A3(new_n14200_), .ZN(new_n20698_));
  NOR2_X1    g17572(.A1(new_n20698_), .A2(new_n14217_), .ZN(new_n20699_));
  NOR4_X1    g17573(.A1(new_n20564_), .A2(new_n20555_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n20700_));
  NOR2_X1    g17574(.A1(new_n20699_), .A2(new_n20700_), .ZN(new_n20701_));
  OAI21_X1   g17575(.A1(new_n12776_), .A2(new_n20561_), .B(new_n20563_), .ZN(new_n20702_));
  OR3_X2     g17576(.A1(new_n20561_), .A2(new_n20563_), .A3(new_n12776_), .Z(new_n20703_));
  NOR2_X1    g17577(.A1(new_n20416_), .A2(new_n14211_), .ZN(new_n20704_));
  AOI21_X1   g17578(.A1(new_n20538_), .A2(new_n14211_), .B(new_n20704_), .ZN(new_n20705_));
  OAI21_X1   g17579(.A1(new_n20416_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n20706_));
  NAND2_X1   g17580(.A1(new_n20705_), .A2(new_n20706_), .ZN(new_n20707_));
  NAND2_X1   g17581(.A1(new_n20545_), .A2(new_n20415_), .ZN(new_n20708_));
  NOR4_X1    g17582(.A1(new_n20708_), .A2(new_n12776_), .A3(new_n20543_), .A4(new_n20551_), .ZN(new_n20709_));
  NAND2_X1   g17583(.A1(new_n20708_), .A2(pi0787), .ZN(new_n20710_));
  NOR3_X1    g17584(.A1(new_n20551_), .A2(new_n12776_), .A3(new_n20543_), .ZN(new_n20711_));
  NOR2_X1    g17585(.A1(new_n20710_), .A2(new_n20711_), .ZN(new_n20712_));
  AOI21_X1   g17586(.A1(new_n20707_), .A2(new_n14815_), .B(pi0644), .ZN(new_n20713_));
  AOI21_X1   g17587(.A1(new_n20703_), .A2(new_n20702_), .B(new_n20713_), .ZN(new_n20714_));
  OAI21_X1   g17588(.A1(new_n20415_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n20715_));
  OAI21_X1   g17589(.A1(new_n20712_), .A2(new_n20709_), .B(new_n20715_), .ZN(new_n20716_));
  NOR2_X1    g17590(.A1(new_n20716_), .A2(new_n20705_), .ZN(new_n20717_));
  OAI21_X1   g17591(.A1(new_n20714_), .A2(pi0790), .B(new_n20717_), .ZN(new_n20718_));
  NOR3_X1    g17592(.A1(new_n20701_), .A2(new_n20718_), .A3(new_n20697_), .ZN(po0336));
  NOR2_X1    g17593(.A1(new_n14428_), .A2(pi0180), .ZN(new_n20720_));
  INV_X1     g17594(.I(new_n20720_), .ZN(new_n20721_));
  NAND2_X1   g17595(.A1(new_n20721_), .A2(new_n13965_), .ZN(new_n20722_));
  NOR2_X1    g17596(.A1(new_n20721_), .A2(new_n13919_), .ZN(new_n20723_));
  INV_X1     g17597(.I(pi0702), .ZN(new_n20724_));
  OAI21_X1   g17598(.A1(new_n13721_), .A2(new_n20724_), .B(new_n5642_), .ZN(new_n20725_));
  NAND2_X1   g17599(.A1(new_n16715_), .A2(new_n5642_), .ZN(new_n20726_));
  NAND4_X1   g17600(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n20725_), .A4(new_n20726_), .ZN(new_n20727_));
  AOI21_X1   g17601(.A1(new_n20727_), .A2(new_n14424_), .B(new_n5642_), .ZN(new_n20728_));
  NAND2_X1   g17602(.A1(new_n20720_), .A2(new_n20728_), .ZN(new_n20729_));
  NAND2_X1   g17603(.A1(new_n20729_), .A2(new_n3290_), .ZN(new_n20730_));
  NAND2_X1   g17604(.A1(new_n20730_), .A2(pi0702), .ZN(new_n20731_));
  NAND2_X1   g17605(.A1(new_n20731_), .A2(pi0625), .ZN(new_n20732_));
  XOR2_X1    g17606(.A1(new_n20732_), .A2(new_n13620_), .Z(new_n20733_));
  NAND2_X1   g17607(.A1(new_n20733_), .A2(new_n20720_), .ZN(new_n20734_));
  NAND2_X1   g17608(.A1(new_n20734_), .A2(pi0778), .ZN(new_n20735_));
  NAND2_X1   g17609(.A1(new_n20731_), .A2(pi1153), .ZN(new_n20736_));
  XOR2_X1    g17610(.A1(new_n20736_), .A2(new_n13620_), .Z(new_n20737_));
  NAND2_X1   g17611(.A1(new_n20737_), .A2(new_n20720_), .ZN(new_n20738_));
  NOR3_X1    g17612(.A1(new_n20738_), .A2(new_n13748_), .A3(new_n20731_), .ZN(new_n20739_));
  XNOR2_X1   g17613(.A1(new_n20739_), .A2(new_n20735_), .ZN(new_n20740_));
  INV_X1     g17614(.I(new_n20740_), .ZN(new_n20741_));
  NAND2_X1   g17615(.A1(new_n20720_), .A2(new_n13803_), .ZN(new_n20742_));
  OAI21_X1   g17616(.A1(new_n20741_), .A2(new_n13803_), .B(new_n20742_), .ZN(new_n20743_));
  NOR2_X1    g17617(.A1(new_n20743_), .A2(new_n13879_), .ZN(new_n20744_));
  AOI21_X1   g17618(.A1(new_n13879_), .A2(new_n20721_), .B(new_n20744_), .ZN(new_n20745_));
  AOI21_X1   g17619(.A1(new_n20745_), .A2(new_n13919_), .B(new_n20723_), .ZN(new_n20746_));
  NAND2_X1   g17620(.A1(new_n20746_), .A2(new_n13966_), .ZN(new_n20747_));
  NAND2_X1   g17621(.A1(new_n20747_), .A2(new_n20722_), .ZN(new_n20748_));
  INV_X1     g17622(.I(new_n20748_), .ZN(new_n20749_));
  AOI21_X1   g17623(.A1(new_n20749_), .A2(pi0628), .B(new_n13971_), .ZN(new_n20750_));
  NOR3_X1    g17624(.A1(new_n20748_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n20751_));
  OAI21_X1   g17625(.A1(new_n20750_), .A2(new_n20751_), .B(new_n20720_), .ZN(new_n20752_));
  NAND2_X1   g17626(.A1(new_n20752_), .A2(pi0792), .ZN(new_n20753_));
  NAND3_X1   g17627(.A1(new_n20748_), .A2(pi0628), .A3(pi1156), .ZN(new_n20754_));
  INV_X1     g17628(.I(new_n20754_), .ZN(new_n20755_));
  NOR3_X1    g17629(.A1(new_n20748_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n20756_));
  NOR2_X1    g17630(.A1(new_n20755_), .A2(new_n20756_), .ZN(new_n20757_));
  NOR4_X1    g17631(.A1(new_n20757_), .A2(new_n12777_), .A3(new_n20721_), .A4(new_n20749_), .ZN(new_n20758_));
  NAND2_X1   g17632(.A1(new_n20758_), .A2(new_n20753_), .ZN(new_n20759_));
  NOR2_X1    g17633(.A1(new_n20758_), .A2(new_n20753_), .ZN(new_n20760_));
  INV_X1     g17634(.I(new_n20760_), .ZN(new_n20761_));
  AOI21_X1   g17635(.A1(new_n20761_), .A2(new_n20759_), .B(new_n14005_), .ZN(new_n20762_));
  NOR2_X1    g17636(.A1(new_n20721_), .A2(pi0647), .ZN(new_n20763_));
  NOR2_X1    g17637(.A1(new_n20763_), .A2(new_n14006_), .ZN(new_n20764_));
  INV_X1     g17638(.I(new_n20764_), .ZN(new_n20765_));
  NOR2_X1    g17639(.A1(new_n20762_), .A2(new_n20765_), .ZN(new_n20766_));
  AOI21_X1   g17640(.A1(new_n20761_), .A2(new_n20759_), .B(pi0647), .ZN(new_n20767_));
  NOR2_X1    g17641(.A1(new_n20721_), .A2(new_n14005_), .ZN(new_n20768_));
  NOR3_X1    g17642(.A1(new_n20767_), .A2(pi1157), .A3(new_n20768_), .ZN(new_n20769_));
  OAI21_X1   g17643(.A1(new_n20769_), .A2(new_n20766_), .B(pi0787), .ZN(new_n20770_));
  NAND3_X1   g17644(.A1(new_n20749_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n20771_));
  AOI21_X1   g17645(.A1(new_n20771_), .A2(new_n20754_), .B(new_n20721_), .ZN(new_n20772_));
  NAND3_X1   g17646(.A1(new_n20772_), .A2(pi0792), .A3(new_n20748_), .ZN(new_n20773_));
  AOI21_X1   g17647(.A1(pi0792), .A2(new_n20752_), .B(new_n20773_), .ZN(new_n20774_));
  NOR3_X1    g17648(.A1(new_n20774_), .A2(pi0787), .A3(new_n20760_), .ZN(new_n20775_));
  INV_X1     g17649(.I(new_n20775_), .ZN(new_n20776_));
  NAND2_X1   g17650(.A1(new_n20721_), .A2(new_n14142_), .ZN(new_n20777_));
  NOR2_X1    g17651(.A1(new_n5642_), .A2(new_n17532_), .ZN(new_n20778_));
  INV_X1     g17652(.I(new_n20778_), .ZN(new_n20779_));
  NAND2_X1   g17653(.A1(new_n14366_), .A2(new_n14389_), .ZN(new_n20780_));
  NAND2_X1   g17654(.A1(new_n20780_), .A2(new_n20779_), .ZN(new_n20781_));
  OAI21_X1   g17655(.A1(new_n14298_), .A2(new_n5642_), .B(new_n3183_), .ZN(new_n20782_));
  AOI21_X1   g17656(.A1(new_n13194_), .A2(pi0753), .B(new_n20782_), .ZN(new_n20783_));
  OAI21_X1   g17657(.A1(new_n20783_), .A2(new_n17532_), .B(pi0180), .ZN(new_n20784_));
  NAND2_X1   g17658(.A1(new_n19327_), .A2(pi0038), .ZN(new_n20785_));
  OAI21_X1   g17659(.A1(new_n20785_), .A2(new_n20784_), .B(new_n3183_), .ZN(new_n20786_));
  AOI21_X1   g17660(.A1(new_n13109_), .A2(new_n5642_), .B(new_n3259_), .ZN(new_n20787_));
  AND3_X2    g17661(.A1(new_n20781_), .A2(new_n20786_), .A3(new_n20787_), .Z(new_n20788_));
  OAI21_X1   g17662(.A1(new_n20788_), .A2(new_n13106_), .B(pi0753), .ZN(new_n20789_));
  INV_X1     g17663(.I(new_n20789_), .ZN(new_n20790_));
  NOR2_X1    g17664(.A1(new_n3289_), .A2(pi0180), .ZN(new_n20791_));
  AOI21_X1   g17665(.A1(new_n20790_), .A2(new_n3289_), .B(new_n20791_), .ZN(new_n20792_));
  NAND2_X1   g17666(.A1(new_n20792_), .A2(new_n13776_), .ZN(new_n20793_));
  NAND2_X1   g17667(.A1(new_n20721_), .A2(new_n13780_), .ZN(new_n20794_));
  NAND2_X1   g17668(.A1(new_n20793_), .A2(new_n20794_), .ZN(new_n20795_));
  NAND2_X1   g17669(.A1(new_n20795_), .A2(pi0609), .ZN(new_n20796_));
  NAND2_X1   g17670(.A1(new_n20796_), .A2(pi0785), .ZN(new_n20797_));
  NAND2_X1   g17671(.A1(new_n20720_), .A2(new_n13775_), .ZN(new_n20798_));
  OAI21_X1   g17672(.A1(new_n20792_), .A2(new_n13775_), .B(new_n20798_), .ZN(new_n20799_));
  AOI21_X1   g17673(.A1(new_n20721_), .A2(new_n14467_), .B(pi0609), .ZN(new_n20800_));
  NOR2_X1    g17674(.A1(new_n20793_), .A2(new_n20800_), .ZN(new_n20801_));
  NAND3_X1   g17675(.A1(new_n20801_), .A2(pi0785), .A3(new_n20799_), .ZN(new_n20802_));
  XNOR2_X1   g17676(.A1(new_n20797_), .A2(new_n20802_), .ZN(new_n20803_));
  INV_X1     g17677(.I(new_n20803_), .ZN(new_n20804_));
  NAND3_X1   g17678(.A1(new_n20804_), .A2(pi0618), .A3(pi1154), .ZN(new_n20805_));
  NAND3_X1   g17679(.A1(new_n20803_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n20806_));
  AOI21_X1   g17680(.A1(new_n20805_), .A2(new_n20806_), .B(new_n20721_), .ZN(new_n20807_));
  NAND3_X1   g17681(.A1(new_n20804_), .A2(pi0618), .A3(pi1154), .ZN(new_n20808_));
  NAND3_X1   g17682(.A1(new_n20803_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n20809_));
  AOI21_X1   g17683(.A1(new_n20808_), .A2(new_n20809_), .B(new_n20721_), .ZN(new_n20810_));
  NAND4_X1   g17684(.A1(new_n20807_), .A2(new_n20810_), .A3(pi0781), .A4(new_n20804_), .ZN(new_n20811_));
  NOR2_X1    g17685(.A1(new_n20807_), .A2(new_n13855_), .ZN(new_n20812_));
  INV_X1     g17686(.I(new_n20810_), .ZN(new_n20813_));
  NAND2_X1   g17687(.A1(new_n20804_), .A2(pi0781), .ZN(new_n20814_));
  OAI21_X1   g17688(.A1(new_n20813_), .A2(new_n20814_), .B(new_n20812_), .ZN(new_n20815_));
  NAND2_X1   g17689(.A1(new_n20815_), .A2(new_n20811_), .ZN(new_n20816_));
  NAND3_X1   g17690(.A1(new_n20816_), .A2(pi0619), .A3(pi1159), .ZN(new_n20817_));
  INV_X1     g17691(.I(new_n20816_), .ZN(new_n20818_));
  NAND3_X1   g17692(.A1(new_n20818_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n20819_));
  AOI21_X1   g17693(.A1(new_n20819_), .A2(new_n20817_), .B(new_n20721_), .ZN(new_n20820_));
  NOR2_X1    g17694(.A1(new_n20820_), .A2(new_n13896_), .ZN(new_n20821_));
  INV_X1     g17695(.I(new_n20821_), .ZN(new_n20822_));
  NOR2_X1    g17696(.A1(new_n20816_), .A2(new_n13868_), .ZN(new_n20823_));
  XOR2_X1    g17697(.A1(new_n20823_), .A2(new_n13903_), .Z(new_n20824_));
  NOR2_X1    g17698(.A1(new_n20818_), .A2(new_n13896_), .ZN(new_n20825_));
  NAND4_X1   g17699(.A1(new_n20822_), .A2(new_n20720_), .A3(new_n20824_), .A4(new_n20825_), .ZN(new_n20826_));
  NAND2_X1   g17700(.A1(new_n20824_), .A2(new_n20720_), .ZN(new_n20827_));
  INV_X1     g17701(.I(new_n20825_), .ZN(new_n20828_));
  OAI21_X1   g17702(.A1(new_n20827_), .A2(new_n20828_), .B(new_n20821_), .ZN(new_n20829_));
  NAND2_X1   g17703(.A1(new_n20826_), .A2(new_n20829_), .ZN(new_n20830_));
  OAI21_X1   g17704(.A1(new_n20830_), .A2(new_n14142_), .B(new_n20777_), .ZN(new_n20831_));
  NOR2_X1    g17705(.A1(new_n20720_), .A2(new_n13994_), .ZN(new_n20832_));
  AOI21_X1   g17706(.A1(new_n20831_), .A2(new_n13994_), .B(new_n20832_), .ZN(new_n20833_));
  NAND2_X1   g17707(.A1(new_n20721_), .A2(new_n14210_), .ZN(new_n20834_));
  OAI21_X1   g17708(.A1(new_n20833_), .A2(new_n14210_), .B(new_n20834_), .ZN(new_n20835_));
  NAND2_X1   g17709(.A1(new_n19370_), .A2(new_n14204_), .ZN(new_n20836_));
  NAND3_X1   g17710(.A1(new_n20835_), .A2(pi0715), .A3(new_n20836_), .ZN(new_n20837_));
  AOI22_X1   g17711(.A1(new_n20770_), .A2(new_n20776_), .B1(new_n14204_), .B2(new_n20837_), .ZN(new_n20838_));
  OAI21_X1   g17712(.A1(new_n20774_), .A2(new_n20760_), .B(new_n14005_), .ZN(new_n20839_));
  INV_X1     g17713(.I(new_n20768_), .ZN(new_n20840_));
  NAND2_X1   g17714(.A1(new_n20839_), .A2(new_n20840_), .ZN(new_n20841_));
  OAI22_X1   g17715(.A1(new_n20841_), .A2(pi1157), .B1(new_n20762_), .B2(new_n20765_), .ZN(new_n20842_));
  AOI21_X1   g17716(.A1(new_n20842_), .A2(pi0787), .B(new_n20775_), .ZN(new_n20843_));
  OAI21_X1   g17717(.A1(new_n20720_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n20844_));
  NAND3_X1   g17718(.A1(new_n20835_), .A2(pi0715), .A3(new_n20844_), .ZN(new_n20845_));
  AOI21_X1   g17719(.A1(new_n20843_), .A2(new_n20845_), .B(new_n14204_), .ZN(new_n20846_));
  OAI21_X1   g17720(.A1(new_n20846_), .A2(new_n20838_), .B(pi0790), .ZN(new_n20847_));
  NAND2_X1   g17721(.A1(new_n20835_), .A2(new_n20836_), .ZN(new_n20848_));
  NAND4_X1   g17722(.A1(new_n20835_), .A2(pi0644), .A3(pi0790), .A4(new_n20844_), .ZN(new_n20849_));
  NAND2_X1   g17723(.A1(new_n20835_), .A2(new_n20844_), .ZN(new_n20850_));
  NAND3_X1   g17724(.A1(new_n20850_), .A2(new_n14204_), .A3(pi0790), .ZN(new_n20851_));
  AOI21_X1   g17725(.A1(new_n20851_), .A2(new_n20849_), .B(new_n20848_), .ZN(new_n20852_));
  NOR2_X1    g17726(.A1(new_n20767_), .A2(new_n20768_), .ZN(new_n20853_));
  NOR4_X1    g17727(.A1(new_n20762_), .A2(pi0630), .A3(new_n14006_), .A4(new_n20763_), .ZN(new_n20854_));
  NOR3_X1    g17728(.A1(new_n20762_), .A2(pi0630), .A3(new_n20765_), .ZN(new_n20855_));
  NOR3_X1    g17729(.A1(new_n20855_), .A2(new_n20853_), .A3(new_n14012_), .ZN(new_n20856_));
  OAI21_X1   g17730(.A1(new_n20856_), .A2(new_n20854_), .B(pi0787), .ZN(new_n20857_));
  AOI21_X1   g17731(.A1(new_n20857_), .A2(new_n20833_), .B(new_n16867_), .ZN(new_n20858_));
  NOR2_X1    g17732(.A1(new_n20858_), .A2(new_n20852_), .ZN(new_n20859_));
  INV_X1     g17733(.I(new_n20743_), .ZN(new_n20860_));
  NAND2_X1   g17734(.A1(new_n13461_), .A2(pi0180), .ZN(new_n20861_));
  XOR2_X1    g17735(.A1(new_n20861_), .A2(new_n20779_), .Z(new_n20862_));
  NAND2_X1   g17736(.A1(new_n20862_), .A2(new_n13521_), .ZN(new_n20863_));
  NAND3_X1   g17737(.A1(new_n14270_), .A2(pi0180), .A3(pi0753), .ZN(new_n20864_));
  NAND3_X1   g17738(.A1(new_n14272_), .A2(new_n5642_), .A3(pi0753), .ZN(new_n20865_));
  AOI21_X1   g17739(.A1(new_n20864_), .A2(new_n20865_), .B(new_n13152_), .ZN(new_n20866_));
  NAND3_X1   g17740(.A1(new_n13198_), .A2(pi0180), .A3(pi0753), .ZN(new_n20867_));
  NAND3_X1   g17741(.A1(new_n13200_), .A2(pi0180), .A3(new_n17532_), .ZN(new_n20868_));
  AOI21_X1   g17742(.A1(new_n20868_), .A2(new_n20867_), .B(new_n13191_), .ZN(new_n20869_));
  OAI21_X1   g17743(.A1(new_n20866_), .A2(new_n3262_), .B(new_n20869_), .ZN(new_n20870_));
  NAND3_X1   g17744(.A1(new_n20863_), .A2(new_n3183_), .A3(new_n20870_), .ZN(new_n20871_));
  NOR2_X1    g17745(.A1(new_n14284_), .A2(new_n17532_), .ZN(new_n20872_));
  XOR2_X1    g17746(.A1(new_n20872_), .A2(new_n20778_), .Z(new_n20873_));
  NAND3_X1   g17747(.A1(new_n20871_), .A2(new_n20873_), .A3(new_n13359_), .ZN(new_n20874_));
  NAND3_X1   g17748(.A1(new_n20874_), .A2(new_n20724_), .A3(new_n3290_), .ZN(new_n20875_));
  OAI21_X1   g17749(.A1(new_n15587_), .A2(new_n5642_), .B(new_n17532_), .ZN(new_n20876_));
  NAND2_X1   g17750(.A1(new_n20876_), .A2(new_n13209_), .ZN(new_n20877_));
  NOR2_X1    g17751(.A1(new_n13105_), .A2(pi0753), .ZN(new_n20878_));
  INV_X1     g17752(.I(new_n20878_), .ZN(new_n20879_));
  NAND2_X1   g17753(.A1(new_n20879_), .A2(new_n16751_), .ZN(new_n20880_));
  NAND4_X1   g17754(.A1(new_n5503_), .A2(new_n20880_), .A3(pi0180), .A4(new_n3290_), .ZN(new_n20881_));
  AOI21_X1   g17755(.A1(new_n20877_), .A2(new_n3259_), .B(new_n20881_), .ZN(new_n20882_));
  NAND2_X1   g17756(.A1(new_n20875_), .A2(new_n20882_), .ZN(new_n20883_));
  AOI21_X1   g17757(.A1(new_n20883_), .A2(new_n20724_), .B(new_n20789_), .ZN(new_n20884_));
  INV_X1     g17758(.I(new_n20738_), .ZN(new_n20885_));
  INV_X1     g17759(.I(new_n20884_), .ZN(new_n20886_));
  NAND2_X1   g17760(.A1(new_n20792_), .A2(pi0625), .ZN(new_n20887_));
  XOR2_X1    g17761(.A1(new_n20887_), .A2(new_n13615_), .Z(new_n20888_));
  OAI21_X1   g17762(.A1(new_n20886_), .A2(new_n20888_), .B(new_n14081_), .ZN(new_n20889_));
  NAND2_X1   g17763(.A1(new_n20792_), .A2(pi1153), .ZN(new_n20890_));
  XOR2_X1    g17764(.A1(new_n20890_), .A2(new_n13620_), .Z(new_n20891_));
  AOI21_X1   g17765(.A1(new_n20884_), .A2(new_n20891_), .B(pi0608), .ZN(new_n20892_));
  OAI21_X1   g17766(.A1(new_n20889_), .A2(new_n20885_), .B(new_n20892_), .ZN(new_n20893_));
  NAND4_X1   g17767(.A1(new_n20893_), .A2(pi0778), .A3(new_n20720_), .A4(new_n20733_), .ZN(new_n20894_));
  OAI21_X1   g17768(.A1(pi0778), .A2(new_n20884_), .B(new_n20894_), .ZN(new_n20895_));
  NAND2_X1   g17769(.A1(new_n20895_), .A2(new_n13801_), .ZN(new_n20896_));
  NOR2_X1    g17770(.A1(new_n20895_), .A2(new_n13778_), .ZN(new_n20897_));
  NOR2_X1    g17771(.A1(new_n20897_), .A2(new_n14694_), .ZN(new_n20898_));
  NAND2_X1   g17772(.A1(new_n20897_), .A2(new_n14694_), .ZN(new_n20899_));
  INV_X1     g17773(.I(new_n20899_), .ZN(new_n20900_));
  OAI21_X1   g17774(.A1(new_n20900_), .A2(new_n20898_), .B(new_n20740_), .ZN(new_n20901_));
  NAND2_X1   g17775(.A1(new_n20796_), .A2(pi0660), .ZN(new_n20902_));
  INV_X1     g17776(.I(new_n20902_), .ZN(new_n20903_));
  NOR2_X1    g17777(.A1(new_n20801_), .A2(pi0660), .ZN(new_n20904_));
  INV_X1     g17778(.I(new_n20904_), .ZN(new_n20905_));
  AOI21_X1   g17779(.A1(new_n20901_), .A2(new_n20903_), .B(new_n20905_), .ZN(new_n20906_));
  NOR2_X1    g17780(.A1(new_n20895_), .A2(new_n13766_), .ZN(new_n20907_));
  XOR2_X1    g17781(.A1(new_n20907_), .A2(new_n14694_), .Z(new_n20908_));
  NAND2_X1   g17782(.A1(new_n20740_), .A2(pi0785), .ZN(new_n20909_));
  NOR2_X1    g17783(.A1(new_n20908_), .A2(new_n20909_), .ZN(new_n20910_));
  INV_X1     g17784(.I(new_n20910_), .ZN(new_n20911_));
  OAI21_X1   g17785(.A1(new_n20911_), .A2(new_n20906_), .B(new_n20896_), .ZN(new_n20912_));
  NAND3_X1   g17786(.A1(new_n20912_), .A2(pi0618), .A3(pi1154), .ZN(new_n20913_));
  INV_X1     g17787(.I(new_n20898_), .ZN(new_n20914_));
  AOI21_X1   g17788(.A1(new_n20914_), .A2(new_n20899_), .B(new_n20741_), .ZN(new_n20915_));
  OAI21_X1   g17789(.A1(new_n20915_), .A2(new_n20902_), .B(new_n20904_), .ZN(new_n20916_));
  AOI22_X1   g17790(.A1(new_n20916_), .A2(new_n20910_), .B1(new_n13801_), .B2(new_n20895_), .ZN(new_n20917_));
  NAND3_X1   g17791(.A1(new_n20917_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n20918_));
  AOI21_X1   g17792(.A1(new_n20918_), .A2(new_n20913_), .B(new_n20860_), .ZN(new_n20919_));
  NOR2_X1    g17793(.A1(new_n20807_), .A2(new_n13823_), .ZN(new_n20920_));
  INV_X1     g17794(.I(new_n20920_), .ZN(new_n20921_));
  OAI21_X1   g17795(.A1(new_n20919_), .A2(new_n20921_), .B(pi0781), .ZN(new_n20922_));
  NAND3_X1   g17796(.A1(new_n20912_), .A2(pi0618), .A3(pi1154), .ZN(new_n20923_));
  NAND3_X1   g17797(.A1(new_n20917_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n20924_));
  NAND2_X1   g17798(.A1(new_n20924_), .A2(new_n20923_), .ZN(new_n20925_));
  NAND3_X1   g17799(.A1(new_n20912_), .A2(new_n19177_), .A3(new_n20813_), .ZN(new_n20926_));
  AOI21_X1   g17800(.A1(new_n20925_), .A2(new_n20743_), .B(new_n20926_), .ZN(new_n20927_));
  NAND2_X1   g17801(.A1(new_n20922_), .A2(new_n20927_), .ZN(new_n20928_));
  AOI21_X1   g17802(.A1(new_n20917_), .A2(pi1154), .B(new_n13819_), .ZN(new_n20929_));
  NOR3_X1    g17803(.A1(new_n20912_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n20930_));
  OAI21_X1   g17804(.A1(new_n20929_), .A2(new_n20930_), .B(new_n20743_), .ZN(new_n20931_));
  AOI21_X1   g17805(.A1(new_n20931_), .A2(new_n20920_), .B(new_n13855_), .ZN(new_n20932_));
  AOI21_X1   g17806(.A1(new_n20917_), .A2(pi0618), .B(new_n13819_), .ZN(new_n20933_));
  NOR3_X1    g17807(.A1(new_n20912_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n20934_));
  OAI21_X1   g17808(.A1(new_n20933_), .A2(new_n20934_), .B(new_n20743_), .ZN(new_n20935_));
  NAND4_X1   g17809(.A1(new_n20935_), .A2(new_n19177_), .A3(new_n20813_), .A4(new_n20912_), .ZN(new_n20936_));
  NAND2_X1   g17810(.A1(new_n20936_), .A2(new_n20932_), .ZN(new_n20937_));
  NAND2_X1   g17811(.A1(new_n20937_), .A2(new_n20928_), .ZN(new_n20938_));
  NAND3_X1   g17812(.A1(new_n20938_), .A2(pi0619), .A3(pi1159), .ZN(new_n20939_));
  NOR2_X1    g17813(.A1(new_n20936_), .A2(new_n20932_), .ZN(new_n20940_));
  NOR2_X1    g17814(.A1(new_n20922_), .A2(new_n20927_), .ZN(new_n20941_));
  NOR2_X1    g17815(.A1(new_n20940_), .A2(new_n20941_), .ZN(new_n20942_));
  NAND3_X1   g17816(.A1(new_n20942_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n20943_));
  AOI21_X1   g17817(.A1(new_n20943_), .A2(new_n20939_), .B(new_n20745_), .ZN(new_n20944_));
  OAI21_X1   g17818(.A1(new_n20944_), .A2(new_n20003_), .B(new_n20820_), .ZN(new_n20945_));
  NAND2_X1   g17819(.A1(new_n20938_), .A2(new_n13896_), .ZN(new_n20946_));
  NAND3_X1   g17820(.A1(new_n20830_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n20947_));
  INV_X1     g17821(.I(new_n20830_), .ZN(new_n20948_));
  NAND3_X1   g17822(.A1(new_n20948_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n20949_));
  AOI21_X1   g17823(.A1(new_n20949_), .A2(new_n20947_), .B(new_n20721_), .ZN(new_n20950_));
  NOR2_X1    g17824(.A1(new_n20746_), .A2(new_n14162_), .ZN(new_n20951_));
  OAI21_X1   g17825(.A1(new_n20950_), .A2(new_n20951_), .B(new_n19204_), .ZN(new_n20952_));
  NOR2_X1    g17826(.A1(new_n20830_), .A2(new_n19208_), .ZN(new_n20953_));
  XNOR2_X1   g17827(.A1(new_n20953_), .A2(new_n19028_), .ZN(new_n20954_));
  NOR2_X1    g17828(.A1(new_n20721_), .A2(new_n15479_), .ZN(new_n20955_));
  NAND4_X1   g17829(.A1(new_n20952_), .A2(new_n20946_), .A3(new_n20954_), .A4(new_n20955_), .ZN(new_n20956_));
  INV_X1     g17830(.I(new_n20745_), .ZN(new_n20957_));
  AOI21_X1   g17831(.A1(new_n20942_), .A2(pi0619), .B(new_n13904_), .ZN(new_n20958_));
  NOR4_X1    g17832(.A1(new_n20940_), .A2(new_n20941_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n20959_));
  OAI21_X1   g17833(.A1(new_n20958_), .A2(new_n20959_), .B(new_n20957_), .ZN(new_n20960_));
  NAND3_X1   g17834(.A1(new_n20960_), .A2(new_n20173_), .A3(new_n20827_), .ZN(new_n20961_));
  AOI21_X1   g17835(.A1(new_n20945_), .A2(new_n20956_), .B(new_n20961_), .ZN(new_n20962_));
  AND2_X2    g17836(.A1(new_n20752_), .A2(pi0629), .Z(new_n20963_));
  NOR2_X1    g17837(.A1(new_n20772_), .A2(pi0629), .ZN(new_n20964_));
  NOR2_X1    g17838(.A1(new_n9992_), .A2(pi0180), .ZN(new_n20965_));
  NOR3_X1    g17839(.A1(new_n13219_), .A2(pi0625), .A3(pi0702), .ZN(new_n20966_));
  INV_X1     g17840(.I(new_n20966_), .ZN(new_n20967_));
  NOR2_X1    g17841(.A1(new_n20965_), .A2(pi1153), .ZN(new_n20968_));
  NAND2_X1   g17842(.A1(new_n20967_), .A2(new_n20968_), .ZN(new_n20969_));
  INV_X1     g17843(.I(new_n20969_), .ZN(new_n20970_));
  NOR2_X1    g17844(.A1(new_n20970_), .A2(new_n13748_), .ZN(new_n20971_));
  AOI21_X1   g17845(.A1(new_n13218_), .A2(new_n20724_), .B(new_n20965_), .ZN(new_n20972_));
  INV_X1     g17846(.I(new_n20972_), .ZN(new_n20973_));
  AOI21_X1   g17847(.A1(new_n20967_), .A2(new_n20973_), .B(new_n13614_), .ZN(new_n20974_));
  INV_X1     g17848(.I(new_n20974_), .ZN(new_n20975_));
  NOR3_X1    g17849(.A1(new_n20975_), .A2(new_n13748_), .A3(new_n20973_), .ZN(new_n20976_));
  XNOR2_X1   g17850(.A1(new_n20976_), .A2(new_n20971_), .ZN(new_n20977_));
  NAND2_X1   g17851(.A1(new_n20977_), .A2(new_n14049_), .ZN(new_n20978_));
  NOR2_X1    g17852(.A1(new_n20978_), .A2(new_n14051_), .ZN(new_n20979_));
  INV_X1     g17853(.I(new_n20979_), .ZN(new_n20980_));
  NOR2_X1    g17854(.A1(new_n20980_), .A2(new_n14163_), .ZN(new_n20981_));
  NOR2_X1    g17855(.A1(new_n20878_), .A2(new_n20965_), .ZN(new_n20982_));
  INV_X1     g17856(.I(new_n20982_), .ZN(new_n20983_));
  NAND3_X1   g17857(.A1(new_n20983_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n20984_));
  AOI21_X1   g17858(.A1(new_n20984_), .A2(new_n16444_), .B(new_n20879_), .ZN(new_n20985_));
  NOR2_X1    g17859(.A1(new_n20985_), .A2(new_n13801_), .ZN(new_n20986_));
  NOR2_X1    g17860(.A1(new_n20965_), .A2(pi1155), .ZN(new_n20987_));
  NOR3_X1    g17861(.A1(new_n20879_), .A2(new_n16444_), .A3(new_n20987_), .ZN(new_n20988_));
  NAND4_X1   g17862(.A1(new_n20988_), .A2(new_n20983_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n20989_));
  XOR2_X1    g17863(.A1(new_n20986_), .A2(new_n20989_), .Z(new_n20990_));
  NOR2_X1    g17864(.A1(new_n20990_), .A2(new_n13817_), .ZN(new_n20991_));
  OAI21_X1   g17865(.A1(new_n20991_), .A2(pi0618), .B(new_n9992_), .ZN(new_n20992_));
  NAND2_X1   g17866(.A1(new_n20992_), .A2(pi0781), .ZN(new_n20993_));
  OAI21_X1   g17867(.A1(new_n20991_), .A2(new_n9992_), .B(pi0618), .ZN(new_n20994_));
  NOR3_X1    g17868(.A1(new_n20994_), .A2(new_n13855_), .A3(new_n20990_), .ZN(new_n20995_));
  XOR2_X1    g17869(.A1(new_n20995_), .A2(new_n20993_), .Z(new_n20996_));
  NOR2_X1    g17870(.A1(new_n20996_), .A2(new_n13868_), .ZN(new_n20997_));
  OAI21_X1   g17871(.A1(new_n20997_), .A2(pi0619), .B(new_n9992_), .ZN(new_n20998_));
  NAND2_X1   g17872(.A1(new_n20998_), .A2(pi0789), .ZN(new_n20999_));
  OAI21_X1   g17873(.A1(new_n20997_), .A2(new_n9992_), .B(pi0619), .ZN(new_n21000_));
  NOR3_X1    g17874(.A1(new_n21000_), .A2(new_n13896_), .A3(new_n20996_), .ZN(new_n21001_));
  XOR2_X1    g17875(.A1(new_n21001_), .A2(new_n20999_), .Z(new_n21002_));
  NAND2_X1   g17876(.A1(new_n21002_), .A2(new_n13962_), .ZN(new_n21003_));
  XOR2_X1    g17877(.A1(new_n21003_), .A2(new_n18976_), .Z(new_n21004_));
  AOI22_X1   g17878(.A1(new_n21004_), .A2(new_n20965_), .B1(new_n16639_), .B2(new_n20981_), .ZN(new_n21005_));
  NOR2_X1    g17879(.A1(new_n20972_), .A2(new_n13203_), .ZN(new_n21006_));
  NAND2_X1   g17880(.A1(new_n21006_), .A2(pi0625), .ZN(new_n21007_));
  NAND3_X1   g17881(.A1(new_n21007_), .A2(pi1153), .A3(new_n20982_), .ZN(new_n21008_));
  NOR2_X1    g17882(.A1(new_n20970_), .A2(new_n14081_), .ZN(new_n21009_));
  AOI21_X1   g17883(.A1(new_n21009_), .A2(new_n21008_), .B(new_n13748_), .ZN(new_n21010_));
  NOR2_X1    g17884(.A1(new_n20983_), .A2(new_n21006_), .ZN(new_n21011_));
  INV_X1     g17885(.I(new_n21007_), .ZN(new_n21012_));
  OAI21_X1   g17886(.A1(new_n21011_), .A2(new_n21012_), .B(new_n20968_), .ZN(new_n21013_));
  NAND4_X1   g17887(.A1(new_n21013_), .A2(new_n13749_), .A3(new_n20975_), .A4(new_n21011_), .ZN(new_n21014_));
  XNOR2_X1   g17888(.A1(new_n21014_), .A2(new_n21010_), .ZN(new_n21015_));
  NAND2_X1   g17889(.A1(new_n21015_), .A2(new_n13801_), .ZN(new_n21016_));
  NOR2_X1    g17890(.A1(new_n20985_), .A2(pi0660), .ZN(new_n21020_));
  NOR2_X1    g17891(.A1(new_n21015_), .A2(new_n13766_), .ZN(new_n21021_));
  XOR2_X1    g17892(.A1(new_n21021_), .A2(new_n14090_), .Z(new_n21022_));
  NOR2_X1    g17893(.A1(new_n20977_), .A2(new_n13801_), .ZN(new_n21023_));
  NAND2_X1   g17894(.A1(new_n21022_), .A2(new_n21023_), .ZN(new_n21024_));
  OAI21_X1   g17895(.A1(new_n21024_), .A2(new_n21020_), .B(new_n21016_), .ZN(new_n21025_));
  NAND2_X1   g17896(.A1(new_n21025_), .A2(new_n13855_), .ZN(new_n21026_));
  INV_X1     g17897(.I(new_n20978_), .ZN(new_n21027_));
  NOR2_X1    g17898(.A1(new_n21025_), .A2(new_n13816_), .ZN(new_n21028_));
  XOR2_X1    g17899(.A1(new_n21028_), .A2(new_n13818_), .Z(new_n21029_));
  NAND2_X1   g17900(.A1(new_n21029_), .A2(new_n21027_), .ZN(new_n21030_));
  NAND3_X1   g17901(.A1(new_n21030_), .A2(new_n13823_), .A3(new_n20994_), .ZN(new_n21031_));
  NAND3_X1   g17902(.A1(new_n21031_), .A2(new_n13823_), .A3(new_n20992_), .ZN(new_n21032_));
  NOR2_X1    g17903(.A1(new_n21025_), .A2(new_n13817_), .ZN(new_n21033_));
  XOR2_X1    g17904(.A1(new_n21033_), .A2(new_n13818_), .Z(new_n21034_));
  NAND4_X1   g17905(.A1(new_n21032_), .A2(pi0781), .A3(new_n21027_), .A4(new_n21034_), .ZN(new_n21035_));
  NAND2_X1   g17906(.A1(new_n21035_), .A2(new_n21026_), .ZN(new_n21036_));
  NOR2_X1    g17907(.A1(new_n21036_), .A2(new_n13860_), .ZN(new_n21037_));
  XOR2_X1    g17908(.A1(new_n21037_), .A2(new_n13904_), .Z(new_n21038_));
  NOR2_X1    g17909(.A1(new_n21038_), .A2(new_n20980_), .ZN(new_n21039_));
  NAND2_X1   g17910(.A1(new_n21000_), .A2(new_n13884_), .ZN(new_n21040_));
  INV_X1     g17911(.I(new_n21036_), .ZN(new_n21041_));
  AOI21_X1   g17912(.A1(new_n21041_), .A2(new_n14143_), .B(pi0789), .ZN(new_n21042_));
  OAI21_X1   g17913(.A1(new_n21039_), .A2(new_n21040_), .B(new_n21042_), .ZN(new_n21043_));
  NOR2_X1    g17914(.A1(new_n21036_), .A2(new_n13868_), .ZN(new_n21044_));
  XOR2_X1    g17915(.A1(new_n21044_), .A2(new_n13903_), .Z(new_n21045_));
  NAND2_X1   g17916(.A1(new_n20998_), .A2(new_n19018_), .ZN(new_n21046_));
  AOI21_X1   g17917(.A1(new_n21045_), .A2(new_n20979_), .B(new_n21046_), .ZN(new_n21047_));
  AOI21_X1   g17918(.A1(new_n21043_), .A2(new_n21047_), .B(new_n21005_), .ZN(new_n21048_));
  NOR3_X1    g17919(.A1(new_n20980_), .A2(new_n14163_), .A3(new_n18928_), .ZN(new_n21049_));
  NAND2_X1   g17920(.A1(new_n21002_), .A2(new_n16372_), .ZN(new_n21050_));
  OAI21_X1   g17921(.A1(new_n16372_), .A2(new_n20965_), .B(new_n21050_), .ZN(new_n21051_));
  NAND2_X1   g17922(.A1(new_n21051_), .A2(new_n21049_), .ZN(new_n21052_));
  NAND2_X1   g17923(.A1(new_n21052_), .A2(new_n19022_), .ZN(new_n21053_));
  NAND2_X1   g17924(.A1(new_n21052_), .A2(new_n16569_), .ZN(new_n21054_));
  XNOR2_X1   g17925(.A1(new_n21054_), .A2(new_n16572_), .ZN(new_n21055_));
  AOI21_X1   g17926(.A1(new_n21055_), .A2(new_n21053_), .B(new_n16574_), .ZN(new_n21056_));
  NAND2_X1   g17927(.A1(new_n21002_), .A2(new_n13963_), .ZN(new_n21057_));
  XNOR2_X1   g17928(.A1(new_n21057_), .A2(new_n19028_), .ZN(new_n21058_));
  NAND2_X1   g17929(.A1(new_n16423_), .A2(new_n20965_), .ZN(new_n21059_));
  NOR4_X1    g17930(.A1(new_n21048_), .A2(new_n21056_), .A3(new_n21058_), .A4(new_n21059_), .ZN(new_n21060_));
  INV_X1     g17931(.I(new_n20965_), .ZN(new_n21061_));
  NAND2_X1   g17932(.A1(new_n21049_), .A2(new_n14061_), .ZN(new_n21062_));
  NAND2_X1   g17933(.A1(new_n20965_), .A2(new_n14005_), .ZN(new_n21063_));
  OAI21_X1   g17934(.A1(new_n21062_), .A2(new_n14005_), .B(new_n21063_), .ZN(new_n21064_));
  NOR2_X1    g17935(.A1(new_n21051_), .A2(new_n13994_), .ZN(new_n21065_));
  XOR2_X1    g17936(.A1(new_n21065_), .A2(new_n19033_), .Z(new_n21066_));
  OAI22_X1   g17937(.A1(new_n21066_), .A2(new_n21061_), .B1(new_n14207_), .B2(new_n21064_), .ZN(new_n21067_));
  NAND2_X1   g17938(.A1(new_n21062_), .A2(pi0647), .ZN(new_n21068_));
  XOR2_X1    g17939(.A1(new_n21068_), .A2(new_n14007_), .Z(new_n21069_));
  NOR3_X1    g17940(.A1(new_n21069_), .A2(new_n14010_), .A3(new_n21061_), .ZN(new_n21070_));
  AOI21_X1   g17941(.A1(new_n21067_), .A2(new_n21070_), .B(new_n12776_), .ZN(new_n21071_));
  NOR2_X1    g17942(.A1(new_n21060_), .A2(new_n21071_), .ZN(new_n21072_));
  NOR2_X1    g17943(.A1(new_n21069_), .A2(new_n21061_), .ZN(new_n21073_));
  OAI21_X1   g17944(.A1(new_n21064_), .A2(new_n14006_), .B(pi0787), .ZN(new_n21074_));
  OAI22_X1   g17945(.A1(new_n21073_), .A2(new_n21074_), .B1(pi0787), .B2(new_n21062_), .ZN(new_n21075_));
  NOR2_X1    g17946(.A1(new_n21072_), .A2(new_n14204_), .ZN(new_n21076_));
  XOR2_X1    g17947(.A1(new_n21076_), .A2(new_n14205_), .Z(new_n21077_));
  NAND2_X1   g17948(.A1(new_n21077_), .A2(new_n21075_), .ZN(new_n21078_));
  NOR2_X1    g17949(.A1(new_n21051_), .A2(new_n18968_), .ZN(new_n21079_));
  NAND2_X1   g17950(.A1(new_n18967_), .A2(new_n20965_), .ZN(new_n21080_));
  XOR2_X1    g17951(.A1(new_n21079_), .A2(new_n21080_), .Z(new_n21081_));
  NAND2_X1   g17952(.A1(new_n21081_), .A2(pi0715), .ZN(new_n21082_));
  XOR2_X1    g17953(.A1(new_n21082_), .A2(new_n14217_), .Z(new_n21083_));
  AOI21_X1   g17954(.A1(new_n21083_), .A2(new_n20965_), .B(pi1160), .ZN(new_n21084_));
  NAND2_X1   g17955(.A1(new_n21081_), .A2(pi0644), .ZN(new_n21085_));
  XOR2_X1    g17956(.A1(new_n21085_), .A2(new_n14205_), .Z(new_n21086_));
  OAI21_X1   g17957(.A1(new_n21086_), .A2(new_n21061_), .B(new_n14203_), .ZN(new_n21087_));
  AOI21_X1   g17958(.A1(new_n21078_), .A2(new_n21084_), .B(new_n21087_), .ZN(new_n21088_));
  NOR2_X1    g17959(.A1(new_n21072_), .A2(new_n14200_), .ZN(new_n21089_));
  XOR2_X1    g17960(.A1(new_n21089_), .A2(new_n14205_), .Z(new_n21090_));
  NAND2_X1   g17961(.A1(new_n21090_), .A2(new_n21075_), .ZN(new_n21091_));
  OAI21_X1   g17962(.A1(new_n21088_), .A2(new_n21091_), .B(pi0832), .ZN(new_n21092_));
  XOR2_X1    g17963(.A1(new_n21092_), .A2(new_n14801_), .Z(new_n21093_));
  NAND2_X1   g17964(.A1(po1038), .A2(new_n5642_), .ZN(new_n21094_));
  NAND4_X1   g17965(.A1(new_n21093_), .A2(new_n14799_), .A3(new_n21072_), .A4(new_n21094_), .ZN(new_n21095_));
  NAND2_X1   g17966(.A1(new_n21095_), .A2(new_n7240_), .ZN(new_n21096_));
  OAI21_X1   g17967(.A1(new_n20963_), .A2(new_n20964_), .B(new_n21096_), .ZN(new_n21097_));
  AOI21_X1   g17968(.A1(new_n16875_), .A2(new_n20831_), .B(new_n21097_), .ZN(new_n21098_));
  OAI21_X1   g17969(.A1(new_n20962_), .A2(pi0792), .B(new_n21098_), .ZN(new_n21099_));
  AOI21_X1   g17970(.A1(new_n20859_), .A2(new_n20847_), .B(new_n21099_), .ZN(po0337));
  NOR2_X1    g17971(.A1(new_n14428_), .A2(pi0181), .ZN(new_n21101_));
  INV_X1     g17972(.I(new_n21101_), .ZN(new_n21102_));
  NAND2_X1   g17973(.A1(new_n21102_), .A2(new_n13965_), .ZN(new_n21103_));
  NOR2_X1    g17974(.A1(new_n21102_), .A2(new_n13919_), .ZN(new_n21104_));
  INV_X1     g17975(.I(pi0709), .ZN(new_n21105_));
  OAI21_X1   g17976(.A1(new_n13721_), .A2(new_n21105_), .B(new_n5643_), .ZN(new_n21106_));
  NAND2_X1   g17977(.A1(new_n16715_), .A2(new_n5643_), .ZN(new_n21107_));
  NAND4_X1   g17978(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n21106_), .A4(new_n21107_), .ZN(new_n21108_));
  AOI21_X1   g17979(.A1(new_n21108_), .A2(new_n14424_), .B(new_n5643_), .ZN(new_n21109_));
  NAND2_X1   g17980(.A1(new_n21101_), .A2(new_n21109_), .ZN(new_n21110_));
  NAND2_X1   g17981(.A1(new_n21110_), .A2(new_n3290_), .ZN(new_n21111_));
  NAND2_X1   g17982(.A1(new_n21111_), .A2(pi0709), .ZN(new_n21112_));
  NAND2_X1   g17983(.A1(new_n21112_), .A2(pi0625), .ZN(new_n21113_));
  XOR2_X1    g17984(.A1(new_n21113_), .A2(new_n13620_), .Z(new_n21114_));
  NAND2_X1   g17985(.A1(new_n21114_), .A2(new_n21101_), .ZN(new_n21115_));
  NAND2_X1   g17986(.A1(new_n21115_), .A2(pi0778), .ZN(new_n21116_));
  NAND2_X1   g17987(.A1(new_n21112_), .A2(pi1153), .ZN(new_n21117_));
  XOR2_X1    g17988(.A1(new_n21117_), .A2(new_n13620_), .Z(new_n21118_));
  NAND2_X1   g17989(.A1(new_n21118_), .A2(new_n21101_), .ZN(new_n21119_));
  NOR3_X1    g17990(.A1(new_n21119_), .A2(new_n13748_), .A3(new_n21112_), .ZN(new_n21120_));
  XNOR2_X1   g17991(.A1(new_n21120_), .A2(new_n21116_), .ZN(new_n21121_));
  INV_X1     g17992(.I(new_n21121_), .ZN(new_n21122_));
  NAND2_X1   g17993(.A1(new_n21101_), .A2(new_n13803_), .ZN(new_n21123_));
  OAI21_X1   g17994(.A1(new_n21122_), .A2(new_n13803_), .B(new_n21123_), .ZN(new_n21124_));
  NOR2_X1    g17995(.A1(new_n21124_), .A2(new_n13879_), .ZN(new_n21125_));
  AOI21_X1   g17996(.A1(new_n13879_), .A2(new_n21102_), .B(new_n21125_), .ZN(new_n21126_));
  AOI21_X1   g17997(.A1(new_n21126_), .A2(new_n13919_), .B(new_n21104_), .ZN(new_n21127_));
  NAND2_X1   g17998(.A1(new_n21127_), .A2(new_n13966_), .ZN(new_n21128_));
  NAND2_X1   g17999(.A1(new_n21128_), .A2(new_n21103_), .ZN(new_n21129_));
  INV_X1     g18000(.I(new_n21129_), .ZN(new_n21130_));
  AOI21_X1   g18001(.A1(new_n21130_), .A2(pi0628), .B(new_n13971_), .ZN(new_n21131_));
  NOR3_X1    g18002(.A1(new_n21129_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n21132_));
  OAI21_X1   g18003(.A1(new_n21131_), .A2(new_n21132_), .B(new_n21101_), .ZN(new_n21133_));
  NAND2_X1   g18004(.A1(new_n21133_), .A2(pi0792), .ZN(new_n21134_));
  NAND3_X1   g18005(.A1(new_n21129_), .A2(pi0628), .A3(pi1156), .ZN(new_n21135_));
  INV_X1     g18006(.I(new_n21135_), .ZN(new_n21136_));
  NOR3_X1    g18007(.A1(new_n21129_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n21137_));
  NOR2_X1    g18008(.A1(new_n21136_), .A2(new_n21137_), .ZN(new_n21138_));
  NOR4_X1    g18009(.A1(new_n21138_), .A2(new_n12777_), .A3(new_n21102_), .A4(new_n21130_), .ZN(new_n21139_));
  NAND2_X1   g18010(.A1(new_n21139_), .A2(new_n21134_), .ZN(new_n21140_));
  NOR2_X1    g18011(.A1(new_n21139_), .A2(new_n21134_), .ZN(new_n21141_));
  INV_X1     g18012(.I(new_n21141_), .ZN(new_n21142_));
  AOI21_X1   g18013(.A1(new_n21142_), .A2(new_n21140_), .B(new_n14005_), .ZN(new_n21143_));
  NOR2_X1    g18014(.A1(new_n21102_), .A2(pi0647), .ZN(new_n21144_));
  NOR2_X1    g18015(.A1(new_n21144_), .A2(new_n14006_), .ZN(new_n21145_));
  INV_X1     g18016(.I(new_n21145_), .ZN(new_n21146_));
  NOR2_X1    g18017(.A1(new_n21143_), .A2(new_n21146_), .ZN(new_n21147_));
  AOI21_X1   g18018(.A1(new_n21142_), .A2(new_n21140_), .B(pi0647), .ZN(new_n21148_));
  NOR2_X1    g18019(.A1(new_n21102_), .A2(new_n14005_), .ZN(new_n21149_));
  NOR3_X1    g18020(.A1(new_n21148_), .A2(pi1157), .A3(new_n21149_), .ZN(new_n21150_));
  OAI21_X1   g18021(.A1(new_n21150_), .A2(new_n21147_), .B(pi0787), .ZN(new_n21151_));
  NAND3_X1   g18022(.A1(new_n21130_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n21152_));
  AOI21_X1   g18023(.A1(new_n21152_), .A2(new_n21135_), .B(new_n21102_), .ZN(new_n21153_));
  NAND3_X1   g18024(.A1(new_n21153_), .A2(pi0792), .A3(new_n21129_), .ZN(new_n21154_));
  AOI21_X1   g18025(.A1(pi0792), .A2(new_n21133_), .B(new_n21154_), .ZN(new_n21155_));
  NOR3_X1    g18026(.A1(new_n21155_), .A2(pi0787), .A3(new_n21141_), .ZN(new_n21156_));
  INV_X1     g18027(.I(new_n21156_), .ZN(new_n21157_));
  NAND2_X1   g18028(.A1(new_n21102_), .A2(new_n14142_), .ZN(new_n21158_));
  NOR2_X1    g18029(.A1(new_n5643_), .A2(new_n17569_), .ZN(new_n21159_));
  INV_X1     g18030(.I(new_n21159_), .ZN(new_n21160_));
  NAND2_X1   g18031(.A1(new_n20780_), .A2(new_n21160_), .ZN(new_n21161_));
  OAI21_X1   g18032(.A1(new_n14298_), .A2(new_n5643_), .B(new_n3183_), .ZN(new_n21162_));
  AOI21_X1   g18033(.A1(new_n13194_), .A2(pi0754), .B(new_n21162_), .ZN(new_n21163_));
  OAI21_X1   g18034(.A1(new_n21163_), .A2(new_n17569_), .B(pi0181), .ZN(new_n21164_));
  OAI21_X1   g18035(.A1(new_n20785_), .A2(new_n21164_), .B(new_n3183_), .ZN(new_n21165_));
  AOI21_X1   g18036(.A1(new_n13109_), .A2(new_n5643_), .B(new_n3259_), .ZN(new_n21166_));
  AND3_X2    g18037(.A1(new_n21161_), .A2(new_n21165_), .A3(new_n21166_), .Z(new_n21167_));
  OAI21_X1   g18038(.A1(new_n21167_), .A2(new_n13106_), .B(pi0754), .ZN(new_n21168_));
  INV_X1     g18039(.I(new_n21168_), .ZN(new_n21169_));
  NOR2_X1    g18040(.A1(new_n3289_), .A2(pi0181), .ZN(new_n21170_));
  AOI21_X1   g18041(.A1(new_n21169_), .A2(new_n3289_), .B(new_n21170_), .ZN(new_n21171_));
  NAND2_X1   g18042(.A1(new_n21171_), .A2(new_n13776_), .ZN(new_n21172_));
  NAND2_X1   g18043(.A1(new_n21102_), .A2(new_n13780_), .ZN(new_n21173_));
  NAND2_X1   g18044(.A1(new_n21172_), .A2(new_n21173_), .ZN(new_n21174_));
  NAND2_X1   g18045(.A1(new_n21174_), .A2(pi0609), .ZN(new_n21175_));
  NAND2_X1   g18046(.A1(new_n21175_), .A2(pi0785), .ZN(new_n21176_));
  NAND2_X1   g18047(.A1(new_n21101_), .A2(new_n13775_), .ZN(new_n21177_));
  OAI21_X1   g18048(.A1(new_n21171_), .A2(new_n13775_), .B(new_n21177_), .ZN(new_n21178_));
  AOI21_X1   g18049(.A1(new_n21102_), .A2(new_n14467_), .B(pi0609), .ZN(new_n21179_));
  NOR2_X1    g18050(.A1(new_n21172_), .A2(new_n21179_), .ZN(new_n21180_));
  NAND3_X1   g18051(.A1(new_n21180_), .A2(pi0785), .A3(new_n21178_), .ZN(new_n21181_));
  XNOR2_X1   g18052(.A1(new_n21176_), .A2(new_n21181_), .ZN(new_n21182_));
  INV_X1     g18053(.I(new_n21182_), .ZN(new_n21183_));
  NAND3_X1   g18054(.A1(new_n21183_), .A2(pi0618), .A3(pi1154), .ZN(new_n21184_));
  NAND3_X1   g18055(.A1(new_n21182_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n21185_));
  AOI21_X1   g18056(.A1(new_n21184_), .A2(new_n21185_), .B(new_n21102_), .ZN(new_n21186_));
  NAND3_X1   g18057(.A1(new_n21183_), .A2(pi0618), .A3(pi1154), .ZN(new_n21187_));
  NAND3_X1   g18058(.A1(new_n21182_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n21188_));
  AOI21_X1   g18059(.A1(new_n21187_), .A2(new_n21188_), .B(new_n21102_), .ZN(new_n21189_));
  NAND4_X1   g18060(.A1(new_n21186_), .A2(new_n21189_), .A3(pi0781), .A4(new_n21183_), .ZN(new_n21190_));
  NOR2_X1    g18061(.A1(new_n21186_), .A2(new_n13855_), .ZN(new_n21191_));
  INV_X1     g18062(.I(new_n21189_), .ZN(new_n21192_));
  NAND2_X1   g18063(.A1(new_n21183_), .A2(pi0781), .ZN(new_n21193_));
  OAI21_X1   g18064(.A1(new_n21192_), .A2(new_n21193_), .B(new_n21191_), .ZN(new_n21194_));
  NAND2_X1   g18065(.A1(new_n21194_), .A2(new_n21190_), .ZN(new_n21195_));
  NAND3_X1   g18066(.A1(new_n21195_), .A2(pi0619), .A3(pi1159), .ZN(new_n21196_));
  INV_X1     g18067(.I(new_n21195_), .ZN(new_n21197_));
  NAND3_X1   g18068(.A1(new_n21197_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n21198_));
  AOI21_X1   g18069(.A1(new_n21198_), .A2(new_n21196_), .B(new_n21102_), .ZN(new_n21199_));
  NOR2_X1    g18070(.A1(new_n21199_), .A2(new_n13896_), .ZN(new_n21200_));
  INV_X1     g18071(.I(new_n21200_), .ZN(new_n21201_));
  NOR2_X1    g18072(.A1(new_n21195_), .A2(new_n13868_), .ZN(new_n21202_));
  XOR2_X1    g18073(.A1(new_n21202_), .A2(new_n13903_), .Z(new_n21203_));
  NOR2_X1    g18074(.A1(new_n21197_), .A2(new_n13896_), .ZN(new_n21204_));
  NAND4_X1   g18075(.A1(new_n21201_), .A2(new_n21101_), .A3(new_n21203_), .A4(new_n21204_), .ZN(new_n21205_));
  NAND2_X1   g18076(.A1(new_n21203_), .A2(new_n21101_), .ZN(new_n21206_));
  INV_X1     g18077(.I(new_n21204_), .ZN(new_n21207_));
  OAI21_X1   g18078(.A1(new_n21206_), .A2(new_n21207_), .B(new_n21200_), .ZN(new_n21208_));
  NAND2_X1   g18079(.A1(new_n21205_), .A2(new_n21208_), .ZN(new_n21209_));
  OAI21_X1   g18080(.A1(new_n21209_), .A2(new_n14142_), .B(new_n21158_), .ZN(new_n21210_));
  NOR2_X1    g18081(.A1(new_n21101_), .A2(new_n13994_), .ZN(new_n21211_));
  AOI21_X1   g18082(.A1(new_n21210_), .A2(new_n13994_), .B(new_n21211_), .ZN(new_n21212_));
  NAND2_X1   g18083(.A1(new_n21102_), .A2(new_n14210_), .ZN(new_n21213_));
  OAI21_X1   g18084(.A1(new_n21212_), .A2(new_n14210_), .B(new_n21213_), .ZN(new_n21214_));
  NAND2_X1   g18085(.A1(new_n19370_), .A2(new_n14204_), .ZN(new_n21215_));
  NAND3_X1   g18086(.A1(new_n21214_), .A2(pi0715), .A3(new_n21215_), .ZN(new_n21216_));
  AOI22_X1   g18087(.A1(new_n21151_), .A2(new_n21157_), .B1(new_n14204_), .B2(new_n21216_), .ZN(new_n21217_));
  OAI21_X1   g18088(.A1(new_n21155_), .A2(new_n21141_), .B(new_n14005_), .ZN(new_n21218_));
  INV_X1     g18089(.I(new_n21149_), .ZN(new_n21219_));
  NAND2_X1   g18090(.A1(new_n21218_), .A2(new_n21219_), .ZN(new_n21220_));
  OAI22_X1   g18091(.A1(new_n21220_), .A2(pi1157), .B1(new_n21143_), .B2(new_n21146_), .ZN(new_n21221_));
  AOI21_X1   g18092(.A1(new_n21221_), .A2(pi0787), .B(new_n21156_), .ZN(new_n21222_));
  OAI21_X1   g18093(.A1(new_n21101_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n21223_));
  NAND3_X1   g18094(.A1(new_n21214_), .A2(pi0715), .A3(new_n21223_), .ZN(new_n21224_));
  AOI21_X1   g18095(.A1(new_n21222_), .A2(new_n21224_), .B(new_n14204_), .ZN(new_n21225_));
  OAI21_X1   g18096(.A1(new_n21225_), .A2(new_n21217_), .B(pi0790), .ZN(new_n21226_));
  NAND2_X1   g18097(.A1(new_n21214_), .A2(new_n21215_), .ZN(new_n21227_));
  NAND4_X1   g18098(.A1(new_n21214_), .A2(pi0644), .A3(pi0790), .A4(new_n21223_), .ZN(new_n21228_));
  NAND2_X1   g18099(.A1(new_n21214_), .A2(new_n21223_), .ZN(new_n21229_));
  NAND3_X1   g18100(.A1(new_n21229_), .A2(new_n14204_), .A3(pi0790), .ZN(new_n21230_));
  AOI21_X1   g18101(.A1(new_n21230_), .A2(new_n21228_), .B(new_n21227_), .ZN(new_n21231_));
  NOR2_X1    g18102(.A1(new_n21148_), .A2(new_n21149_), .ZN(new_n21232_));
  NOR4_X1    g18103(.A1(new_n21143_), .A2(pi0630), .A3(new_n14006_), .A4(new_n21144_), .ZN(new_n21233_));
  NOR3_X1    g18104(.A1(new_n21143_), .A2(pi0630), .A3(new_n21146_), .ZN(new_n21234_));
  NOR3_X1    g18105(.A1(new_n21234_), .A2(new_n21232_), .A3(new_n14012_), .ZN(new_n21235_));
  OAI21_X1   g18106(.A1(new_n21235_), .A2(new_n21233_), .B(pi0787), .ZN(new_n21236_));
  AOI21_X1   g18107(.A1(new_n21236_), .A2(new_n21212_), .B(new_n16867_), .ZN(new_n21237_));
  NOR2_X1    g18108(.A1(new_n21237_), .A2(new_n21231_), .ZN(new_n21238_));
  INV_X1     g18109(.I(new_n21124_), .ZN(new_n21239_));
  NAND2_X1   g18110(.A1(new_n13461_), .A2(pi0181), .ZN(new_n21240_));
  XOR2_X1    g18111(.A1(new_n21240_), .A2(new_n21160_), .Z(new_n21241_));
  NAND2_X1   g18112(.A1(new_n21241_), .A2(new_n13521_), .ZN(new_n21242_));
  NAND3_X1   g18113(.A1(new_n14270_), .A2(pi0181), .A3(pi0754), .ZN(new_n21243_));
  NAND3_X1   g18114(.A1(new_n14272_), .A2(new_n5643_), .A3(pi0754), .ZN(new_n21244_));
  AOI21_X1   g18115(.A1(new_n21243_), .A2(new_n21244_), .B(new_n13152_), .ZN(new_n21245_));
  NAND3_X1   g18116(.A1(new_n13198_), .A2(pi0181), .A3(pi0754), .ZN(new_n21246_));
  NAND3_X1   g18117(.A1(new_n13200_), .A2(pi0181), .A3(new_n17569_), .ZN(new_n21247_));
  AOI21_X1   g18118(.A1(new_n21247_), .A2(new_n21246_), .B(new_n13191_), .ZN(new_n21248_));
  OAI21_X1   g18119(.A1(new_n21245_), .A2(new_n3262_), .B(new_n21248_), .ZN(new_n21249_));
  NAND3_X1   g18120(.A1(new_n21242_), .A2(new_n3183_), .A3(new_n21249_), .ZN(new_n21250_));
  NOR2_X1    g18121(.A1(new_n14284_), .A2(new_n17569_), .ZN(new_n21251_));
  XOR2_X1    g18122(.A1(new_n21251_), .A2(new_n21159_), .Z(new_n21252_));
  NAND3_X1   g18123(.A1(new_n21250_), .A2(new_n21252_), .A3(new_n13359_), .ZN(new_n21253_));
  NAND3_X1   g18124(.A1(new_n21253_), .A2(new_n21105_), .A3(new_n3290_), .ZN(new_n21254_));
  OAI21_X1   g18125(.A1(new_n15587_), .A2(new_n5643_), .B(new_n17569_), .ZN(new_n21255_));
  NAND2_X1   g18126(.A1(new_n21255_), .A2(new_n13209_), .ZN(new_n21256_));
  NOR2_X1    g18127(.A1(new_n13105_), .A2(pi0754), .ZN(new_n21257_));
  INV_X1     g18128(.I(new_n21257_), .ZN(new_n21258_));
  NAND2_X1   g18129(.A1(new_n21258_), .A2(new_n16751_), .ZN(new_n21259_));
  NAND4_X1   g18130(.A1(new_n5503_), .A2(new_n21259_), .A3(pi0181), .A4(new_n3290_), .ZN(new_n21260_));
  AOI21_X1   g18131(.A1(new_n21256_), .A2(new_n3259_), .B(new_n21260_), .ZN(new_n21261_));
  NAND2_X1   g18132(.A1(new_n21254_), .A2(new_n21261_), .ZN(new_n21262_));
  AOI21_X1   g18133(.A1(new_n21262_), .A2(new_n21105_), .B(new_n21168_), .ZN(new_n21263_));
  INV_X1     g18134(.I(new_n21119_), .ZN(new_n21264_));
  INV_X1     g18135(.I(new_n21263_), .ZN(new_n21265_));
  NAND2_X1   g18136(.A1(new_n21171_), .A2(pi0625), .ZN(new_n21266_));
  XOR2_X1    g18137(.A1(new_n21266_), .A2(new_n13615_), .Z(new_n21267_));
  OAI21_X1   g18138(.A1(new_n21265_), .A2(new_n21267_), .B(new_n14081_), .ZN(new_n21268_));
  NAND2_X1   g18139(.A1(new_n21171_), .A2(pi1153), .ZN(new_n21269_));
  XOR2_X1    g18140(.A1(new_n21269_), .A2(new_n13620_), .Z(new_n21270_));
  AOI21_X1   g18141(.A1(new_n21263_), .A2(new_n21270_), .B(pi0608), .ZN(new_n21271_));
  OAI21_X1   g18142(.A1(new_n21268_), .A2(new_n21264_), .B(new_n21271_), .ZN(new_n21272_));
  NAND4_X1   g18143(.A1(new_n21272_), .A2(pi0778), .A3(new_n21101_), .A4(new_n21114_), .ZN(new_n21273_));
  OAI21_X1   g18144(.A1(pi0778), .A2(new_n21263_), .B(new_n21273_), .ZN(new_n21274_));
  NAND2_X1   g18145(.A1(new_n21274_), .A2(new_n13801_), .ZN(new_n21275_));
  NOR2_X1    g18146(.A1(new_n21274_), .A2(new_n13778_), .ZN(new_n21276_));
  NOR2_X1    g18147(.A1(new_n21276_), .A2(new_n14694_), .ZN(new_n21277_));
  NAND2_X1   g18148(.A1(new_n21276_), .A2(new_n14694_), .ZN(new_n21278_));
  INV_X1     g18149(.I(new_n21278_), .ZN(new_n21279_));
  OAI21_X1   g18150(.A1(new_n21279_), .A2(new_n21277_), .B(new_n21121_), .ZN(new_n21280_));
  NAND2_X1   g18151(.A1(new_n21175_), .A2(pi0660), .ZN(new_n21281_));
  INV_X1     g18152(.I(new_n21281_), .ZN(new_n21282_));
  NOR2_X1    g18153(.A1(new_n21180_), .A2(pi0660), .ZN(new_n21283_));
  INV_X1     g18154(.I(new_n21283_), .ZN(new_n21284_));
  AOI21_X1   g18155(.A1(new_n21280_), .A2(new_n21282_), .B(new_n21284_), .ZN(new_n21285_));
  NOR2_X1    g18156(.A1(new_n21274_), .A2(new_n13766_), .ZN(new_n21286_));
  XOR2_X1    g18157(.A1(new_n21286_), .A2(new_n14694_), .Z(new_n21287_));
  NAND2_X1   g18158(.A1(new_n21121_), .A2(pi0785), .ZN(new_n21288_));
  NOR2_X1    g18159(.A1(new_n21287_), .A2(new_n21288_), .ZN(new_n21289_));
  INV_X1     g18160(.I(new_n21289_), .ZN(new_n21290_));
  OAI21_X1   g18161(.A1(new_n21290_), .A2(new_n21285_), .B(new_n21275_), .ZN(new_n21291_));
  NAND3_X1   g18162(.A1(new_n21291_), .A2(pi0618), .A3(pi1154), .ZN(new_n21292_));
  INV_X1     g18163(.I(new_n21277_), .ZN(new_n21293_));
  AOI21_X1   g18164(.A1(new_n21293_), .A2(new_n21278_), .B(new_n21122_), .ZN(new_n21294_));
  OAI21_X1   g18165(.A1(new_n21294_), .A2(new_n21281_), .B(new_n21283_), .ZN(new_n21295_));
  AOI22_X1   g18166(.A1(new_n21295_), .A2(new_n21289_), .B1(new_n13801_), .B2(new_n21274_), .ZN(new_n21296_));
  NAND3_X1   g18167(.A1(new_n21296_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n21297_));
  AOI21_X1   g18168(.A1(new_n21297_), .A2(new_n21292_), .B(new_n21239_), .ZN(new_n21298_));
  NOR2_X1    g18169(.A1(new_n21186_), .A2(new_n13823_), .ZN(new_n21299_));
  INV_X1     g18170(.I(new_n21299_), .ZN(new_n21300_));
  OAI21_X1   g18171(.A1(new_n21298_), .A2(new_n21300_), .B(pi0781), .ZN(new_n21301_));
  NAND3_X1   g18172(.A1(new_n21291_), .A2(pi0618), .A3(pi1154), .ZN(new_n21302_));
  NAND3_X1   g18173(.A1(new_n21296_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n21303_));
  NAND2_X1   g18174(.A1(new_n21303_), .A2(new_n21302_), .ZN(new_n21304_));
  NAND3_X1   g18175(.A1(new_n21291_), .A2(new_n19177_), .A3(new_n21192_), .ZN(new_n21305_));
  AOI21_X1   g18176(.A1(new_n21304_), .A2(new_n21124_), .B(new_n21305_), .ZN(new_n21306_));
  NAND2_X1   g18177(.A1(new_n21301_), .A2(new_n21306_), .ZN(new_n21307_));
  AOI21_X1   g18178(.A1(new_n21296_), .A2(pi1154), .B(new_n13819_), .ZN(new_n21308_));
  NOR3_X1    g18179(.A1(new_n21291_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n21309_));
  OAI21_X1   g18180(.A1(new_n21308_), .A2(new_n21309_), .B(new_n21124_), .ZN(new_n21310_));
  AOI21_X1   g18181(.A1(new_n21310_), .A2(new_n21299_), .B(new_n13855_), .ZN(new_n21311_));
  AOI21_X1   g18182(.A1(new_n21296_), .A2(pi0618), .B(new_n13819_), .ZN(new_n21312_));
  NOR3_X1    g18183(.A1(new_n21291_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n21313_));
  OAI21_X1   g18184(.A1(new_n21312_), .A2(new_n21313_), .B(new_n21124_), .ZN(new_n21314_));
  NAND4_X1   g18185(.A1(new_n21314_), .A2(new_n19177_), .A3(new_n21192_), .A4(new_n21291_), .ZN(new_n21315_));
  NAND2_X1   g18186(.A1(new_n21315_), .A2(new_n21311_), .ZN(new_n21316_));
  NAND2_X1   g18187(.A1(new_n21316_), .A2(new_n21307_), .ZN(new_n21317_));
  NAND3_X1   g18188(.A1(new_n21317_), .A2(pi0619), .A3(pi1159), .ZN(new_n21318_));
  NOR2_X1    g18189(.A1(new_n21315_), .A2(new_n21311_), .ZN(new_n21319_));
  NOR2_X1    g18190(.A1(new_n21301_), .A2(new_n21306_), .ZN(new_n21320_));
  NOR2_X1    g18191(.A1(new_n21319_), .A2(new_n21320_), .ZN(new_n21321_));
  NAND3_X1   g18192(.A1(new_n21321_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n21322_));
  AOI21_X1   g18193(.A1(new_n21322_), .A2(new_n21318_), .B(new_n21126_), .ZN(new_n21323_));
  OAI21_X1   g18194(.A1(new_n21323_), .A2(new_n20003_), .B(new_n21199_), .ZN(new_n21324_));
  NAND2_X1   g18195(.A1(new_n21317_), .A2(new_n13896_), .ZN(new_n21325_));
  NAND3_X1   g18196(.A1(new_n21209_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n21326_));
  INV_X1     g18197(.I(new_n21209_), .ZN(new_n21327_));
  NAND3_X1   g18198(.A1(new_n21327_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n21328_));
  AOI21_X1   g18199(.A1(new_n21328_), .A2(new_n21326_), .B(new_n21102_), .ZN(new_n21329_));
  NOR2_X1    g18200(.A1(new_n21127_), .A2(new_n14162_), .ZN(new_n21330_));
  OAI21_X1   g18201(.A1(new_n21329_), .A2(new_n21330_), .B(new_n19204_), .ZN(new_n21331_));
  NOR2_X1    g18202(.A1(new_n21209_), .A2(new_n19208_), .ZN(new_n21332_));
  XNOR2_X1   g18203(.A1(new_n21332_), .A2(new_n19028_), .ZN(new_n21333_));
  NOR2_X1    g18204(.A1(new_n21102_), .A2(new_n15479_), .ZN(new_n21334_));
  NAND4_X1   g18205(.A1(new_n21331_), .A2(new_n21325_), .A3(new_n21333_), .A4(new_n21334_), .ZN(new_n21335_));
  INV_X1     g18206(.I(new_n21126_), .ZN(new_n21336_));
  AOI21_X1   g18207(.A1(new_n21321_), .A2(pi0619), .B(new_n13904_), .ZN(new_n21337_));
  NOR4_X1    g18208(.A1(new_n21319_), .A2(new_n21320_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n21338_));
  OAI21_X1   g18209(.A1(new_n21337_), .A2(new_n21338_), .B(new_n21336_), .ZN(new_n21339_));
  NAND3_X1   g18210(.A1(new_n21339_), .A2(new_n20173_), .A3(new_n21206_), .ZN(new_n21340_));
  AOI21_X1   g18211(.A1(new_n21324_), .A2(new_n21335_), .B(new_n21340_), .ZN(new_n21341_));
  AND2_X2    g18212(.A1(new_n21133_), .A2(pi0629), .Z(new_n21342_));
  NOR2_X1    g18213(.A1(new_n21153_), .A2(pi0629), .ZN(new_n21343_));
  NOR2_X1    g18214(.A1(new_n9992_), .A2(pi0181), .ZN(new_n21344_));
  NOR3_X1    g18215(.A1(new_n13219_), .A2(pi0625), .A3(pi0709), .ZN(new_n21345_));
  INV_X1     g18216(.I(new_n21345_), .ZN(new_n21346_));
  NOR2_X1    g18217(.A1(new_n21344_), .A2(pi1153), .ZN(new_n21347_));
  NAND2_X1   g18218(.A1(new_n21346_), .A2(new_n21347_), .ZN(new_n21348_));
  INV_X1     g18219(.I(new_n21348_), .ZN(new_n21349_));
  NOR2_X1    g18220(.A1(new_n21349_), .A2(new_n13748_), .ZN(new_n21350_));
  AOI21_X1   g18221(.A1(new_n13218_), .A2(new_n21105_), .B(new_n21344_), .ZN(new_n21351_));
  INV_X1     g18222(.I(new_n21351_), .ZN(new_n21352_));
  AOI21_X1   g18223(.A1(new_n21346_), .A2(new_n21352_), .B(new_n13614_), .ZN(new_n21353_));
  INV_X1     g18224(.I(new_n21353_), .ZN(new_n21354_));
  NOR3_X1    g18225(.A1(new_n21354_), .A2(new_n13748_), .A3(new_n21352_), .ZN(new_n21355_));
  XNOR2_X1   g18226(.A1(new_n21355_), .A2(new_n21350_), .ZN(new_n21356_));
  NAND2_X1   g18227(.A1(new_n21356_), .A2(new_n14049_), .ZN(new_n21357_));
  NOR2_X1    g18228(.A1(new_n21357_), .A2(new_n14051_), .ZN(new_n21358_));
  INV_X1     g18229(.I(new_n21358_), .ZN(new_n21359_));
  NOR2_X1    g18230(.A1(new_n21359_), .A2(new_n14163_), .ZN(new_n21360_));
  NOR2_X1    g18231(.A1(new_n21257_), .A2(new_n21344_), .ZN(new_n21361_));
  INV_X1     g18232(.I(new_n21361_), .ZN(new_n21362_));
  NAND3_X1   g18233(.A1(new_n21362_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n21363_));
  AOI21_X1   g18234(.A1(new_n21363_), .A2(new_n16444_), .B(new_n21258_), .ZN(new_n21364_));
  NOR2_X1    g18235(.A1(new_n21364_), .A2(new_n13801_), .ZN(new_n21365_));
  NOR2_X1    g18236(.A1(new_n21344_), .A2(pi1155), .ZN(new_n21366_));
  NOR3_X1    g18237(.A1(new_n21258_), .A2(new_n16444_), .A3(new_n21366_), .ZN(new_n21367_));
  NAND4_X1   g18238(.A1(new_n21367_), .A2(new_n21362_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n21368_));
  XOR2_X1    g18239(.A1(new_n21365_), .A2(new_n21368_), .Z(new_n21369_));
  NOR2_X1    g18240(.A1(new_n21369_), .A2(new_n13817_), .ZN(new_n21370_));
  OAI21_X1   g18241(.A1(new_n21370_), .A2(pi0618), .B(new_n9992_), .ZN(new_n21371_));
  NAND2_X1   g18242(.A1(new_n21371_), .A2(pi0781), .ZN(new_n21372_));
  OAI21_X1   g18243(.A1(new_n21370_), .A2(new_n9992_), .B(pi0618), .ZN(new_n21373_));
  NOR3_X1    g18244(.A1(new_n21373_), .A2(new_n13855_), .A3(new_n21369_), .ZN(new_n21374_));
  XOR2_X1    g18245(.A1(new_n21374_), .A2(new_n21372_), .Z(new_n21375_));
  NOR2_X1    g18246(.A1(new_n21375_), .A2(new_n13868_), .ZN(new_n21376_));
  OAI21_X1   g18247(.A1(new_n21376_), .A2(pi0619), .B(new_n9992_), .ZN(new_n21377_));
  NAND2_X1   g18248(.A1(new_n21377_), .A2(pi0789), .ZN(new_n21378_));
  OAI21_X1   g18249(.A1(new_n21376_), .A2(new_n9992_), .B(pi0619), .ZN(new_n21379_));
  NOR3_X1    g18250(.A1(new_n21379_), .A2(new_n13896_), .A3(new_n21375_), .ZN(new_n21380_));
  XOR2_X1    g18251(.A1(new_n21380_), .A2(new_n21378_), .Z(new_n21381_));
  NAND2_X1   g18252(.A1(new_n21381_), .A2(new_n13962_), .ZN(new_n21382_));
  XOR2_X1    g18253(.A1(new_n21382_), .A2(new_n18976_), .Z(new_n21383_));
  AOI22_X1   g18254(.A1(new_n21383_), .A2(new_n21344_), .B1(new_n16639_), .B2(new_n21360_), .ZN(new_n21384_));
  NOR2_X1    g18255(.A1(new_n21351_), .A2(new_n13203_), .ZN(new_n21385_));
  NAND2_X1   g18256(.A1(new_n21385_), .A2(pi0625), .ZN(new_n21386_));
  NAND3_X1   g18257(.A1(new_n21386_), .A2(pi1153), .A3(new_n21361_), .ZN(new_n21387_));
  NOR2_X1    g18258(.A1(new_n21349_), .A2(new_n14081_), .ZN(new_n21388_));
  AOI21_X1   g18259(.A1(new_n21388_), .A2(new_n21387_), .B(new_n13748_), .ZN(new_n21389_));
  NOR2_X1    g18260(.A1(new_n21362_), .A2(new_n21385_), .ZN(new_n21390_));
  INV_X1     g18261(.I(new_n21386_), .ZN(new_n21391_));
  OAI21_X1   g18262(.A1(new_n21390_), .A2(new_n21391_), .B(new_n21347_), .ZN(new_n21392_));
  NAND4_X1   g18263(.A1(new_n21392_), .A2(new_n13749_), .A3(new_n21354_), .A4(new_n21390_), .ZN(new_n21393_));
  XNOR2_X1   g18264(.A1(new_n21393_), .A2(new_n21389_), .ZN(new_n21394_));
  NAND2_X1   g18265(.A1(new_n21394_), .A2(new_n13801_), .ZN(new_n21395_));
  NOR2_X1    g18266(.A1(new_n21364_), .A2(pi0660), .ZN(new_n21399_));
  NOR2_X1    g18267(.A1(new_n21394_), .A2(new_n13766_), .ZN(new_n21400_));
  XOR2_X1    g18268(.A1(new_n21400_), .A2(new_n14090_), .Z(new_n21401_));
  NOR2_X1    g18269(.A1(new_n21356_), .A2(new_n13801_), .ZN(new_n21402_));
  NAND2_X1   g18270(.A1(new_n21401_), .A2(new_n21402_), .ZN(new_n21403_));
  OAI21_X1   g18271(.A1(new_n21403_), .A2(new_n21399_), .B(new_n21395_), .ZN(new_n21404_));
  NAND2_X1   g18272(.A1(new_n21404_), .A2(new_n13855_), .ZN(new_n21405_));
  INV_X1     g18273(.I(new_n21357_), .ZN(new_n21406_));
  NOR2_X1    g18274(.A1(new_n21404_), .A2(new_n13816_), .ZN(new_n21407_));
  XOR2_X1    g18275(.A1(new_n21407_), .A2(new_n13818_), .Z(new_n21408_));
  NAND2_X1   g18276(.A1(new_n21408_), .A2(new_n21406_), .ZN(new_n21409_));
  NAND3_X1   g18277(.A1(new_n21409_), .A2(new_n13823_), .A3(new_n21373_), .ZN(new_n21410_));
  NAND3_X1   g18278(.A1(new_n21410_), .A2(new_n13823_), .A3(new_n21371_), .ZN(new_n21411_));
  NOR2_X1    g18279(.A1(new_n21404_), .A2(new_n13817_), .ZN(new_n21412_));
  XOR2_X1    g18280(.A1(new_n21412_), .A2(new_n13818_), .Z(new_n21413_));
  NAND4_X1   g18281(.A1(new_n21411_), .A2(pi0781), .A3(new_n21406_), .A4(new_n21413_), .ZN(new_n21414_));
  NAND2_X1   g18282(.A1(new_n21414_), .A2(new_n21405_), .ZN(new_n21415_));
  NOR2_X1    g18283(.A1(new_n21415_), .A2(new_n13860_), .ZN(new_n21416_));
  XOR2_X1    g18284(.A1(new_n21416_), .A2(new_n13904_), .Z(new_n21417_));
  NOR2_X1    g18285(.A1(new_n21417_), .A2(new_n21359_), .ZN(new_n21418_));
  NAND2_X1   g18286(.A1(new_n21379_), .A2(new_n13884_), .ZN(new_n21419_));
  INV_X1     g18287(.I(new_n21415_), .ZN(new_n21420_));
  AOI21_X1   g18288(.A1(new_n21420_), .A2(new_n14143_), .B(pi0789), .ZN(new_n21421_));
  OAI21_X1   g18289(.A1(new_n21418_), .A2(new_n21419_), .B(new_n21421_), .ZN(new_n21422_));
  NOR2_X1    g18290(.A1(new_n21415_), .A2(new_n13868_), .ZN(new_n21423_));
  XOR2_X1    g18291(.A1(new_n21423_), .A2(new_n13903_), .Z(new_n21424_));
  NAND2_X1   g18292(.A1(new_n21377_), .A2(new_n19018_), .ZN(new_n21425_));
  AOI21_X1   g18293(.A1(new_n21424_), .A2(new_n21358_), .B(new_n21425_), .ZN(new_n21426_));
  AOI21_X1   g18294(.A1(new_n21422_), .A2(new_n21426_), .B(new_n21384_), .ZN(new_n21427_));
  NOR3_X1    g18295(.A1(new_n21359_), .A2(new_n14163_), .A3(new_n18928_), .ZN(new_n21428_));
  NAND2_X1   g18296(.A1(new_n21381_), .A2(new_n16372_), .ZN(new_n21429_));
  OAI21_X1   g18297(.A1(new_n16372_), .A2(new_n21344_), .B(new_n21429_), .ZN(new_n21430_));
  NAND2_X1   g18298(.A1(new_n21430_), .A2(new_n21428_), .ZN(new_n21431_));
  NAND2_X1   g18299(.A1(new_n21431_), .A2(new_n19022_), .ZN(new_n21432_));
  NAND2_X1   g18300(.A1(new_n21431_), .A2(new_n16569_), .ZN(new_n21433_));
  XNOR2_X1   g18301(.A1(new_n21433_), .A2(new_n16572_), .ZN(new_n21434_));
  AOI21_X1   g18302(.A1(new_n21434_), .A2(new_n21432_), .B(new_n16574_), .ZN(new_n21435_));
  NAND2_X1   g18303(.A1(new_n21381_), .A2(new_n13963_), .ZN(new_n21436_));
  XNOR2_X1   g18304(.A1(new_n21436_), .A2(new_n19028_), .ZN(new_n21437_));
  NAND2_X1   g18305(.A1(new_n16423_), .A2(new_n21344_), .ZN(new_n21438_));
  NOR4_X1    g18306(.A1(new_n21427_), .A2(new_n21435_), .A3(new_n21437_), .A4(new_n21438_), .ZN(new_n21439_));
  INV_X1     g18307(.I(new_n21344_), .ZN(new_n21440_));
  NAND2_X1   g18308(.A1(new_n21428_), .A2(new_n14061_), .ZN(new_n21441_));
  NAND2_X1   g18309(.A1(new_n21344_), .A2(new_n14005_), .ZN(new_n21442_));
  OAI21_X1   g18310(.A1(new_n21441_), .A2(new_n14005_), .B(new_n21442_), .ZN(new_n21443_));
  NOR2_X1    g18311(.A1(new_n21430_), .A2(new_n13994_), .ZN(new_n21444_));
  XOR2_X1    g18312(.A1(new_n21444_), .A2(new_n19033_), .Z(new_n21445_));
  OAI22_X1   g18313(.A1(new_n21445_), .A2(new_n21440_), .B1(new_n14207_), .B2(new_n21443_), .ZN(new_n21446_));
  NAND2_X1   g18314(.A1(new_n21441_), .A2(pi0647), .ZN(new_n21447_));
  XOR2_X1    g18315(.A1(new_n21447_), .A2(new_n14007_), .Z(new_n21448_));
  NOR3_X1    g18316(.A1(new_n21448_), .A2(new_n14010_), .A3(new_n21440_), .ZN(new_n21449_));
  AOI21_X1   g18317(.A1(new_n21446_), .A2(new_n21449_), .B(new_n12776_), .ZN(new_n21450_));
  NOR2_X1    g18318(.A1(new_n21439_), .A2(new_n21450_), .ZN(new_n21451_));
  NOR2_X1    g18319(.A1(new_n21448_), .A2(new_n21440_), .ZN(new_n21452_));
  OAI21_X1   g18320(.A1(new_n21443_), .A2(new_n14006_), .B(pi0787), .ZN(new_n21453_));
  OAI22_X1   g18321(.A1(new_n21452_), .A2(new_n21453_), .B1(pi0787), .B2(new_n21441_), .ZN(new_n21454_));
  NOR2_X1    g18322(.A1(new_n21451_), .A2(new_n14204_), .ZN(new_n21455_));
  XOR2_X1    g18323(.A1(new_n21455_), .A2(new_n14205_), .Z(new_n21456_));
  NAND2_X1   g18324(.A1(new_n21456_), .A2(new_n21454_), .ZN(new_n21457_));
  NOR2_X1    g18325(.A1(new_n21430_), .A2(new_n18968_), .ZN(new_n21458_));
  NAND2_X1   g18326(.A1(new_n18967_), .A2(new_n21344_), .ZN(new_n21459_));
  XOR2_X1    g18327(.A1(new_n21458_), .A2(new_n21459_), .Z(new_n21460_));
  NAND2_X1   g18328(.A1(new_n21460_), .A2(pi0715), .ZN(new_n21461_));
  XOR2_X1    g18329(.A1(new_n21461_), .A2(new_n14217_), .Z(new_n21462_));
  AOI21_X1   g18330(.A1(new_n21462_), .A2(new_n21344_), .B(pi1160), .ZN(new_n21463_));
  NAND2_X1   g18331(.A1(new_n21460_), .A2(pi0644), .ZN(new_n21464_));
  XOR2_X1    g18332(.A1(new_n21464_), .A2(new_n14205_), .Z(new_n21465_));
  OAI21_X1   g18333(.A1(new_n21465_), .A2(new_n21440_), .B(new_n14203_), .ZN(new_n21466_));
  AOI21_X1   g18334(.A1(new_n21457_), .A2(new_n21463_), .B(new_n21466_), .ZN(new_n21467_));
  NOR2_X1    g18335(.A1(new_n21451_), .A2(new_n14200_), .ZN(new_n21468_));
  XOR2_X1    g18336(.A1(new_n21468_), .A2(new_n14205_), .Z(new_n21469_));
  NAND2_X1   g18337(.A1(new_n21469_), .A2(new_n21454_), .ZN(new_n21470_));
  OAI21_X1   g18338(.A1(new_n21467_), .A2(new_n21470_), .B(pi0832), .ZN(new_n21471_));
  XOR2_X1    g18339(.A1(new_n21471_), .A2(new_n14801_), .Z(new_n21472_));
  NAND2_X1   g18340(.A1(po1038), .A2(new_n5643_), .ZN(new_n21473_));
  NAND4_X1   g18341(.A1(new_n21472_), .A2(new_n14799_), .A3(new_n21451_), .A4(new_n21473_), .ZN(new_n21474_));
  NAND2_X1   g18342(.A1(new_n21474_), .A2(new_n7240_), .ZN(new_n21475_));
  OAI21_X1   g18343(.A1(new_n21342_), .A2(new_n21343_), .B(new_n21475_), .ZN(new_n21476_));
  AOI21_X1   g18344(.A1(new_n16875_), .A2(new_n21210_), .B(new_n21476_), .ZN(new_n21477_));
  OAI21_X1   g18345(.A1(new_n21341_), .A2(pi0792), .B(new_n21477_), .ZN(new_n21478_));
  AOI21_X1   g18346(.A1(new_n21238_), .A2(new_n21226_), .B(new_n21478_), .ZN(po0338));
  NAND2_X1   g18347(.A1(new_n13627_), .A2(new_n5644_), .ZN(new_n21480_));
  INV_X1     g18348(.I(new_n21480_), .ZN(new_n21481_));
  AOI21_X1   g18349(.A1(new_n5644_), .A2(new_n17609_), .B(pi0038), .ZN(new_n21482_));
  NOR2_X1    g18350(.A1(new_n5644_), .A2(new_n17609_), .ZN(new_n21483_));
  OAI21_X1   g18351(.A1(new_n20007_), .A2(new_n21483_), .B(pi0038), .ZN(new_n21484_));
  INV_X1     g18352(.I(new_n21484_), .ZN(new_n21485_));
  AOI21_X1   g18353(.A1(new_n13097_), .A2(new_n21482_), .B(new_n21485_), .ZN(new_n21486_));
  NOR2_X1    g18354(.A1(new_n3289_), .A2(pi0182), .ZN(new_n21487_));
  AOI21_X1   g18355(.A1(new_n21486_), .A2(new_n3289_), .B(new_n21487_), .ZN(new_n21488_));
  NAND2_X1   g18356(.A1(new_n21488_), .A2(new_n13776_), .ZN(new_n21489_));
  OAI21_X1   g18357(.A1(new_n15147_), .A2(new_n21481_), .B(new_n21489_), .ZN(new_n21490_));
  NAND2_X1   g18358(.A1(new_n21490_), .A2(pi0609), .ZN(new_n21491_));
  NAND2_X1   g18359(.A1(new_n21491_), .A2(pi0785), .ZN(new_n21492_));
  AOI21_X1   g18360(.A1(new_n21480_), .A2(new_n14467_), .B(pi0609), .ZN(new_n21493_));
  NOR2_X1    g18361(.A1(new_n21493_), .A2(new_n21489_), .ZN(new_n21494_));
  NAND2_X1   g18362(.A1(new_n21481_), .A2(new_n13775_), .ZN(new_n21495_));
  OAI21_X1   g18363(.A1(new_n13775_), .A2(new_n21488_), .B(new_n21495_), .ZN(new_n21496_));
  NAND3_X1   g18364(.A1(new_n21496_), .A2(pi0785), .A3(new_n21494_), .ZN(new_n21497_));
  XNOR2_X1   g18365(.A1(new_n21492_), .A2(new_n21497_), .ZN(new_n21498_));
  NAND2_X1   g18366(.A1(new_n21498_), .A2(pi0618), .ZN(new_n21499_));
  XOR2_X1    g18367(.A1(new_n21499_), .A2(new_n13819_), .Z(new_n21500_));
  NAND2_X1   g18368(.A1(new_n21500_), .A2(new_n21481_), .ZN(new_n21501_));
  NAND2_X1   g18369(.A1(new_n21501_), .A2(pi0781), .ZN(new_n21502_));
  NAND2_X1   g18370(.A1(new_n21498_), .A2(pi1154), .ZN(new_n21503_));
  XOR2_X1    g18371(.A1(new_n21503_), .A2(new_n13819_), .Z(new_n21504_));
  NAND2_X1   g18372(.A1(new_n21504_), .A2(new_n21481_), .ZN(new_n21505_));
  NOR3_X1    g18373(.A1(new_n21505_), .A2(new_n13855_), .A3(new_n21498_), .ZN(new_n21506_));
  XNOR2_X1   g18374(.A1(new_n21506_), .A2(new_n21502_), .ZN(new_n21507_));
  NAND3_X1   g18375(.A1(new_n21507_), .A2(pi0619), .A3(pi1159), .ZN(new_n21508_));
  XOR2_X1    g18376(.A1(new_n21506_), .A2(new_n21502_), .Z(new_n21509_));
  NAND3_X1   g18377(.A1(new_n21509_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n21510_));
  AOI21_X1   g18378(.A1(new_n21508_), .A2(new_n21510_), .B(new_n21480_), .ZN(new_n21511_));
  NOR2_X1    g18379(.A1(new_n21481_), .A2(new_n13880_), .ZN(new_n21512_));
  OAI21_X1   g18380(.A1(new_n13721_), .A2(new_n17604_), .B(new_n5644_), .ZN(new_n21513_));
  NAND2_X1   g18381(.A1(new_n16715_), .A2(new_n5644_), .ZN(new_n21514_));
  NAND4_X1   g18382(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n21513_), .A4(new_n21514_), .ZN(new_n21515_));
  NAND2_X1   g18383(.A1(new_n21515_), .A2(new_n14424_), .ZN(new_n21516_));
  NAND2_X1   g18384(.A1(new_n21516_), .A2(pi0182), .ZN(new_n21517_));
  OAI21_X1   g18385(.A1(new_n21517_), .A2(new_n21480_), .B(new_n3290_), .ZN(new_n21518_));
  NAND2_X1   g18386(.A1(new_n21518_), .A2(pi0734), .ZN(new_n21519_));
  NAND2_X1   g18387(.A1(new_n21519_), .A2(pi0625), .ZN(new_n21520_));
  XOR2_X1    g18388(.A1(new_n21520_), .A2(new_n13620_), .Z(new_n21521_));
  NAND2_X1   g18389(.A1(new_n21521_), .A2(new_n21481_), .ZN(new_n21522_));
  NAND2_X1   g18390(.A1(new_n21522_), .A2(pi0778), .ZN(new_n21523_));
  NAND2_X1   g18391(.A1(new_n21519_), .A2(pi1153), .ZN(new_n21524_));
  XOR2_X1    g18392(.A1(new_n21524_), .A2(new_n13620_), .Z(new_n21525_));
  NAND2_X1   g18393(.A1(new_n21525_), .A2(new_n21481_), .ZN(new_n21526_));
  NOR3_X1    g18394(.A1(new_n21526_), .A2(new_n13748_), .A3(new_n21519_), .ZN(new_n21527_));
  XNOR2_X1   g18395(.A1(new_n21527_), .A2(new_n21523_), .ZN(new_n21528_));
  NOR2_X1    g18396(.A1(new_n21480_), .A2(new_n13805_), .ZN(new_n21529_));
  AOI21_X1   g18397(.A1(new_n21528_), .A2(new_n13805_), .B(new_n21529_), .ZN(new_n21530_));
  AOI21_X1   g18398(.A1(new_n21530_), .A2(new_n13880_), .B(new_n21512_), .ZN(new_n21531_));
  NOR2_X1    g18399(.A1(new_n13453_), .A2(new_n5644_), .ZN(new_n21532_));
  XOR2_X1    g18400(.A1(new_n21532_), .A2(new_n21483_), .Z(new_n21533_));
  NAND2_X1   g18401(.A1(new_n21533_), .A2(new_n13521_), .ZN(new_n21534_));
  NAND3_X1   g18402(.A1(new_n14270_), .A2(pi0182), .A3(pi0756), .ZN(new_n21535_));
  NAND3_X1   g18403(.A1(new_n14272_), .A2(new_n5644_), .A3(pi0756), .ZN(new_n21536_));
  AOI21_X1   g18404(.A1(new_n21535_), .A2(new_n21536_), .B(new_n13152_), .ZN(new_n21537_));
  NAND3_X1   g18405(.A1(new_n13198_), .A2(pi0182), .A3(pi0756), .ZN(new_n21538_));
  NAND3_X1   g18406(.A1(new_n13200_), .A2(pi0182), .A3(new_n17609_), .ZN(new_n21539_));
  AOI21_X1   g18407(.A1(new_n21539_), .A2(new_n21538_), .B(new_n13191_), .ZN(new_n21540_));
  OAI21_X1   g18408(.A1(new_n21537_), .A2(new_n3262_), .B(new_n21540_), .ZN(new_n21541_));
  NAND3_X1   g18409(.A1(new_n21534_), .A2(new_n3183_), .A3(new_n21541_), .ZN(new_n21542_));
  NOR2_X1    g18410(.A1(new_n14284_), .A2(new_n17609_), .ZN(new_n21543_));
  XOR2_X1    g18411(.A1(new_n21543_), .A2(new_n21483_), .Z(new_n21544_));
  NAND3_X1   g18412(.A1(new_n21542_), .A2(new_n21544_), .A3(new_n13359_), .ZN(new_n21545_));
  NAND3_X1   g18413(.A1(new_n21545_), .A2(new_n17604_), .A3(new_n3290_), .ZN(new_n21546_));
  OAI21_X1   g18414(.A1(new_n15587_), .A2(new_n5644_), .B(new_n17609_), .ZN(new_n21547_));
  NAND2_X1   g18415(.A1(new_n21547_), .A2(new_n13209_), .ZN(new_n21548_));
  NOR2_X1    g18416(.A1(new_n13105_), .A2(pi0756), .ZN(new_n21549_));
  INV_X1     g18417(.I(new_n21549_), .ZN(new_n21550_));
  NAND2_X1   g18418(.A1(new_n21550_), .A2(new_n16751_), .ZN(new_n21551_));
  NAND4_X1   g18419(.A1(new_n5503_), .A2(new_n21551_), .A3(pi0182), .A4(new_n3290_), .ZN(new_n21552_));
  AOI21_X1   g18420(.A1(new_n21548_), .A2(new_n3259_), .B(new_n21552_), .ZN(new_n21553_));
  AOI21_X1   g18421(.A1(new_n21546_), .A2(new_n21553_), .B(pi0734), .ZN(new_n21554_));
  NOR2_X1    g18422(.A1(new_n21554_), .A2(new_n21486_), .ZN(new_n21555_));
  INV_X1     g18423(.I(new_n21555_), .ZN(new_n21556_));
  INV_X1     g18424(.I(new_n21488_), .ZN(new_n21557_));
  NOR2_X1    g18425(.A1(new_n21555_), .A2(new_n13613_), .ZN(new_n21558_));
  XOR2_X1    g18426(.A1(new_n21558_), .A2(new_n13615_), .Z(new_n21559_));
  NAND2_X1   g18427(.A1(new_n21526_), .A2(new_n14081_), .ZN(new_n21560_));
  AOI21_X1   g18428(.A1(new_n21559_), .A2(new_n21557_), .B(new_n21560_), .ZN(new_n21561_));
  INV_X1     g18429(.I(new_n21561_), .ZN(new_n21562_));
  NOR2_X1    g18430(.A1(new_n21555_), .A2(new_n13614_), .ZN(new_n21563_));
  XOR2_X1    g18431(.A1(new_n21563_), .A2(new_n13615_), .Z(new_n21564_));
  AOI21_X1   g18432(.A1(new_n21564_), .A2(new_n21557_), .B(pi0608), .ZN(new_n21565_));
  NAND2_X1   g18433(.A1(new_n21562_), .A2(new_n21565_), .ZN(new_n21566_));
  NOR2_X1    g18434(.A1(new_n21522_), .A2(new_n13748_), .ZN(new_n21567_));
  AOI22_X1   g18435(.A1(new_n21566_), .A2(new_n21567_), .B1(new_n13748_), .B2(new_n21556_), .ZN(new_n21568_));
  AOI21_X1   g18436(.A1(new_n21568_), .A2(pi1155), .B(new_n14694_), .ZN(new_n21569_));
  INV_X1     g18437(.I(new_n21565_), .ZN(new_n21570_));
  NOR2_X1    g18438(.A1(new_n21570_), .A2(new_n21561_), .ZN(new_n21571_));
  INV_X1     g18439(.I(new_n21567_), .ZN(new_n21572_));
  OAI22_X1   g18440(.A1(new_n21571_), .A2(new_n21572_), .B1(pi0778), .B2(new_n21555_), .ZN(new_n21573_));
  NOR3_X1    g18441(.A1(new_n21573_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n21574_));
  OAI21_X1   g18442(.A1(new_n21574_), .A2(new_n21569_), .B(new_n21528_), .ZN(new_n21575_));
  NAND2_X1   g18443(.A1(new_n21491_), .A2(pi0660), .ZN(new_n21576_));
  INV_X1     g18444(.I(new_n21576_), .ZN(new_n21577_));
  NOR2_X1    g18445(.A1(new_n21494_), .A2(pi0660), .ZN(new_n21578_));
  INV_X1     g18446(.I(new_n21578_), .ZN(new_n21579_));
  AOI21_X1   g18447(.A1(new_n21575_), .A2(new_n21577_), .B(new_n21579_), .ZN(new_n21580_));
  NOR2_X1    g18448(.A1(new_n21573_), .A2(new_n13766_), .ZN(new_n21581_));
  NOR2_X1    g18449(.A1(new_n21581_), .A2(new_n14694_), .ZN(new_n21582_));
  NAND2_X1   g18450(.A1(new_n21581_), .A2(new_n14694_), .ZN(new_n21583_));
  INV_X1     g18451(.I(new_n21583_), .ZN(new_n21584_));
  INV_X1     g18452(.I(new_n21528_), .ZN(new_n21585_));
  NOR2_X1    g18453(.A1(new_n21585_), .A2(new_n13801_), .ZN(new_n21586_));
  OAI21_X1   g18454(.A1(new_n21584_), .A2(new_n21582_), .B(new_n21586_), .ZN(new_n21587_));
  OAI22_X1   g18455(.A1(new_n21587_), .A2(new_n21580_), .B1(pi0785), .B2(new_n21568_), .ZN(new_n21588_));
  NAND3_X1   g18456(.A1(new_n21588_), .A2(pi0618), .A3(pi1154), .ZN(new_n21589_));
  NAND3_X1   g18457(.A1(new_n21573_), .A2(pi0609), .A3(pi1155), .ZN(new_n21590_));
  NAND3_X1   g18458(.A1(new_n21568_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n21591_));
  AOI21_X1   g18459(.A1(new_n21590_), .A2(new_n21591_), .B(new_n21585_), .ZN(new_n21592_));
  OAI21_X1   g18460(.A1(new_n21592_), .A2(new_n21576_), .B(new_n21578_), .ZN(new_n21593_));
  NAND2_X1   g18461(.A1(new_n21568_), .A2(pi0609), .ZN(new_n21594_));
  NAND2_X1   g18462(.A1(new_n21594_), .A2(new_n14090_), .ZN(new_n21595_));
  INV_X1     g18463(.I(new_n21586_), .ZN(new_n21596_));
  AOI21_X1   g18464(.A1(new_n21583_), .A2(new_n21595_), .B(new_n21596_), .ZN(new_n21597_));
  AOI22_X1   g18465(.A1(new_n21593_), .A2(new_n21597_), .B1(new_n13801_), .B2(new_n21573_), .ZN(new_n21598_));
  NAND3_X1   g18466(.A1(new_n21598_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n21599_));
  AOI21_X1   g18467(.A1(new_n21589_), .A2(new_n21599_), .B(new_n21530_), .ZN(new_n21600_));
  NAND2_X1   g18468(.A1(new_n21501_), .A2(pi0627), .ZN(new_n21601_));
  OAI21_X1   g18469(.A1(new_n21600_), .A2(new_n21601_), .B(pi0781), .ZN(new_n21602_));
  INV_X1     g18470(.I(new_n21530_), .ZN(new_n21603_));
  AOI21_X1   g18471(.A1(new_n21598_), .A2(pi0618), .B(new_n13819_), .ZN(new_n21604_));
  NOR3_X1    g18472(.A1(new_n21588_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n21605_));
  OAI21_X1   g18473(.A1(new_n21605_), .A2(new_n21604_), .B(new_n21603_), .ZN(new_n21606_));
  AND3_X2    g18474(.A1(new_n21588_), .A2(new_n19177_), .A3(new_n21505_), .Z(new_n21607_));
  NAND3_X1   g18475(.A1(new_n21602_), .A2(new_n21606_), .A3(new_n21607_), .ZN(new_n21608_));
  AOI21_X1   g18476(.A1(new_n21598_), .A2(pi1154), .B(new_n13819_), .ZN(new_n21609_));
  NOR3_X1    g18477(.A1(new_n21588_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n21610_));
  OAI21_X1   g18478(.A1(new_n21610_), .A2(new_n21609_), .B(new_n21603_), .ZN(new_n21611_));
  INV_X1     g18479(.I(new_n21601_), .ZN(new_n21612_));
  AOI21_X1   g18480(.A1(new_n21611_), .A2(new_n21612_), .B(new_n13855_), .ZN(new_n21613_));
  NAND4_X1   g18481(.A1(new_n21606_), .A2(new_n19177_), .A3(new_n21505_), .A4(new_n21588_), .ZN(new_n21614_));
  NAND2_X1   g18482(.A1(new_n21614_), .A2(new_n21613_), .ZN(new_n21615_));
  NAND2_X1   g18483(.A1(new_n21615_), .A2(new_n21608_), .ZN(new_n21616_));
  NAND3_X1   g18484(.A1(new_n21616_), .A2(pi0619), .A3(pi1159), .ZN(new_n21617_));
  NAND4_X1   g18485(.A1(new_n21615_), .A2(new_n21608_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n21618_));
  AOI21_X1   g18486(.A1(new_n21617_), .A2(new_n21618_), .B(new_n21531_), .ZN(new_n21619_));
  OAI21_X1   g18487(.A1(new_n21619_), .A2(new_n20003_), .B(new_n21511_), .ZN(new_n21620_));
  NAND2_X1   g18488(.A1(new_n21616_), .A2(new_n13896_), .ZN(new_n21621_));
  NOR2_X1    g18489(.A1(new_n21511_), .A2(new_n13896_), .ZN(new_n21622_));
  NAND3_X1   g18490(.A1(new_n21507_), .A2(pi0619), .A3(pi1159), .ZN(new_n21623_));
  NAND3_X1   g18491(.A1(new_n21509_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n21624_));
  NAND2_X1   g18492(.A1(new_n21623_), .A2(new_n21624_), .ZN(new_n21625_));
  NAND4_X1   g18493(.A1(new_n21625_), .A2(pi0789), .A3(new_n21481_), .A4(new_n21507_), .ZN(new_n21626_));
  OR2_X2     g18494(.A1(new_n21626_), .A2(new_n21622_), .Z(new_n21627_));
  NAND2_X1   g18495(.A1(new_n21626_), .A2(new_n21622_), .ZN(new_n21628_));
  NAND2_X1   g18496(.A1(new_n21627_), .A2(new_n21628_), .ZN(new_n21629_));
  NAND3_X1   g18497(.A1(new_n21629_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n21630_));
  NAND4_X1   g18498(.A1(new_n21627_), .A2(new_n13901_), .A3(new_n13962_), .A4(new_n21628_), .ZN(new_n21631_));
  AOI21_X1   g18499(.A1(new_n21630_), .A2(new_n21631_), .B(new_n21480_), .ZN(new_n21632_));
  NOR2_X1    g18500(.A1(new_n21480_), .A2(new_n13919_), .ZN(new_n21633_));
  NAND2_X1   g18501(.A1(new_n21531_), .A2(new_n13919_), .ZN(new_n21634_));
  INV_X1     g18502(.I(new_n21634_), .ZN(new_n21635_));
  NOR2_X1    g18503(.A1(new_n21635_), .A2(new_n21633_), .ZN(new_n21636_));
  NOR2_X1    g18504(.A1(new_n21636_), .A2(new_n14162_), .ZN(new_n21637_));
  OAI21_X1   g18505(.A1(new_n21632_), .A2(new_n21637_), .B(new_n19204_), .ZN(new_n21638_));
  NOR2_X1    g18506(.A1(new_n21629_), .A2(new_n19208_), .ZN(new_n21639_));
  XNOR2_X1   g18507(.A1(new_n21639_), .A2(new_n19028_), .ZN(new_n21640_));
  NOR2_X1    g18508(.A1(new_n21480_), .A2(new_n15479_), .ZN(new_n21641_));
  NAND4_X1   g18509(.A1(new_n21621_), .A2(new_n21638_), .A3(new_n21640_), .A4(new_n21641_), .ZN(new_n21642_));
  NAND2_X1   g18510(.A1(new_n21620_), .A2(new_n21642_), .ZN(new_n21643_));
  INV_X1     g18511(.I(new_n21531_), .ZN(new_n21644_));
  NAND3_X1   g18512(.A1(new_n21615_), .A2(new_n21608_), .A3(pi0619), .ZN(new_n21645_));
  XOR2_X1    g18513(.A1(new_n21645_), .A2(new_n13904_), .Z(new_n21646_));
  NAND2_X1   g18514(.A1(new_n21625_), .A2(new_n21481_), .ZN(new_n21647_));
  NAND2_X1   g18515(.A1(new_n21647_), .A2(new_n20173_), .ZN(new_n21648_));
  AOI21_X1   g18516(.A1(new_n21646_), .A2(new_n21644_), .B(new_n21648_), .ZN(new_n21649_));
  AOI21_X1   g18517(.A1(new_n21643_), .A2(new_n21649_), .B(pi0792), .ZN(new_n21650_));
  NOR2_X1    g18518(.A1(new_n21481_), .A2(new_n13966_), .ZN(new_n21651_));
  NOR3_X1    g18519(.A1(new_n21635_), .A2(new_n13965_), .A3(new_n21633_), .ZN(new_n21652_));
  NOR2_X1    g18520(.A1(new_n21652_), .A2(new_n21651_), .ZN(new_n21653_));
  INV_X1     g18521(.I(new_n21653_), .ZN(new_n21654_));
  NAND3_X1   g18522(.A1(new_n21654_), .A2(pi0628), .A3(pi1156), .ZN(new_n21655_));
  NAND3_X1   g18523(.A1(new_n21653_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n21656_));
  AOI21_X1   g18524(.A1(new_n21655_), .A2(new_n21656_), .B(new_n21480_), .ZN(new_n21657_));
  NOR2_X1    g18525(.A1(new_n21657_), .A2(new_n12777_), .ZN(new_n21658_));
  NAND3_X1   g18526(.A1(new_n21654_), .A2(pi0628), .A3(pi1156), .ZN(new_n21659_));
  NAND3_X1   g18527(.A1(new_n21653_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n21660_));
  AOI21_X1   g18528(.A1(new_n21659_), .A2(new_n21660_), .B(new_n21480_), .ZN(new_n21661_));
  NAND3_X1   g18529(.A1(new_n21661_), .A2(pi0792), .A3(new_n21654_), .ZN(new_n21662_));
  NOR2_X1    g18530(.A1(new_n21662_), .A2(new_n21658_), .ZN(new_n21663_));
  INV_X1     g18531(.I(new_n21663_), .ZN(new_n21664_));
  NAND2_X1   g18532(.A1(new_n21662_), .A2(new_n21658_), .ZN(new_n21665_));
  NAND2_X1   g18533(.A1(new_n21664_), .A2(new_n21665_), .ZN(new_n21666_));
  NAND2_X1   g18534(.A1(new_n21481_), .A2(new_n14005_), .ZN(new_n21667_));
  NAND2_X1   g18535(.A1(new_n21667_), .A2(pi1157), .ZN(new_n21668_));
  AOI21_X1   g18536(.A1(new_n21666_), .A2(pi0647), .B(new_n21668_), .ZN(new_n21669_));
  AOI21_X1   g18537(.A1(new_n21664_), .A2(new_n21665_), .B(pi0647), .ZN(new_n21670_));
  NOR2_X1    g18538(.A1(new_n21480_), .A2(new_n14005_), .ZN(new_n21671_));
  NOR3_X1    g18539(.A1(new_n21670_), .A2(pi1157), .A3(new_n21671_), .ZN(new_n21672_));
  OAI21_X1   g18540(.A1(new_n21672_), .A2(new_n21669_), .B(pi0787), .ZN(new_n21673_));
  OAI21_X1   g18541(.A1(pi0787), .A2(new_n21666_), .B(new_n21673_), .ZN(new_n21674_));
  NOR2_X1    g18542(.A1(new_n21481_), .A2(new_n16372_), .ZN(new_n21675_));
  NOR2_X1    g18543(.A1(new_n21629_), .A2(new_n14142_), .ZN(new_n21676_));
  OAI21_X1   g18544(.A1(new_n21676_), .A2(new_n21675_), .B(new_n13994_), .ZN(new_n21677_));
  NOR2_X1    g18545(.A1(new_n21481_), .A2(new_n13994_), .ZN(new_n21678_));
  INV_X1     g18546(.I(new_n21678_), .ZN(new_n21679_));
  AOI21_X1   g18547(.A1(new_n21677_), .A2(new_n21679_), .B(new_n14210_), .ZN(new_n21680_));
  NOR2_X1    g18548(.A1(new_n21481_), .A2(new_n14211_), .ZN(new_n21681_));
  NOR2_X1    g18549(.A1(new_n21680_), .A2(new_n21681_), .ZN(new_n21682_));
  NOR2_X1    g18550(.A1(new_n14243_), .A2(pi0644), .ZN(new_n21683_));
  NOR2_X1    g18551(.A1(new_n21682_), .A2(new_n21683_), .ZN(new_n21684_));
  NAND2_X1   g18552(.A1(new_n21684_), .A2(pi0715), .ZN(new_n21685_));
  NAND2_X1   g18553(.A1(new_n21685_), .A2(new_n14204_), .ZN(new_n21686_));
  NAND2_X1   g18554(.A1(new_n21674_), .A2(new_n21686_), .ZN(new_n21687_));
  AOI21_X1   g18555(.A1(new_n21481_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n21688_));
  NOR2_X1    g18556(.A1(new_n21688_), .A2(pi0644), .ZN(new_n21689_));
  NOR3_X1    g18557(.A1(new_n21682_), .A2(new_n14200_), .A3(new_n21689_), .ZN(new_n21690_));
  OAI21_X1   g18558(.A1(new_n21674_), .A2(new_n21690_), .B(pi0644), .ZN(new_n21691_));
  AOI21_X1   g18559(.A1(new_n21691_), .A2(new_n21687_), .B(new_n12775_), .ZN(new_n21692_));
  NOR3_X1    g18560(.A1(new_n21682_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n21693_));
  OAI21_X1   g18561(.A1(new_n21682_), .A2(new_n21689_), .B(pi0790), .ZN(new_n21694_));
  NOR2_X1    g18562(.A1(new_n21694_), .A2(new_n19379_), .ZN(new_n21695_));
  OAI21_X1   g18563(.A1(new_n21695_), .A2(new_n21693_), .B(new_n21684_), .ZN(new_n21696_));
  NAND2_X1   g18564(.A1(new_n21677_), .A2(new_n21679_), .ZN(new_n21697_));
  INV_X1     g18565(.I(new_n21665_), .ZN(new_n21698_));
  OAI21_X1   g18566(.A1(new_n21698_), .A2(new_n21663_), .B(pi0647), .ZN(new_n21699_));
  NOR2_X1    g18567(.A1(new_n21698_), .A2(new_n21663_), .ZN(new_n21700_));
  INV_X1     g18568(.I(new_n21671_), .ZN(new_n21701_));
  OAI21_X1   g18569(.A1(new_n21700_), .A2(pi0647), .B(new_n21701_), .ZN(new_n21702_));
  NAND4_X1   g18570(.A1(new_n21699_), .A2(new_n14010_), .A3(pi1157), .A4(new_n21667_), .ZN(new_n21704_));
  NAND4_X1   g18571(.A1(new_n21699_), .A2(new_n14010_), .A3(pi1157), .A4(new_n21667_), .ZN(new_n21705_));
  NAND3_X1   g18572(.A1(new_n21705_), .A2(new_n21702_), .A3(new_n14011_), .ZN(new_n21706_));
  AOI21_X1   g18573(.A1(new_n21706_), .A2(new_n21704_), .B(new_n12776_), .ZN(new_n21707_));
  OAI21_X1   g18574(.A1(new_n21707_), .A2(new_n21697_), .B(new_n16576_), .ZN(new_n21708_));
  NAND2_X1   g18575(.A1(new_n21708_), .A2(new_n21696_), .ZN(new_n21709_));
  NOR2_X1    g18576(.A1(new_n21657_), .A2(new_n13976_), .ZN(new_n21710_));
  NOR2_X1    g18577(.A1(new_n21661_), .A2(pi0629), .ZN(new_n21711_));
  NOR2_X1    g18578(.A1(new_n21710_), .A2(new_n21711_), .ZN(new_n21712_));
  NOR2_X1    g18579(.A1(new_n21676_), .A2(new_n21675_), .ZN(new_n21713_));
  NOR2_X1    g18580(.A1(new_n21713_), .A2(new_n16874_), .ZN(new_n21714_));
  NOR3_X1    g18581(.A1(new_n13219_), .A2(pi0625), .A3(pi0734), .ZN(new_n21715_));
  INV_X1     g18582(.I(new_n21715_), .ZN(new_n21716_));
  NOR2_X1    g18583(.A1(new_n9992_), .A2(pi0182), .ZN(new_n21717_));
  NOR2_X1    g18584(.A1(new_n21717_), .A2(pi1153), .ZN(new_n21718_));
  NAND2_X1   g18585(.A1(new_n21716_), .A2(new_n21718_), .ZN(new_n21719_));
  INV_X1     g18586(.I(new_n21719_), .ZN(new_n21720_));
  NOR2_X1    g18587(.A1(new_n21720_), .A2(new_n13748_), .ZN(new_n21721_));
  AOI21_X1   g18588(.A1(new_n13218_), .A2(new_n17604_), .B(new_n21717_), .ZN(new_n21722_));
  INV_X1     g18589(.I(new_n21722_), .ZN(new_n21723_));
  AOI21_X1   g18590(.A1(new_n21716_), .A2(new_n21723_), .B(new_n13614_), .ZN(new_n21724_));
  INV_X1     g18591(.I(new_n21724_), .ZN(new_n21725_));
  NOR3_X1    g18592(.A1(new_n21725_), .A2(new_n13748_), .A3(new_n21723_), .ZN(new_n21726_));
  XNOR2_X1   g18593(.A1(new_n21726_), .A2(new_n21721_), .ZN(new_n21727_));
  NAND2_X1   g18594(.A1(new_n21727_), .A2(new_n14049_), .ZN(new_n21728_));
  NOR2_X1    g18595(.A1(new_n21728_), .A2(new_n14051_), .ZN(new_n21729_));
  INV_X1     g18596(.I(new_n21729_), .ZN(new_n21730_));
  NOR4_X1    g18597(.A1(new_n21730_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n21731_));
  NOR2_X1    g18598(.A1(new_n21731_), .A2(new_n14005_), .ZN(new_n21732_));
  XOR2_X1    g18599(.A1(new_n21732_), .A2(new_n14007_), .Z(new_n21733_));
  NAND2_X1   g18600(.A1(new_n21733_), .A2(new_n21717_), .ZN(new_n21734_));
  INV_X1     g18601(.I(new_n21717_), .ZN(new_n21735_));
  NOR2_X1    g18602(.A1(new_n21735_), .A2(pi0647), .ZN(new_n21736_));
  AOI21_X1   g18603(.A1(new_n21731_), .A2(pi0647), .B(new_n21736_), .ZN(new_n21737_));
  AOI21_X1   g18604(.A1(new_n21737_), .A2(pi1157), .B(new_n12776_), .ZN(new_n21738_));
  AOI22_X1   g18605(.A1(new_n21734_), .A2(new_n21738_), .B1(new_n12776_), .B2(new_n21731_), .ZN(new_n21739_));
  NOR2_X1    g18606(.A1(new_n21730_), .A2(new_n14163_), .ZN(new_n21740_));
  NOR2_X1    g18607(.A1(new_n21549_), .A2(new_n21717_), .ZN(new_n21741_));
  INV_X1     g18608(.I(new_n21741_), .ZN(new_n21742_));
  NAND3_X1   g18609(.A1(new_n21742_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n21743_));
  AOI21_X1   g18610(.A1(new_n21743_), .A2(new_n16444_), .B(new_n21550_), .ZN(new_n21744_));
  NOR2_X1    g18611(.A1(new_n21744_), .A2(new_n13801_), .ZN(new_n21745_));
  NOR2_X1    g18612(.A1(new_n21717_), .A2(pi1155), .ZN(new_n21746_));
  NOR3_X1    g18613(.A1(new_n21550_), .A2(new_n16444_), .A3(new_n21746_), .ZN(new_n21747_));
  NAND4_X1   g18614(.A1(new_n21747_), .A2(new_n21742_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n21748_));
  XOR2_X1    g18615(.A1(new_n21745_), .A2(new_n21748_), .Z(new_n21749_));
  NOR2_X1    g18616(.A1(new_n21749_), .A2(new_n13817_), .ZN(new_n21750_));
  OAI21_X1   g18617(.A1(new_n21750_), .A2(pi0618), .B(new_n9992_), .ZN(new_n21751_));
  NAND2_X1   g18618(.A1(new_n21751_), .A2(pi0781), .ZN(new_n21752_));
  OAI21_X1   g18619(.A1(new_n21750_), .A2(new_n9992_), .B(pi0618), .ZN(new_n21753_));
  NOR3_X1    g18620(.A1(new_n21753_), .A2(new_n13855_), .A3(new_n21749_), .ZN(new_n21754_));
  XOR2_X1    g18621(.A1(new_n21754_), .A2(new_n21752_), .Z(new_n21755_));
  NOR2_X1    g18622(.A1(new_n21755_), .A2(new_n13868_), .ZN(new_n21756_));
  OAI21_X1   g18623(.A1(new_n21756_), .A2(pi0619), .B(new_n9992_), .ZN(new_n21757_));
  NAND2_X1   g18624(.A1(new_n21757_), .A2(pi0789), .ZN(new_n21758_));
  OAI21_X1   g18625(.A1(new_n21756_), .A2(new_n9992_), .B(pi0619), .ZN(new_n21759_));
  NOR3_X1    g18626(.A1(new_n21759_), .A2(new_n13896_), .A3(new_n21755_), .ZN(new_n21760_));
  XOR2_X1    g18627(.A1(new_n21760_), .A2(new_n21758_), .Z(new_n21761_));
  NAND2_X1   g18628(.A1(new_n21761_), .A2(new_n13962_), .ZN(new_n21762_));
  XOR2_X1    g18629(.A1(new_n21762_), .A2(new_n18976_), .Z(new_n21763_));
  AOI22_X1   g18630(.A1(new_n21763_), .A2(new_n21717_), .B1(new_n16639_), .B2(new_n21740_), .ZN(new_n21764_));
  NOR2_X1    g18631(.A1(new_n21722_), .A2(new_n13203_), .ZN(new_n21765_));
  NAND2_X1   g18632(.A1(new_n21765_), .A2(pi0625), .ZN(new_n21766_));
  NAND3_X1   g18633(.A1(new_n21766_), .A2(pi1153), .A3(new_n21741_), .ZN(new_n21767_));
  NOR2_X1    g18634(.A1(new_n21720_), .A2(new_n14081_), .ZN(new_n21768_));
  AOI21_X1   g18635(.A1(new_n21768_), .A2(new_n21767_), .B(new_n13748_), .ZN(new_n21769_));
  NOR2_X1    g18636(.A1(new_n21742_), .A2(new_n21765_), .ZN(new_n21770_));
  INV_X1     g18637(.I(new_n21766_), .ZN(new_n21771_));
  OAI21_X1   g18638(.A1(new_n21770_), .A2(new_n21771_), .B(new_n21718_), .ZN(new_n21772_));
  NAND4_X1   g18639(.A1(new_n21772_), .A2(new_n13749_), .A3(new_n21725_), .A4(new_n21770_), .ZN(new_n21773_));
  XNOR2_X1   g18640(.A1(new_n21773_), .A2(new_n21769_), .ZN(new_n21774_));
  NAND2_X1   g18641(.A1(new_n21774_), .A2(new_n13801_), .ZN(new_n21775_));
  NOR2_X1    g18642(.A1(new_n21744_), .A2(pi0660), .ZN(new_n21779_));
  NOR2_X1    g18643(.A1(new_n21774_), .A2(new_n13766_), .ZN(new_n21780_));
  XOR2_X1    g18644(.A1(new_n21780_), .A2(new_n14090_), .Z(new_n21781_));
  NOR2_X1    g18645(.A1(new_n21727_), .A2(new_n13801_), .ZN(new_n21782_));
  NAND2_X1   g18646(.A1(new_n21781_), .A2(new_n21782_), .ZN(new_n21783_));
  OAI21_X1   g18647(.A1(new_n21783_), .A2(new_n21779_), .B(new_n21775_), .ZN(new_n21784_));
  NAND2_X1   g18648(.A1(new_n21784_), .A2(new_n13855_), .ZN(new_n21785_));
  INV_X1     g18649(.I(new_n21728_), .ZN(new_n21786_));
  NOR2_X1    g18650(.A1(new_n21784_), .A2(new_n13816_), .ZN(new_n21787_));
  XOR2_X1    g18651(.A1(new_n21787_), .A2(new_n13818_), .Z(new_n21788_));
  NAND2_X1   g18652(.A1(new_n21788_), .A2(new_n21786_), .ZN(new_n21789_));
  NAND3_X1   g18653(.A1(new_n21789_), .A2(new_n13823_), .A3(new_n21753_), .ZN(new_n21790_));
  NAND3_X1   g18654(.A1(new_n21790_), .A2(new_n13823_), .A3(new_n21751_), .ZN(new_n21791_));
  NOR2_X1    g18655(.A1(new_n21784_), .A2(new_n13817_), .ZN(new_n21792_));
  XOR2_X1    g18656(.A1(new_n21792_), .A2(new_n13818_), .Z(new_n21793_));
  NAND4_X1   g18657(.A1(new_n21791_), .A2(pi0781), .A3(new_n21786_), .A4(new_n21793_), .ZN(new_n21794_));
  NAND2_X1   g18658(.A1(new_n21794_), .A2(new_n21785_), .ZN(new_n21795_));
  NOR2_X1    g18659(.A1(new_n21795_), .A2(new_n13860_), .ZN(new_n21796_));
  XOR2_X1    g18660(.A1(new_n21796_), .A2(new_n13904_), .Z(new_n21797_));
  NOR2_X1    g18661(.A1(new_n21797_), .A2(new_n21730_), .ZN(new_n21798_));
  NAND2_X1   g18662(.A1(new_n21759_), .A2(new_n13884_), .ZN(new_n21799_));
  INV_X1     g18663(.I(new_n21795_), .ZN(new_n21800_));
  AOI21_X1   g18664(.A1(new_n21800_), .A2(new_n14143_), .B(pi0789), .ZN(new_n21801_));
  OAI21_X1   g18665(.A1(new_n21798_), .A2(new_n21799_), .B(new_n21801_), .ZN(new_n21802_));
  NOR2_X1    g18666(.A1(new_n21795_), .A2(new_n13868_), .ZN(new_n21803_));
  XOR2_X1    g18667(.A1(new_n21803_), .A2(new_n13903_), .Z(new_n21804_));
  NAND2_X1   g18668(.A1(new_n21757_), .A2(new_n19018_), .ZN(new_n21805_));
  AOI21_X1   g18669(.A1(new_n21804_), .A2(new_n21729_), .B(new_n21805_), .ZN(new_n21806_));
  AOI21_X1   g18670(.A1(new_n21802_), .A2(new_n21806_), .B(new_n21764_), .ZN(new_n21807_));
  NAND2_X1   g18671(.A1(new_n21761_), .A2(new_n16372_), .ZN(new_n21808_));
  OAI21_X1   g18672(.A1(new_n16372_), .A2(new_n21717_), .B(new_n21808_), .ZN(new_n21809_));
  NAND3_X1   g18673(.A1(new_n21809_), .A2(new_n18929_), .A3(new_n21740_), .ZN(new_n21810_));
  NAND2_X1   g18674(.A1(new_n21810_), .A2(new_n16569_), .ZN(new_n21811_));
  XOR2_X1    g18675(.A1(new_n21811_), .A2(new_n16572_), .Z(new_n21812_));
  AOI21_X1   g18676(.A1(new_n19022_), .A2(new_n21810_), .B(new_n21812_), .ZN(new_n21813_));
  NAND2_X1   g18677(.A1(new_n21761_), .A2(new_n13963_), .ZN(new_n21814_));
  XNOR2_X1   g18678(.A1(new_n21814_), .A2(new_n19028_), .ZN(new_n21815_));
  NOR3_X1    g18679(.A1(new_n21815_), .A2(new_n16424_), .A3(new_n21735_), .ZN(new_n21816_));
  OAI21_X1   g18680(.A1(new_n21813_), .A2(new_n16574_), .B(new_n21816_), .ZN(new_n21817_));
  NOR2_X1    g18681(.A1(new_n21809_), .A2(new_n13994_), .ZN(new_n21818_));
  XNOR2_X1   g18682(.A1(new_n21818_), .A2(new_n19033_), .ZN(new_n21819_));
  AOI22_X1   g18683(.A1(new_n21819_), .A2(new_n21717_), .B1(new_n14206_), .B2(new_n21737_), .ZN(new_n21820_));
  NOR3_X1    g18684(.A1(new_n21820_), .A2(new_n14010_), .A3(new_n21734_), .ZN(new_n21821_));
  OAI22_X1   g18685(.A1(new_n21807_), .A2(new_n21817_), .B1(new_n12776_), .B2(new_n21821_), .ZN(new_n21822_));
  NAND2_X1   g18686(.A1(new_n21822_), .A2(pi0644), .ZN(new_n21823_));
  XOR2_X1    g18687(.A1(new_n21823_), .A2(new_n14205_), .Z(new_n21824_));
  NOR2_X1    g18688(.A1(new_n21824_), .A2(new_n21739_), .ZN(new_n21825_));
  NOR2_X1    g18689(.A1(new_n21809_), .A2(new_n18968_), .ZN(new_n21826_));
  NAND2_X1   g18690(.A1(new_n18967_), .A2(new_n21717_), .ZN(new_n21827_));
  XOR2_X1    g18691(.A1(new_n21826_), .A2(new_n21827_), .Z(new_n21828_));
  NAND2_X1   g18692(.A1(new_n21828_), .A2(pi0715), .ZN(new_n21829_));
  XOR2_X1    g18693(.A1(new_n21829_), .A2(new_n14205_), .Z(new_n21830_));
  OAI21_X1   g18694(.A1(new_n21830_), .A2(new_n21735_), .B(new_n14203_), .ZN(new_n21831_));
  NAND2_X1   g18695(.A1(new_n21828_), .A2(pi0644), .ZN(new_n21832_));
  XOR2_X1    g18696(.A1(new_n21832_), .A2(new_n14217_), .Z(new_n21833_));
  AOI21_X1   g18697(.A1(new_n21833_), .A2(new_n21717_), .B(pi1160), .ZN(new_n21834_));
  OAI21_X1   g18698(.A1(new_n21825_), .A2(new_n21831_), .B(new_n21834_), .ZN(new_n21835_));
  NAND2_X1   g18699(.A1(new_n21822_), .A2(pi0715), .ZN(new_n21836_));
  XOR2_X1    g18700(.A1(new_n21836_), .A2(new_n14205_), .Z(new_n21837_));
  NOR2_X1    g18701(.A1(new_n21837_), .A2(new_n21739_), .ZN(new_n21838_));
  AOI21_X1   g18702(.A1(new_n21835_), .A2(new_n21838_), .B(new_n14799_), .ZN(new_n21839_));
  XOR2_X1    g18703(.A1(new_n21839_), .A2(new_n14800_), .Z(new_n21840_));
  OAI21_X1   g18704(.A1(new_n7240_), .A2(pi0182), .B(new_n14799_), .ZN(new_n21841_));
  NOR2_X1    g18705(.A1(new_n21822_), .A2(new_n21841_), .ZN(new_n21842_));
  AOI21_X1   g18706(.A1(new_n21840_), .A2(new_n21842_), .B(po1038), .ZN(new_n21843_));
  NOR3_X1    g18707(.A1(new_n21714_), .A2(new_n21712_), .A3(new_n21843_), .ZN(new_n21844_));
  OAI21_X1   g18708(.A1(new_n21692_), .A2(new_n21709_), .B(new_n21844_), .ZN(new_n21845_));
  NOR2_X1    g18709(.A1(new_n21845_), .A2(new_n21650_), .ZN(po0339));
  NAND2_X1   g18710(.A1(new_n13627_), .A2(new_n7375_), .ZN(new_n21847_));
  INV_X1     g18711(.I(new_n21847_), .ZN(new_n21848_));
  AOI21_X1   g18712(.A1(new_n7375_), .A2(new_n17153_), .B(pi0038), .ZN(new_n21849_));
  NOR2_X1    g18713(.A1(new_n7375_), .A2(new_n17153_), .ZN(new_n21850_));
  OAI21_X1   g18714(.A1(new_n20007_), .A2(new_n21850_), .B(pi0038), .ZN(new_n21851_));
  INV_X1     g18715(.I(new_n21851_), .ZN(new_n21852_));
  AOI21_X1   g18716(.A1(new_n13097_), .A2(new_n21849_), .B(new_n21852_), .ZN(new_n21853_));
  NOR2_X1    g18717(.A1(new_n3289_), .A2(pi0183), .ZN(new_n21854_));
  AOI21_X1   g18718(.A1(new_n21853_), .A2(new_n3289_), .B(new_n21854_), .ZN(new_n21855_));
  NAND2_X1   g18719(.A1(new_n21855_), .A2(new_n13776_), .ZN(new_n21856_));
  OAI21_X1   g18720(.A1(new_n15147_), .A2(new_n21848_), .B(new_n21856_), .ZN(new_n21857_));
  NAND2_X1   g18721(.A1(new_n21857_), .A2(pi0609), .ZN(new_n21858_));
  NAND2_X1   g18722(.A1(new_n21858_), .A2(pi0785), .ZN(new_n21859_));
  AOI21_X1   g18723(.A1(new_n21847_), .A2(new_n14467_), .B(pi0609), .ZN(new_n21860_));
  NOR2_X1    g18724(.A1(new_n21860_), .A2(new_n21856_), .ZN(new_n21861_));
  NAND2_X1   g18725(.A1(new_n21848_), .A2(new_n13775_), .ZN(new_n21862_));
  OAI21_X1   g18726(.A1(new_n13775_), .A2(new_n21855_), .B(new_n21862_), .ZN(new_n21863_));
  NAND3_X1   g18727(.A1(new_n21863_), .A2(pi0785), .A3(new_n21861_), .ZN(new_n21864_));
  XNOR2_X1   g18728(.A1(new_n21859_), .A2(new_n21864_), .ZN(new_n21865_));
  NAND2_X1   g18729(.A1(new_n21865_), .A2(pi0618), .ZN(new_n21866_));
  XOR2_X1    g18730(.A1(new_n21866_), .A2(new_n13819_), .Z(new_n21867_));
  NAND2_X1   g18731(.A1(new_n21867_), .A2(new_n21848_), .ZN(new_n21868_));
  NAND2_X1   g18732(.A1(new_n21868_), .A2(pi0781), .ZN(new_n21869_));
  NAND2_X1   g18733(.A1(new_n21865_), .A2(pi1154), .ZN(new_n21870_));
  XOR2_X1    g18734(.A1(new_n21870_), .A2(new_n13819_), .Z(new_n21871_));
  NAND2_X1   g18735(.A1(new_n21871_), .A2(new_n21848_), .ZN(new_n21872_));
  NOR3_X1    g18736(.A1(new_n21872_), .A2(new_n13855_), .A3(new_n21865_), .ZN(new_n21873_));
  XNOR2_X1   g18737(.A1(new_n21873_), .A2(new_n21869_), .ZN(new_n21874_));
  NAND3_X1   g18738(.A1(new_n21874_), .A2(pi0619), .A3(pi1159), .ZN(new_n21875_));
  XOR2_X1    g18739(.A1(new_n21873_), .A2(new_n21869_), .Z(new_n21876_));
  NAND3_X1   g18740(.A1(new_n21876_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n21877_));
  AOI21_X1   g18741(.A1(new_n21875_), .A2(new_n21877_), .B(new_n21847_), .ZN(new_n21878_));
  NOR2_X1    g18742(.A1(new_n21848_), .A2(new_n13880_), .ZN(new_n21879_));
  OAI21_X1   g18743(.A1(new_n13721_), .A2(new_n17148_), .B(new_n7375_), .ZN(new_n21880_));
  NAND2_X1   g18744(.A1(new_n16715_), .A2(new_n7375_), .ZN(new_n21881_));
  NAND4_X1   g18745(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n21880_), .A4(new_n21881_), .ZN(new_n21882_));
  NAND2_X1   g18746(.A1(new_n21882_), .A2(new_n14424_), .ZN(new_n21883_));
  NAND2_X1   g18747(.A1(new_n21883_), .A2(pi0183), .ZN(new_n21884_));
  OAI21_X1   g18748(.A1(new_n21884_), .A2(new_n21847_), .B(new_n3290_), .ZN(new_n21885_));
  NAND2_X1   g18749(.A1(new_n21885_), .A2(pi0725), .ZN(new_n21886_));
  NAND2_X1   g18750(.A1(new_n21886_), .A2(pi0625), .ZN(new_n21887_));
  XOR2_X1    g18751(.A1(new_n21887_), .A2(new_n13620_), .Z(new_n21888_));
  NAND2_X1   g18752(.A1(new_n21888_), .A2(new_n21848_), .ZN(new_n21889_));
  NAND2_X1   g18753(.A1(new_n21889_), .A2(pi0778), .ZN(new_n21890_));
  NAND2_X1   g18754(.A1(new_n21886_), .A2(pi1153), .ZN(new_n21891_));
  XOR2_X1    g18755(.A1(new_n21891_), .A2(new_n13620_), .Z(new_n21892_));
  NAND2_X1   g18756(.A1(new_n21892_), .A2(new_n21848_), .ZN(new_n21893_));
  NOR3_X1    g18757(.A1(new_n21893_), .A2(new_n13748_), .A3(new_n21886_), .ZN(new_n21894_));
  XNOR2_X1   g18758(.A1(new_n21894_), .A2(new_n21890_), .ZN(new_n21895_));
  NOR2_X1    g18759(.A1(new_n21847_), .A2(new_n13805_), .ZN(new_n21896_));
  AOI21_X1   g18760(.A1(new_n21895_), .A2(new_n13805_), .B(new_n21896_), .ZN(new_n21897_));
  AOI21_X1   g18761(.A1(new_n21897_), .A2(new_n13880_), .B(new_n21879_), .ZN(new_n21898_));
  NOR2_X1    g18762(.A1(new_n13453_), .A2(new_n7375_), .ZN(new_n21899_));
  XOR2_X1    g18763(.A1(new_n21899_), .A2(new_n21850_), .Z(new_n21900_));
  NAND2_X1   g18764(.A1(new_n21900_), .A2(new_n13521_), .ZN(new_n21901_));
  NAND3_X1   g18765(.A1(new_n14270_), .A2(pi0183), .A3(pi0755), .ZN(new_n21902_));
  NAND3_X1   g18766(.A1(new_n14272_), .A2(new_n7375_), .A3(pi0755), .ZN(new_n21903_));
  AOI21_X1   g18767(.A1(new_n21902_), .A2(new_n21903_), .B(new_n13152_), .ZN(new_n21904_));
  NAND3_X1   g18768(.A1(new_n13198_), .A2(pi0183), .A3(pi0755), .ZN(new_n21905_));
  NAND3_X1   g18769(.A1(new_n13200_), .A2(pi0183), .A3(new_n17153_), .ZN(new_n21906_));
  AOI21_X1   g18770(.A1(new_n21906_), .A2(new_n21905_), .B(new_n13191_), .ZN(new_n21907_));
  OAI21_X1   g18771(.A1(new_n21904_), .A2(new_n3262_), .B(new_n21907_), .ZN(new_n21908_));
  NAND3_X1   g18772(.A1(new_n21901_), .A2(new_n3183_), .A3(new_n21908_), .ZN(new_n21909_));
  NOR2_X1    g18773(.A1(new_n14284_), .A2(new_n17153_), .ZN(new_n21910_));
  XOR2_X1    g18774(.A1(new_n21910_), .A2(new_n21850_), .Z(new_n21911_));
  NAND3_X1   g18775(.A1(new_n21909_), .A2(new_n21911_), .A3(new_n13359_), .ZN(new_n21912_));
  NAND3_X1   g18776(.A1(new_n21912_), .A2(new_n17148_), .A3(new_n3290_), .ZN(new_n21913_));
  OAI21_X1   g18777(.A1(new_n15587_), .A2(new_n7375_), .B(new_n17153_), .ZN(new_n21914_));
  NAND2_X1   g18778(.A1(new_n21914_), .A2(new_n13209_), .ZN(new_n21915_));
  NOR2_X1    g18779(.A1(new_n13105_), .A2(pi0755), .ZN(new_n21916_));
  INV_X1     g18780(.I(new_n21916_), .ZN(new_n21917_));
  NAND2_X1   g18781(.A1(new_n21917_), .A2(new_n16751_), .ZN(new_n21918_));
  NAND4_X1   g18782(.A1(new_n5503_), .A2(new_n21918_), .A3(pi0183), .A4(new_n3290_), .ZN(new_n21919_));
  AOI21_X1   g18783(.A1(new_n21915_), .A2(new_n3259_), .B(new_n21919_), .ZN(new_n21920_));
  AOI21_X1   g18784(.A1(new_n21913_), .A2(new_n21920_), .B(pi0725), .ZN(new_n21921_));
  NOR2_X1    g18785(.A1(new_n21921_), .A2(new_n21853_), .ZN(new_n21922_));
  INV_X1     g18786(.I(new_n21922_), .ZN(new_n21923_));
  INV_X1     g18787(.I(new_n21855_), .ZN(new_n21924_));
  NOR2_X1    g18788(.A1(new_n21922_), .A2(new_n13613_), .ZN(new_n21925_));
  XOR2_X1    g18789(.A1(new_n21925_), .A2(new_n13615_), .Z(new_n21926_));
  NAND2_X1   g18790(.A1(new_n21893_), .A2(new_n14081_), .ZN(new_n21927_));
  AOI21_X1   g18791(.A1(new_n21926_), .A2(new_n21924_), .B(new_n21927_), .ZN(new_n21928_));
  INV_X1     g18792(.I(new_n21928_), .ZN(new_n21929_));
  NOR2_X1    g18793(.A1(new_n21922_), .A2(new_n13614_), .ZN(new_n21930_));
  XOR2_X1    g18794(.A1(new_n21930_), .A2(new_n13615_), .Z(new_n21931_));
  AOI21_X1   g18795(.A1(new_n21931_), .A2(new_n21924_), .B(pi0608), .ZN(new_n21932_));
  NAND2_X1   g18796(.A1(new_n21929_), .A2(new_n21932_), .ZN(new_n21933_));
  NOR2_X1    g18797(.A1(new_n21889_), .A2(new_n13748_), .ZN(new_n21934_));
  AOI22_X1   g18798(.A1(new_n21933_), .A2(new_n21934_), .B1(new_n13748_), .B2(new_n21923_), .ZN(new_n21935_));
  AOI21_X1   g18799(.A1(new_n21935_), .A2(pi1155), .B(new_n14694_), .ZN(new_n21936_));
  INV_X1     g18800(.I(new_n21932_), .ZN(new_n21937_));
  NOR2_X1    g18801(.A1(new_n21937_), .A2(new_n21928_), .ZN(new_n21938_));
  INV_X1     g18802(.I(new_n21934_), .ZN(new_n21939_));
  OAI22_X1   g18803(.A1(new_n21938_), .A2(new_n21939_), .B1(pi0778), .B2(new_n21922_), .ZN(new_n21940_));
  NOR3_X1    g18804(.A1(new_n21940_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n21941_));
  OAI21_X1   g18805(.A1(new_n21941_), .A2(new_n21936_), .B(new_n21895_), .ZN(new_n21942_));
  NAND2_X1   g18806(.A1(new_n21858_), .A2(pi0660), .ZN(new_n21943_));
  INV_X1     g18807(.I(new_n21943_), .ZN(new_n21944_));
  NOR2_X1    g18808(.A1(new_n21861_), .A2(pi0660), .ZN(new_n21945_));
  INV_X1     g18809(.I(new_n21945_), .ZN(new_n21946_));
  AOI21_X1   g18810(.A1(new_n21942_), .A2(new_n21944_), .B(new_n21946_), .ZN(new_n21947_));
  NOR2_X1    g18811(.A1(new_n21940_), .A2(new_n13766_), .ZN(new_n21948_));
  NOR2_X1    g18812(.A1(new_n21948_), .A2(new_n14694_), .ZN(new_n21949_));
  NAND2_X1   g18813(.A1(new_n21948_), .A2(new_n14694_), .ZN(new_n21950_));
  INV_X1     g18814(.I(new_n21950_), .ZN(new_n21951_));
  INV_X1     g18815(.I(new_n21895_), .ZN(new_n21952_));
  NOR2_X1    g18816(.A1(new_n21952_), .A2(new_n13801_), .ZN(new_n21953_));
  OAI21_X1   g18817(.A1(new_n21951_), .A2(new_n21949_), .B(new_n21953_), .ZN(new_n21954_));
  OAI22_X1   g18818(.A1(new_n21954_), .A2(new_n21947_), .B1(pi0785), .B2(new_n21935_), .ZN(new_n21955_));
  NAND3_X1   g18819(.A1(new_n21955_), .A2(pi0618), .A3(pi1154), .ZN(new_n21956_));
  NAND3_X1   g18820(.A1(new_n21940_), .A2(pi0609), .A3(pi1155), .ZN(new_n21957_));
  NAND3_X1   g18821(.A1(new_n21935_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n21958_));
  AOI21_X1   g18822(.A1(new_n21957_), .A2(new_n21958_), .B(new_n21952_), .ZN(new_n21959_));
  OAI21_X1   g18823(.A1(new_n21959_), .A2(new_n21943_), .B(new_n21945_), .ZN(new_n21960_));
  NAND2_X1   g18824(.A1(new_n21935_), .A2(pi0609), .ZN(new_n21961_));
  NAND2_X1   g18825(.A1(new_n21961_), .A2(new_n14090_), .ZN(new_n21962_));
  INV_X1     g18826(.I(new_n21953_), .ZN(new_n21963_));
  AOI21_X1   g18827(.A1(new_n21950_), .A2(new_n21962_), .B(new_n21963_), .ZN(new_n21964_));
  AOI22_X1   g18828(.A1(new_n21960_), .A2(new_n21964_), .B1(new_n13801_), .B2(new_n21940_), .ZN(new_n21965_));
  NAND3_X1   g18829(.A1(new_n21965_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n21966_));
  AOI21_X1   g18830(.A1(new_n21956_), .A2(new_n21966_), .B(new_n21897_), .ZN(new_n21967_));
  NAND2_X1   g18831(.A1(new_n21868_), .A2(pi0627), .ZN(new_n21968_));
  OAI21_X1   g18832(.A1(new_n21967_), .A2(new_n21968_), .B(pi0781), .ZN(new_n21969_));
  INV_X1     g18833(.I(new_n21897_), .ZN(new_n21970_));
  AOI21_X1   g18834(.A1(new_n21965_), .A2(pi0618), .B(new_n13819_), .ZN(new_n21971_));
  NOR3_X1    g18835(.A1(new_n21955_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n21972_));
  OAI21_X1   g18836(.A1(new_n21972_), .A2(new_n21971_), .B(new_n21970_), .ZN(new_n21973_));
  AND3_X2    g18837(.A1(new_n21955_), .A2(new_n19177_), .A3(new_n21872_), .Z(new_n21974_));
  NAND3_X1   g18838(.A1(new_n21969_), .A2(new_n21973_), .A3(new_n21974_), .ZN(new_n21975_));
  AOI21_X1   g18839(.A1(new_n21965_), .A2(pi1154), .B(new_n13819_), .ZN(new_n21976_));
  NOR3_X1    g18840(.A1(new_n21955_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n21977_));
  OAI21_X1   g18841(.A1(new_n21977_), .A2(new_n21976_), .B(new_n21970_), .ZN(new_n21978_));
  INV_X1     g18842(.I(new_n21968_), .ZN(new_n21979_));
  AOI21_X1   g18843(.A1(new_n21978_), .A2(new_n21979_), .B(new_n13855_), .ZN(new_n21980_));
  NAND4_X1   g18844(.A1(new_n21973_), .A2(new_n19177_), .A3(new_n21872_), .A4(new_n21955_), .ZN(new_n21981_));
  NAND2_X1   g18845(.A1(new_n21981_), .A2(new_n21980_), .ZN(new_n21982_));
  NAND2_X1   g18846(.A1(new_n21982_), .A2(new_n21975_), .ZN(new_n21983_));
  NAND3_X1   g18847(.A1(new_n21983_), .A2(pi0619), .A3(pi1159), .ZN(new_n21984_));
  NAND4_X1   g18848(.A1(new_n21982_), .A2(new_n21975_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n21985_));
  AOI21_X1   g18849(.A1(new_n21984_), .A2(new_n21985_), .B(new_n21898_), .ZN(new_n21986_));
  OAI21_X1   g18850(.A1(new_n21986_), .A2(new_n20003_), .B(new_n21878_), .ZN(new_n21987_));
  NAND2_X1   g18851(.A1(new_n21983_), .A2(new_n13896_), .ZN(new_n21988_));
  NOR2_X1    g18852(.A1(new_n21878_), .A2(new_n13896_), .ZN(new_n21989_));
  NAND3_X1   g18853(.A1(new_n21874_), .A2(pi0619), .A3(pi1159), .ZN(new_n21990_));
  NAND3_X1   g18854(.A1(new_n21876_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n21991_));
  NAND2_X1   g18855(.A1(new_n21990_), .A2(new_n21991_), .ZN(new_n21992_));
  NAND4_X1   g18856(.A1(new_n21992_), .A2(pi0789), .A3(new_n21848_), .A4(new_n21874_), .ZN(new_n21993_));
  OR2_X2     g18857(.A1(new_n21993_), .A2(new_n21989_), .Z(new_n21994_));
  NAND2_X1   g18858(.A1(new_n21993_), .A2(new_n21989_), .ZN(new_n21995_));
  NAND2_X1   g18859(.A1(new_n21994_), .A2(new_n21995_), .ZN(new_n21996_));
  NAND3_X1   g18860(.A1(new_n21996_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n21997_));
  NAND4_X1   g18861(.A1(new_n21994_), .A2(new_n13901_), .A3(new_n13962_), .A4(new_n21995_), .ZN(new_n21998_));
  AOI21_X1   g18862(.A1(new_n21997_), .A2(new_n21998_), .B(new_n21847_), .ZN(new_n21999_));
  NOR2_X1    g18863(.A1(new_n21847_), .A2(new_n13919_), .ZN(new_n22000_));
  NAND2_X1   g18864(.A1(new_n21898_), .A2(new_n13919_), .ZN(new_n22001_));
  INV_X1     g18865(.I(new_n22001_), .ZN(new_n22002_));
  NOR2_X1    g18866(.A1(new_n22002_), .A2(new_n22000_), .ZN(new_n22003_));
  NOR2_X1    g18867(.A1(new_n22003_), .A2(new_n14162_), .ZN(new_n22004_));
  OAI21_X1   g18868(.A1(new_n21999_), .A2(new_n22004_), .B(new_n19204_), .ZN(new_n22005_));
  NOR2_X1    g18869(.A1(new_n21996_), .A2(new_n19208_), .ZN(new_n22006_));
  XNOR2_X1   g18870(.A1(new_n22006_), .A2(new_n19028_), .ZN(new_n22007_));
  NOR2_X1    g18871(.A1(new_n21847_), .A2(new_n15479_), .ZN(new_n22008_));
  NAND4_X1   g18872(.A1(new_n21988_), .A2(new_n22005_), .A3(new_n22007_), .A4(new_n22008_), .ZN(new_n22009_));
  NAND2_X1   g18873(.A1(new_n21987_), .A2(new_n22009_), .ZN(new_n22010_));
  INV_X1     g18874(.I(new_n21898_), .ZN(new_n22011_));
  NAND3_X1   g18875(.A1(new_n21982_), .A2(new_n21975_), .A3(pi0619), .ZN(new_n22012_));
  XOR2_X1    g18876(.A1(new_n22012_), .A2(new_n13904_), .Z(new_n22013_));
  NAND2_X1   g18877(.A1(new_n21992_), .A2(new_n21848_), .ZN(new_n22014_));
  NAND2_X1   g18878(.A1(new_n22014_), .A2(new_n20173_), .ZN(new_n22015_));
  AOI21_X1   g18879(.A1(new_n22013_), .A2(new_n22011_), .B(new_n22015_), .ZN(new_n22016_));
  AOI21_X1   g18880(.A1(new_n22010_), .A2(new_n22016_), .B(pi0792), .ZN(new_n22017_));
  NOR2_X1    g18881(.A1(new_n21848_), .A2(new_n13966_), .ZN(new_n22018_));
  NOR3_X1    g18882(.A1(new_n22002_), .A2(new_n13965_), .A3(new_n22000_), .ZN(new_n22019_));
  NOR2_X1    g18883(.A1(new_n22019_), .A2(new_n22018_), .ZN(new_n22020_));
  INV_X1     g18884(.I(new_n22020_), .ZN(new_n22021_));
  NAND3_X1   g18885(.A1(new_n22021_), .A2(pi0628), .A3(pi1156), .ZN(new_n22022_));
  NAND3_X1   g18886(.A1(new_n22020_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n22023_));
  AOI21_X1   g18887(.A1(new_n22022_), .A2(new_n22023_), .B(new_n21847_), .ZN(new_n22024_));
  NOR2_X1    g18888(.A1(new_n22024_), .A2(new_n12777_), .ZN(new_n22025_));
  NAND3_X1   g18889(.A1(new_n22021_), .A2(pi0628), .A3(pi1156), .ZN(new_n22026_));
  NAND3_X1   g18890(.A1(new_n22020_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n22027_));
  AOI21_X1   g18891(.A1(new_n22026_), .A2(new_n22027_), .B(new_n21847_), .ZN(new_n22028_));
  NAND3_X1   g18892(.A1(new_n22028_), .A2(pi0792), .A3(new_n22021_), .ZN(new_n22029_));
  NOR2_X1    g18893(.A1(new_n22029_), .A2(new_n22025_), .ZN(new_n22030_));
  INV_X1     g18894(.I(new_n22030_), .ZN(new_n22031_));
  NAND2_X1   g18895(.A1(new_n22029_), .A2(new_n22025_), .ZN(new_n22032_));
  NAND2_X1   g18896(.A1(new_n22031_), .A2(new_n22032_), .ZN(new_n22033_));
  NAND2_X1   g18897(.A1(new_n21848_), .A2(new_n14005_), .ZN(new_n22034_));
  NAND2_X1   g18898(.A1(new_n22034_), .A2(pi1157), .ZN(new_n22035_));
  AOI21_X1   g18899(.A1(new_n22033_), .A2(pi0647), .B(new_n22035_), .ZN(new_n22036_));
  AOI21_X1   g18900(.A1(new_n22031_), .A2(new_n22032_), .B(pi0647), .ZN(new_n22037_));
  NOR2_X1    g18901(.A1(new_n21847_), .A2(new_n14005_), .ZN(new_n22038_));
  NOR3_X1    g18902(.A1(new_n22037_), .A2(pi1157), .A3(new_n22038_), .ZN(new_n22039_));
  OAI21_X1   g18903(.A1(new_n22039_), .A2(new_n22036_), .B(pi0787), .ZN(new_n22040_));
  OAI21_X1   g18904(.A1(pi0787), .A2(new_n22033_), .B(new_n22040_), .ZN(new_n22041_));
  NOR2_X1    g18905(.A1(new_n21848_), .A2(new_n16372_), .ZN(new_n22042_));
  NOR2_X1    g18906(.A1(new_n21996_), .A2(new_n14142_), .ZN(new_n22043_));
  OAI21_X1   g18907(.A1(new_n22043_), .A2(new_n22042_), .B(new_n13994_), .ZN(new_n22044_));
  NOR2_X1    g18908(.A1(new_n21848_), .A2(new_n13994_), .ZN(new_n22045_));
  INV_X1     g18909(.I(new_n22045_), .ZN(new_n22046_));
  AOI21_X1   g18910(.A1(new_n22044_), .A2(new_n22046_), .B(new_n14210_), .ZN(new_n22047_));
  NOR2_X1    g18911(.A1(new_n21848_), .A2(new_n14211_), .ZN(new_n22048_));
  NOR2_X1    g18912(.A1(new_n22047_), .A2(new_n22048_), .ZN(new_n22049_));
  NOR2_X1    g18913(.A1(new_n14243_), .A2(pi0644), .ZN(new_n22050_));
  NOR2_X1    g18914(.A1(new_n22049_), .A2(new_n22050_), .ZN(new_n22051_));
  NAND2_X1   g18915(.A1(new_n22051_), .A2(pi0715), .ZN(new_n22052_));
  NAND2_X1   g18916(.A1(new_n22052_), .A2(new_n14204_), .ZN(new_n22053_));
  NAND2_X1   g18917(.A1(new_n22041_), .A2(new_n22053_), .ZN(new_n22054_));
  AOI21_X1   g18918(.A1(new_n21848_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n22055_));
  NOR2_X1    g18919(.A1(new_n22055_), .A2(pi0644), .ZN(new_n22056_));
  NOR3_X1    g18920(.A1(new_n22049_), .A2(new_n14200_), .A3(new_n22056_), .ZN(new_n22057_));
  OAI21_X1   g18921(.A1(new_n22041_), .A2(new_n22057_), .B(pi0644), .ZN(new_n22058_));
  AOI21_X1   g18922(.A1(new_n22058_), .A2(new_n22054_), .B(new_n12775_), .ZN(new_n22059_));
  NOR3_X1    g18923(.A1(new_n22049_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n22060_));
  OAI21_X1   g18924(.A1(new_n22049_), .A2(new_n22056_), .B(pi0790), .ZN(new_n22061_));
  NOR2_X1    g18925(.A1(new_n22061_), .A2(new_n19379_), .ZN(new_n22062_));
  OAI21_X1   g18926(.A1(new_n22062_), .A2(new_n22060_), .B(new_n22051_), .ZN(new_n22063_));
  NAND2_X1   g18927(.A1(new_n22044_), .A2(new_n22046_), .ZN(new_n22064_));
  INV_X1     g18928(.I(new_n22032_), .ZN(new_n22065_));
  OAI21_X1   g18929(.A1(new_n22065_), .A2(new_n22030_), .B(pi0647), .ZN(new_n22066_));
  NOR2_X1    g18930(.A1(new_n22065_), .A2(new_n22030_), .ZN(new_n22067_));
  INV_X1     g18931(.I(new_n22038_), .ZN(new_n22068_));
  OAI21_X1   g18932(.A1(new_n22067_), .A2(pi0647), .B(new_n22068_), .ZN(new_n22069_));
  NAND4_X1   g18933(.A1(new_n22066_), .A2(new_n14010_), .A3(pi1157), .A4(new_n22034_), .ZN(new_n22071_));
  NAND4_X1   g18934(.A1(new_n22066_), .A2(new_n14010_), .A3(pi1157), .A4(new_n22034_), .ZN(new_n22072_));
  NAND3_X1   g18935(.A1(new_n22072_), .A2(new_n22069_), .A3(new_n14011_), .ZN(new_n22073_));
  AOI21_X1   g18936(.A1(new_n22073_), .A2(new_n22071_), .B(new_n12776_), .ZN(new_n22074_));
  OAI21_X1   g18937(.A1(new_n22074_), .A2(new_n22064_), .B(new_n16576_), .ZN(new_n22075_));
  NAND2_X1   g18938(.A1(new_n22075_), .A2(new_n22063_), .ZN(new_n22076_));
  NOR2_X1    g18939(.A1(new_n22024_), .A2(new_n13976_), .ZN(new_n22077_));
  NOR2_X1    g18940(.A1(new_n22028_), .A2(pi0629), .ZN(new_n22078_));
  NOR2_X1    g18941(.A1(new_n22077_), .A2(new_n22078_), .ZN(new_n22079_));
  NOR2_X1    g18942(.A1(new_n22043_), .A2(new_n22042_), .ZN(new_n22080_));
  NOR2_X1    g18943(.A1(new_n22080_), .A2(new_n16874_), .ZN(new_n22081_));
  NOR3_X1    g18944(.A1(new_n13219_), .A2(pi0625), .A3(pi0725), .ZN(new_n22082_));
  INV_X1     g18945(.I(new_n22082_), .ZN(new_n22083_));
  NOR2_X1    g18946(.A1(new_n9992_), .A2(pi0183), .ZN(new_n22084_));
  NOR2_X1    g18947(.A1(new_n22084_), .A2(pi1153), .ZN(new_n22085_));
  NAND2_X1   g18948(.A1(new_n22083_), .A2(new_n22085_), .ZN(new_n22086_));
  INV_X1     g18949(.I(new_n22086_), .ZN(new_n22087_));
  NOR2_X1    g18950(.A1(new_n22087_), .A2(new_n13748_), .ZN(new_n22088_));
  AOI21_X1   g18951(.A1(new_n13218_), .A2(new_n17148_), .B(new_n22084_), .ZN(new_n22089_));
  INV_X1     g18952(.I(new_n22089_), .ZN(new_n22090_));
  AOI21_X1   g18953(.A1(new_n22083_), .A2(new_n22090_), .B(new_n13614_), .ZN(new_n22091_));
  INV_X1     g18954(.I(new_n22091_), .ZN(new_n22092_));
  NOR3_X1    g18955(.A1(new_n22092_), .A2(new_n13748_), .A3(new_n22090_), .ZN(new_n22093_));
  XNOR2_X1   g18956(.A1(new_n22093_), .A2(new_n22088_), .ZN(new_n22094_));
  NAND2_X1   g18957(.A1(new_n22094_), .A2(new_n14049_), .ZN(new_n22095_));
  NOR2_X1    g18958(.A1(new_n22095_), .A2(new_n14051_), .ZN(new_n22096_));
  INV_X1     g18959(.I(new_n22096_), .ZN(new_n22097_));
  NOR4_X1    g18960(.A1(new_n22097_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n22098_));
  NOR2_X1    g18961(.A1(new_n22098_), .A2(new_n14005_), .ZN(new_n22099_));
  XOR2_X1    g18962(.A1(new_n22099_), .A2(new_n14007_), .Z(new_n22100_));
  NAND2_X1   g18963(.A1(new_n22100_), .A2(new_n22084_), .ZN(new_n22101_));
  INV_X1     g18964(.I(new_n22084_), .ZN(new_n22102_));
  NOR2_X1    g18965(.A1(new_n22102_), .A2(pi0647), .ZN(new_n22103_));
  AOI21_X1   g18966(.A1(new_n22098_), .A2(pi0647), .B(new_n22103_), .ZN(new_n22104_));
  AOI21_X1   g18967(.A1(new_n22104_), .A2(pi1157), .B(new_n12776_), .ZN(new_n22105_));
  AOI22_X1   g18968(.A1(new_n22101_), .A2(new_n22105_), .B1(new_n12776_), .B2(new_n22098_), .ZN(new_n22106_));
  NOR2_X1    g18969(.A1(new_n22097_), .A2(new_n14163_), .ZN(new_n22107_));
  NOR2_X1    g18970(.A1(new_n21916_), .A2(new_n22084_), .ZN(new_n22108_));
  INV_X1     g18971(.I(new_n22108_), .ZN(new_n22109_));
  NAND3_X1   g18972(.A1(new_n22109_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n22110_));
  AOI21_X1   g18973(.A1(new_n22110_), .A2(new_n16444_), .B(new_n21917_), .ZN(new_n22111_));
  NOR2_X1    g18974(.A1(new_n22111_), .A2(new_n13801_), .ZN(new_n22112_));
  NOR2_X1    g18975(.A1(new_n22084_), .A2(pi1155), .ZN(new_n22113_));
  NOR3_X1    g18976(.A1(new_n21917_), .A2(new_n16444_), .A3(new_n22113_), .ZN(new_n22114_));
  NAND4_X1   g18977(.A1(new_n22114_), .A2(new_n22109_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n22115_));
  XOR2_X1    g18978(.A1(new_n22112_), .A2(new_n22115_), .Z(new_n22116_));
  NOR2_X1    g18979(.A1(new_n22116_), .A2(new_n13817_), .ZN(new_n22117_));
  OAI21_X1   g18980(.A1(new_n22117_), .A2(pi0618), .B(new_n9992_), .ZN(new_n22118_));
  NAND2_X1   g18981(.A1(new_n22118_), .A2(pi0781), .ZN(new_n22119_));
  OAI21_X1   g18982(.A1(new_n22117_), .A2(new_n9992_), .B(pi0618), .ZN(new_n22120_));
  NOR3_X1    g18983(.A1(new_n22120_), .A2(new_n13855_), .A3(new_n22116_), .ZN(new_n22121_));
  XOR2_X1    g18984(.A1(new_n22121_), .A2(new_n22119_), .Z(new_n22122_));
  NOR2_X1    g18985(.A1(new_n22122_), .A2(new_n13868_), .ZN(new_n22123_));
  OAI21_X1   g18986(.A1(new_n22123_), .A2(pi0619), .B(new_n9992_), .ZN(new_n22124_));
  NAND2_X1   g18987(.A1(new_n22124_), .A2(pi0789), .ZN(new_n22125_));
  OAI21_X1   g18988(.A1(new_n22123_), .A2(new_n9992_), .B(pi0619), .ZN(new_n22126_));
  NOR3_X1    g18989(.A1(new_n22126_), .A2(new_n13896_), .A3(new_n22122_), .ZN(new_n22127_));
  XOR2_X1    g18990(.A1(new_n22127_), .A2(new_n22125_), .Z(new_n22128_));
  NAND2_X1   g18991(.A1(new_n22128_), .A2(new_n13962_), .ZN(new_n22129_));
  XOR2_X1    g18992(.A1(new_n22129_), .A2(new_n18976_), .Z(new_n22130_));
  AOI22_X1   g18993(.A1(new_n22130_), .A2(new_n22084_), .B1(new_n16639_), .B2(new_n22107_), .ZN(new_n22131_));
  NOR2_X1    g18994(.A1(new_n22089_), .A2(new_n13203_), .ZN(new_n22132_));
  NAND2_X1   g18995(.A1(new_n22132_), .A2(pi0625), .ZN(new_n22133_));
  NAND3_X1   g18996(.A1(new_n22133_), .A2(pi1153), .A3(new_n22108_), .ZN(new_n22134_));
  NOR2_X1    g18997(.A1(new_n22087_), .A2(new_n14081_), .ZN(new_n22135_));
  AOI21_X1   g18998(.A1(new_n22135_), .A2(new_n22134_), .B(new_n13748_), .ZN(new_n22136_));
  NOR2_X1    g18999(.A1(new_n22109_), .A2(new_n22132_), .ZN(new_n22137_));
  INV_X1     g19000(.I(new_n22133_), .ZN(new_n22138_));
  OAI21_X1   g19001(.A1(new_n22137_), .A2(new_n22138_), .B(new_n22085_), .ZN(new_n22139_));
  NAND4_X1   g19002(.A1(new_n22139_), .A2(new_n13749_), .A3(new_n22092_), .A4(new_n22137_), .ZN(new_n22140_));
  XNOR2_X1   g19003(.A1(new_n22140_), .A2(new_n22136_), .ZN(new_n22141_));
  NAND2_X1   g19004(.A1(new_n22141_), .A2(new_n13801_), .ZN(new_n22142_));
  NOR2_X1    g19005(.A1(new_n22111_), .A2(pi0660), .ZN(new_n22146_));
  NOR2_X1    g19006(.A1(new_n22141_), .A2(new_n13766_), .ZN(new_n22147_));
  XOR2_X1    g19007(.A1(new_n22147_), .A2(new_n14090_), .Z(new_n22148_));
  NOR2_X1    g19008(.A1(new_n22094_), .A2(new_n13801_), .ZN(new_n22149_));
  NAND2_X1   g19009(.A1(new_n22148_), .A2(new_n22149_), .ZN(new_n22150_));
  OAI21_X1   g19010(.A1(new_n22150_), .A2(new_n22146_), .B(new_n22142_), .ZN(new_n22151_));
  NAND2_X1   g19011(.A1(new_n22151_), .A2(new_n13855_), .ZN(new_n22152_));
  INV_X1     g19012(.I(new_n22095_), .ZN(new_n22153_));
  NOR2_X1    g19013(.A1(new_n22151_), .A2(new_n13816_), .ZN(new_n22154_));
  XOR2_X1    g19014(.A1(new_n22154_), .A2(new_n13818_), .Z(new_n22155_));
  NAND2_X1   g19015(.A1(new_n22155_), .A2(new_n22153_), .ZN(new_n22156_));
  NAND3_X1   g19016(.A1(new_n22156_), .A2(new_n13823_), .A3(new_n22120_), .ZN(new_n22157_));
  NAND3_X1   g19017(.A1(new_n22157_), .A2(new_n13823_), .A3(new_n22118_), .ZN(new_n22158_));
  NOR2_X1    g19018(.A1(new_n22151_), .A2(new_n13817_), .ZN(new_n22159_));
  XOR2_X1    g19019(.A1(new_n22159_), .A2(new_n13818_), .Z(new_n22160_));
  NAND4_X1   g19020(.A1(new_n22158_), .A2(pi0781), .A3(new_n22153_), .A4(new_n22160_), .ZN(new_n22161_));
  NAND2_X1   g19021(.A1(new_n22161_), .A2(new_n22152_), .ZN(new_n22162_));
  NOR2_X1    g19022(.A1(new_n22162_), .A2(new_n13860_), .ZN(new_n22163_));
  XOR2_X1    g19023(.A1(new_n22163_), .A2(new_n13904_), .Z(new_n22164_));
  NOR2_X1    g19024(.A1(new_n22164_), .A2(new_n22097_), .ZN(new_n22165_));
  NAND2_X1   g19025(.A1(new_n22126_), .A2(new_n13884_), .ZN(new_n22166_));
  INV_X1     g19026(.I(new_n22162_), .ZN(new_n22167_));
  AOI21_X1   g19027(.A1(new_n22167_), .A2(new_n14143_), .B(pi0789), .ZN(new_n22168_));
  OAI21_X1   g19028(.A1(new_n22165_), .A2(new_n22166_), .B(new_n22168_), .ZN(new_n22169_));
  NOR2_X1    g19029(.A1(new_n22162_), .A2(new_n13868_), .ZN(new_n22170_));
  XOR2_X1    g19030(.A1(new_n22170_), .A2(new_n13903_), .Z(new_n22171_));
  NAND2_X1   g19031(.A1(new_n22124_), .A2(new_n19018_), .ZN(new_n22172_));
  AOI21_X1   g19032(.A1(new_n22171_), .A2(new_n22096_), .B(new_n22172_), .ZN(new_n22173_));
  AOI21_X1   g19033(.A1(new_n22169_), .A2(new_n22173_), .B(new_n22131_), .ZN(new_n22174_));
  NAND2_X1   g19034(.A1(new_n22128_), .A2(new_n16372_), .ZN(new_n22175_));
  OAI21_X1   g19035(.A1(new_n16372_), .A2(new_n22084_), .B(new_n22175_), .ZN(new_n22176_));
  NAND3_X1   g19036(.A1(new_n22176_), .A2(new_n18929_), .A3(new_n22107_), .ZN(new_n22177_));
  NAND2_X1   g19037(.A1(new_n22177_), .A2(new_n16569_), .ZN(new_n22178_));
  XOR2_X1    g19038(.A1(new_n22178_), .A2(new_n16572_), .Z(new_n22179_));
  AOI21_X1   g19039(.A1(new_n19022_), .A2(new_n22177_), .B(new_n22179_), .ZN(new_n22180_));
  NAND2_X1   g19040(.A1(new_n22128_), .A2(new_n13963_), .ZN(new_n22181_));
  XNOR2_X1   g19041(.A1(new_n22181_), .A2(new_n19028_), .ZN(new_n22182_));
  NOR3_X1    g19042(.A1(new_n22182_), .A2(new_n16424_), .A3(new_n22102_), .ZN(new_n22183_));
  OAI21_X1   g19043(.A1(new_n22180_), .A2(new_n16574_), .B(new_n22183_), .ZN(new_n22184_));
  NOR2_X1    g19044(.A1(new_n22176_), .A2(new_n13994_), .ZN(new_n22185_));
  XNOR2_X1   g19045(.A1(new_n22185_), .A2(new_n19033_), .ZN(new_n22186_));
  AOI22_X1   g19046(.A1(new_n22186_), .A2(new_n22084_), .B1(new_n14206_), .B2(new_n22104_), .ZN(new_n22187_));
  NOR3_X1    g19047(.A1(new_n22187_), .A2(new_n14010_), .A3(new_n22101_), .ZN(new_n22188_));
  OAI22_X1   g19048(.A1(new_n22174_), .A2(new_n22184_), .B1(new_n12776_), .B2(new_n22188_), .ZN(new_n22189_));
  NAND2_X1   g19049(.A1(new_n22189_), .A2(pi0644), .ZN(new_n22190_));
  XOR2_X1    g19050(.A1(new_n22190_), .A2(new_n14205_), .Z(new_n22191_));
  NOR2_X1    g19051(.A1(new_n22191_), .A2(new_n22106_), .ZN(new_n22192_));
  NOR2_X1    g19052(.A1(new_n22176_), .A2(new_n18968_), .ZN(new_n22193_));
  NAND2_X1   g19053(.A1(new_n18967_), .A2(new_n22084_), .ZN(new_n22194_));
  XOR2_X1    g19054(.A1(new_n22193_), .A2(new_n22194_), .Z(new_n22195_));
  NAND2_X1   g19055(.A1(new_n22195_), .A2(pi0715), .ZN(new_n22196_));
  XOR2_X1    g19056(.A1(new_n22196_), .A2(new_n14205_), .Z(new_n22197_));
  OAI21_X1   g19057(.A1(new_n22197_), .A2(new_n22102_), .B(new_n14203_), .ZN(new_n22198_));
  NAND2_X1   g19058(.A1(new_n22195_), .A2(pi0644), .ZN(new_n22199_));
  XOR2_X1    g19059(.A1(new_n22199_), .A2(new_n14217_), .Z(new_n22200_));
  AOI21_X1   g19060(.A1(new_n22200_), .A2(new_n22084_), .B(pi1160), .ZN(new_n22201_));
  OAI21_X1   g19061(.A1(new_n22192_), .A2(new_n22198_), .B(new_n22201_), .ZN(new_n22202_));
  NAND2_X1   g19062(.A1(new_n22189_), .A2(pi0715), .ZN(new_n22203_));
  XOR2_X1    g19063(.A1(new_n22203_), .A2(new_n14205_), .Z(new_n22204_));
  NOR2_X1    g19064(.A1(new_n22204_), .A2(new_n22106_), .ZN(new_n22205_));
  AOI21_X1   g19065(.A1(new_n22202_), .A2(new_n22205_), .B(new_n14799_), .ZN(new_n22206_));
  XOR2_X1    g19066(.A1(new_n22206_), .A2(new_n14800_), .Z(new_n22207_));
  OAI21_X1   g19067(.A1(new_n7240_), .A2(pi0183), .B(new_n14799_), .ZN(new_n22208_));
  NOR2_X1    g19068(.A1(new_n22189_), .A2(new_n22208_), .ZN(new_n22209_));
  AOI21_X1   g19069(.A1(new_n22207_), .A2(new_n22209_), .B(po1038), .ZN(new_n22210_));
  NOR3_X1    g19070(.A1(new_n22081_), .A2(new_n22079_), .A3(new_n22210_), .ZN(new_n22211_));
  OAI21_X1   g19071(.A1(new_n22059_), .A2(new_n22076_), .B(new_n22211_), .ZN(new_n22212_));
  NOR2_X1    g19072(.A1(new_n22212_), .A2(new_n22017_), .ZN(po0340));
  NAND2_X1   g19073(.A1(new_n13627_), .A2(new_n9471_), .ZN(new_n22214_));
  INV_X1     g19074(.I(new_n22214_), .ZN(new_n22215_));
  AOI21_X1   g19075(.A1(new_n9471_), .A2(new_n17735_), .B(pi0038), .ZN(new_n22216_));
  NOR2_X1    g19076(.A1(new_n9471_), .A2(new_n17735_), .ZN(new_n22217_));
  OAI21_X1   g19077(.A1(new_n20007_), .A2(new_n22217_), .B(pi0038), .ZN(new_n22218_));
  INV_X1     g19078(.I(new_n22218_), .ZN(new_n22219_));
  AOI21_X1   g19079(.A1(new_n13097_), .A2(new_n22216_), .B(new_n22219_), .ZN(new_n22220_));
  NOR2_X1    g19080(.A1(new_n3289_), .A2(pi0184), .ZN(new_n22221_));
  AOI21_X1   g19081(.A1(new_n22220_), .A2(new_n3289_), .B(new_n22221_), .ZN(new_n22222_));
  NAND2_X1   g19082(.A1(new_n22222_), .A2(new_n13776_), .ZN(new_n22223_));
  OAI21_X1   g19083(.A1(new_n15147_), .A2(new_n22215_), .B(new_n22223_), .ZN(new_n22224_));
  NAND2_X1   g19084(.A1(new_n22224_), .A2(pi0609), .ZN(new_n22225_));
  NAND2_X1   g19085(.A1(new_n22225_), .A2(pi0785), .ZN(new_n22226_));
  AOI21_X1   g19086(.A1(new_n22214_), .A2(new_n14467_), .B(pi0609), .ZN(new_n22227_));
  NOR2_X1    g19087(.A1(new_n22227_), .A2(new_n22223_), .ZN(new_n22228_));
  NAND2_X1   g19088(.A1(new_n22215_), .A2(new_n13775_), .ZN(new_n22229_));
  OAI21_X1   g19089(.A1(new_n13775_), .A2(new_n22222_), .B(new_n22229_), .ZN(new_n22230_));
  NAND3_X1   g19090(.A1(new_n22230_), .A2(pi0785), .A3(new_n22228_), .ZN(new_n22231_));
  XNOR2_X1   g19091(.A1(new_n22226_), .A2(new_n22231_), .ZN(new_n22232_));
  NAND2_X1   g19092(.A1(new_n22232_), .A2(pi0618), .ZN(new_n22233_));
  XOR2_X1    g19093(.A1(new_n22233_), .A2(new_n13819_), .Z(new_n22234_));
  NAND2_X1   g19094(.A1(new_n22234_), .A2(new_n22215_), .ZN(new_n22235_));
  NAND2_X1   g19095(.A1(new_n22235_), .A2(pi0781), .ZN(new_n22236_));
  NAND2_X1   g19096(.A1(new_n22232_), .A2(pi1154), .ZN(new_n22237_));
  XOR2_X1    g19097(.A1(new_n22237_), .A2(new_n13819_), .Z(new_n22238_));
  NAND2_X1   g19098(.A1(new_n22238_), .A2(new_n22215_), .ZN(new_n22239_));
  NOR3_X1    g19099(.A1(new_n22239_), .A2(new_n13855_), .A3(new_n22232_), .ZN(new_n22240_));
  XNOR2_X1   g19100(.A1(new_n22240_), .A2(new_n22236_), .ZN(new_n22241_));
  NAND3_X1   g19101(.A1(new_n22241_), .A2(pi0619), .A3(pi1159), .ZN(new_n22242_));
  XOR2_X1    g19102(.A1(new_n22240_), .A2(new_n22236_), .Z(new_n22243_));
  NAND3_X1   g19103(.A1(new_n22243_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n22244_));
  AOI21_X1   g19104(.A1(new_n22242_), .A2(new_n22244_), .B(new_n22214_), .ZN(new_n22245_));
  NOR2_X1    g19105(.A1(new_n22215_), .A2(new_n13880_), .ZN(new_n22246_));
  OAI21_X1   g19106(.A1(new_n13721_), .A2(new_n17730_), .B(new_n9471_), .ZN(new_n22247_));
  NAND2_X1   g19107(.A1(new_n16715_), .A2(new_n9471_), .ZN(new_n22248_));
  NAND4_X1   g19108(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n22247_), .A4(new_n22248_), .ZN(new_n22249_));
  NAND2_X1   g19109(.A1(new_n22249_), .A2(new_n14424_), .ZN(new_n22250_));
  NAND2_X1   g19110(.A1(new_n22250_), .A2(pi0184), .ZN(new_n22251_));
  OAI21_X1   g19111(.A1(new_n22251_), .A2(new_n22214_), .B(new_n3290_), .ZN(new_n22252_));
  NAND2_X1   g19112(.A1(new_n22252_), .A2(pi0737), .ZN(new_n22253_));
  NAND2_X1   g19113(.A1(new_n22253_), .A2(pi0625), .ZN(new_n22254_));
  XOR2_X1    g19114(.A1(new_n22254_), .A2(new_n13620_), .Z(new_n22255_));
  NAND2_X1   g19115(.A1(new_n22255_), .A2(new_n22215_), .ZN(new_n22256_));
  NAND2_X1   g19116(.A1(new_n22256_), .A2(pi0778), .ZN(new_n22257_));
  NAND2_X1   g19117(.A1(new_n22253_), .A2(pi1153), .ZN(new_n22258_));
  XOR2_X1    g19118(.A1(new_n22258_), .A2(new_n13620_), .Z(new_n22259_));
  NAND2_X1   g19119(.A1(new_n22259_), .A2(new_n22215_), .ZN(new_n22260_));
  NOR3_X1    g19120(.A1(new_n22260_), .A2(new_n13748_), .A3(new_n22253_), .ZN(new_n22261_));
  XNOR2_X1   g19121(.A1(new_n22261_), .A2(new_n22257_), .ZN(new_n22262_));
  NOR2_X1    g19122(.A1(new_n22214_), .A2(new_n13805_), .ZN(new_n22263_));
  AOI21_X1   g19123(.A1(new_n22262_), .A2(new_n13805_), .B(new_n22263_), .ZN(new_n22264_));
  AOI21_X1   g19124(.A1(new_n22264_), .A2(new_n13880_), .B(new_n22246_), .ZN(new_n22265_));
  NOR2_X1    g19125(.A1(new_n13453_), .A2(new_n9471_), .ZN(new_n22266_));
  XOR2_X1    g19126(.A1(new_n22266_), .A2(new_n22217_), .Z(new_n22267_));
  NAND2_X1   g19127(.A1(new_n22267_), .A2(new_n13521_), .ZN(new_n22268_));
  NAND3_X1   g19128(.A1(new_n14270_), .A2(pi0184), .A3(pi0777), .ZN(new_n22269_));
  NAND3_X1   g19129(.A1(new_n14272_), .A2(new_n9471_), .A3(pi0777), .ZN(new_n22270_));
  AOI21_X1   g19130(.A1(new_n22269_), .A2(new_n22270_), .B(new_n13152_), .ZN(new_n22271_));
  NAND3_X1   g19131(.A1(new_n13198_), .A2(pi0184), .A3(pi0777), .ZN(new_n22272_));
  NAND3_X1   g19132(.A1(new_n13200_), .A2(pi0184), .A3(new_n17735_), .ZN(new_n22273_));
  AOI21_X1   g19133(.A1(new_n22273_), .A2(new_n22272_), .B(new_n13191_), .ZN(new_n22274_));
  OAI21_X1   g19134(.A1(new_n22271_), .A2(new_n3262_), .B(new_n22274_), .ZN(new_n22275_));
  NAND3_X1   g19135(.A1(new_n22268_), .A2(new_n3183_), .A3(new_n22275_), .ZN(new_n22276_));
  NOR2_X1    g19136(.A1(new_n14284_), .A2(new_n17735_), .ZN(new_n22277_));
  XOR2_X1    g19137(.A1(new_n22277_), .A2(new_n22217_), .Z(new_n22278_));
  NAND3_X1   g19138(.A1(new_n22276_), .A2(new_n22278_), .A3(new_n13359_), .ZN(new_n22279_));
  NAND3_X1   g19139(.A1(new_n22279_), .A2(new_n17730_), .A3(new_n3290_), .ZN(new_n22280_));
  OAI21_X1   g19140(.A1(new_n15587_), .A2(new_n9471_), .B(new_n17735_), .ZN(new_n22281_));
  NAND2_X1   g19141(.A1(new_n22281_), .A2(new_n13209_), .ZN(new_n22282_));
  NOR2_X1    g19142(.A1(new_n13105_), .A2(pi0777), .ZN(new_n22283_));
  INV_X1     g19143(.I(new_n22283_), .ZN(new_n22284_));
  NAND2_X1   g19144(.A1(new_n22284_), .A2(new_n16751_), .ZN(new_n22285_));
  NAND4_X1   g19145(.A1(new_n5503_), .A2(new_n22285_), .A3(pi0184), .A4(new_n3290_), .ZN(new_n22286_));
  AOI21_X1   g19146(.A1(new_n22282_), .A2(new_n3259_), .B(new_n22286_), .ZN(new_n22287_));
  AOI21_X1   g19147(.A1(new_n22280_), .A2(new_n22287_), .B(pi0737), .ZN(new_n22288_));
  NOR2_X1    g19148(.A1(new_n22288_), .A2(new_n22220_), .ZN(new_n22289_));
  INV_X1     g19149(.I(new_n22289_), .ZN(new_n22290_));
  INV_X1     g19150(.I(new_n22222_), .ZN(new_n22291_));
  NOR2_X1    g19151(.A1(new_n22289_), .A2(new_n13613_), .ZN(new_n22292_));
  XOR2_X1    g19152(.A1(new_n22292_), .A2(new_n13615_), .Z(new_n22293_));
  NAND2_X1   g19153(.A1(new_n22260_), .A2(new_n14081_), .ZN(new_n22294_));
  AOI21_X1   g19154(.A1(new_n22293_), .A2(new_n22291_), .B(new_n22294_), .ZN(new_n22295_));
  INV_X1     g19155(.I(new_n22295_), .ZN(new_n22296_));
  NOR2_X1    g19156(.A1(new_n22289_), .A2(new_n13614_), .ZN(new_n22297_));
  XOR2_X1    g19157(.A1(new_n22297_), .A2(new_n13615_), .Z(new_n22298_));
  AOI21_X1   g19158(.A1(new_n22298_), .A2(new_n22291_), .B(pi0608), .ZN(new_n22299_));
  NAND2_X1   g19159(.A1(new_n22296_), .A2(new_n22299_), .ZN(new_n22300_));
  NOR2_X1    g19160(.A1(new_n22256_), .A2(new_n13748_), .ZN(new_n22301_));
  AOI22_X1   g19161(.A1(new_n22300_), .A2(new_n22301_), .B1(new_n13748_), .B2(new_n22290_), .ZN(new_n22302_));
  AOI21_X1   g19162(.A1(new_n22302_), .A2(pi1155), .B(new_n14694_), .ZN(new_n22303_));
  INV_X1     g19163(.I(new_n22299_), .ZN(new_n22304_));
  NOR2_X1    g19164(.A1(new_n22304_), .A2(new_n22295_), .ZN(new_n22305_));
  INV_X1     g19165(.I(new_n22301_), .ZN(new_n22306_));
  OAI22_X1   g19166(.A1(new_n22305_), .A2(new_n22306_), .B1(pi0778), .B2(new_n22289_), .ZN(new_n22307_));
  NOR3_X1    g19167(.A1(new_n22307_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n22308_));
  OAI21_X1   g19168(.A1(new_n22308_), .A2(new_n22303_), .B(new_n22262_), .ZN(new_n22309_));
  NAND2_X1   g19169(.A1(new_n22225_), .A2(pi0660), .ZN(new_n22310_));
  INV_X1     g19170(.I(new_n22310_), .ZN(new_n22311_));
  NOR2_X1    g19171(.A1(new_n22228_), .A2(pi0660), .ZN(new_n22312_));
  INV_X1     g19172(.I(new_n22312_), .ZN(new_n22313_));
  AOI21_X1   g19173(.A1(new_n22309_), .A2(new_n22311_), .B(new_n22313_), .ZN(new_n22314_));
  NOR2_X1    g19174(.A1(new_n22307_), .A2(new_n13766_), .ZN(new_n22315_));
  NOR2_X1    g19175(.A1(new_n22315_), .A2(new_n14694_), .ZN(new_n22316_));
  NAND2_X1   g19176(.A1(new_n22315_), .A2(new_n14694_), .ZN(new_n22317_));
  INV_X1     g19177(.I(new_n22317_), .ZN(new_n22318_));
  INV_X1     g19178(.I(new_n22262_), .ZN(new_n22319_));
  NOR2_X1    g19179(.A1(new_n22319_), .A2(new_n13801_), .ZN(new_n22320_));
  OAI21_X1   g19180(.A1(new_n22318_), .A2(new_n22316_), .B(new_n22320_), .ZN(new_n22321_));
  OAI22_X1   g19181(.A1(new_n22321_), .A2(new_n22314_), .B1(pi0785), .B2(new_n22302_), .ZN(new_n22322_));
  NAND3_X1   g19182(.A1(new_n22322_), .A2(pi0618), .A3(pi1154), .ZN(new_n22323_));
  NAND3_X1   g19183(.A1(new_n22307_), .A2(pi0609), .A3(pi1155), .ZN(new_n22324_));
  NAND3_X1   g19184(.A1(new_n22302_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n22325_));
  AOI21_X1   g19185(.A1(new_n22324_), .A2(new_n22325_), .B(new_n22319_), .ZN(new_n22326_));
  OAI21_X1   g19186(.A1(new_n22326_), .A2(new_n22310_), .B(new_n22312_), .ZN(new_n22327_));
  NAND2_X1   g19187(.A1(new_n22302_), .A2(pi0609), .ZN(new_n22328_));
  NAND2_X1   g19188(.A1(new_n22328_), .A2(new_n14090_), .ZN(new_n22329_));
  INV_X1     g19189(.I(new_n22320_), .ZN(new_n22330_));
  AOI21_X1   g19190(.A1(new_n22317_), .A2(new_n22329_), .B(new_n22330_), .ZN(new_n22331_));
  AOI22_X1   g19191(.A1(new_n22327_), .A2(new_n22331_), .B1(new_n13801_), .B2(new_n22307_), .ZN(new_n22332_));
  NAND3_X1   g19192(.A1(new_n22332_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n22333_));
  AOI21_X1   g19193(.A1(new_n22323_), .A2(new_n22333_), .B(new_n22264_), .ZN(new_n22334_));
  NAND2_X1   g19194(.A1(new_n22235_), .A2(pi0627), .ZN(new_n22335_));
  OAI21_X1   g19195(.A1(new_n22334_), .A2(new_n22335_), .B(pi0781), .ZN(new_n22336_));
  INV_X1     g19196(.I(new_n22264_), .ZN(new_n22337_));
  AOI21_X1   g19197(.A1(new_n22332_), .A2(pi0618), .B(new_n13819_), .ZN(new_n22338_));
  NOR3_X1    g19198(.A1(new_n22322_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n22339_));
  OAI21_X1   g19199(.A1(new_n22339_), .A2(new_n22338_), .B(new_n22337_), .ZN(new_n22340_));
  AND3_X2    g19200(.A1(new_n22322_), .A2(new_n19177_), .A3(new_n22239_), .Z(new_n22341_));
  NAND3_X1   g19201(.A1(new_n22336_), .A2(new_n22340_), .A3(new_n22341_), .ZN(new_n22342_));
  AOI21_X1   g19202(.A1(new_n22332_), .A2(pi1154), .B(new_n13819_), .ZN(new_n22343_));
  NOR3_X1    g19203(.A1(new_n22322_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n22344_));
  OAI21_X1   g19204(.A1(new_n22344_), .A2(new_n22343_), .B(new_n22337_), .ZN(new_n22345_));
  INV_X1     g19205(.I(new_n22335_), .ZN(new_n22346_));
  AOI21_X1   g19206(.A1(new_n22345_), .A2(new_n22346_), .B(new_n13855_), .ZN(new_n22347_));
  NAND4_X1   g19207(.A1(new_n22340_), .A2(new_n19177_), .A3(new_n22239_), .A4(new_n22322_), .ZN(new_n22348_));
  NAND2_X1   g19208(.A1(new_n22348_), .A2(new_n22347_), .ZN(new_n22349_));
  NAND2_X1   g19209(.A1(new_n22349_), .A2(new_n22342_), .ZN(new_n22350_));
  NAND3_X1   g19210(.A1(new_n22350_), .A2(pi0619), .A3(pi1159), .ZN(new_n22351_));
  NAND4_X1   g19211(.A1(new_n22349_), .A2(new_n22342_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n22352_));
  AOI21_X1   g19212(.A1(new_n22351_), .A2(new_n22352_), .B(new_n22265_), .ZN(new_n22353_));
  OAI21_X1   g19213(.A1(new_n22353_), .A2(new_n20003_), .B(new_n22245_), .ZN(new_n22354_));
  NAND2_X1   g19214(.A1(new_n22350_), .A2(new_n13896_), .ZN(new_n22355_));
  NOR2_X1    g19215(.A1(new_n22245_), .A2(new_n13896_), .ZN(new_n22356_));
  NAND3_X1   g19216(.A1(new_n22241_), .A2(pi0619), .A3(pi1159), .ZN(new_n22357_));
  NAND3_X1   g19217(.A1(new_n22243_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n22358_));
  NAND2_X1   g19218(.A1(new_n22357_), .A2(new_n22358_), .ZN(new_n22359_));
  NAND4_X1   g19219(.A1(new_n22359_), .A2(pi0789), .A3(new_n22215_), .A4(new_n22241_), .ZN(new_n22360_));
  OR2_X2     g19220(.A1(new_n22360_), .A2(new_n22356_), .Z(new_n22361_));
  NAND2_X1   g19221(.A1(new_n22360_), .A2(new_n22356_), .ZN(new_n22362_));
  NAND2_X1   g19222(.A1(new_n22361_), .A2(new_n22362_), .ZN(new_n22363_));
  NAND3_X1   g19223(.A1(new_n22363_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n22364_));
  NAND4_X1   g19224(.A1(new_n22361_), .A2(new_n13901_), .A3(new_n13962_), .A4(new_n22362_), .ZN(new_n22365_));
  AOI21_X1   g19225(.A1(new_n22364_), .A2(new_n22365_), .B(new_n22214_), .ZN(new_n22366_));
  NOR2_X1    g19226(.A1(new_n22214_), .A2(new_n13919_), .ZN(new_n22367_));
  NAND2_X1   g19227(.A1(new_n22265_), .A2(new_n13919_), .ZN(new_n22368_));
  INV_X1     g19228(.I(new_n22368_), .ZN(new_n22369_));
  NOR2_X1    g19229(.A1(new_n22369_), .A2(new_n22367_), .ZN(new_n22370_));
  NOR2_X1    g19230(.A1(new_n22370_), .A2(new_n14162_), .ZN(new_n22371_));
  OAI21_X1   g19231(.A1(new_n22366_), .A2(new_n22371_), .B(new_n19204_), .ZN(new_n22372_));
  NOR2_X1    g19232(.A1(new_n22363_), .A2(new_n19208_), .ZN(new_n22373_));
  XNOR2_X1   g19233(.A1(new_n22373_), .A2(new_n19028_), .ZN(new_n22374_));
  NOR2_X1    g19234(.A1(new_n22214_), .A2(new_n15479_), .ZN(new_n22375_));
  NAND4_X1   g19235(.A1(new_n22355_), .A2(new_n22372_), .A3(new_n22374_), .A4(new_n22375_), .ZN(new_n22376_));
  NAND2_X1   g19236(.A1(new_n22354_), .A2(new_n22376_), .ZN(new_n22377_));
  INV_X1     g19237(.I(new_n22265_), .ZN(new_n22378_));
  NAND3_X1   g19238(.A1(new_n22349_), .A2(new_n22342_), .A3(pi0619), .ZN(new_n22379_));
  XOR2_X1    g19239(.A1(new_n22379_), .A2(new_n13904_), .Z(new_n22380_));
  NAND2_X1   g19240(.A1(new_n22359_), .A2(new_n22215_), .ZN(new_n22381_));
  NAND2_X1   g19241(.A1(new_n22381_), .A2(new_n20173_), .ZN(new_n22382_));
  AOI21_X1   g19242(.A1(new_n22380_), .A2(new_n22378_), .B(new_n22382_), .ZN(new_n22383_));
  AOI21_X1   g19243(.A1(new_n22377_), .A2(new_n22383_), .B(pi0792), .ZN(new_n22384_));
  NOR2_X1    g19244(.A1(new_n22215_), .A2(new_n13966_), .ZN(new_n22385_));
  NOR3_X1    g19245(.A1(new_n22369_), .A2(new_n13965_), .A3(new_n22367_), .ZN(new_n22386_));
  NOR2_X1    g19246(.A1(new_n22386_), .A2(new_n22385_), .ZN(new_n22387_));
  INV_X1     g19247(.I(new_n22387_), .ZN(new_n22388_));
  NAND3_X1   g19248(.A1(new_n22388_), .A2(pi0628), .A3(pi1156), .ZN(new_n22389_));
  NAND3_X1   g19249(.A1(new_n22387_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n22390_));
  AOI21_X1   g19250(.A1(new_n22389_), .A2(new_n22390_), .B(new_n22214_), .ZN(new_n22391_));
  NOR2_X1    g19251(.A1(new_n22391_), .A2(new_n12777_), .ZN(new_n22392_));
  NAND3_X1   g19252(.A1(new_n22388_), .A2(pi0628), .A3(pi1156), .ZN(new_n22393_));
  NAND3_X1   g19253(.A1(new_n22387_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n22394_));
  AOI21_X1   g19254(.A1(new_n22393_), .A2(new_n22394_), .B(new_n22214_), .ZN(new_n22395_));
  NAND3_X1   g19255(.A1(new_n22395_), .A2(pi0792), .A3(new_n22388_), .ZN(new_n22396_));
  NOR2_X1    g19256(.A1(new_n22396_), .A2(new_n22392_), .ZN(new_n22397_));
  INV_X1     g19257(.I(new_n22397_), .ZN(new_n22398_));
  NAND2_X1   g19258(.A1(new_n22396_), .A2(new_n22392_), .ZN(new_n22399_));
  NAND2_X1   g19259(.A1(new_n22398_), .A2(new_n22399_), .ZN(new_n22400_));
  NAND2_X1   g19260(.A1(new_n22215_), .A2(new_n14005_), .ZN(new_n22401_));
  NAND2_X1   g19261(.A1(new_n22401_), .A2(pi1157), .ZN(new_n22402_));
  AOI21_X1   g19262(.A1(new_n22400_), .A2(pi0647), .B(new_n22402_), .ZN(new_n22403_));
  AOI21_X1   g19263(.A1(new_n22398_), .A2(new_n22399_), .B(pi0647), .ZN(new_n22404_));
  NOR2_X1    g19264(.A1(new_n22214_), .A2(new_n14005_), .ZN(new_n22405_));
  NOR3_X1    g19265(.A1(new_n22404_), .A2(pi1157), .A3(new_n22405_), .ZN(new_n22406_));
  OAI21_X1   g19266(.A1(new_n22406_), .A2(new_n22403_), .B(pi0787), .ZN(new_n22407_));
  OAI21_X1   g19267(.A1(pi0787), .A2(new_n22400_), .B(new_n22407_), .ZN(new_n22408_));
  NOR2_X1    g19268(.A1(new_n22215_), .A2(new_n16372_), .ZN(new_n22409_));
  NOR2_X1    g19269(.A1(new_n22363_), .A2(new_n14142_), .ZN(new_n22410_));
  OAI21_X1   g19270(.A1(new_n22410_), .A2(new_n22409_), .B(new_n13994_), .ZN(new_n22411_));
  NOR2_X1    g19271(.A1(new_n22215_), .A2(new_n13994_), .ZN(new_n22412_));
  INV_X1     g19272(.I(new_n22412_), .ZN(new_n22413_));
  AOI21_X1   g19273(.A1(new_n22411_), .A2(new_n22413_), .B(new_n14210_), .ZN(new_n22414_));
  NOR2_X1    g19274(.A1(new_n22215_), .A2(new_n14211_), .ZN(new_n22415_));
  NOR2_X1    g19275(.A1(new_n22414_), .A2(new_n22415_), .ZN(new_n22416_));
  NOR2_X1    g19276(.A1(new_n14243_), .A2(pi0644), .ZN(new_n22417_));
  NOR2_X1    g19277(.A1(new_n22416_), .A2(new_n22417_), .ZN(new_n22418_));
  NAND2_X1   g19278(.A1(new_n22418_), .A2(pi0715), .ZN(new_n22419_));
  NAND2_X1   g19279(.A1(new_n22419_), .A2(new_n14204_), .ZN(new_n22420_));
  NAND2_X1   g19280(.A1(new_n22408_), .A2(new_n22420_), .ZN(new_n22421_));
  AOI21_X1   g19281(.A1(new_n22215_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n22422_));
  NOR2_X1    g19282(.A1(new_n22422_), .A2(pi0644), .ZN(new_n22423_));
  NOR3_X1    g19283(.A1(new_n22416_), .A2(new_n14200_), .A3(new_n22423_), .ZN(new_n22424_));
  OAI21_X1   g19284(.A1(new_n22408_), .A2(new_n22424_), .B(pi0644), .ZN(new_n22425_));
  AOI21_X1   g19285(.A1(new_n22425_), .A2(new_n22421_), .B(new_n12775_), .ZN(new_n22426_));
  NOR3_X1    g19286(.A1(new_n22416_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n22427_));
  OAI21_X1   g19287(.A1(new_n22416_), .A2(new_n22423_), .B(pi0790), .ZN(new_n22428_));
  NOR2_X1    g19288(.A1(new_n22428_), .A2(new_n19379_), .ZN(new_n22429_));
  OAI21_X1   g19289(.A1(new_n22429_), .A2(new_n22427_), .B(new_n22418_), .ZN(new_n22430_));
  NAND2_X1   g19290(.A1(new_n22411_), .A2(new_n22413_), .ZN(new_n22431_));
  INV_X1     g19291(.I(new_n22399_), .ZN(new_n22432_));
  OAI21_X1   g19292(.A1(new_n22432_), .A2(new_n22397_), .B(pi0647), .ZN(new_n22433_));
  NOR2_X1    g19293(.A1(new_n22432_), .A2(new_n22397_), .ZN(new_n22434_));
  INV_X1     g19294(.I(new_n22405_), .ZN(new_n22435_));
  OAI21_X1   g19295(.A1(new_n22434_), .A2(pi0647), .B(new_n22435_), .ZN(new_n22436_));
  NAND4_X1   g19296(.A1(new_n22433_), .A2(new_n14010_), .A3(pi1157), .A4(new_n22401_), .ZN(new_n22438_));
  NAND4_X1   g19297(.A1(new_n22433_), .A2(new_n14010_), .A3(pi1157), .A4(new_n22401_), .ZN(new_n22439_));
  NAND3_X1   g19298(.A1(new_n22439_), .A2(new_n22436_), .A3(new_n14011_), .ZN(new_n22440_));
  AOI21_X1   g19299(.A1(new_n22440_), .A2(new_n22438_), .B(new_n12776_), .ZN(new_n22441_));
  OAI21_X1   g19300(.A1(new_n22441_), .A2(new_n22431_), .B(new_n16576_), .ZN(new_n22442_));
  NAND2_X1   g19301(.A1(new_n22442_), .A2(new_n22430_), .ZN(new_n22443_));
  NOR2_X1    g19302(.A1(new_n22391_), .A2(new_n13976_), .ZN(new_n22444_));
  NOR2_X1    g19303(.A1(new_n22395_), .A2(pi0629), .ZN(new_n22445_));
  NOR2_X1    g19304(.A1(new_n22444_), .A2(new_n22445_), .ZN(new_n22446_));
  NOR2_X1    g19305(.A1(new_n22410_), .A2(new_n22409_), .ZN(new_n22447_));
  NOR2_X1    g19306(.A1(new_n22447_), .A2(new_n16874_), .ZN(new_n22448_));
  NOR3_X1    g19307(.A1(new_n13219_), .A2(pi0625), .A3(pi0737), .ZN(new_n22449_));
  INV_X1     g19308(.I(new_n22449_), .ZN(new_n22450_));
  NOR2_X1    g19309(.A1(new_n9992_), .A2(pi0184), .ZN(new_n22451_));
  NOR2_X1    g19310(.A1(new_n22451_), .A2(pi1153), .ZN(new_n22452_));
  NAND2_X1   g19311(.A1(new_n22450_), .A2(new_n22452_), .ZN(new_n22453_));
  INV_X1     g19312(.I(new_n22453_), .ZN(new_n22454_));
  NOR2_X1    g19313(.A1(new_n22454_), .A2(new_n13748_), .ZN(new_n22455_));
  AOI21_X1   g19314(.A1(new_n13218_), .A2(new_n17730_), .B(new_n22451_), .ZN(new_n22456_));
  INV_X1     g19315(.I(new_n22456_), .ZN(new_n22457_));
  AOI21_X1   g19316(.A1(new_n22450_), .A2(new_n22457_), .B(new_n13614_), .ZN(new_n22458_));
  INV_X1     g19317(.I(new_n22458_), .ZN(new_n22459_));
  NOR3_X1    g19318(.A1(new_n22459_), .A2(new_n13748_), .A3(new_n22457_), .ZN(new_n22460_));
  XNOR2_X1   g19319(.A1(new_n22460_), .A2(new_n22455_), .ZN(new_n22461_));
  NAND2_X1   g19320(.A1(new_n22461_), .A2(new_n14049_), .ZN(new_n22462_));
  NOR2_X1    g19321(.A1(new_n22462_), .A2(new_n14051_), .ZN(new_n22463_));
  INV_X1     g19322(.I(new_n22463_), .ZN(new_n22464_));
  NOR4_X1    g19323(.A1(new_n22464_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n22465_));
  NOR2_X1    g19324(.A1(new_n22465_), .A2(new_n14005_), .ZN(new_n22466_));
  XOR2_X1    g19325(.A1(new_n22466_), .A2(new_n14007_), .Z(new_n22467_));
  NAND2_X1   g19326(.A1(new_n22467_), .A2(new_n22451_), .ZN(new_n22468_));
  INV_X1     g19327(.I(new_n22451_), .ZN(new_n22469_));
  NOR2_X1    g19328(.A1(new_n22469_), .A2(pi0647), .ZN(new_n22470_));
  AOI21_X1   g19329(.A1(new_n22465_), .A2(pi0647), .B(new_n22470_), .ZN(new_n22471_));
  AOI21_X1   g19330(.A1(new_n22471_), .A2(pi1157), .B(new_n12776_), .ZN(new_n22472_));
  AOI22_X1   g19331(.A1(new_n22468_), .A2(new_n22472_), .B1(new_n12776_), .B2(new_n22465_), .ZN(new_n22473_));
  NOR2_X1    g19332(.A1(new_n22464_), .A2(new_n14163_), .ZN(new_n22474_));
  NOR2_X1    g19333(.A1(new_n22283_), .A2(new_n22451_), .ZN(new_n22475_));
  INV_X1     g19334(.I(new_n22475_), .ZN(new_n22476_));
  NAND3_X1   g19335(.A1(new_n22476_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n22477_));
  AOI21_X1   g19336(.A1(new_n22477_), .A2(new_n16444_), .B(new_n22284_), .ZN(new_n22478_));
  NOR2_X1    g19337(.A1(new_n22478_), .A2(new_n13801_), .ZN(new_n22479_));
  NOR2_X1    g19338(.A1(new_n22451_), .A2(pi1155), .ZN(new_n22480_));
  NOR3_X1    g19339(.A1(new_n22284_), .A2(new_n16444_), .A3(new_n22480_), .ZN(new_n22481_));
  NAND4_X1   g19340(.A1(new_n22481_), .A2(new_n22476_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n22482_));
  XOR2_X1    g19341(.A1(new_n22479_), .A2(new_n22482_), .Z(new_n22483_));
  NOR2_X1    g19342(.A1(new_n22483_), .A2(new_n13817_), .ZN(new_n22484_));
  OAI21_X1   g19343(.A1(new_n22484_), .A2(pi0618), .B(new_n9992_), .ZN(new_n22485_));
  NAND2_X1   g19344(.A1(new_n22485_), .A2(pi0781), .ZN(new_n22486_));
  OAI21_X1   g19345(.A1(new_n22484_), .A2(new_n9992_), .B(pi0618), .ZN(new_n22487_));
  NOR3_X1    g19346(.A1(new_n22487_), .A2(new_n13855_), .A3(new_n22483_), .ZN(new_n22488_));
  XOR2_X1    g19347(.A1(new_n22488_), .A2(new_n22486_), .Z(new_n22489_));
  NOR2_X1    g19348(.A1(new_n22489_), .A2(new_n13868_), .ZN(new_n22490_));
  OAI21_X1   g19349(.A1(new_n22490_), .A2(pi0619), .B(new_n9992_), .ZN(new_n22491_));
  NAND2_X1   g19350(.A1(new_n22491_), .A2(pi0789), .ZN(new_n22492_));
  OAI21_X1   g19351(.A1(new_n22490_), .A2(new_n9992_), .B(pi0619), .ZN(new_n22493_));
  NOR3_X1    g19352(.A1(new_n22493_), .A2(new_n13896_), .A3(new_n22489_), .ZN(new_n22494_));
  XOR2_X1    g19353(.A1(new_n22494_), .A2(new_n22492_), .Z(new_n22495_));
  NAND2_X1   g19354(.A1(new_n22495_), .A2(new_n13962_), .ZN(new_n22496_));
  XOR2_X1    g19355(.A1(new_n22496_), .A2(new_n18976_), .Z(new_n22497_));
  AOI22_X1   g19356(.A1(new_n22497_), .A2(new_n22451_), .B1(new_n16639_), .B2(new_n22474_), .ZN(new_n22498_));
  NOR2_X1    g19357(.A1(new_n22456_), .A2(new_n13203_), .ZN(new_n22499_));
  NAND2_X1   g19358(.A1(new_n22499_), .A2(pi0625), .ZN(new_n22500_));
  NAND3_X1   g19359(.A1(new_n22500_), .A2(pi1153), .A3(new_n22475_), .ZN(new_n22501_));
  NOR2_X1    g19360(.A1(new_n22454_), .A2(new_n14081_), .ZN(new_n22502_));
  AOI21_X1   g19361(.A1(new_n22502_), .A2(new_n22501_), .B(new_n13748_), .ZN(new_n22503_));
  NOR2_X1    g19362(.A1(new_n22476_), .A2(new_n22499_), .ZN(new_n22504_));
  INV_X1     g19363(.I(new_n22500_), .ZN(new_n22505_));
  OAI21_X1   g19364(.A1(new_n22504_), .A2(new_n22505_), .B(new_n22452_), .ZN(new_n22506_));
  NAND4_X1   g19365(.A1(new_n22506_), .A2(new_n13749_), .A3(new_n22459_), .A4(new_n22504_), .ZN(new_n22507_));
  XNOR2_X1   g19366(.A1(new_n22507_), .A2(new_n22503_), .ZN(new_n22508_));
  NAND2_X1   g19367(.A1(new_n22508_), .A2(new_n13801_), .ZN(new_n22509_));
  NOR2_X1    g19368(.A1(new_n22478_), .A2(pi0660), .ZN(new_n22513_));
  NOR2_X1    g19369(.A1(new_n22508_), .A2(new_n13766_), .ZN(new_n22514_));
  XOR2_X1    g19370(.A1(new_n22514_), .A2(new_n14090_), .Z(new_n22515_));
  NOR2_X1    g19371(.A1(new_n22461_), .A2(new_n13801_), .ZN(new_n22516_));
  NAND2_X1   g19372(.A1(new_n22515_), .A2(new_n22516_), .ZN(new_n22517_));
  OAI21_X1   g19373(.A1(new_n22517_), .A2(new_n22513_), .B(new_n22509_), .ZN(new_n22518_));
  NAND2_X1   g19374(.A1(new_n22518_), .A2(new_n13855_), .ZN(new_n22519_));
  INV_X1     g19375(.I(new_n22462_), .ZN(new_n22520_));
  NOR2_X1    g19376(.A1(new_n22518_), .A2(new_n13816_), .ZN(new_n22521_));
  XOR2_X1    g19377(.A1(new_n22521_), .A2(new_n13818_), .Z(new_n22522_));
  NAND2_X1   g19378(.A1(new_n22522_), .A2(new_n22520_), .ZN(new_n22523_));
  NAND3_X1   g19379(.A1(new_n22523_), .A2(new_n13823_), .A3(new_n22487_), .ZN(new_n22524_));
  NAND3_X1   g19380(.A1(new_n22524_), .A2(new_n13823_), .A3(new_n22485_), .ZN(new_n22525_));
  NOR2_X1    g19381(.A1(new_n22518_), .A2(new_n13817_), .ZN(new_n22526_));
  XOR2_X1    g19382(.A1(new_n22526_), .A2(new_n13818_), .Z(new_n22527_));
  NAND4_X1   g19383(.A1(new_n22525_), .A2(pi0781), .A3(new_n22520_), .A4(new_n22527_), .ZN(new_n22528_));
  NAND2_X1   g19384(.A1(new_n22528_), .A2(new_n22519_), .ZN(new_n22529_));
  NOR2_X1    g19385(.A1(new_n22529_), .A2(new_n13860_), .ZN(new_n22530_));
  XOR2_X1    g19386(.A1(new_n22530_), .A2(new_n13904_), .Z(new_n22531_));
  NOR2_X1    g19387(.A1(new_n22531_), .A2(new_n22464_), .ZN(new_n22532_));
  NAND2_X1   g19388(.A1(new_n22493_), .A2(new_n13884_), .ZN(new_n22533_));
  INV_X1     g19389(.I(new_n22529_), .ZN(new_n22534_));
  AOI21_X1   g19390(.A1(new_n22534_), .A2(new_n14143_), .B(pi0789), .ZN(new_n22535_));
  OAI21_X1   g19391(.A1(new_n22532_), .A2(new_n22533_), .B(new_n22535_), .ZN(new_n22536_));
  NOR2_X1    g19392(.A1(new_n22529_), .A2(new_n13868_), .ZN(new_n22537_));
  XOR2_X1    g19393(.A1(new_n22537_), .A2(new_n13903_), .Z(new_n22538_));
  NAND2_X1   g19394(.A1(new_n22491_), .A2(new_n19018_), .ZN(new_n22539_));
  AOI21_X1   g19395(.A1(new_n22538_), .A2(new_n22463_), .B(new_n22539_), .ZN(new_n22540_));
  AOI21_X1   g19396(.A1(new_n22536_), .A2(new_n22540_), .B(new_n22498_), .ZN(new_n22541_));
  NAND2_X1   g19397(.A1(new_n22495_), .A2(new_n16372_), .ZN(new_n22542_));
  OAI21_X1   g19398(.A1(new_n16372_), .A2(new_n22451_), .B(new_n22542_), .ZN(new_n22543_));
  NAND3_X1   g19399(.A1(new_n22543_), .A2(new_n18929_), .A3(new_n22474_), .ZN(new_n22544_));
  NAND2_X1   g19400(.A1(new_n22544_), .A2(new_n16569_), .ZN(new_n22545_));
  XOR2_X1    g19401(.A1(new_n22545_), .A2(new_n16572_), .Z(new_n22546_));
  AOI21_X1   g19402(.A1(new_n19022_), .A2(new_n22544_), .B(new_n22546_), .ZN(new_n22547_));
  NAND2_X1   g19403(.A1(new_n22495_), .A2(new_n13963_), .ZN(new_n22548_));
  XNOR2_X1   g19404(.A1(new_n22548_), .A2(new_n19028_), .ZN(new_n22549_));
  NOR3_X1    g19405(.A1(new_n22549_), .A2(new_n16424_), .A3(new_n22469_), .ZN(new_n22550_));
  OAI21_X1   g19406(.A1(new_n22547_), .A2(new_n16574_), .B(new_n22550_), .ZN(new_n22551_));
  NOR2_X1    g19407(.A1(new_n22543_), .A2(new_n13994_), .ZN(new_n22552_));
  XNOR2_X1   g19408(.A1(new_n22552_), .A2(new_n19033_), .ZN(new_n22553_));
  AOI22_X1   g19409(.A1(new_n22553_), .A2(new_n22451_), .B1(new_n14206_), .B2(new_n22471_), .ZN(new_n22554_));
  NOR3_X1    g19410(.A1(new_n22554_), .A2(new_n14010_), .A3(new_n22468_), .ZN(new_n22555_));
  OAI22_X1   g19411(.A1(new_n22541_), .A2(new_n22551_), .B1(new_n12776_), .B2(new_n22555_), .ZN(new_n22556_));
  NAND2_X1   g19412(.A1(new_n22556_), .A2(pi0644), .ZN(new_n22557_));
  XOR2_X1    g19413(.A1(new_n22557_), .A2(new_n14205_), .Z(new_n22558_));
  NOR2_X1    g19414(.A1(new_n22558_), .A2(new_n22473_), .ZN(new_n22559_));
  NOR2_X1    g19415(.A1(new_n22543_), .A2(new_n18968_), .ZN(new_n22560_));
  NAND2_X1   g19416(.A1(new_n18967_), .A2(new_n22451_), .ZN(new_n22561_));
  XOR2_X1    g19417(.A1(new_n22560_), .A2(new_n22561_), .Z(new_n22562_));
  NAND2_X1   g19418(.A1(new_n22562_), .A2(pi0715), .ZN(new_n22563_));
  XOR2_X1    g19419(.A1(new_n22563_), .A2(new_n14205_), .Z(new_n22564_));
  OAI21_X1   g19420(.A1(new_n22564_), .A2(new_n22469_), .B(new_n14203_), .ZN(new_n22565_));
  NAND2_X1   g19421(.A1(new_n22562_), .A2(pi0644), .ZN(new_n22566_));
  XOR2_X1    g19422(.A1(new_n22566_), .A2(new_n14217_), .Z(new_n22567_));
  AOI21_X1   g19423(.A1(new_n22567_), .A2(new_n22451_), .B(pi1160), .ZN(new_n22568_));
  OAI21_X1   g19424(.A1(new_n22559_), .A2(new_n22565_), .B(new_n22568_), .ZN(new_n22569_));
  NAND2_X1   g19425(.A1(new_n22556_), .A2(pi0715), .ZN(new_n22570_));
  XOR2_X1    g19426(.A1(new_n22570_), .A2(new_n14205_), .Z(new_n22571_));
  NOR2_X1    g19427(.A1(new_n22571_), .A2(new_n22473_), .ZN(new_n22572_));
  AOI21_X1   g19428(.A1(new_n22569_), .A2(new_n22572_), .B(new_n14799_), .ZN(new_n22573_));
  XOR2_X1    g19429(.A1(new_n22573_), .A2(new_n14800_), .Z(new_n22574_));
  OAI21_X1   g19430(.A1(new_n7240_), .A2(pi0184), .B(new_n14799_), .ZN(new_n22575_));
  NOR2_X1    g19431(.A1(new_n22556_), .A2(new_n22575_), .ZN(new_n22576_));
  AOI21_X1   g19432(.A1(new_n22574_), .A2(new_n22576_), .B(po1038), .ZN(new_n22577_));
  NOR3_X1    g19433(.A1(new_n22448_), .A2(new_n22446_), .A3(new_n22577_), .ZN(new_n22578_));
  OAI21_X1   g19434(.A1(new_n22426_), .A2(new_n22443_), .B(new_n22578_), .ZN(new_n22579_));
  NOR2_X1    g19435(.A1(new_n22579_), .A2(new_n22384_), .ZN(po0341));
  NOR2_X1    g19436(.A1(new_n14428_), .A2(pi0185), .ZN(new_n22581_));
  INV_X1     g19437(.I(new_n22581_), .ZN(new_n22582_));
  NAND2_X1   g19438(.A1(new_n22582_), .A2(new_n13965_), .ZN(new_n22583_));
  NOR2_X1    g19439(.A1(new_n22582_), .A2(new_n13919_), .ZN(new_n22584_));
  INV_X1     g19440(.I(pi0701), .ZN(new_n22585_));
  OAI21_X1   g19441(.A1(new_n13721_), .A2(new_n22585_), .B(new_n10659_), .ZN(new_n22586_));
  NAND2_X1   g19442(.A1(new_n16715_), .A2(new_n10659_), .ZN(new_n22587_));
  NAND4_X1   g19443(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n22586_), .A4(new_n22587_), .ZN(new_n22588_));
  AOI21_X1   g19444(.A1(new_n22588_), .A2(new_n14424_), .B(new_n10659_), .ZN(new_n22589_));
  NAND2_X1   g19445(.A1(new_n22581_), .A2(new_n22589_), .ZN(new_n22590_));
  NAND2_X1   g19446(.A1(new_n22590_), .A2(new_n3290_), .ZN(new_n22591_));
  NAND2_X1   g19447(.A1(new_n22591_), .A2(pi0701), .ZN(new_n22592_));
  NAND2_X1   g19448(.A1(new_n22592_), .A2(pi0625), .ZN(new_n22593_));
  XOR2_X1    g19449(.A1(new_n22593_), .A2(new_n13620_), .Z(new_n22594_));
  NAND2_X1   g19450(.A1(new_n22594_), .A2(new_n22581_), .ZN(new_n22595_));
  NAND2_X1   g19451(.A1(new_n22595_), .A2(pi0778), .ZN(new_n22596_));
  NAND2_X1   g19452(.A1(new_n22592_), .A2(pi1153), .ZN(new_n22597_));
  XOR2_X1    g19453(.A1(new_n22597_), .A2(new_n13620_), .Z(new_n22598_));
  NAND2_X1   g19454(.A1(new_n22598_), .A2(new_n22581_), .ZN(new_n22599_));
  NOR3_X1    g19455(.A1(new_n22599_), .A2(new_n13748_), .A3(new_n22592_), .ZN(new_n22600_));
  XNOR2_X1   g19456(.A1(new_n22600_), .A2(new_n22596_), .ZN(new_n22601_));
  INV_X1     g19457(.I(new_n22601_), .ZN(new_n22602_));
  NAND2_X1   g19458(.A1(new_n22581_), .A2(new_n13803_), .ZN(new_n22603_));
  OAI21_X1   g19459(.A1(new_n22602_), .A2(new_n13803_), .B(new_n22603_), .ZN(new_n22604_));
  NOR2_X1    g19460(.A1(new_n22604_), .A2(new_n13879_), .ZN(new_n22605_));
  AOI21_X1   g19461(.A1(new_n13879_), .A2(new_n22582_), .B(new_n22605_), .ZN(new_n22606_));
  AOI21_X1   g19462(.A1(new_n22606_), .A2(new_n13919_), .B(new_n22584_), .ZN(new_n22607_));
  NAND2_X1   g19463(.A1(new_n22607_), .A2(new_n13966_), .ZN(new_n22608_));
  NAND2_X1   g19464(.A1(new_n22608_), .A2(new_n22583_), .ZN(new_n22609_));
  INV_X1     g19465(.I(new_n22609_), .ZN(new_n22610_));
  AOI21_X1   g19466(.A1(new_n22610_), .A2(pi0628), .B(new_n13971_), .ZN(new_n22611_));
  NOR3_X1    g19467(.A1(new_n22609_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n22612_));
  OAI21_X1   g19468(.A1(new_n22611_), .A2(new_n22612_), .B(new_n22581_), .ZN(new_n22613_));
  NAND2_X1   g19469(.A1(new_n22613_), .A2(pi0792), .ZN(new_n22614_));
  NAND3_X1   g19470(.A1(new_n22609_), .A2(pi0628), .A3(pi1156), .ZN(new_n22615_));
  INV_X1     g19471(.I(new_n22615_), .ZN(new_n22616_));
  NOR3_X1    g19472(.A1(new_n22609_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n22617_));
  NOR2_X1    g19473(.A1(new_n22616_), .A2(new_n22617_), .ZN(new_n22618_));
  NOR4_X1    g19474(.A1(new_n22618_), .A2(new_n12777_), .A3(new_n22582_), .A4(new_n22610_), .ZN(new_n22619_));
  NAND2_X1   g19475(.A1(new_n22619_), .A2(new_n22614_), .ZN(new_n22620_));
  NOR2_X1    g19476(.A1(new_n22619_), .A2(new_n22614_), .ZN(new_n22621_));
  INV_X1     g19477(.I(new_n22621_), .ZN(new_n22622_));
  AOI21_X1   g19478(.A1(new_n22622_), .A2(new_n22620_), .B(new_n14005_), .ZN(new_n22623_));
  NOR2_X1    g19479(.A1(new_n22582_), .A2(pi0647), .ZN(new_n22624_));
  NOR2_X1    g19480(.A1(new_n22624_), .A2(new_n14006_), .ZN(new_n22625_));
  INV_X1     g19481(.I(new_n22625_), .ZN(new_n22626_));
  NOR2_X1    g19482(.A1(new_n22623_), .A2(new_n22626_), .ZN(new_n22627_));
  AOI21_X1   g19483(.A1(new_n22622_), .A2(new_n22620_), .B(pi0647), .ZN(new_n22628_));
  NOR2_X1    g19484(.A1(new_n22582_), .A2(new_n14005_), .ZN(new_n22629_));
  NOR3_X1    g19485(.A1(new_n22628_), .A2(pi1157), .A3(new_n22629_), .ZN(new_n22630_));
  OAI21_X1   g19486(.A1(new_n22630_), .A2(new_n22627_), .B(pi0787), .ZN(new_n22631_));
  NAND3_X1   g19487(.A1(new_n22610_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n22632_));
  AOI21_X1   g19488(.A1(new_n22632_), .A2(new_n22615_), .B(new_n22582_), .ZN(new_n22633_));
  NAND3_X1   g19489(.A1(new_n22633_), .A2(pi0792), .A3(new_n22609_), .ZN(new_n22634_));
  AOI21_X1   g19490(.A1(pi0792), .A2(new_n22613_), .B(new_n22634_), .ZN(new_n22635_));
  NOR3_X1    g19491(.A1(new_n22635_), .A2(pi0787), .A3(new_n22621_), .ZN(new_n22636_));
  INV_X1     g19492(.I(new_n22636_), .ZN(new_n22637_));
  NAND2_X1   g19493(.A1(new_n22582_), .A2(new_n14142_), .ZN(new_n22638_));
  NOR2_X1    g19494(.A1(new_n10659_), .A2(new_n17192_), .ZN(new_n22639_));
  INV_X1     g19495(.I(new_n22639_), .ZN(new_n22640_));
  NAND2_X1   g19496(.A1(new_n20780_), .A2(new_n22640_), .ZN(new_n22641_));
  OAI21_X1   g19497(.A1(new_n14298_), .A2(new_n10659_), .B(new_n3183_), .ZN(new_n22642_));
  AOI21_X1   g19498(.A1(new_n13194_), .A2(pi0751), .B(new_n22642_), .ZN(new_n22643_));
  OAI21_X1   g19499(.A1(new_n22643_), .A2(new_n17192_), .B(pi0185), .ZN(new_n22644_));
  OAI21_X1   g19500(.A1(new_n20785_), .A2(new_n22644_), .B(new_n3183_), .ZN(new_n22645_));
  AOI21_X1   g19501(.A1(new_n13109_), .A2(new_n10659_), .B(new_n3259_), .ZN(new_n22646_));
  AND3_X2    g19502(.A1(new_n22641_), .A2(new_n22645_), .A3(new_n22646_), .Z(new_n22647_));
  OAI21_X1   g19503(.A1(new_n22647_), .A2(new_n13106_), .B(pi0751), .ZN(new_n22648_));
  INV_X1     g19504(.I(new_n22648_), .ZN(new_n22649_));
  NOR2_X1    g19505(.A1(new_n3289_), .A2(pi0185), .ZN(new_n22650_));
  AOI21_X1   g19506(.A1(new_n22649_), .A2(new_n3289_), .B(new_n22650_), .ZN(new_n22651_));
  NAND2_X1   g19507(.A1(new_n22651_), .A2(new_n13776_), .ZN(new_n22652_));
  NAND2_X1   g19508(.A1(new_n22582_), .A2(new_n13780_), .ZN(new_n22653_));
  NAND2_X1   g19509(.A1(new_n22652_), .A2(new_n22653_), .ZN(new_n22654_));
  NAND2_X1   g19510(.A1(new_n22654_), .A2(pi0609), .ZN(new_n22655_));
  NAND2_X1   g19511(.A1(new_n22655_), .A2(pi0785), .ZN(new_n22656_));
  NAND2_X1   g19512(.A1(new_n22581_), .A2(new_n13775_), .ZN(new_n22657_));
  OAI21_X1   g19513(.A1(new_n22651_), .A2(new_n13775_), .B(new_n22657_), .ZN(new_n22658_));
  AOI21_X1   g19514(.A1(new_n22582_), .A2(new_n14467_), .B(pi0609), .ZN(new_n22659_));
  NOR2_X1    g19515(.A1(new_n22652_), .A2(new_n22659_), .ZN(new_n22660_));
  NAND3_X1   g19516(.A1(new_n22660_), .A2(pi0785), .A3(new_n22658_), .ZN(new_n22661_));
  XNOR2_X1   g19517(.A1(new_n22656_), .A2(new_n22661_), .ZN(new_n22662_));
  INV_X1     g19518(.I(new_n22662_), .ZN(new_n22663_));
  NAND3_X1   g19519(.A1(new_n22663_), .A2(pi0618), .A3(pi1154), .ZN(new_n22664_));
  NAND3_X1   g19520(.A1(new_n22662_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n22665_));
  AOI21_X1   g19521(.A1(new_n22664_), .A2(new_n22665_), .B(new_n22582_), .ZN(new_n22666_));
  NAND3_X1   g19522(.A1(new_n22663_), .A2(pi0618), .A3(pi1154), .ZN(new_n22667_));
  NAND3_X1   g19523(.A1(new_n22662_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n22668_));
  AOI21_X1   g19524(.A1(new_n22667_), .A2(new_n22668_), .B(new_n22582_), .ZN(new_n22669_));
  NAND4_X1   g19525(.A1(new_n22666_), .A2(new_n22669_), .A3(pi0781), .A4(new_n22663_), .ZN(new_n22670_));
  NOR2_X1    g19526(.A1(new_n22666_), .A2(new_n13855_), .ZN(new_n22671_));
  INV_X1     g19527(.I(new_n22669_), .ZN(new_n22672_));
  NAND2_X1   g19528(.A1(new_n22663_), .A2(pi0781), .ZN(new_n22673_));
  OAI21_X1   g19529(.A1(new_n22672_), .A2(new_n22673_), .B(new_n22671_), .ZN(new_n22674_));
  NAND2_X1   g19530(.A1(new_n22674_), .A2(new_n22670_), .ZN(new_n22675_));
  NAND3_X1   g19531(.A1(new_n22675_), .A2(pi0619), .A3(pi1159), .ZN(new_n22676_));
  INV_X1     g19532(.I(new_n22675_), .ZN(new_n22677_));
  NAND3_X1   g19533(.A1(new_n22677_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n22678_));
  AOI21_X1   g19534(.A1(new_n22678_), .A2(new_n22676_), .B(new_n22582_), .ZN(new_n22679_));
  NOR2_X1    g19535(.A1(new_n22679_), .A2(new_n13896_), .ZN(new_n22680_));
  INV_X1     g19536(.I(new_n22680_), .ZN(new_n22681_));
  NOR2_X1    g19537(.A1(new_n22675_), .A2(new_n13868_), .ZN(new_n22682_));
  XOR2_X1    g19538(.A1(new_n22682_), .A2(new_n13903_), .Z(new_n22683_));
  NOR2_X1    g19539(.A1(new_n22677_), .A2(new_n13896_), .ZN(new_n22684_));
  NAND4_X1   g19540(.A1(new_n22681_), .A2(new_n22581_), .A3(new_n22683_), .A4(new_n22684_), .ZN(new_n22685_));
  NAND2_X1   g19541(.A1(new_n22683_), .A2(new_n22581_), .ZN(new_n22686_));
  INV_X1     g19542(.I(new_n22684_), .ZN(new_n22687_));
  OAI21_X1   g19543(.A1(new_n22686_), .A2(new_n22687_), .B(new_n22680_), .ZN(new_n22688_));
  NAND2_X1   g19544(.A1(new_n22685_), .A2(new_n22688_), .ZN(new_n22689_));
  OAI21_X1   g19545(.A1(new_n22689_), .A2(new_n14142_), .B(new_n22638_), .ZN(new_n22690_));
  NOR2_X1    g19546(.A1(new_n22581_), .A2(new_n13994_), .ZN(new_n22691_));
  AOI21_X1   g19547(.A1(new_n22690_), .A2(new_n13994_), .B(new_n22691_), .ZN(new_n22692_));
  NAND2_X1   g19548(.A1(new_n22582_), .A2(new_n14210_), .ZN(new_n22693_));
  OAI21_X1   g19549(.A1(new_n22692_), .A2(new_n14210_), .B(new_n22693_), .ZN(new_n22694_));
  NAND2_X1   g19550(.A1(new_n19370_), .A2(new_n14204_), .ZN(new_n22695_));
  NAND3_X1   g19551(.A1(new_n22694_), .A2(pi0715), .A3(new_n22695_), .ZN(new_n22696_));
  AOI22_X1   g19552(.A1(new_n22631_), .A2(new_n22637_), .B1(new_n14204_), .B2(new_n22696_), .ZN(new_n22697_));
  OAI21_X1   g19553(.A1(new_n22635_), .A2(new_n22621_), .B(new_n14005_), .ZN(new_n22698_));
  INV_X1     g19554(.I(new_n22629_), .ZN(new_n22699_));
  NAND2_X1   g19555(.A1(new_n22698_), .A2(new_n22699_), .ZN(new_n22700_));
  OAI22_X1   g19556(.A1(new_n22700_), .A2(pi1157), .B1(new_n22623_), .B2(new_n22626_), .ZN(new_n22701_));
  AOI21_X1   g19557(.A1(new_n22701_), .A2(pi0787), .B(new_n22636_), .ZN(new_n22702_));
  OAI21_X1   g19558(.A1(new_n22581_), .A2(new_n14255_), .B(new_n14204_), .ZN(new_n22703_));
  NAND3_X1   g19559(.A1(new_n22694_), .A2(pi0715), .A3(new_n22703_), .ZN(new_n22704_));
  AOI21_X1   g19560(.A1(new_n22702_), .A2(new_n22704_), .B(new_n14204_), .ZN(new_n22705_));
  OAI21_X1   g19561(.A1(new_n22705_), .A2(new_n22697_), .B(pi0790), .ZN(new_n22706_));
  NAND2_X1   g19562(.A1(new_n22694_), .A2(new_n22695_), .ZN(new_n22707_));
  NAND4_X1   g19563(.A1(new_n22694_), .A2(pi0644), .A3(pi0790), .A4(new_n22703_), .ZN(new_n22708_));
  NAND2_X1   g19564(.A1(new_n22694_), .A2(new_n22703_), .ZN(new_n22709_));
  NAND3_X1   g19565(.A1(new_n22709_), .A2(new_n14204_), .A3(pi0790), .ZN(new_n22710_));
  AOI21_X1   g19566(.A1(new_n22710_), .A2(new_n22708_), .B(new_n22707_), .ZN(new_n22711_));
  NOR2_X1    g19567(.A1(new_n22628_), .A2(new_n22629_), .ZN(new_n22712_));
  NOR4_X1    g19568(.A1(new_n22623_), .A2(pi0630), .A3(new_n14006_), .A4(new_n22624_), .ZN(new_n22713_));
  NOR3_X1    g19569(.A1(new_n22623_), .A2(pi0630), .A3(new_n22626_), .ZN(new_n22714_));
  NOR3_X1    g19570(.A1(new_n22714_), .A2(new_n22712_), .A3(new_n14012_), .ZN(new_n22715_));
  OAI21_X1   g19571(.A1(new_n22715_), .A2(new_n22713_), .B(pi0787), .ZN(new_n22716_));
  AOI21_X1   g19572(.A1(new_n22716_), .A2(new_n22692_), .B(new_n16867_), .ZN(new_n22717_));
  NOR2_X1    g19573(.A1(new_n22717_), .A2(new_n22711_), .ZN(new_n22718_));
  INV_X1     g19574(.I(new_n22604_), .ZN(new_n22719_));
  NAND2_X1   g19575(.A1(new_n13461_), .A2(pi0185), .ZN(new_n22720_));
  XOR2_X1    g19576(.A1(new_n22720_), .A2(new_n22640_), .Z(new_n22721_));
  NAND2_X1   g19577(.A1(new_n22721_), .A2(new_n13521_), .ZN(new_n22722_));
  NAND3_X1   g19578(.A1(new_n14270_), .A2(pi0185), .A3(pi0751), .ZN(new_n22723_));
  NAND3_X1   g19579(.A1(new_n14272_), .A2(new_n10659_), .A3(pi0751), .ZN(new_n22724_));
  AOI21_X1   g19580(.A1(new_n22723_), .A2(new_n22724_), .B(new_n13152_), .ZN(new_n22725_));
  NAND3_X1   g19581(.A1(new_n13198_), .A2(pi0185), .A3(pi0751), .ZN(new_n22726_));
  NAND3_X1   g19582(.A1(new_n13200_), .A2(pi0185), .A3(new_n17192_), .ZN(new_n22727_));
  AOI21_X1   g19583(.A1(new_n22727_), .A2(new_n22726_), .B(new_n13191_), .ZN(new_n22728_));
  OAI21_X1   g19584(.A1(new_n22725_), .A2(new_n3262_), .B(new_n22728_), .ZN(new_n22729_));
  NAND3_X1   g19585(.A1(new_n22722_), .A2(new_n3183_), .A3(new_n22729_), .ZN(new_n22730_));
  NOR2_X1    g19586(.A1(new_n14284_), .A2(new_n17192_), .ZN(new_n22731_));
  XOR2_X1    g19587(.A1(new_n22731_), .A2(new_n22639_), .Z(new_n22732_));
  NAND3_X1   g19588(.A1(new_n22730_), .A2(new_n22732_), .A3(new_n13359_), .ZN(new_n22733_));
  NAND3_X1   g19589(.A1(new_n22733_), .A2(new_n22585_), .A3(new_n3290_), .ZN(new_n22734_));
  OAI21_X1   g19590(.A1(new_n15587_), .A2(new_n10659_), .B(new_n17192_), .ZN(new_n22735_));
  NAND2_X1   g19591(.A1(new_n22735_), .A2(new_n13209_), .ZN(new_n22736_));
  NOR2_X1    g19592(.A1(new_n13105_), .A2(pi0751), .ZN(new_n22737_));
  INV_X1     g19593(.I(new_n22737_), .ZN(new_n22738_));
  NAND2_X1   g19594(.A1(new_n22738_), .A2(new_n16751_), .ZN(new_n22739_));
  NAND4_X1   g19595(.A1(new_n5503_), .A2(new_n22739_), .A3(pi0185), .A4(new_n3290_), .ZN(new_n22740_));
  AOI21_X1   g19596(.A1(new_n22736_), .A2(new_n3259_), .B(new_n22740_), .ZN(new_n22741_));
  NAND2_X1   g19597(.A1(new_n22734_), .A2(new_n22741_), .ZN(new_n22742_));
  AOI21_X1   g19598(.A1(new_n22742_), .A2(new_n22585_), .B(new_n22648_), .ZN(new_n22743_));
  INV_X1     g19599(.I(new_n22599_), .ZN(new_n22744_));
  INV_X1     g19600(.I(new_n22743_), .ZN(new_n22745_));
  NAND2_X1   g19601(.A1(new_n22651_), .A2(pi0625), .ZN(new_n22746_));
  XOR2_X1    g19602(.A1(new_n22746_), .A2(new_n13615_), .Z(new_n22747_));
  OAI21_X1   g19603(.A1(new_n22745_), .A2(new_n22747_), .B(new_n14081_), .ZN(new_n22748_));
  NAND2_X1   g19604(.A1(new_n22651_), .A2(pi1153), .ZN(new_n22749_));
  XOR2_X1    g19605(.A1(new_n22749_), .A2(new_n13620_), .Z(new_n22750_));
  AOI21_X1   g19606(.A1(new_n22743_), .A2(new_n22750_), .B(pi0608), .ZN(new_n22751_));
  OAI21_X1   g19607(.A1(new_n22748_), .A2(new_n22744_), .B(new_n22751_), .ZN(new_n22752_));
  NAND4_X1   g19608(.A1(new_n22752_), .A2(pi0778), .A3(new_n22581_), .A4(new_n22594_), .ZN(new_n22753_));
  OAI21_X1   g19609(.A1(pi0778), .A2(new_n22743_), .B(new_n22753_), .ZN(new_n22754_));
  NAND2_X1   g19610(.A1(new_n22754_), .A2(new_n13801_), .ZN(new_n22755_));
  NOR2_X1    g19611(.A1(new_n22754_), .A2(new_n13778_), .ZN(new_n22756_));
  NOR2_X1    g19612(.A1(new_n22756_), .A2(new_n14694_), .ZN(new_n22757_));
  NAND2_X1   g19613(.A1(new_n22756_), .A2(new_n14694_), .ZN(new_n22758_));
  INV_X1     g19614(.I(new_n22758_), .ZN(new_n22759_));
  OAI21_X1   g19615(.A1(new_n22759_), .A2(new_n22757_), .B(new_n22601_), .ZN(new_n22760_));
  NAND2_X1   g19616(.A1(new_n22655_), .A2(pi0660), .ZN(new_n22761_));
  INV_X1     g19617(.I(new_n22761_), .ZN(new_n22762_));
  NOR2_X1    g19618(.A1(new_n22660_), .A2(pi0660), .ZN(new_n22763_));
  INV_X1     g19619(.I(new_n22763_), .ZN(new_n22764_));
  AOI21_X1   g19620(.A1(new_n22760_), .A2(new_n22762_), .B(new_n22764_), .ZN(new_n22765_));
  NOR2_X1    g19621(.A1(new_n22754_), .A2(new_n13766_), .ZN(new_n22766_));
  XOR2_X1    g19622(.A1(new_n22766_), .A2(new_n14694_), .Z(new_n22767_));
  NAND2_X1   g19623(.A1(new_n22601_), .A2(pi0785), .ZN(new_n22768_));
  NOR2_X1    g19624(.A1(new_n22767_), .A2(new_n22768_), .ZN(new_n22769_));
  INV_X1     g19625(.I(new_n22769_), .ZN(new_n22770_));
  OAI21_X1   g19626(.A1(new_n22770_), .A2(new_n22765_), .B(new_n22755_), .ZN(new_n22771_));
  NAND3_X1   g19627(.A1(new_n22771_), .A2(pi0618), .A3(pi1154), .ZN(new_n22772_));
  INV_X1     g19628(.I(new_n22757_), .ZN(new_n22773_));
  AOI21_X1   g19629(.A1(new_n22773_), .A2(new_n22758_), .B(new_n22602_), .ZN(new_n22774_));
  OAI21_X1   g19630(.A1(new_n22774_), .A2(new_n22761_), .B(new_n22763_), .ZN(new_n22775_));
  AOI22_X1   g19631(.A1(new_n22775_), .A2(new_n22769_), .B1(new_n13801_), .B2(new_n22754_), .ZN(new_n22776_));
  NAND3_X1   g19632(.A1(new_n22776_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n22777_));
  AOI21_X1   g19633(.A1(new_n22777_), .A2(new_n22772_), .B(new_n22719_), .ZN(new_n22778_));
  NOR2_X1    g19634(.A1(new_n22666_), .A2(new_n13823_), .ZN(new_n22779_));
  INV_X1     g19635(.I(new_n22779_), .ZN(new_n22780_));
  OAI21_X1   g19636(.A1(new_n22778_), .A2(new_n22780_), .B(pi0781), .ZN(new_n22781_));
  NAND3_X1   g19637(.A1(new_n22771_), .A2(pi0618), .A3(pi1154), .ZN(new_n22782_));
  NAND3_X1   g19638(.A1(new_n22776_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n22783_));
  NAND2_X1   g19639(.A1(new_n22783_), .A2(new_n22782_), .ZN(new_n22784_));
  NAND3_X1   g19640(.A1(new_n22771_), .A2(new_n19177_), .A3(new_n22672_), .ZN(new_n22785_));
  AOI21_X1   g19641(.A1(new_n22784_), .A2(new_n22604_), .B(new_n22785_), .ZN(new_n22786_));
  NAND2_X1   g19642(.A1(new_n22781_), .A2(new_n22786_), .ZN(new_n22787_));
  AOI21_X1   g19643(.A1(new_n22776_), .A2(pi1154), .B(new_n13819_), .ZN(new_n22788_));
  NOR3_X1    g19644(.A1(new_n22771_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n22789_));
  OAI21_X1   g19645(.A1(new_n22788_), .A2(new_n22789_), .B(new_n22604_), .ZN(new_n22790_));
  AOI21_X1   g19646(.A1(new_n22790_), .A2(new_n22779_), .B(new_n13855_), .ZN(new_n22791_));
  AOI21_X1   g19647(.A1(new_n22776_), .A2(pi0618), .B(new_n13819_), .ZN(new_n22792_));
  NOR3_X1    g19648(.A1(new_n22771_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n22793_));
  OAI21_X1   g19649(.A1(new_n22792_), .A2(new_n22793_), .B(new_n22604_), .ZN(new_n22794_));
  NAND4_X1   g19650(.A1(new_n22794_), .A2(new_n19177_), .A3(new_n22672_), .A4(new_n22771_), .ZN(new_n22795_));
  NAND2_X1   g19651(.A1(new_n22795_), .A2(new_n22791_), .ZN(new_n22796_));
  NAND2_X1   g19652(.A1(new_n22796_), .A2(new_n22787_), .ZN(new_n22797_));
  NAND3_X1   g19653(.A1(new_n22797_), .A2(pi0619), .A3(pi1159), .ZN(new_n22798_));
  NOR2_X1    g19654(.A1(new_n22795_), .A2(new_n22791_), .ZN(new_n22799_));
  NOR2_X1    g19655(.A1(new_n22781_), .A2(new_n22786_), .ZN(new_n22800_));
  NOR2_X1    g19656(.A1(new_n22799_), .A2(new_n22800_), .ZN(new_n22801_));
  NAND3_X1   g19657(.A1(new_n22801_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n22802_));
  AOI21_X1   g19658(.A1(new_n22802_), .A2(new_n22798_), .B(new_n22606_), .ZN(new_n22803_));
  OAI21_X1   g19659(.A1(new_n22803_), .A2(new_n20003_), .B(new_n22679_), .ZN(new_n22804_));
  NAND2_X1   g19660(.A1(new_n22797_), .A2(new_n13896_), .ZN(new_n22805_));
  NAND3_X1   g19661(.A1(new_n22689_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n22806_));
  INV_X1     g19662(.I(new_n22689_), .ZN(new_n22807_));
  NAND3_X1   g19663(.A1(new_n22807_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n22808_));
  AOI21_X1   g19664(.A1(new_n22808_), .A2(new_n22806_), .B(new_n22582_), .ZN(new_n22809_));
  NOR2_X1    g19665(.A1(new_n22607_), .A2(new_n14162_), .ZN(new_n22810_));
  OAI21_X1   g19666(.A1(new_n22809_), .A2(new_n22810_), .B(new_n19204_), .ZN(new_n22811_));
  NOR2_X1    g19667(.A1(new_n22689_), .A2(new_n19208_), .ZN(new_n22812_));
  XNOR2_X1   g19668(.A1(new_n22812_), .A2(new_n19028_), .ZN(new_n22813_));
  NOR2_X1    g19669(.A1(new_n22582_), .A2(new_n15479_), .ZN(new_n22814_));
  NAND4_X1   g19670(.A1(new_n22811_), .A2(new_n22805_), .A3(new_n22813_), .A4(new_n22814_), .ZN(new_n22815_));
  INV_X1     g19671(.I(new_n22606_), .ZN(new_n22816_));
  AOI21_X1   g19672(.A1(new_n22801_), .A2(pi0619), .B(new_n13904_), .ZN(new_n22817_));
  NOR4_X1    g19673(.A1(new_n22799_), .A2(new_n22800_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n22818_));
  OAI21_X1   g19674(.A1(new_n22817_), .A2(new_n22818_), .B(new_n22816_), .ZN(new_n22819_));
  NAND3_X1   g19675(.A1(new_n22819_), .A2(new_n20173_), .A3(new_n22686_), .ZN(new_n22820_));
  AOI21_X1   g19676(.A1(new_n22804_), .A2(new_n22815_), .B(new_n22820_), .ZN(new_n22821_));
  AND2_X2    g19677(.A1(new_n22613_), .A2(pi0629), .Z(new_n22822_));
  NOR2_X1    g19678(.A1(new_n22633_), .A2(pi0629), .ZN(new_n22823_));
  NOR2_X1    g19679(.A1(new_n9992_), .A2(pi0185), .ZN(new_n22824_));
  NOR3_X1    g19680(.A1(new_n13219_), .A2(pi0625), .A3(pi0701), .ZN(new_n22825_));
  INV_X1     g19681(.I(new_n22825_), .ZN(new_n22826_));
  NOR2_X1    g19682(.A1(new_n22824_), .A2(pi1153), .ZN(new_n22827_));
  NAND2_X1   g19683(.A1(new_n22826_), .A2(new_n22827_), .ZN(new_n22828_));
  INV_X1     g19684(.I(new_n22828_), .ZN(new_n22829_));
  NOR2_X1    g19685(.A1(new_n22829_), .A2(new_n13748_), .ZN(new_n22830_));
  AOI21_X1   g19686(.A1(new_n13218_), .A2(new_n22585_), .B(new_n22824_), .ZN(new_n22831_));
  INV_X1     g19687(.I(new_n22831_), .ZN(new_n22832_));
  AOI21_X1   g19688(.A1(new_n22826_), .A2(new_n22832_), .B(new_n13614_), .ZN(new_n22833_));
  INV_X1     g19689(.I(new_n22833_), .ZN(new_n22834_));
  NOR3_X1    g19690(.A1(new_n22834_), .A2(new_n13748_), .A3(new_n22832_), .ZN(new_n22835_));
  XNOR2_X1   g19691(.A1(new_n22835_), .A2(new_n22830_), .ZN(new_n22836_));
  NAND2_X1   g19692(.A1(new_n22836_), .A2(new_n14049_), .ZN(new_n22837_));
  NOR2_X1    g19693(.A1(new_n22837_), .A2(new_n14051_), .ZN(new_n22838_));
  INV_X1     g19694(.I(new_n22838_), .ZN(new_n22839_));
  NOR2_X1    g19695(.A1(new_n22839_), .A2(new_n14163_), .ZN(new_n22840_));
  NOR2_X1    g19696(.A1(new_n22737_), .A2(new_n22824_), .ZN(new_n22841_));
  INV_X1     g19697(.I(new_n22841_), .ZN(new_n22842_));
  NAND3_X1   g19698(.A1(new_n22842_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n22843_));
  AOI21_X1   g19699(.A1(new_n22843_), .A2(new_n16444_), .B(new_n22738_), .ZN(new_n22844_));
  NOR2_X1    g19700(.A1(new_n22844_), .A2(new_n13801_), .ZN(new_n22845_));
  NOR2_X1    g19701(.A1(new_n22824_), .A2(pi1155), .ZN(new_n22846_));
  NOR3_X1    g19702(.A1(new_n22738_), .A2(new_n16444_), .A3(new_n22846_), .ZN(new_n22847_));
  NAND4_X1   g19703(.A1(new_n22847_), .A2(new_n22842_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n22848_));
  XOR2_X1    g19704(.A1(new_n22845_), .A2(new_n22848_), .Z(new_n22849_));
  NOR2_X1    g19705(.A1(new_n22849_), .A2(new_n13817_), .ZN(new_n22850_));
  OAI21_X1   g19706(.A1(new_n22850_), .A2(pi0618), .B(new_n9992_), .ZN(new_n22851_));
  NAND2_X1   g19707(.A1(new_n22851_), .A2(pi0781), .ZN(new_n22852_));
  OAI21_X1   g19708(.A1(new_n22850_), .A2(new_n9992_), .B(pi0618), .ZN(new_n22853_));
  NOR3_X1    g19709(.A1(new_n22853_), .A2(new_n13855_), .A3(new_n22849_), .ZN(new_n22854_));
  XOR2_X1    g19710(.A1(new_n22854_), .A2(new_n22852_), .Z(new_n22855_));
  NOR2_X1    g19711(.A1(new_n22855_), .A2(new_n13868_), .ZN(new_n22856_));
  OAI21_X1   g19712(.A1(new_n22856_), .A2(pi0619), .B(new_n9992_), .ZN(new_n22857_));
  NAND2_X1   g19713(.A1(new_n22857_), .A2(pi0789), .ZN(new_n22858_));
  OAI21_X1   g19714(.A1(new_n22856_), .A2(new_n9992_), .B(pi0619), .ZN(new_n22859_));
  NOR3_X1    g19715(.A1(new_n22859_), .A2(new_n13896_), .A3(new_n22855_), .ZN(new_n22860_));
  XOR2_X1    g19716(.A1(new_n22860_), .A2(new_n22858_), .Z(new_n22861_));
  NAND2_X1   g19717(.A1(new_n22861_), .A2(new_n13962_), .ZN(new_n22862_));
  XOR2_X1    g19718(.A1(new_n22862_), .A2(new_n18976_), .Z(new_n22863_));
  AOI22_X1   g19719(.A1(new_n22863_), .A2(new_n22824_), .B1(new_n16639_), .B2(new_n22840_), .ZN(new_n22864_));
  NOR2_X1    g19720(.A1(new_n22831_), .A2(new_n13203_), .ZN(new_n22865_));
  NAND2_X1   g19721(.A1(new_n22865_), .A2(pi0625), .ZN(new_n22866_));
  NAND3_X1   g19722(.A1(new_n22866_), .A2(pi1153), .A3(new_n22841_), .ZN(new_n22867_));
  NOR2_X1    g19723(.A1(new_n22829_), .A2(new_n14081_), .ZN(new_n22868_));
  AOI21_X1   g19724(.A1(new_n22868_), .A2(new_n22867_), .B(new_n13748_), .ZN(new_n22869_));
  NOR2_X1    g19725(.A1(new_n22842_), .A2(new_n22865_), .ZN(new_n22870_));
  INV_X1     g19726(.I(new_n22866_), .ZN(new_n22871_));
  OAI21_X1   g19727(.A1(new_n22870_), .A2(new_n22871_), .B(new_n22827_), .ZN(new_n22872_));
  NAND4_X1   g19728(.A1(new_n22872_), .A2(new_n13749_), .A3(new_n22834_), .A4(new_n22870_), .ZN(new_n22873_));
  XNOR2_X1   g19729(.A1(new_n22873_), .A2(new_n22869_), .ZN(new_n22874_));
  NAND2_X1   g19730(.A1(new_n22874_), .A2(new_n13801_), .ZN(new_n22875_));
  NOR2_X1    g19731(.A1(new_n22844_), .A2(pi0660), .ZN(new_n22879_));
  NOR2_X1    g19732(.A1(new_n22874_), .A2(new_n13766_), .ZN(new_n22880_));
  XOR2_X1    g19733(.A1(new_n22880_), .A2(new_n14090_), .Z(new_n22881_));
  NOR2_X1    g19734(.A1(new_n22836_), .A2(new_n13801_), .ZN(new_n22882_));
  NAND2_X1   g19735(.A1(new_n22881_), .A2(new_n22882_), .ZN(new_n22883_));
  OAI21_X1   g19736(.A1(new_n22883_), .A2(new_n22879_), .B(new_n22875_), .ZN(new_n22884_));
  NAND2_X1   g19737(.A1(new_n22884_), .A2(new_n13855_), .ZN(new_n22885_));
  INV_X1     g19738(.I(new_n22837_), .ZN(new_n22886_));
  NOR2_X1    g19739(.A1(new_n22884_), .A2(new_n13816_), .ZN(new_n22887_));
  XOR2_X1    g19740(.A1(new_n22887_), .A2(new_n13818_), .Z(new_n22888_));
  NAND2_X1   g19741(.A1(new_n22888_), .A2(new_n22886_), .ZN(new_n22889_));
  NAND3_X1   g19742(.A1(new_n22889_), .A2(new_n13823_), .A3(new_n22853_), .ZN(new_n22890_));
  NAND3_X1   g19743(.A1(new_n22890_), .A2(new_n13823_), .A3(new_n22851_), .ZN(new_n22891_));
  NOR2_X1    g19744(.A1(new_n22884_), .A2(new_n13817_), .ZN(new_n22892_));
  XOR2_X1    g19745(.A1(new_n22892_), .A2(new_n13818_), .Z(new_n22893_));
  NAND4_X1   g19746(.A1(new_n22891_), .A2(pi0781), .A3(new_n22886_), .A4(new_n22893_), .ZN(new_n22894_));
  NAND2_X1   g19747(.A1(new_n22894_), .A2(new_n22885_), .ZN(new_n22895_));
  NOR2_X1    g19748(.A1(new_n22895_), .A2(new_n13860_), .ZN(new_n22896_));
  XOR2_X1    g19749(.A1(new_n22896_), .A2(new_n13904_), .Z(new_n22897_));
  NOR2_X1    g19750(.A1(new_n22897_), .A2(new_n22839_), .ZN(new_n22898_));
  NAND2_X1   g19751(.A1(new_n22859_), .A2(new_n13884_), .ZN(new_n22899_));
  INV_X1     g19752(.I(new_n22895_), .ZN(new_n22900_));
  AOI21_X1   g19753(.A1(new_n22900_), .A2(new_n14143_), .B(pi0789), .ZN(new_n22901_));
  OAI21_X1   g19754(.A1(new_n22898_), .A2(new_n22899_), .B(new_n22901_), .ZN(new_n22902_));
  NOR2_X1    g19755(.A1(new_n22895_), .A2(new_n13868_), .ZN(new_n22903_));
  XOR2_X1    g19756(.A1(new_n22903_), .A2(new_n13903_), .Z(new_n22904_));
  NAND2_X1   g19757(.A1(new_n22857_), .A2(new_n19018_), .ZN(new_n22905_));
  AOI21_X1   g19758(.A1(new_n22904_), .A2(new_n22838_), .B(new_n22905_), .ZN(new_n22906_));
  AOI21_X1   g19759(.A1(new_n22902_), .A2(new_n22906_), .B(new_n22864_), .ZN(new_n22907_));
  NOR3_X1    g19760(.A1(new_n22839_), .A2(new_n14163_), .A3(new_n18928_), .ZN(new_n22908_));
  NAND2_X1   g19761(.A1(new_n22861_), .A2(new_n16372_), .ZN(new_n22909_));
  OAI21_X1   g19762(.A1(new_n16372_), .A2(new_n22824_), .B(new_n22909_), .ZN(new_n22910_));
  NAND2_X1   g19763(.A1(new_n22910_), .A2(new_n22908_), .ZN(new_n22911_));
  NAND2_X1   g19764(.A1(new_n22911_), .A2(new_n19022_), .ZN(new_n22912_));
  NAND2_X1   g19765(.A1(new_n22911_), .A2(new_n16569_), .ZN(new_n22913_));
  XNOR2_X1   g19766(.A1(new_n22913_), .A2(new_n16572_), .ZN(new_n22914_));
  AOI21_X1   g19767(.A1(new_n22914_), .A2(new_n22912_), .B(new_n16574_), .ZN(new_n22915_));
  NAND2_X1   g19768(.A1(new_n22861_), .A2(new_n13963_), .ZN(new_n22916_));
  XNOR2_X1   g19769(.A1(new_n22916_), .A2(new_n19028_), .ZN(new_n22917_));
  NAND2_X1   g19770(.A1(new_n16423_), .A2(new_n22824_), .ZN(new_n22918_));
  NOR4_X1    g19771(.A1(new_n22907_), .A2(new_n22915_), .A3(new_n22917_), .A4(new_n22918_), .ZN(new_n22919_));
  INV_X1     g19772(.I(new_n22824_), .ZN(new_n22920_));
  NAND2_X1   g19773(.A1(new_n22908_), .A2(new_n14061_), .ZN(new_n22921_));
  NAND2_X1   g19774(.A1(new_n22824_), .A2(new_n14005_), .ZN(new_n22922_));
  OAI21_X1   g19775(.A1(new_n22921_), .A2(new_n14005_), .B(new_n22922_), .ZN(new_n22923_));
  NOR2_X1    g19776(.A1(new_n22910_), .A2(new_n13994_), .ZN(new_n22924_));
  XOR2_X1    g19777(.A1(new_n22924_), .A2(new_n19033_), .Z(new_n22925_));
  OAI22_X1   g19778(.A1(new_n22925_), .A2(new_n22920_), .B1(new_n14207_), .B2(new_n22923_), .ZN(new_n22926_));
  NAND2_X1   g19779(.A1(new_n22921_), .A2(pi0647), .ZN(new_n22927_));
  XOR2_X1    g19780(.A1(new_n22927_), .A2(new_n14007_), .Z(new_n22928_));
  NOR3_X1    g19781(.A1(new_n22928_), .A2(new_n14010_), .A3(new_n22920_), .ZN(new_n22929_));
  AOI21_X1   g19782(.A1(new_n22926_), .A2(new_n22929_), .B(new_n12776_), .ZN(new_n22930_));
  NOR2_X1    g19783(.A1(new_n22919_), .A2(new_n22930_), .ZN(new_n22931_));
  NOR2_X1    g19784(.A1(new_n22928_), .A2(new_n22920_), .ZN(new_n22932_));
  OAI21_X1   g19785(.A1(new_n22923_), .A2(new_n14006_), .B(pi0787), .ZN(new_n22933_));
  OAI22_X1   g19786(.A1(new_n22932_), .A2(new_n22933_), .B1(pi0787), .B2(new_n22921_), .ZN(new_n22934_));
  NOR2_X1    g19787(.A1(new_n22931_), .A2(new_n14204_), .ZN(new_n22935_));
  XOR2_X1    g19788(.A1(new_n22935_), .A2(new_n14205_), .Z(new_n22936_));
  NAND2_X1   g19789(.A1(new_n22936_), .A2(new_n22934_), .ZN(new_n22937_));
  NOR2_X1    g19790(.A1(new_n22910_), .A2(new_n18968_), .ZN(new_n22938_));
  NAND2_X1   g19791(.A1(new_n18967_), .A2(new_n22824_), .ZN(new_n22939_));
  XOR2_X1    g19792(.A1(new_n22938_), .A2(new_n22939_), .Z(new_n22940_));
  NAND2_X1   g19793(.A1(new_n22940_), .A2(pi0715), .ZN(new_n22941_));
  XOR2_X1    g19794(.A1(new_n22941_), .A2(new_n14217_), .Z(new_n22942_));
  AOI21_X1   g19795(.A1(new_n22942_), .A2(new_n22824_), .B(pi1160), .ZN(new_n22943_));
  NAND2_X1   g19796(.A1(new_n22940_), .A2(pi0644), .ZN(new_n22944_));
  XOR2_X1    g19797(.A1(new_n22944_), .A2(new_n14205_), .Z(new_n22945_));
  OAI21_X1   g19798(.A1(new_n22945_), .A2(new_n22920_), .B(new_n14203_), .ZN(new_n22946_));
  AOI21_X1   g19799(.A1(new_n22937_), .A2(new_n22943_), .B(new_n22946_), .ZN(new_n22947_));
  NOR2_X1    g19800(.A1(new_n22931_), .A2(new_n14200_), .ZN(new_n22948_));
  XOR2_X1    g19801(.A1(new_n22948_), .A2(new_n14205_), .Z(new_n22949_));
  NAND2_X1   g19802(.A1(new_n22949_), .A2(new_n22934_), .ZN(new_n22950_));
  OAI21_X1   g19803(.A1(new_n22947_), .A2(new_n22950_), .B(pi0832), .ZN(new_n22951_));
  XOR2_X1    g19804(.A1(new_n22951_), .A2(new_n14801_), .Z(new_n22952_));
  NAND2_X1   g19805(.A1(po1038), .A2(new_n10659_), .ZN(new_n22953_));
  NAND4_X1   g19806(.A1(new_n22952_), .A2(new_n14799_), .A3(new_n22931_), .A4(new_n22953_), .ZN(new_n22954_));
  NAND2_X1   g19807(.A1(new_n22954_), .A2(new_n7240_), .ZN(new_n22955_));
  OAI21_X1   g19808(.A1(new_n22822_), .A2(new_n22823_), .B(new_n22955_), .ZN(new_n22956_));
  AOI21_X1   g19809(.A1(new_n16875_), .A2(new_n22690_), .B(new_n22956_), .ZN(new_n22957_));
  OAI21_X1   g19810(.A1(new_n22821_), .A2(pi0792), .B(new_n22957_), .ZN(new_n22958_));
  AOI21_X1   g19811(.A1(new_n22718_), .A2(new_n22706_), .B(new_n22958_), .ZN(po0342));
  NOR2_X1    g19812(.A1(new_n13097_), .A2(new_n3259_), .ZN(new_n22960_));
  NOR2_X1    g19813(.A1(new_n3259_), .A2(new_n7489_), .ZN(new_n22961_));
  XOR2_X1    g19814(.A1(new_n22960_), .A2(new_n22961_), .Z(new_n22962_));
  NAND2_X1   g19815(.A1(new_n22962_), .A2(new_n13624_), .ZN(new_n22963_));
  NAND2_X1   g19816(.A1(new_n19642_), .A2(pi0186), .ZN(new_n22964_));
  OAI22_X1   g19817(.A1(new_n19637_), .A2(new_n22964_), .B1(pi0186), .B2(pi0752), .ZN(new_n22965_));
  NAND2_X1   g19818(.A1(new_n22965_), .A2(new_n15556_), .ZN(new_n22966_));
  NAND2_X1   g19819(.A1(new_n22966_), .A2(new_n3289_), .ZN(new_n22967_));
  AOI21_X1   g19820(.A1(new_n22963_), .A2(pi0752), .B(new_n22967_), .ZN(new_n22968_));
  NOR2_X1    g19821(.A1(new_n3289_), .A2(pi0186), .ZN(new_n22969_));
  NOR2_X1    g19822(.A1(new_n22968_), .A2(new_n22969_), .ZN(new_n22970_));
  INV_X1     g19823(.I(new_n22963_), .ZN(new_n22971_));
  AOI21_X1   g19824(.A1(new_n22966_), .A2(new_n17777_), .B(new_n17769_), .ZN(new_n22972_));
  AOI21_X1   g19825(.A1(new_n22971_), .A2(new_n22972_), .B(new_n3290_), .ZN(new_n22973_));
  INV_X1     g19826(.I(new_n15607_), .ZN(new_n22974_));
  NAND2_X1   g19827(.A1(new_n17769_), .A2(pi0703), .ZN(new_n22975_));
  OAI21_X1   g19828(.A1(new_n22974_), .A2(new_n22975_), .B(new_n7489_), .ZN(new_n22976_));
  AOI21_X1   g19829(.A1(new_n15630_), .A2(new_n17769_), .B(new_n7489_), .ZN(new_n22977_));
  NAND4_X1   g19830(.A1(new_n22976_), .A2(new_n15615_), .A3(new_n15628_), .A4(new_n22977_), .ZN(new_n22978_));
  NAND2_X1   g19831(.A1(new_n22978_), .A2(new_n15595_), .ZN(new_n22979_));
  NOR2_X1    g19832(.A1(new_n3290_), .A2(new_n7489_), .ZN(new_n22980_));
  NAND2_X1   g19833(.A1(new_n22979_), .A2(new_n22980_), .ZN(new_n22981_));
  NOR2_X1    g19834(.A1(new_n22973_), .A2(new_n22981_), .ZN(new_n22982_));
  INV_X1     g19835(.I(new_n22982_), .ZN(new_n22983_));
  NAND2_X1   g19836(.A1(new_n22973_), .A2(new_n22981_), .ZN(new_n22984_));
  NAND3_X1   g19837(.A1(new_n22983_), .A2(pi1153), .A3(new_n22984_), .ZN(new_n22985_));
  NAND2_X1   g19838(.A1(new_n22985_), .A2(new_n13615_), .ZN(new_n22986_));
  INV_X1     g19839(.I(new_n22984_), .ZN(new_n22987_));
  NOR3_X1    g19840(.A1(new_n22987_), .A2(new_n13614_), .A3(new_n22982_), .ZN(new_n22988_));
  NAND2_X1   g19841(.A1(new_n22988_), .A2(new_n13620_), .ZN(new_n22989_));
  AOI21_X1   g19842(.A1(new_n22989_), .A2(new_n22986_), .B(new_n22970_), .ZN(new_n22990_));
  NOR2_X1    g19843(.A1(new_n14428_), .A2(pi0186), .ZN(new_n22991_));
  NAND3_X1   g19844(.A1(new_n14422_), .A2(pi0038), .A3(pi0186), .ZN(new_n22992_));
  NAND3_X1   g19845(.A1(new_n14424_), .A2(new_n3259_), .A3(pi0186), .ZN(new_n22993_));
  AOI21_X1   g19846(.A1(new_n22993_), .A2(new_n22992_), .B(new_n14404_), .ZN(new_n22994_));
  OAI21_X1   g19847(.A1(new_n13721_), .A2(new_n17777_), .B(new_n7489_), .ZN(new_n22995_));
  NAND2_X1   g19848(.A1(new_n22995_), .A2(new_n13108_), .ZN(new_n22996_));
  OAI21_X1   g19849(.A1(new_n22994_), .A2(new_n22996_), .B(new_n3289_), .ZN(new_n22997_));
  NAND3_X1   g19850(.A1(new_n3289_), .A2(pi0186), .A3(new_n17777_), .ZN(new_n22998_));
  NOR2_X1    g19851(.A1(new_n22963_), .A2(new_n22998_), .ZN(new_n22999_));
  NAND2_X1   g19852(.A1(new_n22999_), .A2(new_n22997_), .ZN(new_n23000_));
  INV_X1     g19853(.I(new_n22997_), .ZN(new_n23001_));
  OAI21_X1   g19854(.A1(new_n22963_), .A2(new_n22998_), .B(new_n23001_), .ZN(new_n23002_));
  NAND2_X1   g19855(.A1(new_n23002_), .A2(new_n23000_), .ZN(new_n23003_));
  NAND3_X1   g19856(.A1(new_n23003_), .A2(pi0625), .A3(pi1153), .ZN(new_n23004_));
  INV_X1     g19857(.I(new_n23004_), .ZN(new_n23005_));
  NOR3_X1    g19858(.A1(new_n23003_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n23006_));
  OAI21_X1   g19859(.A1(new_n23005_), .A2(new_n23006_), .B(new_n22991_), .ZN(new_n23007_));
  NAND2_X1   g19860(.A1(new_n23007_), .A2(pi0608), .ZN(new_n23008_));
  OAI21_X1   g19861(.A1(new_n22990_), .A2(new_n23008_), .B(pi0778), .ZN(new_n23009_));
  NAND3_X1   g19862(.A1(new_n22983_), .A2(pi0625), .A3(new_n22984_), .ZN(new_n23010_));
  NAND2_X1   g19863(.A1(new_n23010_), .A2(new_n13615_), .ZN(new_n23011_));
  NOR2_X1    g19864(.A1(new_n22987_), .A2(new_n22982_), .ZN(new_n23012_));
  NAND3_X1   g19865(.A1(new_n23012_), .A2(pi0625), .A3(new_n13620_), .ZN(new_n23013_));
  AOI21_X1   g19866(.A1(new_n23013_), .A2(new_n23011_), .B(new_n22970_), .ZN(new_n23014_));
  INV_X1     g19867(.I(new_n22991_), .ZN(new_n23015_));
  NAND3_X1   g19868(.A1(new_n23003_), .A2(pi0625), .A3(pi1153), .ZN(new_n23016_));
  NAND4_X1   g19869(.A1(new_n23002_), .A2(new_n23000_), .A3(new_n13613_), .A4(pi1153), .ZN(new_n23017_));
  AOI21_X1   g19870(.A1(new_n23016_), .A2(new_n23017_), .B(new_n23015_), .ZN(new_n23018_));
  NOR3_X1    g19871(.A1(new_n23018_), .A2(new_n13750_), .A3(new_n23012_), .ZN(new_n23019_));
  INV_X1     g19872(.I(new_n23019_), .ZN(new_n23020_));
  NOR2_X1    g19873(.A1(new_n23020_), .A2(new_n23014_), .ZN(new_n23021_));
  NAND2_X1   g19874(.A1(new_n23009_), .A2(new_n23021_), .ZN(new_n23022_));
  INV_X1     g19875(.I(new_n22970_), .ZN(new_n23023_));
  NOR2_X1    g19876(.A1(new_n22988_), .A2(new_n13620_), .ZN(new_n23024_));
  NOR2_X1    g19877(.A1(new_n22985_), .A2(new_n13615_), .ZN(new_n23025_));
  OAI21_X1   g19878(.A1(new_n23024_), .A2(new_n23025_), .B(new_n23023_), .ZN(new_n23026_));
  INV_X1     g19879(.I(new_n23006_), .ZN(new_n23027_));
  AOI21_X1   g19880(.A1(new_n23027_), .A2(new_n23004_), .B(new_n23015_), .ZN(new_n23028_));
  NOR2_X1    g19881(.A1(new_n23028_), .A2(new_n14081_), .ZN(new_n23029_));
  AOI21_X1   g19882(.A1(new_n23026_), .A2(new_n23029_), .B(new_n13748_), .ZN(new_n23030_));
  XOR2_X1    g19883(.A1(new_n23010_), .A2(new_n13615_), .Z(new_n23031_));
  OAI21_X1   g19884(.A1(new_n23031_), .A2(new_n22970_), .B(new_n23019_), .ZN(new_n23032_));
  NAND2_X1   g19885(.A1(new_n23032_), .A2(new_n23030_), .ZN(new_n23033_));
  NAND2_X1   g19886(.A1(new_n23033_), .A2(new_n23022_), .ZN(new_n23034_));
  NAND4_X1   g19887(.A1(new_n23028_), .A2(new_n23018_), .A3(pi0778), .A4(new_n23003_), .ZN(new_n23035_));
  NAND3_X1   g19888(.A1(new_n23018_), .A2(pi0778), .A3(new_n23003_), .ZN(new_n23036_));
  NAND3_X1   g19889(.A1(new_n23036_), .A2(pi0778), .A3(new_n23007_), .ZN(new_n23037_));
  NAND2_X1   g19890(.A1(new_n23037_), .A2(new_n23035_), .ZN(new_n23038_));
  NAND2_X1   g19891(.A1(new_n22970_), .A2(new_n13776_), .ZN(new_n23039_));
  NOR2_X1    g19892(.A1(new_n22991_), .A2(new_n15147_), .ZN(new_n23041_));
  OAI21_X1   g19893(.A1(new_n23038_), .A2(new_n13785_), .B(new_n13766_), .ZN(new_n23042_));
  AOI21_X1   g19894(.A1(new_n23037_), .A2(new_n23035_), .B(new_n13766_), .ZN(new_n23043_));
  OAI21_X1   g19895(.A1(new_n22991_), .A2(new_n15707_), .B(new_n13766_), .ZN(new_n23044_));
  INV_X1     g19896(.I(new_n23044_), .ZN(new_n23045_));
  NOR2_X1    g19897(.A1(new_n23039_), .A2(new_n23045_), .ZN(new_n23046_));
  NOR2_X1    g19898(.A1(new_n23046_), .A2(new_n14465_), .ZN(new_n23047_));
  INV_X1     g19899(.I(new_n23047_), .ZN(new_n23048_));
  OAI21_X1   g19900(.A1(new_n23043_), .A2(new_n23048_), .B(new_n13766_), .ZN(new_n23049_));
  NAND4_X1   g19901(.A1(new_n23034_), .A2(new_n23049_), .A3(new_n23042_), .A4(pi0785), .ZN(new_n23050_));
  NAND2_X1   g19902(.A1(new_n23034_), .A2(new_n23042_), .ZN(new_n23051_));
  NAND3_X1   g19903(.A1(new_n23034_), .A2(new_n23049_), .A3(pi0785), .ZN(new_n23052_));
  NAND3_X1   g19904(.A1(new_n23052_), .A2(new_n23051_), .A3(pi0785), .ZN(new_n23053_));
  NAND2_X1   g19905(.A1(new_n23053_), .A2(new_n23050_), .ZN(new_n23054_));
  AOI21_X1   g19906(.A1(new_n22970_), .A2(new_n13776_), .B(new_n23041_), .ZN(new_n23055_));
  OAI21_X1   g19907(.A1(new_n23055_), .A2(new_n13766_), .B(pi0785), .ZN(new_n23056_));
  NAND2_X1   g19908(.A1(new_n22991_), .A2(new_n13775_), .ZN(new_n23057_));
  OAI21_X1   g19909(.A1(new_n22970_), .A2(new_n13775_), .B(new_n23057_), .ZN(new_n23058_));
  NAND3_X1   g19910(.A1(new_n23046_), .A2(pi0785), .A3(new_n23058_), .ZN(new_n23059_));
  XOR2_X1    g19911(.A1(new_n23059_), .A2(new_n23056_), .Z(new_n23060_));
  NAND3_X1   g19912(.A1(new_n23060_), .A2(pi0618), .A3(pi1154), .ZN(new_n23061_));
  XNOR2_X1   g19913(.A1(new_n23059_), .A2(new_n23056_), .ZN(new_n23062_));
  NAND3_X1   g19914(.A1(new_n23062_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n23063_));
  AOI21_X1   g19915(.A1(new_n23063_), .A2(new_n23061_), .B(new_n23015_), .ZN(new_n23064_));
  AOI21_X1   g19916(.A1(new_n23037_), .A2(new_n23035_), .B(new_n13803_), .ZN(new_n23065_));
  NOR2_X1    g19917(.A1(new_n23015_), .A2(new_n13805_), .ZN(new_n23066_));
  NOR2_X1    g19918(.A1(new_n23065_), .A2(new_n23066_), .ZN(new_n23067_));
  OAI21_X1   g19919(.A1(new_n23067_), .A2(pi0618), .B(new_n13824_), .ZN(new_n23068_));
  OAI21_X1   g19920(.A1(new_n23068_), .A2(new_n23064_), .B(new_n13816_), .ZN(new_n23069_));
  AOI21_X1   g19921(.A1(new_n23062_), .A2(pi1154), .B(new_n13819_), .ZN(new_n23070_));
  NOR3_X1    g19922(.A1(new_n23060_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n23071_));
  OAI21_X1   g19923(.A1(new_n23070_), .A2(new_n23071_), .B(new_n22991_), .ZN(new_n23072_));
  OAI21_X1   g19924(.A1(new_n23065_), .A2(new_n23066_), .B(pi0618), .ZN(new_n23073_));
  NAND3_X1   g19925(.A1(new_n23072_), .A2(new_n23073_), .A3(new_n13836_), .ZN(new_n23074_));
  NAND2_X1   g19926(.A1(new_n23074_), .A2(new_n13816_), .ZN(new_n23075_));
  NAND4_X1   g19927(.A1(new_n23054_), .A2(pi0781), .A3(new_n23069_), .A4(new_n23075_), .ZN(new_n23076_));
  INV_X1     g19928(.I(new_n23050_), .ZN(new_n23077_));
  NOR2_X1    g19929(.A1(new_n23032_), .A2(new_n23030_), .ZN(new_n23078_));
  NOR2_X1    g19930(.A1(new_n23009_), .A2(new_n23021_), .ZN(new_n23079_));
  NOR2_X1    g19931(.A1(new_n23078_), .A2(new_n23079_), .ZN(new_n23080_));
  INV_X1     g19932(.I(new_n23042_), .ZN(new_n23081_));
  OAI21_X1   g19933(.A1(new_n23080_), .A2(new_n23081_), .B(pi0785), .ZN(new_n23082_));
  INV_X1     g19934(.I(new_n23049_), .ZN(new_n23083_));
  NOR3_X1    g19935(.A1(new_n23083_), .A2(new_n23080_), .A3(new_n13801_), .ZN(new_n23084_));
  NOR2_X1    g19936(.A1(new_n23084_), .A2(new_n23082_), .ZN(new_n23085_));
  OAI21_X1   g19937(.A1(new_n23085_), .A2(new_n23077_), .B(new_n23069_), .ZN(new_n23086_));
  AOI21_X1   g19938(.A1(new_n23074_), .A2(new_n13816_), .B(new_n13855_), .ZN(new_n23087_));
  OAI21_X1   g19939(.A1(new_n23085_), .A2(new_n23077_), .B(new_n23087_), .ZN(new_n23088_));
  NAND3_X1   g19940(.A1(new_n23088_), .A2(new_n23086_), .A3(pi0781), .ZN(new_n23089_));
  NAND2_X1   g19941(.A1(new_n23089_), .A2(new_n23076_), .ZN(new_n23090_));
  NAND3_X1   g19942(.A1(new_n23060_), .A2(pi0618), .A3(pi1154), .ZN(new_n23091_));
  NAND3_X1   g19943(.A1(new_n23062_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n23092_));
  AOI21_X1   g19944(.A1(new_n23092_), .A2(new_n23091_), .B(new_n23015_), .ZN(new_n23093_));
  NAND4_X1   g19945(.A1(new_n23064_), .A2(new_n23093_), .A3(pi0781), .A4(new_n23060_), .ZN(new_n23094_));
  NOR2_X1    g19946(.A1(new_n23064_), .A2(new_n13855_), .ZN(new_n23095_));
  NAND3_X1   g19947(.A1(new_n23093_), .A2(pi0781), .A3(new_n23060_), .ZN(new_n23096_));
  NAND2_X1   g19948(.A1(new_n23096_), .A2(new_n23095_), .ZN(new_n23097_));
  NAND2_X1   g19949(.A1(new_n23097_), .A2(new_n23094_), .ZN(new_n23098_));
  NAND3_X1   g19950(.A1(new_n23098_), .A2(pi0619), .A3(pi1159), .ZN(new_n23099_));
  NAND4_X1   g19951(.A1(new_n23097_), .A2(pi0619), .A3(new_n13868_), .A4(new_n23094_), .ZN(new_n23100_));
  AOI21_X1   g19952(.A1(new_n23099_), .A2(new_n23100_), .B(new_n23015_), .ZN(new_n23101_));
  NOR2_X1    g19953(.A1(new_n22991_), .A2(new_n13880_), .ZN(new_n23102_));
  AOI21_X1   g19954(.A1(new_n23067_), .A2(new_n13880_), .B(new_n23102_), .ZN(new_n23103_));
  AOI21_X1   g19955(.A1(new_n23103_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n23104_));
  INV_X1     g19956(.I(new_n23104_), .ZN(new_n23105_));
  OAI21_X1   g19957(.A1(new_n23101_), .A2(new_n23105_), .B(new_n13860_), .ZN(new_n23106_));
  NAND3_X1   g19958(.A1(new_n23098_), .A2(pi0619), .A3(pi1159), .ZN(new_n23107_));
  NAND4_X1   g19959(.A1(new_n23097_), .A2(new_n13860_), .A3(pi1159), .A4(new_n23094_), .ZN(new_n23108_));
  AOI21_X1   g19960(.A1(new_n23107_), .A2(new_n23108_), .B(new_n23015_), .ZN(new_n23109_));
  AOI21_X1   g19961(.A1(new_n23103_), .A2(pi0619), .B(new_n15217_), .ZN(new_n23110_));
  INV_X1     g19962(.I(new_n23110_), .ZN(new_n23111_));
  OAI21_X1   g19963(.A1(new_n23109_), .A2(new_n23111_), .B(new_n13860_), .ZN(new_n23112_));
  NAND4_X1   g19964(.A1(new_n23106_), .A2(new_n23112_), .A3(new_n23090_), .A4(pi0789), .ZN(new_n23113_));
  NAND2_X1   g19965(.A1(new_n23106_), .A2(new_n23090_), .ZN(new_n23114_));
  NAND3_X1   g19966(.A1(new_n23112_), .A2(new_n23090_), .A3(pi0789), .ZN(new_n23115_));
  NAND3_X1   g19967(.A1(new_n23115_), .A2(new_n23114_), .A3(pi0789), .ZN(new_n23116_));
  NAND2_X1   g19968(.A1(new_n23116_), .A2(new_n23113_), .ZN(new_n23117_));
  NAND4_X1   g19969(.A1(new_n23101_), .A2(new_n23109_), .A3(pi0789), .A4(new_n23098_), .ZN(new_n23118_));
  XOR2_X1    g19970(.A1(new_n23096_), .A2(new_n23095_), .Z(new_n23119_));
  AOI21_X1   g19971(.A1(new_n23119_), .A2(pi0619), .B(new_n13904_), .ZN(new_n23120_));
  INV_X1     g19972(.I(new_n23100_), .ZN(new_n23121_));
  OAI21_X1   g19973(.A1(new_n23120_), .A2(new_n23121_), .B(new_n22991_), .ZN(new_n23122_));
  NAND3_X1   g19974(.A1(new_n23109_), .A2(pi0789), .A3(new_n23098_), .ZN(new_n23123_));
  NAND3_X1   g19975(.A1(new_n23123_), .A2(pi0789), .A3(new_n23122_), .ZN(new_n23124_));
  NOR2_X1    g19976(.A1(new_n23015_), .A2(new_n13919_), .ZN(new_n23125_));
  AOI21_X1   g19977(.A1(new_n23103_), .A2(new_n13919_), .B(new_n23125_), .ZN(new_n23126_));
  NOR2_X1    g19978(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n23127_));
  INV_X1     g19979(.I(new_n23127_), .ZN(new_n23128_));
  AOI21_X1   g19980(.A1(new_n23124_), .A2(new_n23118_), .B(new_n23128_), .ZN(new_n23129_));
  NAND3_X1   g19981(.A1(new_n23117_), .A2(pi0626), .A3(pi0788), .ZN(new_n23134_));
  INV_X1     g19982(.I(new_n23134_), .ZN(new_n23135_));
  INV_X1     g19983(.I(new_n23118_), .ZN(new_n23136_));
  NAND2_X1   g19984(.A1(new_n23122_), .A2(pi0789), .ZN(new_n23137_));
  AOI21_X1   g19985(.A1(new_n23119_), .A2(pi1159), .B(new_n13904_), .ZN(new_n23138_));
  INV_X1     g19986(.I(new_n23108_), .ZN(new_n23139_));
  OAI21_X1   g19987(.A1(new_n23138_), .A2(new_n23139_), .B(new_n22991_), .ZN(new_n23140_));
  NOR3_X1    g19988(.A1(new_n23140_), .A2(new_n13896_), .A3(new_n23119_), .ZN(new_n23141_));
  NOR2_X1    g19989(.A1(new_n23141_), .A2(new_n23137_), .ZN(new_n23142_));
  OAI21_X1   g19990(.A1(new_n23142_), .A2(new_n23136_), .B(new_n23127_), .ZN(new_n23143_));
  AOI22_X1   g19991(.A1(new_n23143_), .A2(new_n13901_), .B1(new_n23116_), .B2(new_n23113_), .ZN(new_n23144_));
  AOI21_X1   g19992(.A1(new_n23116_), .A2(new_n23113_), .B(new_n15258_), .ZN(new_n23145_));
  NOR3_X1    g19993(.A1(new_n23144_), .A2(new_n13937_), .A3(new_n23145_), .ZN(new_n23146_));
  NOR2_X1    g19994(.A1(new_n23146_), .A2(new_n23135_), .ZN(new_n23147_));
  NOR2_X1    g19995(.A1(new_n22991_), .A2(new_n16372_), .ZN(new_n23148_));
  INV_X1     g19996(.I(new_n23148_), .ZN(new_n23149_));
  NAND3_X1   g19997(.A1(new_n23124_), .A2(new_n16372_), .A3(new_n23118_), .ZN(new_n23150_));
  NAND2_X1   g19998(.A1(new_n23150_), .A2(new_n23149_), .ZN(new_n23151_));
  NOR2_X1    g19999(.A1(new_n22991_), .A2(new_n13966_), .ZN(new_n23153_));
  AOI21_X1   g20000(.A1(new_n23126_), .A2(new_n13966_), .B(new_n23153_), .ZN(new_n23154_));
  AOI21_X1   g20001(.A1(new_n23154_), .A2(pi0628), .B(new_n13971_), .ZN(new_n23155_));
  INV_X1     g20002(.I(new_n23155_), .ZN(new_n23156_));
  NAND3_X1   g20003(.A1(new_n23154_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n23157_));
  AOI21_X1   g20004(.A1(new_n23156_), .A2(new_n23157_), .B(new_n23015_), .ZN(new_n23158_));
  NOR2_X1    g20005(.A1(new_n23158_), .A2(new_n15270_), .ZN(new_n23159_));
  AOI21_X1   g20006(.A1(new_n23154_), .A2(pi1156), .B(new_n13971_), .ZN(new_n23162_));
  INV_X1     g20007(.I(new_n23162_), .ZN(new_n23163_));
  NAND3_X1   g20008(.A1(new_n23154_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n23164_));
  AOI21_X1   g20009(.A1(new_n23163_), .A2(new_n23164_), .B(new_n23015_), .ZN(new_n23165_));
  NOR3_X1    g20010(.A1(new_n23147_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n23169_));
  INV_X1     g20011(.I(new_n23113_), .ZN(new_n23170_));
  AOI21_X1   g20012(.A1(pi0781), .A2(new_n23086_), .B(new_n23088_), .ZN(new_n23171_));
  INV_X1     g20013(.I(new_n23069_), .ZN(new_n23172_));
  AOI21_X1   g20014(.A1(new_n23050_), .A2(new_n23053_), .B(new_n23172_), .ZN(new_n23173_));
  NAND2_X1   g20015(.A1(new_n23073_), .A2(new_n13836_), .ZN(new_n23174_));
  NOR2_X1    g20016(.A1(new_n23174_), .A2(new_n23093_), .ZN(new_n23175_));
  OAI21_X1   g20017(.A1(new_n23175_), .A2(pi0618), .B(pi0781), .ZN(new_n23176_));
  AOI21_X1   g20018(.A1(new_n23050_), .A2(new_n23053_), .B(new_n23176_), .ZN(new_n23177_));
  NOR3_X1    g20019(.A1(new_n23177_), .A2(new_n23173_), .A3(new_n13855_), .ZN(new_n23178_));
  NOR2_X1    g20020(.A1(new_n23178_), .A2(new_n23171_), .ZN(new_n23179_));
  AOI21_X1   g20021(.A1(new_n23122_), .A2(new_n23104_), .B(pi0619), .ZN(new_n23180_));
  OAI21_X1   g20022(.A1(new_n23180_), .A2(new_n23179_), .B(pi0789), .ZN(new_n23181_));
  AOI21_X1   g20023(.A1(new_n23140_), .A2(new_n23110_), .B(pi0619), .ZN(new_n23182_));
  OAI21_X1   g20024(.A1(new_n23178_), .A2(new_n23171_), .B(pi0789), .ZN(new_n23183_));
  NOR2_X1    g20025(.A1(new_n23182_), .A2(new_n23183_), .ZN(new_n23184_));
  NOR2_X1    g20026(.A1(new_n23181_), .A2(new_n23184_), .ZN(new_n23185_));
  OAI22_X1   g20027(.A1(new_n23185_), .A2(new_n23170_), .B1(new_n23129_), .B2(pi0626), .ZN(new_n23186_));
  OAI21_X1   g20028(.A1(new_n23185_), .A2(new_n23170_), .B(new_n14577_), .ZN(new_n23187_));
  NAND3_X1   g20029(.A1(new_n23186_), .A2(new_n23187_), .A3(pi0788), .ZN(new_n23188_));
  AOI21_X1   g20030(.A1(new_n23151_), .A2(new_n23159_), .B(pi0628), .ZN(new_n23189_));
  AOI21_X1   g20031(.A1(new_n23188_), .A2(new_n23134_), .B(new_n23189_), .ZN(new_n23190_));
  AOI21_X1   g20032(.A1(new_n23188_), .A2(new_n23134_), .B(new_n15296_), .ZN(new_n23191_));
  NOR3_X1    g20033(.A1(new_n23190_), .A2(new_n23191_), .A3(new_n12777_), .ZN(new_n23192_));
  NOR2_X1    g20034(.A1(new_n23192_), .A2(new_n23169_), .ZN(new_n23193_));
  INV_X1     g20035(.I(new_n23154_), .ZN(new_n23194_));
  NAND4_X1   g20036(.A1(new_n23158_), .A2(new_n23165_), .A3(pi0792), .A4(new_n23194_), .ZN(new_n23195_));
  INV_X1     g20037(.I(new_n23157_), .ZN(new_n23196_));
  OAI21_X1   g20038(.A1(new_n23196_), .A2(new_n23155_), .B(new_n22991_), .ZN(new_n23197_));
  NOR2_X1    g20039(.A1(new_n23154_), .A2(new_n12777_), .ZN(new_n23198_));
  NAND2_X1   g20040(.A1(new_n23165_), .A2(new_n23198_), .ZN(new_n23199_));
  NAND3_X1   g20041(.A1(new_n23199_), .A2(pi0792), .A3(new_n23197_), .ZN(new_n23200_));
  NAND2_X1   g20042(.A1(new_n23200_), .A2(new_n23195_), .ZN(new_n23201_));
  NAND3_X1   g20043(.A1(new_n23201_), .A2(pi0647), .A3(pi1157), .ZN(new_n23202_));
  INV_X1     g20044(.I(new_n23202_), .ZN(new_n23203_));
  NOR3_X1    g20045(.A1(new_n23201_), .A2(new_n14005_), .A3(pi1157), .ZN(new_n23204_));
  OAI21_X1   g20046(.A1(new_n23203_), .A2(new_n23204_), .B(new_n22991_), .ZN(new_n23205_));
  AOI21_X1   g20047(.A1(new_n23150_), .A2(new_n23149_), .B(new_n13993_), .ZN(new_n23206_));
  NOR2_X1    g20048(.A1(new_n22991_), .A2(new_n13994_), .ZN(new_n23207_));
  NOR2_X1    g20049(.A1(new_n23206_), .A2(new_n23207_), .ZN(new_n23208_));
  AOI21_X1   g20050(.A1(new_n23208_), .A2(new_n14005_), .B(new_n14012_), .ZN(new_n23209_));
  AOI21_X1   g20051(.A1(new_n23205_), .A2(new_n23209_), .B(pi0647), .ZN(new_n23210_));
  NAND3_X1   g20052(.A1(new_n23201_), .A2(pi0647), .A3(pi1157), .ZN(new_n23211_));
  NAND4_X1   g20053(.A1(new_n23200_), .A2(new_n23195_), .A3(new_n14005_), .A4(pi1157), .ZN(new_n23212_));
  AOI21_X1   g20054(.A1(new_n23211_), .A2(new_n23212_), .B(new_n23015_), .ZN(new_n23213_));
  NOR3_X1    g20055(.A1(new_n23206_), .A2(new_n14005_), .A3(new_n23207_), .ZN(new_n23214_));
  NOR3_X1    g20056(.A1(new_n23213_), .A2(new_n23214_), .A3(new_n16329_), .ZN(new_n23215_));
  NOR2_X1    g20057(.A1(new_n23215_), .A2(pi0647), .ZN(new_n23216_));
  NOR4_X1    g20058(.A1(new_n23193_), .A2(new_n12776_), .A3(new_n23210_), .A4(new_n23216_), .ZN(new_n23217_));
  NAND2_X1   g20059(.A1(new_n23188_), .A2(new_n23134_), .ZN(new_n23218_));
  NAND3_X1   g20060(.A1(new_n23218_), .A2(pi0628), .A3(pi0792), .ZN(new_n23219_));
  INV_X1     g20061(.I(new_n23189_), .ZN(new_n23220_));
  OAI21_X1   g20062(.A1(new_n23146_), .A2(new_n23135_), .B(new_n23220_), .ZN(new_n23221_));
  OAI21_X1   g20063(.A1(new_n23146_), .A2(new_n23135_), .B(new_n14606_), .ZN(new_n23222_));
  NAND3_X1   g20064(.A1(new_n23221_), .A2(new_n23222_), .A3(pi0792), .ZN(new_n23223_));
  AOI21_X1   g20065(.A1(new_n23223_), .A2(new_n23219_), .B(new_n23210_), .ZN(new_n23224_));
  OAI21_X1   g20066(.A1(new_n23215_), .A2(pi0647), .B(pi0787), .ZN(new_n23225_));
  AOI21_X1   g20067(.A1(new_n23223_), .A2(new_n23219_), .B(new_n23225_), .ZN(new_n23226_));
  NOR3_X1    g20068(.A1(new_n23226_), .A2(new_n23224_), .A3(new_n12776_), .ZN(new_n23227_));
  OAI21_X1   g20069(.A1(new_n23227_), .A2(new_n23217_), .B(new_n12775_), .ZN(new_n23228_));
  NOR2_X1    g20070(.A1(new_n9992_), .A2(pi0186), .ZN(new_n23229_));
  NOR2_X1    g20071(.A1(new_n14652_), .A2(new_n17777_), .ZN(new_n23230_));
  AOI21_X1   g20072(.A1(new_n13218_), .A2(pi0703), .B(new_n23229_), .ZN(new_n23231_));
  INV_X1     g20073(.I(new_n23231_), .ZN(new_n23232_));
  NAND3_X1   g20074(.A1(new_n23232_), .A2(new_n23230_), .A3(new_n23229_), .ZN(new_n23233_));
  NOR3_X1    g20075(.A1(new_n23230_), .A2(new_n13614_), .A3(new_n23231_), .ZN(new_n23234_));
  XNOR2_X1   g20076(.A1(new_n23233_), .A2(new_n23234_), .ZN(new_n23235_));
  NAND2_X1   g20077(.A1(new_n23235_), .A2(pi0778), .ZN(new_n23236_));
  NAND2_X1   g20078(.A1(new_n23232_), .A2(new_n13748_), .ZN(new_n23237_));
  NAND2_X1   g20079(.A1(new_n23236_), .A2(new_n23237_), .ZN(new_n23238_));
  INV_X1     g20080(.I(new_n23238_), .ZN(new_n23239_));
  NOR2_X1    g20081(.A1(new_n23239_), .A2(new_n14048_), .ZN(new_n23240_));
  INV_X1     g20082(.I(new_n23240_), .ZN(new_n23241_));
  NOR2_X1    g20083(.A1(new_n23241_), .A2(new_n14051_), .ZN(new_n23242_));
  INV_X1     g20084(.I(new_n23242_), .ZN(new_n23243_));
  NOR2_X1    g20085(.A1(new_n23243_), .A2(new_n14163_), .ZN(new_n23244_));
  AOI21_X1   g20086(.A1(new_n13104_), .A2(new_n17769_), .B(new_n23229_), .ZN(new_n23245_));
  NOR2_X1    g20087(.A1(new_n14096_), .A2(new_n23245_), .ZN(new_n23246_));
  AOI21_X1   g20088(.A1(new_n23246_), .A2(new_n14094_), .B(pi1155), .ZN(new_n23247_));
  NOR2_X1    g20089(.A1(new_n23247_), .A2(new_n13801_), .ZN(new_n23248_));
  AOI21_X1   g20090(.A1(new_n23245_), .A2(pi1155), .B(new_n9992_), .ZN(new_n23249_));
  NOR2_X1    g20091(.A1(new_n23249_), .A2(new_n14102_), .ZN(new_n23250_));
  NAND3_X1   g20092(.A1(new_n23250_), .A2(new_n23246_), .A3(pi0785), .ZN(new_n23251_));
  XOR2_X1    g20093(.A1(new_n23248_), .A2(new_n23251_), .Z(new_n23252_));
  NOR2_X1    g20094(.A1(new_n23252_), .A2(new_n13817_), .ZN(new_n23253_));
  OAI21_X1   g20095(.A1(new_n23253_), .A2(pi0618), .B(new_n9992_), .ZN(new_n23254_));
  NAND2_X1   g20096(.A1(new_n23254_), .A2(pi0781), .ZN(new_n23255_));
  OAI21_X1   g20097(.A1(new_n23253_), .A2(new_n9992_), .B(pi0618), .ZN(new_n23256_));
  NOR3_X1    g20098(.A1(new_n23256_), .A2(new_n13855_), .A3(new_n23252_), .ZN(new_n23257_));
  XOR2_X1    g20099(.A1(new_n23257_), .A2(new_n23255_), .Z(new_n23258_));
  NAND2_X1   g20100(.A1(new_n23258_), .A2(pi0619), .ZN(new_n23259_));
  XOR2_X1    g20101(.A1(new_n23259_), .A2(new_n13904_), .Z(new_n23260_));
  NAND2_X1   g20102(.A1(new_n23260_), .A2(new_n23229_), .ZN(new_n23261_));
  NAND2_X1   g20103(.A1(new_n23261_), .A2(pi0789), .ZN(new_n23262_));
  NAND2_X1   g20104(.A1(new_n23258_), .A2(pi1159), .ZN(new_n23263_));
  XOR2_X1    g20105(.A1(new_n23263_), .A2(new_n13904_), .Z(new_n23264_));
  NAND2_X1   g20106(.A1(new_n23264_), .A2(new_n23229_), .ZN(new_n23265_));
  NOR3_X1    g20107(.A1(new_n23265_), .A2(new_n13896_), .A3(new_n23258_), .ZN(new_n23266_));
  XOR2_X1    g20108(.A1(new_n23266_), .A2(new_n23262_), .Z(new_n23267_));
  NAND2_X1   g20109(.A1(new_n23267_), .A2(new_n13962_), .ZN(new_n23268_));
  XOR2_X1    g20110(.A1(new_n23268_), .A2(new_n18976_), .Z(new_n23269_));
  AOI22_X1   g20111(.A1(new_n23269_), .A2(new_n23229_), .B1(new_n16639_), .B2(new_n23244_), .ZN(new_n23270_));
  NOR2_X1    g20112(.A1(new_n23231_), .A2(new_n13203_), .ZN(new_n23271_));
  INV_X1     g20113(.I(new_n23271_), .ZN(new_n23272_));
  NOR2_X1    g20114(.A1(new_n23272_), .A2(new_n13613_), .ZN(new_n23273_));
  NOR2_X1    g20115(.A1(new_n23229_), .A2(pi1153), .ZN(new_n23274_));
  INV_X1     g20116(.I(new_n23274_), .ZN(new_n23275_));
  OAI21_X1   g20117(.A1(new_n23230_), .A2(new_n23275_), .B(pi0608), .ZN(new_n23276_));
  NOR2_X1    g20118(.A1(new_n23245_), .A2(pi1153), .ZN(new_n23277_));
  NAND2_X1   g20119(.A1(new_n23276_), .A2(new_n23277_), .ZN(new_n23278_));
  AOI21_X1   g20120(.A1(new_n23278_), .A2(new_n23273_), .B(new_n13748_), .ZN(new_n23279_));
  NOR2_X1    g20121(.A1(new_n23231_), .A2(new_n14082_), .ZN(new_n23280_));
  NAND2_X1   g20122(.A1(new_n23230_), .A2(new_n23274_), .ZN(new_n23281_));
  OAI22_X1   g20123(.A1(new_n23272_), .A2(new_n13613_), .B1(new_n23281_), .B2(new_n23280_), .ZN(new_n23282_));
  NAND4_X1   g20124(.A1(new_n23282_), .A2(pi0778), .A3(new_n23245_), .A4(new_n23272_), .ZN(new_n23283_));
  XNOR2_X1   g20125(.A1(new_n23283_), .A2(new_n23279_), .ZN(new_n23284_));
  NAND2_X1   g20126(.A1(new_n23284_), .A2(new_n13801_), .ZN(new_n23285_));
  NOR2_X1    g20127(.A1(new_n23284_), .A2(new_n13778_), .ZN(new_n23286_));
  XOR2_X1    g20128(.A1(new_n23286_), .A2(new_n14694_), .Z(new_n23287_));
  NOR2_X1    g20129(.A1(new_n23287_), .A2(new_n23239_), .ZN(new_n23288_));
  NOR3_X1    g20130(.A1(new_n23288_), .A2(new_n13783_), .A3(new_n23247_), .ZN(new_n23289_));
  NOR3_X1    g20131(.A1(new_n23289_), .A2(pi0660), .A3(new_n23250_), .ZN(new_n23290_));
  NOR2_X1    g20132(.A1(new_n23284_), .A2(new_n13766_), .ZN(new_n23291_));
  XOR2_X1    g20133(.A1(new_n23291_), .A2(new_n14090_), .Z(new_n23292_));
  NAND3_X1   g20134(.A1(new_n23292_), .A2(pi0785), .A3(new_n23238_), .ZN(new_n23293_));
  OAI21_X1   g20135(.A1(new_n23290_), .A2(new_n23293_), .B(new_n23285_), .ZN(new_n23294_));
  NAND2_X1   g20136(.A1(new_n23294_), .A2(new_n13855_), .ZN(new_n23295_));
  NOR2_X1    g20137(.A1(new_n23294_), .A2(new_n13816_), .ZN(new_n23296_));
  XOR2_X1    g20138(.A1(new_n23296_), .A2(new_n13818_), .Z(new_n23297_));
  NAND2_X1   g20139(.A1(new_n23297_), .A2(new_n23240_), .ZN(new_n23298_));
  NAND3_X1   g20140(.A1(new_n23298_), .A2(new_n13823_), .A3(new_n23256_), .ZN(new_n23299_));
  AND3_X2    g20141(.A1(new_n23299_), .A2(new_n13823_), .A3(new_n23254_), .Z(new_n23300_));
  NOR2_X1    g20142(.A1(new_n23294_), .A2(new_n13817_), .ZN(new_n23301_));
  XOR2_X1    g20143(.A1(new_n23301_), .A2(new_n13819_), .Z(new_n23302_));
  NOR3_X1    g20144(.A1(new_n23302_), .A2(new_n13855_), .A3(new_n23241_), .ZN(new_n23303_));
  INV_X1     g20145(.I(new_n23303_), .ZN(new_n23304_));
  OAI21_X1   g20146(.A1(new_n23300_), .A2(new_n23304_), .B(new_n23295_), .ZN(new_n23305_));
  NOR2_X1    g20147(.A1(new_n23305_), .A2(new_n13860_), .ZN(new_n23306_));
  XOR2_X1    g20148(.A1(new_n23306_), .A2(new_n13904_), .Z(new_n23307_));
  NOR2_X1    g20149(.A1(new_n23307_), .A2(new_n23243_), .ZN(new_n23308_));
  NAND2_X1   g20150(.A1(new_n23265_), .A2(new_n13884_), .ZN(new_n23309_));
  INV_X1     g20151(.I(new_n23305_), .ZN(new_n23310_));
  AOI21_X1   g20152(.A1(new_n23310_), .A2(new_n14143_), .B(pi0789), .ZN(new_n23311_));
  OAI21_X1   g20153(.A1(new_n23308_), .A2(new_n23309_), .B(new_n23311_), .ZN(new_n23312_));
  NOR2_X1    g20154(.A1(new_n23305_), .A2(new_n13868_), .ZN(new_n23313_));
  XOR2_X1    g20155(.A1(new_n23313_), .A2(new_n13903_), .Z(new_n23314_));
  NAND2_X1   g20156(.A1(new_n23261_), .A2(new_n19018_), .ZN(new_n23315_));
  AOI21_X1   g20157(.A1(new_n23314_), .A2(new_n23242_), .B(new_n23315_), .ZN(new_n23316_));
  AOI21_X1   g20158(.A1(new_n23312_), .A2(new_n23316_), .B(new_n23270_), .ZN(new_n23317_));
  NAND2_X1   g20159(.A1(new_n23267_), .A2(new_n16372_), .ZN(new_n23318_));
  OAI21_X1   g20160(.A1(new_n16372_), .A2(new_n23229_), .B(new_n23318_), .ZN(new_n23319_));
  NAND3_X1   g20161(.A1(new_n23319_), .A2(new_n18929_), .A3(new_n23244_), .ZN(new_n23320_));
  NAND2_X1   g20162(.A1(new_n23320_), .A2(new_n16569_), .ZN(new_n23321_));
  XOR2_X1    g20163(.A1(new_n23321_), .A2(new_n16572_), .Z(new_n23322_));
  AOI21_X1   g20164(.A1(new_n19022_), .A2(new_n23320_), .B(new_n23322_), .ZN(new_n23323_));
  INV_X1     g20165(.I(new_n23229_), .ZN(new_n23324_));
  NAND2_X1   g20166(.A1(new_n23267_), .A2(new_n13963_), .ZN(new_n23325_));
  XNOR2_X1   g20167(.A1(new_n23325_), .A2(new_n19028_), .ZN(new_n23326_));
  NOR3_X1    g20168(.A1(new_n23326_), .A2(new_n16424_), .A3(new_n23324_), .ZN(new_n23327_));
  OAI21_X1   g20169(.A1(new_n23323_), .A2(new_n16574_), .B(new_n23327_), .ZN(new_n23328_));
  NOR4_X1    g20170(.A1(new_n23243_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n23329_));
  NOR2_X1    g20171(.A1(new_n23329_), .A2(new_n14005_), .ZN(new_n23330_));
  XOR2_X1    g20172(.A1(new_n23330_), .A2(new_n14007_), .Z(new_n23331_));
  NAND2_X1   g20173(.A1(new_n23331_), .A2(new_n23229_), .ZN(new_n23332_));
  NOR2_X1    g20174(.A1(new_n23324_), .A2(pi0647), .ZN(new_n23333_));
  AOI21_X1   g20175(.A1(new_n23329_), .A2(pi0647), .B(new_n23333_), .ZN(new_n23334_));
  NOR2_X1    g20176(.A1(new_n23319_), .A2(new_n13994_), .ZN(new_n23335_));
  XNOR2_X1   g20177(.A1(new_n23335_), .A2(new_n19033_), .ZN(new_n23336_));
  AOI22_X1   g20178(.A1(new_n23336_), .A2(new_n23229_), .B1(new_n14206_), .B2(new_n23334_), .ZN(new_n23337_));
  NOR3_X1    g20179(.A1(new_n23337_), .A2(new_n14010_), .A3(new_n23332_), .ZN(new_n23338_));
  OAI22_X1   g20180(.A1(new_n23317_), .A2(new_n23328_), .B1(new_n12776_), .B2(new_n23338_), .ZN(new_n23339_));
  AOI21_X1   g20181(.A1(new_n23334_), .A2(pi1157), .B(new_n12776_), .ZN(new_n23340_));
  AOI22_X1   g20182(.A1(new_n23332_), .A2(new_n23340_), .B1(new_n12776_), .B2(new_n23329_), .ZN(new_n23341_));
  NAND2_X1   g20183(.A1(new_n23339_), .A2(pi0644), .ZN(new_n23342_));
  XOR2_X1    g20184(.A1(new_n23342_), .A2(new_n14205_), .Z(new_n23343_));
  NOR2_X1    g20185(.A1(new_n23343_), .A2(new_n23341_), .ZN(new_n23344_));
  NOR2_X1    g20186(.A1(new_n23319_), .A2(new_n18968_), .ZN(new_n23345_));
  NAND2_X1   g20187(.A1(new_n18967_), .A2(new_n23229_), .ZN(new_n23346_));
  XOR2_X1    g20188(.A1(new_n23345_), .A2(new_n23346_), .Z(new_n23347_));
  NAND2_X1   g20189(.A1(new_n23347_), .A2(pi0715), .ZN(new_n23348_));
  XOR2_X1    g20190(.A1(new_n23348_), .A2(new_n14205_), .Z(new_n23349_));
  OAI21_X1   g20191(.A1(new_n23349_), .A2(new_n23324_), .B(new_n14203_), .ZN(new_n23350_));
  NAND2_X1   g20192(.A1(new_n23347_), .A2(pi0644), .ZN(new_n23351_));
  XOR2_X1    g20193(.A1(new_n23351_), .A2(new_n14217_), .Z(new_n23352_));
  AOI21_X1   g20194(.A1(new_n23352_), .A2(new_n23229_), .B(pi1160), .ZN(new_n23353_));
  OAI21_X1   g20195(.A1(new_n23344_), .A2(new_n23350_), .B(new_n23353_), .ZN(new_n23354_));
  NAND2_X1   g20196(.A1(new_n23339_), .A2(pi0715), .ZN(new_n23355_));
  XOR2_X1    g20197(.A1(new_n23355_), .A2(new_n14205_), .Z(new_n23356_));
  NOR2_X1    g20198(.A1(new_n23356_), .A2(new_n23341_), .ZN(new_n23357_));
  AOI21_X1   g20199(.A1(new_n23354_), .A2(new_n23357_), .B(new_n14799_), .ZN(new_n23358_));
  XOR2_X1    g20200(.A1(new_n23358_), .A2(new_n14801_), .Z(new_n23359_));
  NOR2_X1    g20201(.A1(new_n7240_), .A2(pi0186), .ZN(new_n23360_));
  NOR4_X1    g20202(.A1(new_n23359_), .A2(pi0832), .A3(new_n23339_), .A4(new_n23360_), .ZN(new_n23361_));
  AOI21_X1   g20203(.A1(new_n23228_), .A2(new_n7240_), .B(new_n23361_), .ZN(new_n23362_));
  NOR3_X1    g20204(.A1(new_n23227_), .A2(new_n23217_), .A3(new_n14200_), .ZN(new_n23363_));
  NOR2_X1    g20205(.A1(new_n23363_), .A2(new_n14217_), .ZN(new_n23364_));
  NOR4_X1    g20206(.A1(new_n23227_), .A2(new_n23217_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n23365_));
  NOR2_X1    g20207(.A1(new_n23364_), .A2(new_n23365_), .ZN(new_n23366_));
  NAND2_X1   g20208(.A1(new_n23223_), .A2(new_n23219_), .ZN(new_n23367_));
  INV_X1     g20209(.I(new_n23204_), .ZN(new_n23368_));
  AOI21_X1   g20210(.A1(new_n23368_), .A2(new_n23202_), .B(new_n23015_), .ZN(new_n23369_));
  INV_X1     g20211(.I(new_n23209_), .ZN(new_n23370_));
  OAI21_X1   g20212(.A1(new_n23370_), .A2(new_n23369_), .B(new_n14005_), .ZN(new_n23371_));
  INV_X1     g20213(.I(new_n23216_), .ZN(new_n23372_));
  NAND4_X1   g20214(.A1(new_n23367_), .A2(pi0787), .A3(new_n23371_), .A4(new_n23372_), .ZN(new_n23373_));
  OAI21_X1   g20215(.A1(new_n23192_), .A2(new_n23169_), .B(new_n23371_), .ZN(new_n23374_));
  INV_X1     g20216(.I(new_n23195_), .ZN(new_n23375_));
  NAND2_X1   g20217(.A1(new_n23197_), .A2(pi0792), .ZN(new_n23376_));
  AOI21_X1   g20218(.A1(new_n23165_), .A2(new_n23198_), .B(new_n23376_), .ZN(new_n23377_));
  NOR2_X1    g20219(.A1(new_n23377_), .A2(new_n23375_), .ZN(new_n23378_));
  AOI21_X1   g20220(.A1(new_n23378_), .A2(pi1157), .B(new_n14008_), .ZN(new_n23379_));
  INV_X1     g20221(.I(new_n23212_), .ZN(new_n23380_));
  OAI21_X1   g20222(.A1(new_n23379_), .A2(new_n23380_), .B(new_n22991_), .ZN(new_n23381_));
  NOR2_X1    g20223(.A1(new_n23214_), .A2(new_n16329_), .ZN(new_n23382_));
  NAND2_X1   g20224(.A1(new_n23382_), .A2(new_n23381_), .ZN(new_n23383_));
  AOI21_X1   g20225(.A1(new_n23383_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n23384_));
  OAI21_X1   g20226(.A1(new_n23192_), .A2(new_n23169_), .B(new_n23384_), .ZN(new_n23385_));
  NAND3_X1   g20227(.A1(new_n23385_), .A2(new_n23374_), .A3(pi0787), .ZN(new_n23386_));
  NAND2_X1   g20228(.A1(new_n23205_), .A2(pi0787), .ZN(new_n23387_));
  NOR3_X1    g20229(.A1(new_n23381_), .A2(new_n12776_), .A3(new_n23378_), .ZN(new_n23388_));
  XOR2_X1    g20230(.A1(new_n23387_), .A2(new_n23388_), .Z(new_n23389_));
  NOR2_X1    g20231(.A1(new_n23015_), .A2(new_n14211_), .ZN(new_n23390_));
  AOI21_X1   g20232(.A1(new_n23208_), .A2(new_n14211_), .B(new_n23390_), .ZN(new_n23391_));
  OAI21_X1   g20233(.A1(new_n23015_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n23392_));
  NAND2_X1   g20234(.A1(new_n23391_), .A2(new_n23392_), .ZN(new_n23393_));
  NAND4_X1   g20235(.A1(new_n23389_), .A2(pi0644), .A3(new_n14200_), .A4(new_n23393_), .ZN(new_n23394_));
  AOI22_X1   g20236(.A1(new_n23394_), .A2(new_n14204_), .B1(new_n23386_), .B2(new_n23373_), .ZN(new_n23395_));
  AOI21_X1   g20237(.A1(new_n23015_), .A2(new_n14254_), .B(pi0644), .ZN(new_n23396_));
  NOR3_X1    g20238(.A1(new_n23389_), .A2(new_n23391_), .A3(new_n23396_), .ZN(new_n23397_));
  OAI21_X1   g20239(.A1(new_n23395_), .A2(pi0790), .B(new_n23397_), .ZN(new_n23398_));
  NOR3_X1    g20240(.A1(new_n23366_), .A2(new_n23398_), .A3(new_n23362_), .ZN(po0343));
  NOR3_X1    g20241(.A1(new_n13632_), .A2(new_n3259_), .A3(new_n17019_), .ZN(new_n23400_));
  NOR3_X1    g20242(.A1(new_n13097_), .A2(pi0038), .A3(new_n17019_), .ZN(new_n23401_));
  OAI21_X1   g20243(.A1(new_n23400_), .A2(new_n23401_), .B(new_n13624_), .ZN(new_n23402_));
  NAND2_X1   g20244(.A1(new_n19637_), .A2(pi0187), .ZN(new_n23404_));
  NAND2_X1   g20245(.A1(new_n19329_), .A2(new_n17019_), .ZN(new_n23405_));
  AOI21_X1   g20246(.A1(new_n23402_), .A2(new_n23404_), .B(new_n23405_), .ZN(new_n23406_));
  NAND2_X1   g20247(.A1(new_n16962_), .A2(pi0187), .ZN(new_n23407_));
  OAI21_X1   g20248(.A1(new_n23406_), .A2(new_n23407_), .B(new_n3289_), .ZN(new_n23408_));
  NOR2_X1    g20249(.A1(new_n23406_), .A2(new_n3290_), .ZN(new_n23409_));
  AOI21_X1   g20250(.A1(new_n9528_), .A2(new_n3290_), .B(new_n23409_), .ZN(new_n23410_));
  OAI21_X1   g20251(.A1(new_n13721_), .A2(new_n16962_), .B(new_n9528_), .ZN(new_n23411_));
  NAND2_X1   g20252(.A1(new_n23411_), .A2(new_n13108_), .ZN(new_n23412_));
  NAND2_X1   g20253(.A1(new_n9528_), .A2(new_n16962_), .ZN(new_n23413_));
  NAND4_X1   g20254(.A1(new_n13634_), .A2(pi0187), .A3(new_n3290_), .A4(new_n23413_), .ZN(new_n23414_));
  NOR3_X1    g20255(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n9528_), .ZN(new_n23415_));
  NOR3_X1    g20256(.A1(new_n14422_), .A2(pi0038), .A3(new_n9528_), .ZN(new_n23416_));
  OAI21_X1   g20257(.A1(new_n23415_), .A2(new_n23416_), .B(new_n15655_), .ZN(new_n23417_));
  AOI21_X1   g20258(.A1(new_n23412_), .A2(new_n23414_), .B(new_n23417_), .ZN(new_n23418_));
  NOR3_X1    g20259(.A1(new_n14431_), .A2(new_n9528_), .A3(new_n14081_), .ZN(new_n23419_));
  NOR2_X1    g20260(.A1(new_n23418_), .A2(new_n23419_), .ZN(new_n23420_));
  NOR2_X1    g20261(.A1(new_n23420_), .A2(new_n13620_), .ZN(new_n23421_));
  AOI21_X1   g20262(.A1(new_n23421_), .A2(new_n23410_), .B(pi0625), .ZN(new_n23422_));
  OAI21_X1   g20263(.A1(new_n23422_), .A2(new_n23408_), .B(pi0778), .ZN(new_n23423_));
  NOR3_X1    g20264(.A1(new_n23408_), .A2(new_n13613_), .A3(new_n13748_), .ZN(new_n23427_));
  XOR2_X1    g20265(.A1(new_n23423_), .A2(new_n23427_), .Z(new_n23428_));
  NAND2_X1   g20266(.A1(new_n23410_), .A2(new_n13776_), .ZN(new_n23429_));
  NOR2_X1    g20267(.A1(new_n14428_), .A2(pi0187), .ZN(new_n23430_));
  INV_X1     g20268(.I(new_n23430_), .ZN(new_n23431_));
  NAND2_X1   g20269(.A1(new_n23431_), .A2(new_n13780_), .ZN(new_n23432_));
  AOI21_X1   g20270(.A1(new_n23429_), .A2(new_n23432_), .B(new_n13766_), .ZN(new_n23433_));
  INV_X1     g20271(.I(new_n23433_), .ZN(new_n23434_));
  NAND2_X1   g20272(.A1(new_n23418_), .A2(new_n13748_), .ZN(new_n23435_));
  NOR2_X1    g20273(.A1(new_n23418_), .A2(new_n14452_), .ZN(new_n23436_));
  NOR2_X1    g20274(.A1(new_n23431_), .A2(new_n14452_), .ZN(new_n23437_));
  XNOR2_X1   g20275(.A1(new_n23436_), .A2(new_n23437_), .ZN(new_n23438_));
  OAI21_X1   g20276(.A1(new_n23438_), .A2(new_n13748_), .B(new_n23435_), .ZN(new_n23439_));
  AOI21_X1   g20277(.A1(new_n23439_), .A2(new_n13766_), .B(new_n13785_), .ZN(new_n23440_));
  AOI21_X1   g20278(.A1(new_n23440_), .A2(new_n23434_), .B(pi0609), .ZN(new_n23441_));
  OAI21_X1   g20279(.A1(new_n23441_), .A2(new_n23428_), .B(pi0785), .ZN(new_n23442_));
  NAND2_X1   g20280(.A1(new_n23439_), .A2(pi0609), .ZN(new_n23443_));
  AOI21_X1   g20281(.A1(new_n23431_), .A2(new_n14467_), .B(pi0609), .ZN(new_n23444_));
  NOR2_X1    g20282(.A1(new_n23429_), .A2(new_n23444_), .ZN(new_n23445_));
  NOR2_X1    g20283(.A1(new_n23445_), .A2(new_n14465_), .ZN(new_n23446_));
  AOI21_X1   g20284(.A1(new_n23443_), .A2(new_n23446_), .B(pi0609), .ZN(new_n23447_));
  NOR3_X1    g20285(.A1(new_n23447_), .A2(new_n23428_), .A3(new_n13801_), .ZN(new_n23448_));
  XOR2_X1    g20286(.A1(new_n23442_), .A2(new_n23448_), .Z(new_n23449_));
  NAND2_X1   g20287(.A1(new_n23430_), .A2(new_n13775_), .ZN(new_n23450_));
  OAI21_X1   g20288(.A1(new_n23410_), .A2(new_n13775_), .B(new_n23450_), .ZN(new_n23451_));
  NAND4_X1   g20289(.A1(new_n23433_), .A2(new_n23445_), .A3(pi0785), .A4(new_n23451_), .ZN(new_n23452_));
  NAND3_X1   g20290(.A1(new_n23445_), .A2(pi0785), .A3(new_n23451_), .ZN(new_n23453_));
  NAND3_X1   g20291(.A1(new_n23453_), .A2(new_n23434_), .A3(pi0785), .ZN(new_n23454_));
  NAND2_X1   g20292(.A1(new_n23454_), .A2(new_n23452_), .ZN(new_n23455_));
  NOR2_X1    g20293(.A1(new_n23455_), .A2(new_n13816_), .ZN(new_n23456_));
  NOR2_X1    g20294(.A1(new_n23456_), .A2(new_n13819_), .ZN(new_n23457_));
  NOR3_X1    g20295(.A1(new_n23455_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n23458_));
  OAI21_X1   g20296(.A1(new_n23457_), .A2(new_n23458_), .B(new_n23430_), .ZN(new_n23459_));
  NOR2_X1    g20297(.A1(new_n23431_), .A2(new_n13805_), .ZN(new_n23460_));
  AOI21_X1   g20298(.A1(new_n23439_), .A2(new_n13805_), .B(new_n23460_), .ZN(new_n23461_));
  INV_X1     g20299(.I(new_n23461_), .ZN(new_n23462_));
  AOI21_X1   g20300(.A1(new_n23462_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n23463_));
  AOI21_X1   g20301(.A1(new_n23459_), .A2(new_n23463_), .B(pi0618), .ZN(new_n23464_));
  OR2_X2     g20302(.A1(new_n23464_), .A2(new_n23449_), .Z(new_n23465_));
  NAND3_X1   g20303(.A1(new_n23455_), .A2(pi0618), .A3(pi1154), .ZN(new_n23466_));
  NAND4_X1   g20304(.A1(new_n23454_), .A2(new_n13816_), .A3(pi1154), .A4(new_n23452_), .ZN(new_n23467_));
  AOI21_X1   g20305(.A1(new_n23466_), .A2(new_n23467_), .B(new_n23431_), .ZN(new_n23468_));
  INV_X1     g20306(.I(new_n23468_), .ZN(new_n23469_));
  AOI21_X1   g20307(.A1(new_n23462_), .A2(pi0618), .B(new_n13837_), .ZN(new_n23470_));
  AOI21_X1   g20308(.A1(new_n23469_), .A2(new_n23470_), .B(pi0618), .ZN(new_n23471_));
  OR3_X2     g20309(.A1(new_n23471_), .A2(new_n13855_), .A3(new_n23449_), .Z(new_n23472_));
  AOI21_X1   g20310(.A1(pi0781), .A2(new_n23465_), .B(new_n23472_), .ZN(new_n23473_));
  AND3_X2    g20311(.A1(new_n23472_), .A2(new_n23465_), .A3(pi0781), .Z(new_n23474_));
  NOR2_X1    g20312(.A1(new_n23474_), .A2(new_n23473_), .ZN(new_n23475_));
  INV_X1     g20313(.I(new_n23475_), .ZN(new_n23476_));
  NAND2_X1   g20314(.A1(new_n23459_), .A2(pi0781), .ZN(new_n23477_));
  NAND3_X1   g20315(.A1(new_n23468_), .A2(pi0781), .A3(new_n23455_), .ZN(new_n23478_));
  INV_X1     g20316(.I(new_n23478_), .ZN(new_n23479_));
  NAND2_X1   g20317(.A1(new_n23479_), .A2(new_n23477_), .ZN(new_n23480_));
  NAND3_X1   g20318(.A1(new_n23478_), .A2(new_n23459_), .A3(pi0781), .ZN(new_n23481_));
  NAND2_X1   g20319(.A1(new_n23480_), .A2(new_n23481_), .ZN(new_n23482_));
  NAND3_X1   g20320(.A1(new_n23482_), .A2(pi0619), .A3(pi1159), .ZN(new_n23483_));
  NAND4_X1   g20321(.A1(new_n23480_), .A2(pi0619), .A3(new_n13868_), .A4(new_n23481_), .ZN(new_n23484_));
  AOI21_X1   g20322(.A1(new_n23483_), .A2(new_n23484_), .B(new_n23431_), .ZN(new_n23485_));
  NOR2_X1    g20323(.A1(new_n23430_), .A2(new_n13880_), .ZN(new_n23486_));
  AOI21_X1   g20324(.A1(new_n23461_), .A2(new_n13880_), .B(new_n23486_), .ZN(new_n23487_));
  AOI21_X1   g20325(.A1(new_n23487_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n23488_));
  INV_X1     g20326(.I(new_n23488_), .ZN(new_n23489_));
  OAI21_X1   g20327(.A1(new_n23485_), .A2(new_n23489_), .B(new_n13860_), .ZN(new_n23490_));
  NAND3_X1   g20328(.A1(new_n23482_), .A2(pi0619), .A3(pi1159), .ZN(new_n23491_));
  NAND4_X1   g20329(.A1(new_n23480_), .A2(new_n13860_), .A3(pi1159), .A4(new_n23481_), .ZN(new_n23492_));
  AOI21_X1   g20330(.A1(new_n23491_), .A2(new_n23492_), .B(new_n23431_), .ZN(new_n23493_));
  AOI21_X1   g20331(.A1(new_n23487_), .A2(pi0619), .B(new_n15217_), .ZN(new_n23494_));
  INV_X1     g20332(.I(new_n23494_), .ZN(new_n23495_));
  OAI21_X1   g20333(.A1(new_n23493_), .A2(new_n23495_), .B(new_n13860_), .ZN(new_n23496_));
  NAND4_X1   g20334(.A1(new_n23476_), .A2(new_n23490_), .A3(new_n23496_), .A4(pi0789), .ZN(new_n23497_));
  AOI21_X1   g20335(.A1(new_n23476_), .A2(new_n23490_), .B(new_n13896_), .ZN(new_n23498_));
  NAND3_X1   g20336(.A1(new_n23476_), .A2(new_n23496_), .A3(pi0789), .ZN(new_n23499_));
  NAND2_X1   g20337(.A1(new_n23498_), .A2(new_n23499_), .ZN(new_n23500_));
  NAND2_X1   g20338(.A1(new_n23500_), .A2(new_n23497_), .ZN(new_n23501_));
  NAND4_X1   g20339(.A1(new_n23485_), .A2(new_n23493_), .A3(pi0789), .A4(new_n23482_), .ZN(new_n23502_));
  NAND2_X1   g20340(.A1(new_n23483_), .A2(new_n23484_), .ZN(new_n23503_));
  NAND2_X1   g20341(.A1(new_n23503_), .A2(new_n23430_), .ZN(new_n23504_));
  NAND3_X1   g20342(.A1(new_n23493_), .A2(pi0789), .A3(new_n23482_), .ZN(new_n23505_));
  NAND3_X1   g20343(.A1(new_n23505_), .A2(new_n23504_), .A3(pi0789), .ZN(new_n23506_));
  NOR2_X1    g20344(.A1(new_n23431_), .A2(new_n13919_), .ZN(new_n23507_));
  AOI21_X1   g20345(.A1(new_n23487_), .A2(new_n13919_), .B(new_n23507_), .ZN(new_n23508_));
  NOR2_X1    g20346(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n23509_));
  INV_X1     g20347(.I(new_n23509_), .ZN(new_n23510_));
  AOI21_X1   g20348(.A1(new_n23506_), .A2(new_n23502_), .B(new_n23510_), .ZN(new_n23511_));
  INV_X1     g20349(.I(new_n23502_), .ZN(new_n23512_));
  NOR2_X1    g20350(.A1(new_n23485_), .A2(new_n13896_), .ZN(new_n23513_));
  AND2_X2    g20351(.A1(new_n23505_), .A2(new_n23513_), .Z(new_n23514_));
  NOR2_X1    g20352(.A1(new_n23514_), .A2(new_n23512_), .ZN(new_n23515_));
  NAND3_X1   g20353(.A1(new_n23501_), .A2(pi0626), .A3(pi0788), .ZN(new_n23520_));
  INV_X1     g20354(.I(new_n23520_), .ZN(new_n23521_));
  OAI21_X1   g20355(.A1(new_n23514_), .A2(new_n23512_), .B(new_n23509_), .ZN(new_n23522_));
  AOI22_X1   g20356(.A1(new_n23522_), .A2(new_n13901_), .B1(new_n23497_), .B2(new_n23500_), .ZN(new_n23523_));
  AOI21_X1   g20357(.A1(new_n23500_), .A2(new_n23497_), .B(new_n15258_), .ZN(new_n23524_));
  NOR3_X1    g20358(.A1(new_n23523_), .A2(new_n13937_), .A3(new_n23524_), .ZN(new_n23525_));
  NOR2_X1    g20359(.A1(new_n23525_), .A2(new_n23521_), .ZN(new_n23526_));
  NOR2_X1    g20360(.A1(new_n23430_), .A2(new_n16372_), .ZN(new_n23527_));
  AOI21_X1   g20361(.A1(new_n23515_), .A2(new_n16372_), .B(new_n23527_), .ZN(new_n23528_));
  NOR2_X1    g20362(.A1(new_n23430_), .A2(new_n13966_), .ZN(new_n23529_));
  AOI21_X1   g20363(.A1(new_n23508_), .A2(new_n13966_), .B(new_n23529_), .ZN(new_n23530_));
  NAND2_X1   g20364(.A1(new_n23530_), .A2(pi0628), .ZN(new_n23531_));
  NAND2_X1   g20365(.A1(new_n23531_), .A2(new_n13970_), .ZN(new_n23532_));
  NAND3_X1   g20366(.A1(new_n23530_), .A2(pi0628), .A3(new_n13971_), .ZN(new_n23533_));
  AOI21_X1   g20367(.A1(new_n23532_), .A2(new_n23533_), .B(new_n23431_), .ZN(new_n23534_));
  NOR2_X1    g20368(.A1(new_n23534_), .A2(new_n15270_), .ZN(new_n23535_));
  INV_X1     g20369(.I(new_n23535_), .ZN(new_n23536_));
  NAND2_X1   g20370(.A1(new_n23530_), .A2(pi1156), .ZN(new_n23538_));
  XOR2_X1    g20371(.A1(new_n23538_), .A2(new_n13971_), .Z(new_n23539_));
  NAND2_X1   g20372(.A1(new_n23539_), .A2(new_n23430_), .ZN(new_n23540_));
  NOR3_X1    g20373(.A1(new_n23526_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n23543_));
  INV_X1     g20374(.I(new_n23497_), .ZN(new_n23544_));
  AOI21_X1   g20375(.A1(new_n23504_), .A2(new_n23488_), .B(pi0619), .ZN(new_n23545_));
  OAI21_X1   g20376(.A1(new_n23545_), .A2(new_n23475_), .B(pi0789), .ZN(new_n23546_));
  OR2_X2     g20377(.A1(new_n23493_), .A2(new_n23495_), .Z(new_n23547_));
  OAI21_X1   g20378(.A1(new_n23474_), .A2(new_n23473_), .B(pi0789), .ZN(new_n23548_));
  AOI21_X1   g20379(.A1(new_n23547_), .A2(new_n13860_), .B(new_n23548_), .ZN(new_n23549_));
  NOR2_X1    g20380(.A1(new_n23546_), .A2(new_n23549_), .ZN(new_n23550_));
  OAI22_X1   g20381(.A1(new_n23550_), .A2(new_n23544_), .B1(pi0626), .B2(new_n23511_), .ZN(new_n23551_));
  OAI21_X1   g20382(.A1(new_n23550_), .A2(new_n23544_), .B(new_n14577_), .ZN(new_n23552_));
  NAND3_X1   g20383(.A1(new_n23551_), .A2(new_n23552_), .A3(pi0788), .ZN(new_n23553_));
  NAND3_X1   g20384(.A1(new_n23506_), .A2(new_n16372_), .A3(new_n23502_), .ZN(new_n23554_));
  OAI21_X1   g20385(.A1(new_n16372_), .A2(new_n23430_), .B(new_n23554_), .ZN(new_n23555_));
  AOI21_X1   g20386(.A1(new_n23555_), .A2(new_n23535_), .B(pi0628), .ZN(new_n23556_));
  AOI21_X1   g20387(.A1(new_n23553_), .A2(new_n23520_), .B(new_n23556_), .ZN(new_n23557_));
  AOI21_X1   g20388(.A1(new_n23553_), .A2(new_n23520_), .B(new_n15296_), .ZN(new_n23558_));
  NOR3_X1    g20389(.A1(new_n23557_), .A2(new_n23558_), .A3(new_n12777_), .ZN(new_n23559_));
  NOR2_X1    g20390(.A1(new_n23559_), .A2(new_n23543_), .ZN(new_n23560_));
  NOR2_X1    g20391(.A1(new_n23430_), .A2(new_n13994_), .ZN(new_n23561_));
  AOI21_X1   g20392(.A1(new_n23555_), .A2(new_n13994_), .B(new_n23561_), .ZN(new_n23562_));
  INV_X1     g20393(.I(new_n23562_), .ZN(new_n23563_));
  NOR2_X1    g20394(.A1(new_n23534_), .A2(new_n12777_), .ZN(new_n23564_));
  NOR4_X1    g20395(.A1(new_n23540_), .A2(new_n12777_), .A3(new_n23564_), .A4(new_n23530_), .ZN(new_n23565_));
  NOR3_X1    g20396(.A1(new_n23540_), .A2(new_n12777_), .A3(new_n23530_), .ZN(new_n23566_));
  NOR3_X1    g20397(.A1(new_n23566_), .A2(new_n12777_), .A3(new_n23534_), .ZN(new_n23567_));
  NOR2_X1    g20398(.A1(new_n23567_), .A2(new_n23565_), .ZN(new_n23568_));
  NAND2_X1   g20399(.A1(new_n23568_), .A2(pi0647), .ZN(new_n23569_));
  XOR2_X1    g20400(.A1(new_n23569_), .A2(new_n14008_), .Z(new_n23570_));
  AOI21_X1   g20401(.A1(new_n23570_), .A2(new_n23430_), .B(new_n14012_), .ZN(new_n23571_));
  AOI21_X1   g20402(.A1(new_n23563_), .A2(new_n23571_), .B(pi0647), .ZN(new_n23572_));
  AOI21_X1   g20403(.A1(new_n23568_), .A2(pi1157), .B(new_n14008_), .ZN(new_n23573_));
  NOR4_X1    g20404(.A1(new_n23567_), .A2(new_n23565_), .A3(pi0647), .A4(new_n14006_), .ZN(new_n23574_));
  OAI21_X1   g20405(.A1(new_n23573_), .A2(new_n23574_), .B(new_n23430_), .ZN(new_n23575_));
  NAND2_X1   g20406(.A1(new_n23575_), .A2(new_n14027_), .ZN(new_n23576_));
  AOI21_X1   g20407(.A1(new_n23562_), .A2(pi0647), .B(new_n23576_), .ZN(new_n23577_));
  NOR2_X1    g20408(.A1(new_n23577_), .A2(pi0647), .ZN(new_n23578_));
  NOR4_X1    g20409(.A1(new_n23560_), .A2(new_n12776_), .A3(new_n23572_), .A4(new_n23578_), .ZN(new_n23579_));
  NAND2_X1   g20410(.A1(new_n23553_), .A2(new_n23520_), .ZN(new_n23580_));
  NAND3_X1   g20411(.A1(new_n23580_), .A2(pi0628), .A3(pi0792), .ZN(new_n23581_));
  OAI21_X1   g20412(.A1(new_n23528_), .A2(new_n23536_), .B(new_n13942_), .ZN(new_n23582_));
  OAI21_X1   g20413(.A1(new_n23525_), .A2(new_n23521_), .B(new_n23582_), .ZN(new_n23583_));
  OAI21_X1   g20414(.A1(new_n23525_), .A2(new_n23521_), .B(new_n14606_), .ZN(new_n23584_));
  NAND3_X1   g20415(.A1(new_n23583_), .A2(new_n23584_), .A3(pi0792), .ZN(new_n23585_));
  AOI21_X1   g20416(.A1(new_n23585_), .A2(new_n23581_), .B(new_n23572_), .ZN(new_n23586_));
  OAI21_X1   g20417(.A1(new_n23577_), .A2(pi0647), .B(pi0787), .ZN(new_n23587_));
  AOI21_X1   g20418(.A1(new_n23585_), .A2(new_n23581_), .B(new_n23587_), .ZN(new_n23588_));
  NOR3_X1    g20419(.A1(new_n23586_), .A2(new_n23588_), .A3(new_n12776_), .ZN(new_n23589_));
  OAI21_X1   g20420(.A1(new_n23589_), .A2(new_n23579_), .B(new_n12775_), .ZN(new_n23590_));
  NOR2_X1    g20421(.A1(new_n9992_), .A2(pi0187), .ZN(new_n23591_));
  NOR2_X1    g20422(.A1(new_n14652_), .A2(new_n16962_), .ZN(new_n23592_));
  AOI21_X1   g20423(.A1(new_n13218_), .A2(pi0726), .B(new_n23591_), .ZN(new_n23593_));
  INV_X1     g20424(.I(new_n23593_), .ZN(new_n23594_));
  NAND3_X1   g20425(.A1(new_n23594_), .A2(new_n23592_), .A3(new_n23591_), .ZN(new_n23595_));
  NOR3_X1    g20426(.A1(new_n23592_), .A2(new_n13614_), .A3(new_n23593_), .ZN(new_n23596_));
  XNOR2_X1   g20427(.A1(new_n23595_), .A2(new_n23596_), .ZN(new_n23597_));
  NAND2_X1   g20428(.A1(new_n23597_), .A2(pi0778), .ZN(new_n23598_));
  NAND2_X1   g20429(.A1(new_n23594_), .A2(new_n13748_), .ZN(new_n23599_));
  NAND2_X1   g20430(.A1(new_n23598_), .A2(new_n23599_), .ZN(new_n23600_));
  INV_X1     g20431(.I(new_n23600_), .ZN(new_n23601_));
  NOR2_X1    g20432(.A1(new_n23601_), .A2(new_n14048_), .ZN(new_n23602_));
  INV_X1     g20433(.I(new_n23602_), .ZN(new_n23603_));
  NOR2_X1    g20434(.A1(new_n23603_), .A2(new_n14051_), .ZN(new_n23604_));
  INV_X1     g20435(.I(new_n23604_), .ZN(new_n23605_));
  NOR2_X1    g20436(.A1(new_n23605_), .A2(new_n14163_), .ZN(new_n23606_));
  AOI21_X1   g20437(.A1(new_n13104_), .A2(new_n17019_), .B(new_n23591_), .ZN(new_n23607_));
  NOR2_X1    g20438(.A1(new_n14096_), .A2(new_n23607_), .ZN(new_n23608_));
  AOI21_X1   g20439(.A1(new_n23608_), .A2(new_n14094_), .B(pi1155), .ZN(new_n23609_));
  NOR2_X1    g20440(.A1(new_n23609_), .A2(new_n13801_), .ZN(new_n23610_));
  AOI21_X1   g20441(.A1(new_n23607_), .A2(pi1155), .B(new_n9992_), .ZN(new_n23611_));
  NOR2_X1    g20442(.A1(new_n23611_), .A2(new_n14102_), .ZN(new_n23612_));
  NAND3_X1   g20443(.A1(new_n23612_), .A2(new_n23608_), .A3(pi0785), .ZN(new_n23613_));
  XOR2_X1    g20444(.A1(new_n23610_), .A2(new_n23613_), .Z(new_n23614_));
  NOR2_X1    g20445(.A1(new_n23614_), .A2(new_n13817_), .ZN(new_n23615_));
  OAI21_X1   g20446(.A1(new_n23615_), .A2(pi0618), .B(new_n9992_), .ZN(new_n23616_));
  NAND2_X1   g20447(.A1(new_n23616_), .A2(pi0781), .ZN(new_n23617_));
  OAI21_X1   g20448(.A1(new_n23615_), .A2(new_n9992_), .B(pi0618), .ZN(new_n23618_));
  NOR3_X1    g20449(.A1(new_n23618_), .A2(new_n13855_), .A3(new_n23614_), .ZN(new_n23619_));
  XOR2_X1    g20450(.A1(new_n23619_), .A2(new_n23617_), .Z(new_n23620_));
  NAND2_X1   g20451(.A1(new_n23620_), .A2(pi0619), .ZN(new_n23621_));
  XOR2_X1    g20452(.A1(new_n23621_), .A2(new_n13904_), .Z(new_n23622_));
  NAND2_X1   g20453(.A1(new_n23622_), .A2(new_n23591_), .ZN(new_n23623_));
  NAND2_X1   g20454(.A1(new_n23623_), .A2(pi0789), .ZN(new_n23624_));
  NAND2_X1   g20455(.A1(new_n23620_), .A2(pi1159), .ZN(new_n23625_));
  XOR2_X1    g20456(.A1(new_n23625_), .A2(new_n13904_), .Z(new_n23626_));
  NAND2_X1   g20457(.A1(new_n23626_), .A2(new_n23591_), .ZN(new_n23627_));
  NOR3_X1    g20458(.A1(new_n23627_), .A2(new_n13896_), .A3(new_n23620_), .ZN(new_n23628_));
  XOR2_X1    g20459(.A1(new_n23628_), .A2(new_n23624_), .Z(new_n23629_));
  NAND2_X1   g20460(.A1(new_n23629_), .A2(new_n13962_), .ZN(new_n23630_));
  XOR2_X1    g20461(.A1(new_n23630_), .A2(new_n18976_), .Z(new_n23631_));
  AOI22_X1   g20462(.A1(new_n23631_), .A2(new_n23591_), .B1(new_n16639_), .B2(new_n23606_), .ZN(new_n23632_));
  NOR2_X1    g20463(.A1(new_n23593_), .A2(new_n13203_), .ZN(new_n23633_));
  INV_X1     g20464(.I(new_n23633_), .ZN(new_n23634_));
  NOR2_X1    g20465(.A1(new_n23634_), .A2(new_n13613_), .ZN(new_n23635_));
  NOR2_X1    g20466(.A1(new_n23591_), .A2(pi1153), .ZN(new_n23636_));
  INV_X1     g20467(.I(new_n23636_), .ZN(new_n23637_));
  OAI21_X1   g20468(.A1(new_n23592_), .A2(new_n23637_), .B(pi0608), .ZN(new_n23638_));
  NOR2_X1    g20469(.A1(new_n23607_), .A2(pi1153), .ZN(new_n23639_));
  NAND2_X1   g20470(.A1(new_n23638_), .A2(new_n23639_), .ZN(new_n23640_));
  AOI21_X1   g20471(.A1(new_n23640_), .A2(new_n23635_), .B(new_n13748_), .ZN(new_n23641_));
  NOR2_X1    g20472(.A1(new_n23593_), .A2(new_n14082_), .ZN(new_n23642_));
  NAND2_X1   g20473(.A1(new_n23592_), .A2(new_n23636_), .ZN(new_n23643_));
  OAI22_X1   g20474(.A1(new_n23634_), .A2(new_n13613_), .B1(new_n23643_), .B2(new_n23642_), .ZN(new_n23644_));
  NAND4_X1   g20475(.A1(new_n23644_), .A2(pi0778), .A3(new_n23607_), .A4(new_n23634_), .ZN(new_n23645_));
  XNOR2_X1   g20476(.A1(new_n23645_), .A2(new_n23641_), .ZN(new_n23646_));
  NAND2_X1   g20477(.A1(new_n23646_), .A2(new_n13801_), .ZN(new_n23647_));
  NOR2_X1    g20478(.A1(new_n23646_), .A2(new_n13778_), .ZN(new_n23648_));
  XOR2_X1    g20479(.A1(new_n23648_), .A2(new_n14694_), .Z(new_n23649_));
  NOR2_X1    g20480(.A1(new_n23649_), .A2(new_n23601_), .ZN(new_n23650_));
  NOR3_X1    g20481(.A1(new_n23650_), .A2(new_n13783_), .A3(new_n23609_), .ZN(new_n23651_));
  NOR3_X1    g20482(.A1(new_n23651_), .A2(pi0660), .A3(new_n23612_), .ZN(new_n23652_));
  NOR2_X1    g20483(.A1(new_n23646_), .A2(new_n13766_), .ZN(new_n23653_));
  XOR2_X1    g20484(.A1(new_n23653_), .A2(new_n14090_), .Z(new_n23654_));
  NAND3_X1   g20485(.A1(new_n23654_), .A2(pi0785), .A3(new_n23600_), .ZN(new_n23655_));
  OAI21_X1   g20486(.A1(new_n23652_), .A2(new_n23655_), .B(new_n23647_), .ZN(new_n23656_));
  NAND2_X1   g20487(.A1(new_n23656_), .A2(new_n13855_), .ZN(new_n23657_));
  NOR2_X1    g20488(.A1(new_n23656_), .A2(new_n13816_), .ZN(new_n23658_));
  XOR2_X1    g20489(.A1(new_n23658_), .A2(new_n13818_), .Z(new_n23659_));
  NAND2_X1   g20490(.A1(new_n23659_), .A2(new_n23602_), .ZN(new_n23660_));
  NAND3_X1   g20491(.A1(new_n23660_), .A2(new_n13823_), .A3(new_n23618_), .ZN(new_n23661_));
  AND3_X2    g20492(.A1(new_n23661_), .A2(new_n13823_), .A3(new_n23616_), .Z(new_n23662_));
  NOR2_X1    g20493(.A1(new_n23656_), .A2(new_n13817_), .ZN(new_n23663_));
  XOR2_X1    g20494(.A1(new_n23663_), .A2(new_n13819_), .Z(new_n23664_));
  NOR3_X1    g20495(.A1(new_n23664_), .A2(new_n13855_), .A3(new_n23603_), .ZN(new_n23665_));
  INV_X1     g20496(.I(new_n23665_), .ZN(new_n23666_));
  OAI21_X1   g20497(.A1(new_n23662_), .A2(new_n23666_), .B(new_n23657_), .ZN(new_n23667_));
  NOR2_X1    g20498(.A1(new_n23667_), .A2(new_n13860_), .ZN(new_n23668_));
  XOR2_X1    g20499(.A1(new_n23668_), .A2(new_n13904_), .Z(new_n23669_));
  NOR2_X1    g20500(.A1(new_n23669_), .A2(new_n23605_), .ZN(new_n23670_));
  NAND2_X1   g20501(.A1(new_n23627_), .A2(new_n13884_), .ZN(new_n23671_));
  INV_X1     g20502(.I(new_n23667_), .ZN(new_n23672_));
  AOI21_X1   g20503(.A1(new_n23672_), .A2(new_n14143_), .B(pi0789), .ZN(new_n23673_));
  OAI21_X1   g20504(.A1(new_n23670_), .A2(new_n23671_), .B(new_n23673_), .ZN(new_n23674_));
  NOR2_X1    g20505(.A1(new_n23667_), .A2(new_n13868_), .ZN(new_n23675_));
  XOR2_X1    g20506(.A1(new_n23675_), .A2(new_n13903_), .Z(new_n23676_));
  NAND2_X1   g20507(.A1(new_n23623_), .A2(new_n19018_), .ZN(new_n23677_));
  AOI21_X1   g20508(.A1(new_n23676_), .A2(new_n23604_), .B(new_n23677_), .ZN(new_n23678_));
  AOI21_X1   g20509(.A1(new_n23674_), .A2(new_n23678_), .B(new_n23632_), .ZN(new_n23679_));
  NAND2_X1   g20510(.A1(new_n23629_), .A2(new_n16372_), .ZN(new_n23680_));
  OAI21_X1   g20511(.A1(new_n16372_), .A2(new_n23591_), .B(new_n23680_), .ZN(new_n23681_));
  NAND3_X1   g20512(.A1(new_n23681_), .A2(new_n18929_), .A3(new_n23606_), .ZN(new_n23682_));
  NAND2_X1   g20513(.A1(new_n23682_), .A2(new_n16569_), .ZN(new_n23683_));
  XOR2_X1    g20514(.A1(new_n23683_), .A2(new_n16572_), .Z(new_n23684_));
  AOI21_X1   g20515(.A1(new_n19022_), .A2(new_n23682_), .B(new_n23684_), .ZN(new_n23685_));
  INV_X1     g20516(.I(new_n23591_), .ZN(new_n23686_));
  NAND2_X1   g20517(.A1(new_n23629_), .A2(new_n13963_), .ZN(new_n23687_));
  XNOR2_X1   g20518(.A1(new_n23687_), .A2(new_n19028_), .ZN(new_n23688_));
  NOR3_X1    g20519(.A1(new_n23688_), .A2(new_n16424_), .A3(new_n23686_), .ZN(new_n23689_));
  OAI21_X1   g20520(.A1(new_n23685_), .A2(new_n16574_), .B(new_n23689_), .ZN(new_n23690_));
  NOR4_X1    g20521(.A1(new_n23605_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n23691_));
  NOR2_X1    g20522(.A1(new_n23691_), .A2(new_n14005_), .ZN(new_n23692_));
  XOR2_X1    g20523(.A1(new_n23692_), .A2(new_n14007_), .Z(new_n23693_));
  NAND2_X1   g20524(.A1(new_n23693_), .A2(new_n23591_), .ZN(new_n23694_));
  NOR2_X1    g20525(.A1(new_n23686_), .A2(pi0647), .ZN(new_n23695_));
  AOI21_X1   g20526(.A1(new_n23691_), .A2(pi0647), .B(new_n23695_), .ZN(new_n23696_));
  NOR2_X1    g20527(.A1(new_n23681_), .A2(new_n13994_), .ZN(new_n23697_));
  XNOR2_X1   g20528(.A1(new_n23697_), .A2(new_n19033_), .ZN(new_n23698_));
  AOI22_X1   g20529(.A1(new_n23698_), .A2(new_n23591_), .B1(new_n14206_), .B2(new_n23696_), .ZN(new_n23699_));
  NOR3_X1    g20530(.A1(new_n23699_), .A2(new_n14010_), .A3(new_n23694_), .ZN(new_n23700_));
  OAI22_X1   g20531(.A1(new_n23679_), .A2(new_n23690_), .B1(new_n12776_), .B2(new_n23700_), .ZN(new_n23701_));
  AOI21_X1   g20532(.A1(new_n23696_), .A2(pi1157), .B(new_n12776_), .ZN(new_n23702_));
  AOI22_X1   g20533(.A1(new_n23694_), .A2(new_n23702_), .B1(new_n12776_), .B2(new_n23691_), .ZN(new_n23703_));
  NAND2_X1   g20534(.A1(new_n23701_), .A2(pi0644), .ZN(new_n23704_));
  XOR2_X1    g20535(.A1(new_n23704_), .A2(new_n14205_), .Z(new_n23705_));
  NOR2_X1    g20536(.A1(new_n23705_), .A2(new_n23703_), .ZN(new_n23706_));
  NOR2_X1    g20537(.A1(new_n23681_), .A2(new_n18968_), .ZN(new_n23707_));
  NAND2_X1   g20538(.A1(new_n18967_), .A2(new_n23591_), .ZN(new_n23708_));
  XOR2_X1    g20539(.A1(new_n23707_), .A2(new_n23708_), .Z(new_n23709_));
  NAND2_X1   g20540(.A1(new_n23709_), .A2(pi0715), .ZN(new_n23710_));
  XOR2_X1    g20541(.A1(new_n23710_), .A2(new_n14205_), .Z(new_n23711_));
  OAI21_X1   g20542(.A1(new_n23711_), .A2(new_n23686_), .B(new_n14203_), .ZN(new_n23712_));
  NAND2_X1   g20543(.A1(new_n23709_), .A2(pi0644), .ZN(new_n23713_));
  XOR2_X1    g20544(.A1(new_n23713_), .A2(new_n14217_), .Z(new_n23714_));
  AOI21_X1   g20545(.A1(new_n23714_), .A2(new_n23591_), .B(pi1160), .ZN(new_n23715_));
  OAI21_X1   g20546(.A1(new_n23706_), .A2(new_n23712_), .B(new_n23715_), .ZN(new_n23716_));
  NAND2_X1   g20547(.A1(new_n23701_), .A2(pi0715), .ZN(new_n23717_));
  XOR2_X1    g20548(.A1(new_n23717_), .A2(new_n14205_), .Z(new_n23718_));
  NOR2_X1    g20549(.A1(new_n23718_), .A2(new_n23703_), .ZN(new_n23719_));
  AOI21_X1   g20550(.A1(new_n23716_), .A2(new_n23719_), .B(new_n14799_), .ZN(new_n23720_));
  XOR2_X1    g20551(.A1(new_n23720_), .A2(new_n14801_), .Z(new_n23721_));
  NOR2_X1    g20552(.A1(new_n7240_), .A2(pi0187), .ZN(new_n23722_));
  NOR4_X1    g20553(.A1(new_n23721_), .A2(pi0832), .A3(new_n23701_), .A4(new_n23722_), .ZN(new_n23723_));
  AOI21_X1   g20554(.A1(new_n23590_), .A2(new_n7240_), .B(new_n23723_), .ZN(new_n23724_));
  NOR3_X1    g20555(.A1(new_n23589_), .A2(new_n23579_), .A3(new_n14200_), .ZN(new_n23725_));
  NOR2_X1    g20556(.A1(new_n23725_), .A2(new_n14217_), .ZN(new_n23726_));
  NOR4_X1    g20557(.A1(new_n23589_), .A2(new_n23579_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n23727_));
  NOR2_X1    g20558(.A1(new_n23726_), .A2(new_n23727_), .ZN(new_n23728_));
  OAI21_X1   g20559(.A1(new_n12776_), .A2(new_n23586_), .B(new_n23588_), .ZN(new_n23729_));
  INV_X1     g20560(.I(new_n23572_), .ZN(new_n23730_));
  OAI21_X1   g20561(.A1(new_n23543_), .A2(new_n23559_), .B(new_n23730_), .ZN(new_n23731_));
  INV_X1     g20562(.I(new_n23587_), .ZN(new_n23732_));
  OAI21_X1   g20563(.A1(new_n23543_), .A2(new_n23559_), .B(new_n23732_), .ZN(new_n23733_));
  NAND3_X1   g20564(.A1(new_n23733_), .A2(new_n23731_), .A3(pi0787), .ZN(new_n23734_));
  NOR2_X1    g20565(.A1(new_n23431_), .A2(new_n14211_), .ZN(new_n23735_));
  AOI21_X1   g20566(.A1(new_n23562_), .A2(new_n14211_), .B(new_n23735_), .ZN(new_n23736_));
  OAI21_X1   g20567(.A1(new_n23431_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n23737_));
  NAND2_X1   g20568(.A1(new_n23736_), .A2(new_n23737_), .ZN(new_n23738_));
  AOI21_X1   g20569(.A1(new_n23570_), .A2(new_n23430_), .B(new_n12776_), .ZN(new_n23739_));
  NOR3_X1    g20570(.A1(new_n23575_), .A2(new_n12776_), .A3(new_n23568_), .ZN(new_n23740_));
  XNOR2_X1   g20571(.A1(new_n23739_), .A2(new_n23740_), .ZN(new_n23741_));
  AOI21_X1   g20572(.A1(new_n23738_), .A2(new_n14815_), .B(pi0644), .ZN(new_n23742_));
  AOI21_X1   g20573(.A1(new_n23734_), .A2(new_n23729_), .B(new_n23742_), .ZN(new_n23743_));
  AOI21_X1   g20574(.A1(new_n23431_), .A2(new_n14254_), .B(pi0644), .ZN(new_n23744_));
  NOR3_X1    g20575(.A1(new_n23741_), .A2(new_n23736_), .A3(new_n23744_), .ZN(new_n23745_));
  OAI21_X1   g20576(.A1(new_n23743_), .A2(pi0790), .B(new_n23745_), .ZN(new_n23746_));
  NOR3_X1    g20577(.A1(new_n23728_), .A2(new_n23724_), .A3(new_n23746_), .ZN(po0344));
  NAND2_X1   g20578(.A1(new_n19637_), .A2(pi0188), .ZN(new_n23749_));
  NAND2_X1   g20579(.A1(new_n19329_), .A2(new_n17881_), .ZN(new_n23750_));
  AOI21_X1   g20580(.A1(new_n17895_), .A2(new_n23749_), .B(new_n23750_), .ZN(new_n23751_));
  NAND2_X1   g20581(.A1(new_n17880_), .A2(pi0188), .ZN(new_n23752_));
  OAI21_X1   g20582(.A1(new_n23751_), .A2(new_n23752_), .B(new_n3289_), .ZN(new_n23753_));
  NOR2_X1    g20583(.A1(new_n23751_), .A2(new_n3290_), .ZN(new_n23754_));
  AOI21_X1   g20584(.A1(new_n8000_), .A2(new_n3290_), .B(new_n23754_), .ZN(new_n23755_));
  OAI21_X1   g20585(.A1(new_n13721_), .A2(new_n17880_), .B(new_n8000_), .ZN(new_n23756_));
  NAND2_X1   g20586(.A1(new_n23756_), .A2(new_n13108_), .ZN(new_n23757_));
  NAND2_X1   g20587(.A1(new_n8000_), .A2(new_n17880_), .ZN(new_n23758_));
  NAND4_X1   g20588(.A1(new_n13634_), .A2(pi0188), .A3(new_n3290_), .A4(new_n23758_), .ZN(new_n23759_));
  NOR3_X1    g20589(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n8000_), .ZN(new_n23760_));
  NOR3_X1    g20590(.A1(new_n14422_), .A2(pi0038), .A3(new_n8000_), .ZN(new_n23761_));
  OAI21_X1   g20591(.A1(new_n23760_), .A2(new_n23761_), .B(new_n15655_), .ZN(new_n23762_));
  AOI21_X1   g20592(.A1(new_n23757_), .A2(new_n23759_), .B(new_n23762_), .ZN(new_n23763_));
  NOR3_X1    g20593(.A1(new_n14431_), .A2(new_n8000_), .A3(new_n14081_), .ZN(new_n23764_));
  NOR2_X1    g20594(.A1(new_n23763_), .A2(new_n23764_), .ZN(new_n23765_));
  NOR2_X1    g20595(.A1(new_n23765_), .A2(new_n13620_), .ZN(new_n23766_));
  AOI21_X1   g20596(.A1(new_n23766_), .A2(new_n23755_), .B(pi0625), .ZN(new_n23767_));
  OAI21_X1   g20597(.A1(new_n23767_), .A2(new_n23753_), .B(pi0778), .ZN(new_n23768_));
  NOR3_X1    g20598(.A1(new_n23753_), .A2(new_n13613_), .A3(new_n13748_), .ZN(new_n23772_));
  XOR2_X1    g20599(.A1(new_n23768_), .A2(new_n23772_), .Z(new_n23773_));
  NAND2_X1   g20600(.A1(new_n23755_), .A2(new_n13776_), .ZN(new_n23774_));
  NOR2_X1    g20601(.A1(new_n14428_), .A2(pi0188), .ZN(new_n23775_));
  INV_X1     g20602(.I(new_n23775_), .ZN(new_n23776_));
  NAND2_X1   g20603(.A1(new_n23776_), .A2(new_n13780_), .ZN(new_n23777_));
  AOI21_X1   g20604(.A1(new_n23774_), .A2(new_n23777_), .B(new_n13766_), .ZN(new_n23778_));
  INV_X1     g20605(.I(new_n23778_), .ZN(new_n23779_));
  NAND2_X1   g20606(.A1(new_n23763_), .A2(new_n13748_), .ZN(new_n23780_));
  NOR2_X1    g20607(.A1(new_n23763_), .A2(new_n14452_), .ZN(new_n23781_));
  NOR2_X1    g20608(.A1(new_n23776_), .A2(new_n14452_), .ZN(new_n23782_));
  XNOR2_X1   g20609(.A1(new_n23781_), .A2(new_n23782_), .ZN(new_n23783_));
  OAI21_X1   g20610(.A1(new_n23783_), .A2(new_n13748_), .B(new_n23780_), .ZN(new_n23784_));
  AOI21_X1   g20611(.A1(new_n23784_), .A2(new_n13766_), .B(new_n13785_), .ZN(new_n23785_));
  AOI21_X1   g20612(.A1(new_n23785_), .A2(new_n23779_), .B(pi0609), .ZN(new_n23786_));
  OAI21_X1   g20613(.A1(new_n23786_), .A2(new_n23773_), .B(pi0785), .ZN(new_n23787_));
  NAND2_X1   g20614(.A1(new_n23784_), .A2(pi0609), .ZN(new_n23788_));
  AOI21_X1   g20615(.A1(new_n23776_), .A2(new_n14467_), .B(pi0609), .ZN(new_n23789_));
  NOR2_X1    g20616(.A1(new_n23774_), .A2(new_n23789_), .ZN(new_n23790_));
  NOR2_X1    g20617(.A1(new_n23790_), .A2(new_n14465_), .ZN(new_n23791_));
  AOI21_X1   g20618(.A1(new_n23788_), .A2(new_n23791_), .B(pi0609), .ZN(new_n23792_));
  NOR3_X1    g20619(.A1(new_n23792_), .A2(new_n23773_), .A3(new_n13801_), .ZN(new_n23793_));
  XOR2_X1    g20620(.A1(new_n23787_), .A2(new_n23793_), .Z(new_n23794_));
  NAND2_X1   g20621(.A1(new_n23775_), .A2(new_n13775_), .ZN(new_n23795_));
  OAI21_X1   g20622(.A1(new_n23755_), .A2(new_n13775_), .B(new_n23795_), .ZN(new_n23796_));
  NAND4_X1   g20623(.A1(new_n23778_), .A2(new_n23790_), .A3(pi0785), .A4(new_n23796_), .ZN(new_n23797_));
  NAND3_X1   g20624(.A1(new_n23790_), .A2(pi0785), .A3(new_n23796_), .ZN(new_n23798_));
  NAND3_X1   g20625(.A1(new_n23798_), .A2(new_n23779_), .A3(pi0785), .ZN(new_n23799_));
  NAND2_X1   g20626(.A1(new_n23799_), .A2(new_n23797_), .ZN(new_n23800_));
  NOR2_X1    g20627(.A1(new_n23800_), .A2(new_n13816_), .ZN(new_n23801_));
  NOR2_X1    g20628(.A1(new_n23801_), .A2(new_n13819_), .ZN(new_n23802_));
  NOR3_X1    g20629(.A1(new_n23800_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n23803_));
  OAI21_X1   g20630(.A1(new_n23802_), .A2(new_n23803_), .B(new_n23775_), .ZN(new_n23804_));
  NOR2_X1    g20631(.A1(new_n23776_), .A2(new_n13805_), .ZN(new_n23805_));
  AOI21_X1   g20632(.A1(new_n23784_), .A2(new_n13805_), .B(new_n23805_), .ZN(new_n23806_));
  INV_X1     g20633(.I(new_n23806_), .ZN(new_n23807_));
  AOI21_X1   g20634(.A1(new_n23807_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n23808_));
  AOI21_X1   g20635(.A1(new_n23804_), .A2(new_n23808_), .B(pi0618), .ZN(new_n23809_));
  OR2_X2     g20636(.A1(new_n23809_), .A2(new_n23794_), .Z(new_n23810_));
  NAND3_X1   g20637(.A1(new_n23800_), .A2(pi0618), .A3(pi1154), .ZN(new_n23811_));
  NAND4_X1   g20638(.A1(new_n23799_), .A2(new_n13816_), .A3(pi1154), .A4(new_n23797_), .ZN(new_n23812_));
  AOI21_X1   g20639(.A1(new_n23811_), .A2(new_n23812_), .B(new_n23776_), .ZN(new_n23813_));
  INV_X1     g20640(.I(new_n23813_), .ZN(new_n23814_));
  AOI21_X1   g20641(.A1(new_n23807_), .A2(pi0618), .B(new_n13837_), .ZN(new_n23815_));
  AOI21_X1   g20642(.A1(new_n23814_), .A2(new_n23815_), .B(pi0618), .ZN(new_n23816_));
  OR3_X2     g20643(.A1(new_n23816_), .A2(new_n13855_), .A3(new_n23794_), .Z(new_n23817_));
  AOI21_X1   g20644(.A1(pi0781), .A2(new_n23810_), .B(new_n23817_), .ZN(new_n23818_));
  AND3_X2    g20645(.A1(new_n23817_), .A2(new_n23810_), .A3(pi0781), .Z(new_n23819_));
  NOR2_X1    g20646(.A1(new_n23819_), .A2(new_n23818_), .ZN(new_n23820_));
  INV_X1     g20647(.I(new_n23820_), .ZN(new_n23821_));
  NAND2_X1   g20648(.A1(new_n23804_), .A2(pi0781), .ZN(new_n23822_));
  NAND3_X1   g20649(.A1(new_n23813_), .A2(pi0781), .A3(new_n23800_), .ZN(new_n23823_));
  INV_X1     g20650(.I(new_n23823_), .ZN(new_n23824_));
  NAND2_X1   g20651(.A1(new_n23824_), .A2(new_n23822_), .ZN(new_n23825_));
  NAND3_X1   g20652(.A1(new_n23823_), .A2(new_n23804_), .A3(pi0781), .ZN(new_n23826_));
  NAND2_X1   g20653(.A1(new_n23825_), .A2(new_n23826_), .ZN(new_n23827_));
  NAND3_X1   g20654(.A1(new_n23827_), .A2(pi0619), .A3(pi1159), .ZN(new_n23828_));
  NAND4_X1   g20655(.A1(new_n23825_), .A2(pi0619), .A3(new_n13868_), .A4(new_n23826_), .ZN(new_n23829_));
  AOI21_X1   g20656(.A1(new_n23828_), .A2(new_n23829_), .B(new_n23776_), .ZN(new_n23830_));
  NOR2_X1    g20657(.A1(new_n23775_), .A2(new_n13880_), .ZN(new_n23831_));
  AOI21_X1   g20658(.A1(new_n23806_), .A2(new_n13880_), .B(new_n23831_), .ZN(new_n23832_));
  AOI21_X1   g20659(.A1(new_n23832_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n23833_));
  INV_X1     g20660(.I(new_n23833_), .ZN(new_n23834_));
  OAI21_X1   g20661(.A1(new_n23830_), .A2(new_n23834_), .B(new_n13860_), .ZN(new_n23835_));
  NAND3_X1   g20662(.A1(new_n23827_), .A2(pi0619), .A3(pi1159), .ZN(new_n23836_));
  NAND4_X1   g20663(.A1(new_n23825_), .A2(new_n13860_), .A3(pi1159), .A4(new_n23826_), .ZN(new_n23837_));
  AOI21_X1   g20664(.A1(new_n23836_), .A2(new_n23837_), .B(new_n23776_), .ZN(new_n23838_));
  AOI21_X1   g20665(.A1(new_n23832_), .A2(pi0619), .B(new_n15217_), .ZN(new_n23839_));
  INV_X1     g20666(.I(new_n23839_), .ZN(new_n23840_));
  OAI21_X1   g20667(.A1(new_n23838_), .A2(new_n23840_), .B(new_n13860_), .ZN(new_n23841_));
  NAND4_X1   g20668(.A1(new_n23821_), .A2(new_n23835_), .A3(new_n23841_), .A4(pi0789), .ZN(new_n23842_));
  AOI21_X1   g20669(.A1(new_n23821_), .A2(new_n23835_), .B(new_n13896_), .ZN(new_n23843_));
  NAND3_X1   g20670(.A1(new_n23821_), .A2(new_n23841_), .A3(pi0789), .ZN(new_n23844_));
  NAND2_X1   g20671(.A1(new_n23843_), .A2(new_n23844_), .ZN(new_n23845_));
  NAND2_X1   g20672(.A1(new_n23845_), .A2(new_n23842_), .ZN(new_n23846_));
  NAND4_X1   g20673(.A1(new_n23830_), .A2(new_n23838_), .A3(pi0789), .A4(new_n23827_), .ZN(new_n23847_));
  NAND2_X1   g20674(.A1(new_n23828_), .A2(new_n23829_), .ZN(new_n23848_));
  NAND2_X1   g20675(.A1(new_n23848_), .A2(new_n23775_), .ZN(new_n23849_));
  NAND3_X1   g20676(.A1(new_n23838_), .A2(pi0789), .A3(new_n23827_), .ZN(new_n23850_));
  NAND3_X1   g20677(.A1(new_n23850_), .A2(new_n23849_), .A3(pi0789), .ZN(new_n23851_));
  NOR2_X1    g20678(.A1(new_n23776_), .A2(new_n13919_), .ZN(new_n23852_));
  AOI21_X1   g20679(.A1(new_n23832_), .A2(new_n13919_), .B(new_n23852_), .ZN(new_n23853_));
  NOR2_X1    g20680(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n23854_));
  INV_X1     g20681(.I(new_n23854_), .ZN(new_n23855_));
  AOI21_X1   g20682(.A1(new_n23851_), .A2(new_n23847_), .B(new_n23855_), .ZN(new_n23856_));
  INV_X1     g20683(.I(new_n23847_), .ZN(new_n23857_));
  NOR2_X1    g20684(.A1(new_n23830_), .A2(new_n13896_), .ZN(new_n23858_));
  AND2_X2    g20685(.A1(new_n23850_), .A2(new_n23858_), .Z(new_n23859_));
  NOR2_X1    g20686(.A1(new_n23859_), .A2(new_n23857_), .ZN(new_n23860_));
  NAND3_X1   g20687(.A1(new_n23846_), .A2(pi0626), .A3(pi0788), .ZN(new_n23865_));
  INV_X1     g20688(.I(new_n23865_), .ZN(new_n23866_));
  OAI21_X1   g20689(.A1(new_n23859_), .A2(new_n23857_), .B(new_n23854_), .ZN(new_n23867_));
  AOI22_X1   g20690(.A1(new_n23867_), .A2(new_n13901_), .B1(new_n23842_), .B2(new_n23845_), .ZN(new_n23868_));
  AOI21_X1   g20691(.A1(new_n23845_), .A2(new_n23842_), .B(new_n15258_), .ZN(new_n23869_));
  NOR3_X1    g20692(.A1(new_n23868_), .A2(new_n13937_), .A3(new_n23869_), .ZN(new_n23870_));
  NOR2_X1    g20693(.A1(new_n23870_), .A2(new_n23866_), .ZN(new_n23871_));
  NOR2_X1    g20694(.A1(new_n23775_), .A2(new_n16372_), .ZN(new_n23872_));
  AOI21_X1   g20695(.A1(new_n23860_), .A2(new_n16372_), .B(new_n23872_), .ZN(new_n23873_));
  NOR2_X1    g20696(.A1(new_n23775_), .A2(new_n13966_), .ZN(new_n23874_));
  AOI21_X1   g20697(.A1(new_n23853_), .A2(new_n13966_), .B(new_n23874_), .ZN(new_n23875_));
  NAND2_X1   g20698(.A1(new_n23875_), .A2(pi0628), .ZN(new_n23876_));
  NAND2_X1   g20699(.A1(new_n23876_), .A2(new_n13970_), .ZN(new_n23877_));
  NAND3_X1   g20700(.A1(new_n23875_), .A2(pi0628), .A3(new_n13971_), .ZN(new_n23878_));
  AOI21_X1   g20701(.A1(new_n23877_), .A2(new_n23878_), .B(new_n23776_), .ZN(new_n23879_));
  NOR2_X1    g20702(.A1(new_n23879_), .A2(new_n15270_), .ZN(new_n23880_));
  INV_X1     g20703(.I(new_n23880_), .ZN(new_n23881_));
  NAND2_X1   g20704(.A1(new_n23875_), .A2(pi1156), .ZN(new_n23883_));
  XOR2_X1    g20705(.A1(new_n23883_), .A2(new_n13971_), .Z(new_n23884_));
  NAND2_X1   g20706(.A1(new_n23884_), .A2(new_n23775_), .ZN(new_n23885_));
  NOR3_X1    g20707(.A1(new_n23871_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n23888_));
  INV_X1     g20708(.I(new_n23842_), .ZN(new_n23889_));
  AOI21_X1   g20709(.A1(new_n23849_), .A2(new_n23833_), .B(pi0619), .ZN(new_n23890_));
  OAI21_X1   g20710(.A1(new_n23890_), .A2(new_n23820_), .B(pi0789), .ZN(new_n23891_));
  OR2_X2     g20711(.A1(new_n23838_), .A2(new_n23840_), .Z(new_n23892_));
  OAI21_X1   g20712(.A1(new_n23819_), .A2(new_n23818_), .B(pi0789), .ZN(new_n23893_));
  AOI21_X1   g20713(.A1(new_n23892_), .A2(new_n13860_), .B(new_n23893_), .ZN(new_n23894_));
  NOR2_X1    g20714(.A1(new_n23891_), .A2(new_n23894_), .ZN(new_n23895_));
  OAI22_X1   g20715(.A1(new_n23895_), .A2(new_n23889_), .B1(pi0626), .B2(new_n23856_), .ZN(new_n23896_));
  OAI21_X1   g20716(.A1(new_n23895_), .A2(new_n23889_), .B(new_n14577_), .ZN(new_n23897_));
  NAND3_X1   g20717(.A1(new_n23896_), .A2(new_n23897_), .A3(pi0788), .ZN(new_n23898_));
  NAND3_X1   g20718(.A1(new_n23851_), .A2(new_n16372_), .A3(new_n23847_), .ZN(new_n23899_));
  OAI21_X1   g20719(.A1(new_n16372_), .A2(new_n23775_), .B(new_n23899_), .ZN(new_n23900_));
  AOI21_X1   g20720(.A1(new_n23900_), .A2(new_n23880_), .B(pi0628), .ZN(new_n23901_));
  AOI21_X1   g20721(.A1(new_n23898_), .A2(new_n23865_), .B(new_n23901_), .ZN(new_n23902_));
  AOI21_X1   g20722(.A1(new_n23898_), .A2(new_n23865_), .B(new_n15296_), .ZN(new_n23903_));
  NOR3_X1    g20723(.A1(new_n23902_), .A2(new_n23903_), .A3(new_n12777_), .ZN(new_n23904_));
  NOR2_X1    g20724(.A1(new_n23904_), .A2(new_n23888_), .ZN(new_n23905_));
  NOR2_X1    g20725(.A1(new_n23775_), .A2(new_n13994_), .ZN(new_n23906_));
  AOI21_X1   g20726(.A1(new_n23900_), .A2(new_n13994_), .B(new_n23906_), .ZN(new_n23907_));
  INV_X1     g20727(.I(new_n23907_), .ZN(new_n23908_));
  NOR2_X1    g20728(.A1(new_n23879_), .A2(new_n12777_), .ZN(new_n23909_));
  NOR4_X1    g20729(.A1(new_n23885_), .A2(new_n12777_), .A3(new_n23909_), .A4(new_n23875_), .ZN(new_n23910_));
  NOR3_X1    g20730(.A1(new_n23885_), .A2(new_n12777_), .A3(new_n23875_), .ZN(new_n23911_));
  NOR3_X1    g20731(.A1(new_n23911_), .A2(new_n12777_), .A3(new_n23879_), .ZN(new_n23912_));
  NOR2_X1    g20732(.A1(new_n23912_), .A2(new_n23910_), .ZN(new_n23913_));
  NAND2_X1   g20733(.A1(new_n23913_), .A2(pi0647), .ZN(new_n23914_));
  XOR2_X1    g20734(.A1(new_n23914_), .A2(new_n14008_), .Z(new_n23915_));
  AOI21_X1   g20735(.A1(new_n23915_), .A2(new_n23775_), .B(new_n14012_), .ZN(new_n23916_));
  AOI21_X1   g20736(.A1(new_n23908_), .A2(new_n23916_), .B(pi0647), .ZN(new_n23917_));
  AOI21_X1   g20737(.A1(new_n23913_), .A2(pi1157), .B(new_n14008_), .ZN(new_n23918_));
  NOR4_X1    g20738(.A1(new_n23912_), .A2(new_n23910_), .A3(pi0647), .A4(new_n14006_), .ZN(new_n23919_));
  OAI21_X1   g20739(.A1(new_n23918_), .A2(new_n23919_), .B(new_n23775_), .ZN(new_n23920_));
  NAND2_X1   g20740(.A1(new_n23920_), .A2(new_n14027_), .ZN(new_n23921_));
  AOI21_X1   g20741(.A1(new_n23907_), .A2(pi0647), .B(new_n23921_), .ZN(new_n23922_));
  NOR2_X1    g20742(.A1(new_n23922_), .A2(pi0647), .ZN(new_n23923_));
  NOR4_X1    g20743(.A1(new_n23905_), .A2(new_n12776_), .A3(new_n23917_), .A4(new_n23923_), .ZN(new_n23924_));
  NAND2_X1   g20744(.A1(new_n23898_), .A2(new_n23865_), .ZN(new_n23925_));
  NAND3_X1   g20745(.A1(new_n23925_), .A2(pi0628), .A3(pi0792), .ZN(new_n23926_));
  OAI21_X1   g20746(.A1(new_n23873_), .A2(new_n23881_), .B(new_n13942_), .ZN(new_n23927_));
  OAI21_X1   g20747(.A1(new_n23870_), .A2(new_n23866_), .B(new_n23927_), .ZN(new_n23928_));
  OAI21_X1   g20748(.A1(new_n23870_), .A2(new_n23866_), .B(new_n14606_), .ZN(new_n23929_));
  NAND3_X1   g20749(.A1(new_n23928_), .A2(new_n23929_), .A3(pi0792), .ZN(new_n23930_));
  AOI21_X1   g20750(.A1(new_n23930_), .A2(new_n23926_), .B(new_n23917_), .ZN(new_n23931_));
  OAI21_X1   g20751(.A1(new_n23922_), .A2(pi0647), .B(pi0787), .ZN(new_n23932_));
  AOI21_X1   g20752(.A1(new_n23930_), .A2(new_n23926_), .B(new_n23932_), .ZN(new_n23933_));
  NOR3_X1    g20753(.A1(new_n23931_), .A2(new_n23933_), .A3(new_n12776_), .ZN(new_n23934_));
  OAI21_X1   g20754(.A1(new_n23934_), .A2(new_n23924_), .B(new_n12775_), .ZN(new_n23935_));
  NOR2_X1    g20755(.A1(new_n9992_), .A2(pi0188), .ZN(new_n23936_));
  NOR2_X1    g20756(.A1(new_n14652_), .A2(new_n17880_), .ZN(new_n23937_));
  AOI21_X1   g20757(.A1(new_n13218_), .A2(pi0705), .B(new_n23936_), .ZN(new_n23938_));
  INV_X1     g20758(.I(new_n23938_), .ZN(new_n23939_));
  NAND3_X1   g20759(.A1(new_n23939_), .A2(new_n23937_), .A3(new_n23936_), .ZN(new_n23940_));
  NOR3_X1    g20760(.A1(new_n23937_), .A2(new_n13614_), .A3(new_n23938_), .ZN(new_n23941_));
  XNOR2_X1   g20761(.A1(new_n23940_), .A2(new_n23941_), .ZN(new_n23942_));
  NAND2_X1   g20762(.A1(new_n23942_), .A2(pi0778), .ZN(new_n23943_));
  NAND2_X1   g20763(.A1(new_n23939_), .A2(new_n13748_), .ZN(new_n23944_));
  NAND2_X1   g20764(.A1(new_n23943_), .A2(new_n23944_), .ZN(new_n23945_));
  INV_X1     g20765(.I(new_n23945_), .ZN(new_n23946_));
  NOR2_X1    g20766(.A1(new_n23946_), .A2(new_n14048_), .ZN(new_n23947_));
  INV_X1     g20767(.I(new_n23947_), .ZN(new_n23948_));
  NOR2_X1    g20768(.A1(new_n23948_), .A2(new_n14051_), .ZN(new_n23949_));
  INV_X1     g20769(.I(new_n23949_), .ZN(new_n23950_));
  NOR2_X1    g20770(.A1(new_n23950_), .A2(new_n14163_), .ZN(new_n23951_));
  AOI21_X1   g20771(.A1(new_n13104_), .A2(new_n17881_), .B(new_n23936_), .ZN(new_n23952_));
  NOR2_X1    g20772(.A1(new_n14096_), .A2(new_n23952_), .ZN(new_n23953_));
  AOI21_X1   g20773(.A1(new_n23953_), .A2(new_n14094_), .B(pi1155), .ZN(new_n23954_));
  NOR2_X1    g20774(.A1(new_n23954_), .A2(new_n13801_), .ZN(new_n23955_));
  AOI21_X1   g20775(.A1(new_n23952_), .A2(pi1155), .B(new_n9992_), .ZN(new_n23956_));
  NOR2_X1    g20776(.A1(new_n23956_), .A2(new_n14102_), .ZN(new_n23957_));
  NAND3_X1   g20777(.A1(new_n23957_), .A2(new_n23953_), .A3(pi0785), .ZN(new_n23958_));
  XOR2_X1    g20778(.A1(new_n23955_), .A2(new_n23958_), .Z(new_n23959_));
  NOR2_X1    g20779(.A1(new_n23959_), .A2(new_n13817_), .ZN(new_n23960_));
  OAI21_X1   g20780(.A1(new_n23960_), .A2(pi0618), .B(new_n9992_), .ZN(new_n23961_));
  NAND2_X1   g20781(.A1(new_n23961_), .A2(pi0781), .ZN(new_n23962_));
  OAI21_X1   g20782(.A1(new_n23960_), .A2(new_n9992_), .B(pi0618), .ZN(new_n23963_));
  NOR3_X1    g20783(.A1(new_n23963_), .A2(new_n13855_), .A3(new_n23959_), .ZN(new_n23964_));
  XOR2_X1    g20784(.A1(new_n23964_), .A2(new_n23962_), .Z(new_n23965_));
  NAND2_X1   g20785(.A1(new_n23965_), .A2(pi0619), .ZN(new_n23966_));
  XOR2_X1    g20786(.A1(new_n23966_), .A2(new_n13904_), .Z(new_n23967_));
  NAND2_X1   g20787(.A1(new_n23967_), .A2(new_n23936_), .ZN(new_n23968_));
  NAND2_X1   g20788(.A1(new_n23968_), .A2(pi0789), .ZN(new_n23969_));
  NAND2_X1   g20789(.A1(new_n23965_), .A2(pi1159), .ZN(new_n23970_));
  XOR2_X1    g20790(.A1(new_n23970_), .A2(new_n13904_), .Z(new_n23971_));
  NAND2_X1   g20791(.A1(new_n23971_), .A2(new_n23936_), .ZN(new_n23972_));
  NOR3_X1    g20792(.A1(new_n23972_), .A2(new_n13896_), .A3(new_n23965_), .ZN(new_n23973_));
  XOR2_X1    g20793(.A1(new_n23973_), .A2(new_n23969_), .Z(new_n23974_));
  NAND2_X1   g20794(.A1(new_n23974_), .A2(new_n13962_), .ZN(new_n23975_));
  XOR2_X1    g20795(.A1(new_n23975_), .A2(new_n18976_), .Z(new_n23976_));
  AOI22_X1   g20796(.A1(new_n23976_), .A2(new_n23936_), .B1(new_n16639_), .B2(new_n23951_), .ZN(new_n23977_));
  NOR2_X1    g20797(.A1(new_n23938_), .A2(new_n13203_), .ZN(new_n23978_));
  INV_X1     g20798(.I(new_n23978_), .ZN(new_n23979_));
  NOR2_X1    g20799(.A1(new_n23979_), .A2(new_n13613_), .ZN(new_n23980_));
  NOR2_X1    g20800(.A1(new_n23936_), .A2(pi1153), .ZN(new_n23981_));
  INV_X1     g20801(.I(new_n23981_), .ZN(new_n23982_));
  OAI21_X1   g20802(.A1(new_n23937_), .A2(new_n23982_), .B(pi0608), .ZN(new_n23983_));
  NOR2_X1    g20803(.A1(new_n23952_), .A2(pi1153), .ZN(new_n23984_));
  NAND2_X1   g20804(.A1(new_n23983_), .A2(new_n23984_), .ZN(new_n23985_));
  AOI21_X1   g20805(.A1(new_n23985_), .A2(new_n23980_), .B(new_n13748_), .ZN(new_n23986_));
  NOR2_X1    g20806(.A1(new_n23938_), .A2(new_n14082_), .ZN(new_n23987_));
  NAND2_X1   g20807(.A1(new_n23937_), .A2(new_n23981_), .ZN(new_n23988_));
  OAI22_X1   g20808(.A1(new_n23979_), .A2(new_n13613_), .B1(new_n23988_), .B2(new_n23987_), .ZN(new_n23989_));
  NAND4_X1   g20809(.A1(new_n23989_), .A2(pi0778), .A3(new_n23952_), .A4(new_n23979_), .ZN(new_n23990_));
  XNOR2_X1   g20810(.A1(new_n23990_), .A2(new_n23986_), .ZN(new_n23991_));
  NAND2_X1   g20811(.A1(new_n23991_), .A2(new_n13801_), .ZN(new_n23992_));
  NOR2_X1    g20812(.A1(new_n23991_), .A2(new_n13778_), .ZN(new_n23993_));
  XOR2_X1    g20813(.A1(new_n23993_), .A2(new_n14694_), .Z(new_n23994_));
  NOR2_X1    g20814(.A1(new_n23994_), .A2(new_n23946_), .ZN(new_n23995_));
  NOR3_X1    g20815(.A1(new_n23995_), .A2(new_n13783_), .A3(new_n23954_), .ZN(new_n23996_));
  NOR3_X1    g20816(.A1(new_n23996_), .A2(pi0660), .A3(new_n23957_), .ZN(new_n23997_));
  NOR2_X1    g20817(.A1(new_n23991_), .A2(new_n13766_), .ZN(new_n23998_));
  XOR2_X1    g20818(.A1(new_n23998_), .A2(new_n14090_), .Z(new_n23999_));
  NAND3_X1   g20819(.A1(new_n23999_), .A2(pi0785), .A3(new_n23945_), .ZN(new_n24000_));
  OAI21_X1   g20820(.A1(new_n23997_), .A2(new_n24000_), .B(new_n23992_), .ZN(new_n24001_));
  NAND2_X1   g20821(.A1(new_n24001_), .A2(new_n13855_), .ZN(new_n24002_));
  NOR2_X1    g20822(.A1(new_n24001_), .A2(new_n13816_), .ZN(new_n24003_));
  XOR2_X1    g20823(.A1(new_n24003_), .A2(new_n13818_), .Z(new_n24004_));
  NAND2_X1   g20824(.A1(new_n24004_), .A2(new_n23947_), .ZN(new_n24005_));
  NAND3_X1   g20825(.A1(new_n24005_), .A2(new_n13823_), .A3(new_n23963_), .ZN(new_n24006_));
  AND3_X2    g20826(.A1(new_n24006_), .A2(new_n13823_), .A3(new_n23961_), .Z(new_n24007_));
  NOR2_X1    g20827(.A1(new_n24001_), .A2(new_n13817_), .ZN(new_n24008_));
  XOR2_X1    g20828(.A1(new_n24008_), .A2(new_n13819_), .Z(new_n24009_));
  NOR3_X1    g20829(.A1(new_n24009_), .A2(new_n13855_), .A3(new_n23948_), .ZN(new_n24010_));
  INV_X1     g20830(.I(new_n24010_), .ZN(new_n24011_));
  OAI21_X1   g20831(.A1(new_n24007_), .A2(new_n24011_), .B(new_n24002_), .ZN(new_n24012_));
  NOR2_X1    g20832(.A1(new_n24012_), .A2(new_n13860_), .ZN(new_n24013_));
  XOR2_X1    g20833(.A1(new_n24013_), .A2(new_n13904_), .Z(new_n24014_));
  NOR2_X1    g20834(.A1(new_n24014_), .A2(new_n23950_), .ZN(new_n24015_));
  NAND2_X1   g20835(.A1(new_n23972_), .A2(new_n13884_), .ZN(new_n24016_));
  INV_X1     g20836(.I(new_n24012_), .ZN(new_n24017_));
  AOI21_X1   g20837(.A1(new_n24017_), .A2(new_n14143_), .B(pi0789), .ZN(new_n24018_));
  OAI21_X1   g20838(.A1(new_n24015_), .A2(new_n24016_), .B(new_n24018_), .ZN(new_n24019_));
  NOR2_X1    g20839(.A1(new_n24012_), .A2(new_n13868_), .ZN(new_n24020_));
  XOR2_X1    g20840(.A1(new_n24020_), .A2(new_n13903_), .Z(new_n24021_));
  NAND2_X1   g20841(.A1(new_n23968_), .A2(new_n19018_), .ZN(new_n24022_));
  AOI21_X1   g20842(.A1(new_n24021_), .A2(new_n23949_), .B(new_n24022_), .ZN(new_n24023_));
  AOI21_X1   g20843(.A1(new_n24019_), .A2(new_n24023_), .B(new_n23977_), .ZN(new_n24024_));
  NAND2_X1   g20844(.A1(new_n23974_), .A2(new_n16372_), .ZN(new_n24025_));
  OAI21_X1   g20845(.A1(new_n16372_), .A2(new_n23936_), .B(new_n24025_), .ZN(new_n24026_));
  NAND3_X1   g20846(.A1(new_n24026_), .A2(new_n18929_), .A3(new_n23951_), .ZN(new_n24027_));
  NAND2_X1   g20847(.A1(new_n24027_), .A2(new_n16569_), .ZN(new_n24028_));
  XOR2_X1    g20848(.A1(new_n24028_), .A2(new_n16572_), .Z(new_n24029_));
  AOI21_X1   g20849(.A1(new_n19022_), .A2(new_n24027_), .B(new_n24029_), .ZN(new_n24030_));
  INV_X1     g20850(.I(new_n23936_), .ZN(new_n24031_));
  NAND2_X1   g20851(.A1(new_n23974_), .A2(new_n13963_), .ZN(new_n24032_));
  XNOR2_X1   g20852(.A1(new_n24032_), .A2(new_n19028_), .ZN(new_n24033_));
  NOR3_X1    g20853(.A1(new_n24033_), .A2(new_n16424_), .A3(new_n24031_), .ZN(new_n24034_));
  OAI21_X1   g20854(.A1(new_n24030_), .A2(new_n16574_), .B(new_n24034_), .ZN(new_n24035_));
  NOR4_X1    g20855(.A1(new_n23950_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n24036_));
  NOR2_X1    g20856(.A1(new_n24036_), .A2(new_n14005_), .ZN(new_n24037_));
  XOR2_X1    g20857(.A1(new_n24037_), .A2(new_n14007_), .Z(new_n24038_));
  NAND2_X1   g20858(.A1(new_n24038_), .A2(new_n23936_), .ZN(new_n24039_));
  NOR2_X1    g20859(.A1(new_n24031_), .A2(pi0647), .ZN(new_n24040_));
  AOI21_X1   g20860(.A1(new_n24036_), .A2(pi0647), .B(new_n24040_), .ZN(new_n24041_));
  NOR2_X1    g20861(.A1(new_n24026_), .A2(new_n13994_), .ZN(new_n24042_));
  XNOR2_X1   g20862(.A1(new_n24042_), .A2(new_n19033_), .ZN(new_n24043_));
  AOI22_X1   g20863(.A1(new_n24043_), .A2(new_n23936_), .B1(new_n14206_), .B2(new_n24041_), .ZN(new_n24044_));
  NOR3_X1    g20864(.A1(new_n24044_), .A2(new_n14010_), .A3(new_n24039_), .ZN(new_n24045_));
  OAI22_X1   g20865(.A1(new_n24024_), .A2(new_n24035_), .B1(new_n12776_), .B2(new_n24045_), .ZN(new_n24046_));
  AOI21_X1   g20866(.A1(new_n24041_), .A2(pi1157), .B(new_n12776_), .ZN(new_n24047_));
  AOI22_X1   g20867(.A1(new_n24039_), .A2(new_n24047_), .B1(new_n12776_), .B2(new_n24036_), .ZN(new_n24048_));
  NAND2_X1   g20868(.A1(new_n24046_), .A2(pi0644), .ZN(new_n24049_));
  XOR2_X1    g20869(.A1(new_n24049_), .A2(new_n14205_), .Z(new_n24050_));
  NOR2_X1    g20870(.A1(new_n24050_), .A2(new_n24048_), .ZN(new_n24051_));
  NOR2_X1    g20871(.A1(new_n24026_), .A2(new_n18968_), .ZN(new_n24052_));
  NAND2_X1   g20872(.A1(new_n18967_), .A2(new_n23936_), .ZN(new_n24053_));
  XOR2_X1    g20873(.A1(new_n24052_), .A2(new_n24053_), .Z(new_n24054_));
  NAND2_X1   g20874(.A1(new_n24054_), .A2(pi0715), .ZN(new_n24055_));
  XOR2_X1    g20875(.A1(new_n24055_), .A2(new_n14205_), .Z(new_n24056_));
  OAI21_X1   g20876(.A1(new_n24056_), .A2(new_n24031_), .B(new_n14203_), .ZN(new_n24057_));
  NAND2_X1   g20877(.A1(new_n24054_), .A2(pi0644), .ZN(new_n24058_));
  XOR2_X1    g20878(.A1(new_n24058_), .A2(new_n14217_), .Z(new_n24059_));
  AOI21_X1   g20879(.A1(new_n24059_), .A2(new_n23936_), .B(pi1160), .ZN(new_n24060_));
  OAI21_X1   g20880(.A1(new_n24051_), .A2(new_n24057_), .B(new_n24060_), .ZN(new_n24061_));
  NAND2_X1   g20881(.A1(new_n24046_), .A2(pi0715), .ZN(new_n24062_));
  XOR2_X1    g20882(.A1(new_n24062_), .A2(new_n14205_), .Z(new_n24063_));
  NOR2_X1    g20883(.A1(new_n24063_), .A2(new_n24048_), .ZN(new_n24064_));
  AOI21_X1   g20884(.A1(new_n24061_), .A2(new_n24064_), .B(new_n14799_), .ZN(new_n24065_));
  XOR2_X1    g20885(.A1(new_n24065_), .A2(new_n14801_), .Z(new_n24066_));
  NOR2_X1    g20886(.A1(new_n7240_), .A2(pi0188), .ZN(new_n24067_));
  NOR4_X1    g20887(.A1(new_n24066_), .A2(pi0832), .A3(new_n24046_), .A4(new_n24067_), .ZN(new_n24068_));
  AOI21_X1   g20888(.A1(new_n23935_), .A2(new_n7240_), .B(new_n24068_), .ZN(new_n24069_));
  NOR3_X1    g20889(.A1(new_n23934_), .A2(new_n23924_), .A3(new_n14200_), .ZN(new_n24070_));
  NOR2_X1    g20890(.A1(new_n24070_), .A2(new_n14217_), .ZN(new_n24071_));
  NOR4_X1    g20891(.A1(new_n23934_), .A2(new_n23924_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n24072_));
  NOR2_X1    g20892(.A1(new_n24071_), .A2(new_n24072_), .ZN(new_n24073_));
  OAI21_X1   g20893(.A1(new_n12776_), .A2(new_n23931_), .B(new_n23933_), .ZN(new_n24074_));
  INV_X1     g20894(.I(new_n23917_), .ZN(new_n24075_));
  OAI21_X1   g20895(.A1(new_n23888_), .A2(new_n23904_), .B(new_n24075_), .ZN(new_n24076_));
  INV_X1     g20896(.I(new_n23932_), .ZN(new_n24077_));
  OAI21_X1   g20897(.A1(new_n23888_), .A2(new_n23904_), .B(new_n24077_), .ZN(new_n24078_));
  NAND3_X1   g20898(.A1(new_n24078_), .A2(new_n24076_), .A3(pi0787), .ZN(new_n24079_));
  NOR2_X1    g20899(.A1(new_n23776_), .A2(new_n14211_), .ZN(new_n24080_));
  AOI21_X1   g20900(.A1(new_n23907_), .A2(new_n14211_), .B(new_n24080_), .ZN(new_n24081_));
  OAI21_X1   g20901(.A1(new_n23776_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n24082_));
  NAND2_X1   g20902(.A1(new_n24081_), .A2(new_n24082_), .ZN(new_n24083_));
  AOI21_X1   g20903(.A1(new_n23915_), .A2(new_n23775_), .B(new_n12776_), .ZN(new_n24084_));
  NOR3_X1    g20904(.A1(new_n23920_), .A2(new_n12776_), .A3(new_n23913_), .ZN(new_n24085_));
  XNOR2_X1   g20905(.A1(new_n24084_), .A2(new_n24085_), .ZN(new_n24086_));
  AOI21_X1   g20906(.A1(new_n24083_), .A2(new_n14815_), .B(pi0644), .ZN(new_n24087_));
  AOI21_X1   g20907(.A1(new_n24079_), .A2(new_n24074_), .B(new_n24087_), .ZN(new_n24088_));
  AOI21_X1   g20908(.A1(new_n23776_), .A2(new_n14254_), .B(pi0644), .ZN(new_n24089_));
  NOR3_X1    g20909(.A1(new_n24086_), .A2(new_n24081_), .A3(new_n24089_), .ZN(new_n24090_));
  OAI21_X1   g20910(.A1(new_n24088_), .A2(pi0790), .B(new_n24090_), .ZN(new_n24091_));
  NOR3_X1    g20911(.A1(new_n24073_), .A2(new_n24069_), .A3(new_n24091_), .ZN(po0345));
  NOR3_X1    g20912(.A1(new_n13085_), .A2(new_n16088_), .A3(new_n17845_), .ZN(new_n24093_));
  NOR3_X1    g20913(.A1(new_n12977_), .A2(new_n16086_), .A3(new_n17845_), .ZN(new_n24094_));
  NAND3_X1   g20914(.A1(new_n14356_), .A2(pi0039), .A3(pi0772), .ZN(new_n24095_));
  NAND3_X1   g20915(.A1(new_n14338_), .A2(new_n3183_), .A3(pi0772), .ZN(new_n24096_));
  NAND2_X1   g20916(.A1(new_n14874_), .A2(pi0189), .ZN(new_n24097_));
  AOI21_X1   g20917(.A1(new_n24095_), .A2(new_n24096_), .B(new_n24097_), .ZN(new_n24098_));
  OAI22_X1   g20918(.A1(new_n24094_), .A2(new_n24093_), .B1(pi0039), .B2(new_n24098_), .ZN(new_n24099_));
  AOI21_X1   g20919(.A1(new_n13203_), .A2(pi0772), .B(new_n3259_), .ZN(new_n24100_));
  XOR2_X1    g20920(.A1(new_n13723_), .A2(new_n24100_), .Z(new_n24101_));
  NAND2_X1   g20921(.A1(new_n24101_), .A2(pi0189), .ZN(new_n24102_));
  OAI21_X1   g20922(.A1(new_n3259_), .A2(new_n24102_), .B(new_n24099_), .ZN(new_n24103_));
  NAND4_X1   g20923(.A1(new_n24103_), .A2(new_n8642_), .A3(pi0772), .A4(new_n16114_), .ZN(new_n24104_));
  NOR2_X1    g20924(.A1(new_n24104_), .A2(new_n3290_), .ZN(new_n24105_));
  NOR2_X1    g20925(.A1(new_n3289_), .A2(pi0189), .ZN(new_n24106_));
  OR2_X2     g20926(.A1(new_n24105_), .A2(new_n24106_), .Z(new_n24107_));
  NAND3_X1   g20927(.A1(new_n14270_), .A2(pi0189), .A3(pi0772), .ZN(new_n24108_));
  NAND3_X1   g20928(.A1(new_n14272_), .A2(pi0189), .A3(new_n17845_), .ZN(new_n24109_));
  NAND2_X1   g20929(.A1(new_n24109_), .A2(new_n24108_), .ZN(new_n24110_));
  AOI21_X1   g20930(.A1(new_n14269_), .A2(new_n24110_), .B(new_n3212_), .ZN(new_n24111_));
  NOR3_X1    g20931(.A1(new_n13200_), .A2(new_n8642_), .A3(new_n17845_), .ZN(new_n24112_));
  NOR3_X1    g20932(.A1(new_n13198_), .A2(pi0189), .A3(new_n17845_), .ZN(new_n24113_));
  OAI21_X1   g20933(.A1(new_n24112_), .A2(new_n24113_), .B(new_n13190_), .ZN(new_n24114_));
  NOR2_X1    g20934(.A1(new_n3290_), .A2(new_n17866_), .ZN(new_n24115_));
  NAND3_X1   g20935(.A1(new_n24102_), .A2(new_n15630_), .A3(new_n24115_), .ZN(new_n24116_));
  OAI21_X1   g20936(.A1(new_n24111_), .A2(new_n24114_), .B(new_n24116_), .ZN(new_n24117_));
  NAND4_X1   g20937(.A1(new_n24117_), .A2(pi0189), .A3(new_n3290_), .A4(new_n14284_), .ZN(new_n24122_));
  AOI21_X1   g20938(.A1(new_n24122_), .A2(new_n24104_), .B(new_n17866_), .ZN(new_n24123_));
  NAND3_X1   g20939(.A1(new_n24123_), .A2(pi0625), .A3(pi1153), .ZN(new_n24124_));
  INV_X1     g20940(.I(new_n24123_), .ZN(new_n24125_));
  NAND3_X1   g20941(.A1(new_n24125_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n24126_));
  NAND2_X1   g20942(.A1(new_n24126_), .A2(new_n24124_), .ZN(new_n24127_));
  NAND3_X1   g20943(.A1(new_n14422_), .A2(pi0038), .A3(pi0189), .ZN(new_n24128_));
  NAND3_X1   g20944(.A1(new_n14424_), .A2(new_n3259_), .A3(pi0189), .ZN(new_n24129_));
  AOI21_X1   g20945(.A1(new_n24129_), .A2(new_n24128_), .B(new_n14404_), .ZN(new_n24130_));
  OAI21_X1   g20946(.A1(new_n16149_), .A2(new_n8642_), .B(new_n24115_), .ZN(new_n24131_));
  NOR2_X1    g20947(.A1(new_n24130_), .A2(new_n24131_), .ZN(new_n24132_));
  NOR2_X1    g20948(.A1(new_n24132_), .A2(pi0189), .ZN(new_n24133_));
  NOR2_X1    g20949(.A1(new_n24133_), .A2(new_n13627_), .ZN(new_n24134_));
  NOR2_X1    g20950(.A1(new_n14428_), .A2(new_n8642_), .ZN(new_n24135_));
  NOR2_X1    g20951(.A1(new_n24135_), .A2(new_n13613_), .ZN(new_n24136_));
  XOR2_X1    g20952(.A1(new_n24136_), .A2(new_n13615_), .Z(new_n24137_));
  NAND2_X1   g20953(.A1(new_n24137_), .A2(new_n24134_), .ZN(new_n24138_));
  NAND2_X1   g20954(.A1(new_n24138_), .A2(pi0608), .ZN(new_n24139_));
  AOI21_X1   g20955(.A1(new_n24127_), .A2(new_n24107_), .B(new_n24139_), .ZN(new_n24140_));
  NOR2_X1    g20956(.A1(new_n24140_), .A2(new_n13748_), .ZN(new_n24141_));
  INV_X1     g20957(.I(new_n24107_), .ZN(new_n24142_));
  NAND3_X1   g20958(.A1(new_n24123_), .A2(pi0625), .A3(pi1153), .ZN(new_n24143_));
  NAND3_X1   g20959(.A1(new_n24125_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n24144_));
  AOI21_X1   g20960(.A1(new_n24144_), .A2(new_n24143_), .B(new_n24142_), .ZN(new_n24145_));
  NOR2_X1    g20961(.A1(new_n24135_), .A2(new_n13614_), .ZN(new_n24146_));
  XOR2_X1    g20962(.A1(new_n24146_), .A2(new_n13615_), .Z(new_n24147_));
  AND2_X2    g20963(.A1(new_n24147_), .A2(new_n24134_), .Z(new_n24148_));
  NOR4_X1    g20964(.A1(new_n24145_), .A2(new_n13750_), .A3(new_n24125_), .A4(new_n24148_), .ZN(new_n24149_));
  XOR2_X1    g20965(.A1(new_n24141_), .A2(new_n24149_), .Z(new_n24150_));
  INV_X1     g20966(.I(new_n24150_), .ZN(new_n24151_));
  NAND2_X1   g20967(.A1(new_n24138_), .A2(pi0778), .ZN(new_n24152_));
  NAND3_X1   g20968(.A1(new_n24147_), .A2(pi0778), .A3(new_n24134_), .ZN(new_n24153_));
  XNOR2_X1   g20969(.A1(new_n24152_), .A2(new_n24153_), .ZN(new_n24154_));
  INV_X1     g20970(.I(new_n24135_), .ZN(new_n24155_));
  NAND2_X1   g20971(.A1(new_n24135_), .A2(new_n13775_), .ZN(new_n24156_));
  OAI21_X1   g20972(.A1(new_n24107_), .A2(new_n13775_), .B(new_n24156_), .ZN(new_n24157_));
  NAND3_X1   g20973(.A1(new_n24157_), .A2(pi0609), .A3(pi1155), .ZN(new_n24158_));
  INV_X1     g20974(.I(new_n24157_), .ZN(new_n24159_));
  NAND3_X1   g20975(.A1(new_n24159_), .A2(pi0609), .A3(new_n14694_), .ZN(new_n24160_));
  AOI21_X1   g20976(.A1(new_n24160_), .A2(new_n24158_), .B(new_n24155_), .ZN(new_n24161_));
  NOR2_X1    g20977(.A1(new_n24161_), .A2(new_n13785_), .ZN(new_n24162_));
  AOI21_X1   g20978(.A1(new_n24162_), .A2(new_n24154_), .B(pi0609), .ZN(new_n24163_));
  OAI21_X1   g20979(.A1(new_n24151_), .A2(new_n24163_), .B(pi0785), .ZN(new_n24164_));
  NOR2_X1    g20980(.A1(new_n24154_), .A2(new_n13766_), .ZN(new_n24165_));
  NAND3_X1   g20981(.A1(new_n24157_), .A2(pi0609), .A3(pi1155), .ZN(new_n24166_));
  INV_X1     g20982(.I(new_n24166_), .ZN(new_n24167_));
  NOR3_X1    g20983(.A1(new_n24157_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n24168_));
  OAI21_X1   g20984(.A1(new_n24167_), .A2(new_n24168_), .B(new_n24135_), .ZN(new_n24169_));
  NAND2_X1   g20985(.A1(new_n24169_), .A2(new_n13793_), .ZN(new_n24170_));
  OAI21_X1   g20986(.A1(new_n24165_), .A2(new_n24170_), .B(new_n13766_), .ZN(new_n24171_));
  NAND3_X1   g20987(.A1(new_n24150_), .A2(new_n24171_), .A3(pi0785), .ZN(new_n24172_));
  XNOR2_X1   g20988(.A1(new_n24164_), .A2(new_n24172_), .ZN(new_n24173_));
  INV_X1     g20989(.I(new_n24168_), .ZN(new_n24174_));
  AOI21_X1   g20990(.A1(new_n24174_), .A2(new_n24166_), .B(new_n24155_), .ZN(new_n24175_));
  NAND4_X1   g20991(.A1(new_n24175_), .A2(new_n24161_), .A3(pi0785), .A4(new_n24157_), .ZN(new_n24176_));
  INV_X1     g20992(.I(new_n24176_), .ZN(new_n24177_));
  NOR3_X1    g20993(.A1(new_n24169_), .A2(new_n13801_), .A3(new_n24159_), .ZN(new_n24178_));
  NOR3_X1    g20994(.A1(new_n24178_), .A2(new_n13801_), .A3(new_n24161_), .ZN(new_n24179_));
  NOR2_X1    g20995(.A1(new_n24179_), .A2(new_n24177_), .ZN(new_n24180_));
  AOI21_X1   g20996(.A1(new_n24180_), .A2(pi0618), .B(new_n13819_), .ZN(new_n24181_));
  NOR2_X1    g20997(.A1(new_n24161_), .A2(new_n13801_), .ZN(new_n24182_));
  NOR2_X1    g20998(.A1(new_n24159_), .A2(new_n13801_), .ZN(new_n24183_));
  NAND2_X1   g20999(.A1(new_n24175_), .A2(new_n24183_), .ZN(new_n24184_));
  NAND2_X1   g21000(.A1(new_n24184_), .A2(new_n24182_), .ZN(new_n24185_));
  NAND2_X1   g21001(.A1(new_n24185_), .A2(new_n24176_), .ZN(new_n24186_));
  NOR3_X1    g21002(.A1(new_n24186_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n24187_));
  OAI21_X1   g21003(.A1(new_n24181_), .A2(new_n24187_), .B(new_n24135_), .ZN(new_n24188_));
  NOR2_X1    g21004(.A1(new_n24155_), .A2(new_n13805_), .ZN(new_n24189_));
  AOI21_X1   g21005(.A1(new_n24154_), .A2(new_n13805_), .B(new_n24189_), .ZN(new_n24190_));
  AOI21_X1   g21006(.A1(new_n24190_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n24191_));
  AOI21_X1   g21007(.A1(new_n24188_), .A2(new_n24191_), .B(pi0618), .ZN(new_n24192_));
  OAI21_X1   g21008(.A1(new_n24173_), .A2(new_n24192_), .B(pi0781), .ZN(new_n24193_));
  XOR2_X1    g21009(.A1(new_n24164_), .A2(new_n24172_), .Z(new_n24194_));
  NAND3_X1   g21010(.A1(new_n24186_), .A2(pi0618), .A3(pi1154), .ZN(new_n24195_));
  NAND4_X1   g21011(.A1(new_n24185_), .A2(new_n13816_), .A3(pi1154), .A4(new_n24176_), .ZN(new_n24196_));
  AOI21_X1   g21012(.A1(new_n24195_), .A2(new_n24196_), .B(new_n24155_), .ZN(new_n24197_));
  NAND2_X1   g21013(.A1(new_n24190_), .A2(pi0618), .ZN(new_n24198_));
  NAND2_X1   g21014(.A1(new_n24198_), .A2(new_n13836_), .ZN(new_n24199_));
  OAI21_X1   g21015(.A1(new_n24197_), .A2(new_n24199_), .B(new_n13816_), .ZN(new_n24200_));
  NAND3_X1   g21016(.A1(new_n24194_), .A2(new_n24200_), .A3(pi0781), .ZN(new_n24201_));
  XOR2_X1    g21017(.A1(new_n24193_), .A2(new_n24201_), .Z(new_n24202_));
  NAND3_X1   g21018(.A1(new_n24186_), .A2(pi0618), .A3(pi1154), .ZN(new_n24203_));
  NAND3_X1   g21019(.A1(new_n24180_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n24204_));
  AOI21_X1   g21020(.A1(new_n24204_), .A2(new_n24203_), .B(new_n24155_), .ZN(new_n24205_));
  NAND4_X1   g21021(.A1(new_n24205_), .A2(new_n24197_), .A3(pi0781), .A4(new_n24186_), .ZN(new_n24206_));
  NOR2_X1    g21022(.A1(new_n24180_), .A2(new_n13855_), .ZN(new_n24207_));
  NAND2_X1   g21023(.A1(new_n24197_), .A2(new_n24207_), .ZN(new_n24208_));
  NAND3_X1   g21024(.A1(new_n24208_), .A2(pi0781), .A3(new_n24188_), .ZN(new_n24209_));
  NAND2_X1   g21025(.A1(new_n24209_), .A2(new_n24206_), .ZN(new_n24210_));
  NAND3_X1   g21026(.A1(new_n24210_), .A2(pi0619), .A3(pi1159), .ZN(new_n24211_));
  NAND4_X1   g21027(.A1(new_n24209_), .A2(pi0619), .A3(new_n13868_), .A4(new_n24206_), .ZN(new_n24212_));
  AOI21_X1   g21028(.A1(new_n24211_), .A2(new_n24212_), .B(new_n24155_), .ZN(new_n24213_));
  NOR2_X1    g21029(.A1(new_n24135_), .A2(new_n13880_), .ZN(new_n24214_));
  AOI21_X1   g21030(.A1(new_n24190_), .A2(new_n13880_), .B(new_n24214_), .ZN(new_n24215_));
  INV_X1     g21031(.I(new_n24215_), .ZN(new_n24216_));
  AOI21_X1   g21032(.A1(new_n24216_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n24217_));
  INV_X1     g21033(.I(new_n24217_), .ZN(new_n24218_));
  OAI21_X1   g21034(.A1(new_n24213_), .A2(new_n24218_), .B(new_n13860_), .ZN(new_n24219_));
  NAND3_X1   g21035(.A1(new_n24210_), .A2(pi0619), .A3(pi1159), .ZN(new_n24220_));
  NAND4_X1   g21036(.A1(new_n24209_), .A2(new_n13860_), .A3(pi1159), .A4(new_n24206_), .ZN(new_n24221_));
  AOI21_X1   g21037(.A1(new_n24220_), .A2(new_n24221_), .B(new_n24155_), .ZN(new_n24222_));
  AOI21_X1   g21038(.A1(new_n24216_), .A2(pi0619), .B(new_n15217_), .ZN(new_n24223_));
  INV_X1     g21039(.I(new_n24223_), .ZN(new_n24224_));
  OAI21_X1   g21040(.A1(new_n24222_), .A2(new_n24224_), .B(new_n13860_), .ZN(new_n24225_));
  NAND4_X1   g21041(.A1(new_n24219_), .A2(new_n24225_), .A3(pi0789), .A4(new_n24202_), .ZN(new_n24226_));
  NAND2_X1   g21042(.A1(new_n24219_), .A2(new_n24202_), .ZN(new_n24227_));
  NAND3_X1   g21043(.A1(new_n24225_), .A2(pi0789), .A3(new_n24202_), .ZN(new_n24228_));
  NAND3_X1   g21044(.A1(new_n24228_), .A2(new_n24227_), .A3(pi0789), .ZN(new_n24229_));
  NAND2_X1   g21045(.A1(new_n24229_), .A2(new_n24226_), .ZN(new_n24230_));
  NAND4_X1   g21046(.A1(new_n24213_), .A2(new_n24222_), .A3(pi0789), .A4(new_n24210_), .ZN(new_n24231_));
  AOI21_X1   g21047(.A1(new_n24180_), .A2(pi1154), .B(new_n13819_), .ZN(new_n24232_));
  INV_X1     g21048(.I(new_n24196_), .ZN(new_n24233_));
  OAI21_X1   g21049(.A1(new_n24232_), .A2(new_n24233_), .B(new_n24135_), .ZN(new_n24234_));
  NOR4_X1    g21050(.A1(new_n24188_), .A2(new_n24234_), .A3(new_n13855_), .A4(new_n24180_), .ZN(new_n24235_));
  NAND2_X1   g21051(.A1(new_n24188_), .A2(pi0781), .ZN(new_n24236_));
  NOR3_X1    g21052(.A1(new_n24234_), .A2(new_n13855_), .A3(new_n24180_), .ZN(new_n24237_));
  NOR2_X1    g21053(.A1(new_n24237_), .A2(new_n24236_), .ZN(new_n24238_));
  NOR2_X1    g21054(.A1(new_n24238_), .A2(new_n24235_), .ZN(new_n24239_));
  AOI21_X1   g21055(.A1(new_n24239_), .A2(pi0619), .B(new_n13904_), .ZN(new_n24240_));
  INV_X1     g21056(.I(new_n24212_), .ZN(new_n24241_));
  OAI21_X1   g21057(.A1(new_n24240_), .A2(new_n24241_), .B(new_n24135_), .ZN(new_n24242_));
  NOR2_X1    g21058(.A1(new_n24239_), .A2(new_n13896_), .ZN(new_n24243_));
  NAND2_X1   g21059(.A1(new_n24222_), .A2(new_n24243_), .ZN(new_n24244_));
  NAND3_X1   g21060(.A1(new_n24244_), .A2(pi0789), .A3(new_n24242_), .ZN(new_n24245_));
  NOR2_X1    g21061(.A1(new_n24155_), .A2(new_n13919_), .ZN(new_n24246_));
  AOI21_X1   g21062(.A1(new_n24215_), .A2(new_n13919_), .B(new_n24246_), .ZN(new_n24247_));
  NOR2_X1    g21063(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n24248_));
  INV_X1     g21064(.I(new_n24248_), .ZN(new_n24249_));
  AOI21_X1   g21065(.A1(new_n24245_), .A2(new_n24231_), .B(new_n24249_), .ZN(new_n24250_));
  AND3_X2    g21066(.A1(new_n24230_), .A2(pi0626), .A3(pi0788), .Z(new_n24254_));
  INV_X1     g21067(.I(new_n24231_), .ZN(new_n24255_));
  NAND2_X1   g21068(.A1(new_n24242_), .A2(pi0789), .ZN(new_n24256_));
  AOI21_X1   g21069(.A1(new_n24239_), .A2(pi1159), .B(new_n13904_), .ZN(new_n24257_));
  INV_X1     g21070(.I(new_n24221_), .ZN(new_n24258_));
  OAI21_X1   g21071(.A1(new_n24257_), .A2(new_n24258_), .B(new_n24135_), .ZN(new_n24259_));
  NOR3_X1    g21072(.A1(new_n24259_), .A2(new_n13896_), .A3(new_n24239_), .ZN(new_n24260_));
  NOR2_X1    g21073(.A1(new_n24260_), .A2(new_n24256_), .ZN(new_n24261_));
  OAI21_X1   g21074(.A1(new_n24261_), .A2(new_n24255_), .B(new_n24248_), .ZN(new_n24262_));
  AOI22_X1   g21075(.A1(new_n24262_), .A2(new_n13901_), .B1(new_n24226_), .B2(new_n24229_), .ZN(new_n24263_));
  AOI21_X1   g21076(.A1(new_n24229_), .A2(new_n24226_), .B(new_n15258_), .ZN(new_n24264_));
  NOR3_X1    g21077(.A1(new_n24263_), .A2(new_n13937_), .A3(new_n24264_), .ZN(new_n24265_));
  NOR2_X1    g21078(.A1(new_n24265_), .A2(new_n24254_), .ZN(new_n24266_));
  NAND2_X1   g21079(.A1(new_n24245_), .A2(new_n24231_), .ZN(new_n24267_));
  NOR2_X1    g21080(.A1(new_n24135_), .A2(new_n16372_), .ZN(new_n24268_));
  AOI21_X1   g21081(.A1(new_n24267_), .A2(new_n16372_), .B(new_n24268_), .ZN(new_n24269_));
  NOR2_X1    g21082(.A1(new_n24135_), .A2(new_n13966_), .ZN(new_n24271_));
  AOI21_X1   g21083(.A1(new_n24247_), .A2(new_n13966_), .B(new_n24271_), .ZN(new_n24272_));
  AOI21_X1   g21084(.A1(new_n24272_), .A2(pi0628), .B(new_n13971_), .ZN(new_n24273_));
  INV_X1     g21085(.I(new_n24272_), .ZN(new_n24274_));
  NOR3_X1    g21086(.A1(new_n24274_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n24275_));
  OAI21_X1   g21087(.A1(new_n24275_), .A2(new_n24273_), .B(new_n24135_), .ZN(new_n24276_));
  INV_X1     g21088(.I(new_n24276_), .ZN(new_n24277_));
  NOR2_X1    g21089(.A1(new_n24277_), .A2(new_n15270_), .ZN(new_n24278_));
  AOI21_X1   g21090(.A1(new_n24272_), .A2(pi1156), .B(new_n13971_), .ZN(new_n24281_));
  NOR3_X1    g21091(.A1(new_n24274_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n24282_));
  OAI21_X1   g21092(.A1(new_n24282_), .A2(new_n24281_), .B(new_n24135_), .ZN(new_n24283_));
  NOR3_X1    g21093(.A1(new_n24266_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n24286_));
  NAND3_X1   g21094(.A1(new_n24230_), .A2(pi0626), .A3(pi0788), .ZN(new_n24287_));
  INV_X1     g21095(.I(new_n24226_), .ZN(new_n24288_));
  INV_X1     g21096(.I(new_n24202_), .ZN(new_n24289_));
  AOI21_X1   g21097(.A1(new_n24242_), .A2(new_n24217_), .B(pi0619), .ZN(new_n24290_));
  OAI21_X1   g21098(.A1(new_n24290_), .A2(new_n24289_), .B(pi0789), .ZN(new_n24291_));
  AOI21_X1   g21099(.A1(new_n24259_), .A2(new_n24223_), .B(pi0619), .ZN(new_n24292_));
  INV_X1     g21100(.I(new_n24192_), .ZN(new_n24293_));
  AOI21_X1   g21101(.A1(new_n24194_), .A2(new_n24293_), .B(new_n13855_), .ZN(new_n24294_));
  NOR2_X1    g21102(.A1(new_n24294_), .A2(new_n24201_), .ZN(new_n24295_));
  NAND2_X1   g21103(.A1(new_n24294_), .A2(new_n24201_), .ZN(new_n24296_));
  INV_X1     g21104(.I(new_n24296_), .ZN(new_n24297_));
  OAI21_X1   g21105(.A1(new_n24297_), .A2(new_n24295_), .B(pi0789), .ZN(new_n24298_));
  NOR2_X1    g21106(.A1(new_n24292_), .A2(new_n24298_), .ZN(new_n24299_));
  NOR2_X1    g21107(.A1(new_n24291_), .A2(new_n24299_), .ZN(new_n24300_));
  OAI22_X1   g21108(.A1(new_n24300_), .A2(new_n24288_), .B1(pi0626), .B2(new_n24250_), .ZN(new_n24301_));
  OAI21_X1   g21109(.A1(new_n24300_), .A2(new_n24288_), .B(new_n14577_), .ZN(new_n24302_));
  NAND3_X1   g21110(.A1(new_n24301_), .A2(new_n24302_), .A3(pi0788), .ZN(new_n24303_));
  AOI21_X1   g21111(.A1(new_n24269_), .A2(new_n24278_), .B(pi0628), .ZN(new_n24304_));
  AOI21_X1   g21112(.A1(new_n24303_), .A2(new_n24287_), .B(new_n24304_), .ZN(new_n24305_));
  AOI21_X1   g21113(.A1(new_n24303_), .A2(new_n24287_), .B(new_n15296_), .ZN(new_n24306_));
  NOR3_X1    g21114(.A1(new_n24305_), .A2(new_n24306_), .A3(new_n12777_), .ZN(new_n24307_));
  NOR2_X1    g21115(.A1(new_n24307_), .A2(new_n24286_), .ZN(new_n24308_));
  NOR2_X1    g21116(.A1(new_n24135_), .A2(new_n13994_), .ZN(new_n24309_));
  INV_X1     g21117(.I(new_n24309_), .ZN(new_n24310_));
  OAI21_X1   g21118(.A1(new_n24269_), .A2(new_n13993_), .B(new_n24310_), .ZN(new_n24311_));
  NOR2_X1    g21119(.A1(new_n24277_), .A2(new_n12777_), .ZN(new_n24312_));
  NOR3_X1    g21120(.A1(new_n24283_), .A2(new_n12777_), .A3(new_n24272_), .ZN(new_n24313_));
  INV_X1     g21121(.I(new_n24313_), .ZN(new_n24314_));
  NOR2_X1    g21122(.A1(new_n24314_), .A2(new_n24312_), .ZN(new_n24315_));
  NAND2_X1   g21123(.A1(new_n24314_), .A2(new_n24312_), .ZN(new_n24316_));
  INV_X1     g21124(.I(new_n24316_), .ZN(new_n24317_));
  NOR2_X1    g21125(.A1(new_n24317_), .A2(new_n24315_), .ZN(new_n24318_));
  AOI21_X1   g21126(.A1(new_n24318_), .A2(pi0647), .B(new_n14008_), .ZN(new_n24319_));
  INV_X1     g21127(.I(new_n24315_), .ZN(new_n24320_));
  NAND2_X1   g21128(.A1(new_n24320_), .A2(new_n24316_), .ZN(new_n24321_));
  NOR3_X1    g21129(.A1(new_n24321_), .A2(new_n14005_), .A3(new_n14007_), .ZN(new_n24322_));
  OAI21_X1   g21130(.A1(new_n24322_), .A2(new_n24319_), .B(new_n24135_), .ZN(new_n24323_));
  NAND2_X1   g21131(.A1(new_n24323_), .A2(new_n14011_), .ZN(new_n24324_));
  OAI21_X1   g21132(.A1(new_n24324_), .A2(new_n24311_), .B(new_n14005_), .ZN(new_n24325_));
  INV_X1     g21133(.I(new_n24325_), .ZN(new_n24326_));
  AOI21_X1   g21134(.A1(new_n24318_), .A2(pi1157), .B(new_n14008_), .ZN(new_n24327_));
  NAND4_X1   g21135(.A1(new_n24320_), .A2(new_n24316_), .A3(new_n14005_), .A4(pi1157), .ZN(new_n24328_));
  INV_X1     g21136(.I(new_n24328_), .ZN(new_n24329_));
  OAI21_X1   g21137(.A1(new_n24327_), .A2(new_n24329_), .B(new_n24135_), .ZN(new_n24330_));
  NAND2_X1   g21138(.A1(new_n24330_), .A2(new_n14027_), .ZN(new_n24331_));
  AOI21_X1   g21139(.A1(pi0647), .A2(new_n24311_), .B(new_n24331_), .ZN(new_n24332_));
  NOR2_X1    g21140(.A1(new_n24332_), .A2(pi0647), .ZN(new_n24333_));
  NOR4_X1    g21141(.A1(new_n24308_), .A2(new_n12776_), .A3(new_n24326_), .A4(new_n24333_), .ZN(new_n24334_));
  NAND2_X1   g21142(.A1(new_n24303_), .A2(new_n24287_), .ZN(new_n24335_));
  NAND3_X1   g21143(.A1(new_n24335_), .A2(pi0628), .A3(pi0792), .ZN(new_n24336_));
  INV_X1     g21144(.I(new_n24304_), .ZN(new_n24337_));
  OAI21_X1   g21145(.A1(new_n24265_), .A2(new_n24254_), .B(new_n24337_), .ZN(new_n24338_));
  OAI21_X1   g21146(.A1(new_n24265_), .A2(new_n24254_), .B(new_n14606_), .ZN(new_n24339_));
  NAND3_X1   g21147(.A1(new_n24338_), .A2(new_n24339_), .A3(pi0792), .ZN(new_n24340_));
  AOI21_X1   g21148(.A1(new_n24340_), .A2(new_n24336_), .B(new_n24326_), .ZN(new_n24341_));
  OAI21_X1   g21149(.A1(new_n24332_), .A2(pi0647), .B(pi0787), .ZN(new_n24342_));
  AOI21_X1   g21150(.A1(new_n24340_), .A2(new_n24336_), .B(new_n24342_), .ZN(new_n24343_));
  NOR3_X1    g21151(.A1(new_n24343_), .A2(new_n24341_), .A3(new_n12776_), .ZN(new_n24344_));
  OAI21_X1   g21152(.A1(new_n24344_), .A2(new_n24334_), .B(new_n12775_), .ZN(new_n24345_));
  NAND2_X1   g21153(.A1(new_n24345_), .A2(new_n5787_), .ZN(new_n24346_));
  NAND2_X1   g21154(.A1(new_n24340_), .A2(new_n24336_), .ZN(new_n24347_));
  INV_X1     g21155(.I(new_n24333_), .ZN(new_n24348_));
  NAND4_X1   g21156(.A1(new_n24347_), .A2(pi0787), .A3(new_n24325_), .A4(new_n24348_), .ZN(new_n24349_));
  OAI21_X1   g21157(.A1(new_n24307_), .A2(new_n24286_), .B(new_n24325_), .ZN(new_n24350_));
  NAND2_X1   g21158(.A1(new_n24311_), .A2(pi0647), .ZN(new_n24351_));
  NAND3_X1   g21159(.A1(new_n24321_), .A2(pi0647), .A3(pi1157), .ZN(new_n24352_));
  NAND2_X1   g21160(.A1(new_n24352_), .A2(new_n24328_), .ZN(new_n24353_));
  AOI21_X1   g21161(.A1(new_n24353_), .A2(new_n24135_), .B(new_n16329_), .ZN(new_n24354_));
  NAND2_X1   g21162(.A1(new_n24351_), .A2(new_n24354_), .ZN(new_n24355_));
  AOI21_X1   g21163(.A1(new_n24355_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n24356_));
  OAI21_X1   g21164(.A1(new_n24307_), .A2(new_n24286_), .B(new_n24356_), .ZN(new_n24357_));
  NAND3_X1   g21165(.A1(new_n24350_), .A2(new_n24357_), .A3(pi0787), .ZN(new_n24358_));
  NAND2_X1   g21166(.A1(new_n24358_), .A2(new_n24349_), .ZN(new_n24359_));
  NOR4_X1    g21167(.A1(new_n24323_), .A2(new_n24330_), .A3(new_n12776_), .A4(new_n24318_), .ZN(new_n24360_));
  NAND2_X1   g21168(.A1(new_n24323_), .A2(pi0787), .ZN(new_n24361_));
  NOR3_X1    g21169(.A1(new_n24330_), .A2(new_n12776_), .A3(new_n24318_), .ZN(new_n24362_));
  NOR2_X1    g21170(.A1(new_n24362_), .A2(new_n24361_), .ZN(new_n24363_));
  OR2_X2     g21171(.A1(new_n24363_), .A2(new_n24360_), .Z(new_n24364_));
  NAND2_X1   g21172(.A1(new_n24135_), .A2(new_n14210_), .ZN(new_n24365_));
  OAI21_X1   g21173(.A1(new_n24311_), .A2(new_n14210_), .B(new_n24365_), .ZN(new_n24366_));
  NOR2_X1    g21174(.A1(new_n14204_), .A2(new_n14200_), .ZN(new_n24367_));
  NAND2_X1   g21175(.A1(new_n24366_), .A2(new_n24367_), .ZN(new_n24368_));
  OAI21_X1   g21176(.A1(new_n24364_), .A2(new_n24368_), .B(new_n14204_), .ZN(new_n24369_));
  AOI21_X1   g21177(.A1(new_n24359_), .A2(new_n24369_), .B(pi0790), .ZN(new_n24370_));
  OAI21_X1   g21178(.A1(new_n24363_), .A2(new_n24360_), .B(pi0644), .ZN(new_n24371_));
  NOR2_X1    g21179(.A1(new_n14204_), .A2(pi0715), .ZN(new_n24372_));
  NAND3_X1   g21180(.A1(new_n24371_), .A2(new_n24366_), .A3(new_n24372_), .ZN(new_n24373_));
  NAND2_X1   g21181(.A1(new_n5788_), .A2(new_n8642_), .ZN(new_n24374_));
  NOR2_X1    g21182(.A1(new_n13105_), .A2(new_n17845_), .ZN(new_n24375_));
  INV_X1     g21183(.I(new_n24375_), .ZN(new_n24376_));
  NOR2_X1    g21184(.A1(new_n24376_), .A2(new_n16376_), .ZN(new_n24377_));
  INV_X1     g21185(.I(new_n24377_), .ZN(new_n24378_));
  NOR2_X1    g21186(.A1(new_n16388_), .A2(new_n24378_), .ZN(new_n24379_));
  NOR2_X1    g21187(.A1(new_n9992_), .A2(new_n8642_), .ZN(new_n24380_));
  NOR2_X1    g21188(.A1(new_n24380_), .A2(pi0715), .ZN(new_n24381_));
  NOR4_X1    g21189(.A1(new_n18968_), .A2(new_n14204_), .A3(new_n16372_), .A4(new_n24381_), .ZN(new_n24382_));
  NAND2_X1   g21190(.A1(new_n24379_), .A2(new_n24382_), .ZN(new_n24383_));
  NOR2_X1    g21191(.A1(new_n13219_), .A2(new_n17866_), .ZN(new_n24384_));
  INV_X1     g21192(.I(new_n24380_), .ZN(new_n24385_));
  AOI21_X1   g21193(.A1(new_n24385_), .A2(new_n13614_), .B(new_n13613_), .ZN(new_n24386_));
  AOI21_X1   g21194(.A1(new_n24386_), .A2(new_n24384_), .B(new_n13748_), .ZN(new_n24387_));
  NOR4_X1    g21195(.A1(new_n13219_), .A2(new_n13613_), .A3(new_n17866_), .A4(new_n13614_), .ZN(new_n24388_));
  NOR4_X1    g21196(.A1(new_n13219_), .A2(pi0625), .A3(new_n17866_), .A4(pi1153), .ZN(new_n24389_));
  OAI21_X1   g21197(.A1(new_n24388_), .A2(new_n24389_), .B(new_n24380_), .ZN(new_n24390_));
  NOR4_X1    g21198(.A1(new_n24390_), .A2(new_n13748_), .A3(new_n24380_), .A4(new_n24384_), .ZN(new_n24391_));
  XNOR2_X1   g21199(.A1(new_n24391_), .A2(new_n24387_), .ZN(new_n24392_));
  NOR2_X1    g21200(.A1(new_n24392_), .A2(new_n15396_), .ZN(new_n24393_));
  INV_X1     g21201(.I(new_n24393_), .ZN(new_n24394_));
  NOR2_X1    g21202(.A1(new_n24394_), .A2(new_n14058_), .ZN(new_n24395_));
  AOI21_X1   g21203(.A1(new_n24395_), .A2(new_n15402_), .B(new_n24380_), .ZN(new_n24396_));
  NOR2_X1    g21204(.A1(new_n16435_), .A2(new_n17866_), .ZN(new_n24397_));
  NAND4_X1   g21205(.A1(new_n24397_), .A2(pi1153), .A3(new_n24375_), .A4(new_n24380_), .ZN(new_n24398_));
  NAND3_X1   g21206(.A1(new_n24398_), .A2(pi0608), .A3(new_n24390_), .ZN(new_n24399_));
  NAND2_X1   g21207(.A1(new_n24399_), .A2(pi0778), .ZN(new_n24400_));
  NOR2_X1    g21208(.A1(new_n24400_), .A2(pi0785), .ZN(new_n24401_));
  NAND2_X1   g21209(.A1(new_n24400_), .A2(pi1155), .ZN(new_n24402_));
  XOR2_X1    g21210(.A1(new_n24402_), .A2(new_n14090_), .Z(new_n24403_));
  NOR2_X1    g21211(.A1(new_n24380_), .A2(pi1155), .ZN(new_n24404_));
  NOR2_X1    g21212(.A1(new_n16444_), .A2(new_n24404_), .ZN(new_n24405_));
  AOI21_X1   g21213(.A1(new_n24405_), .A2(new_n24375_), .B(new_n13783_), .ZN(new_n24406_));
  OAI21_X1   g21214(.A1(new_n24403_), .A2(new_n24392_), .B(new_n24406_), .ZN(new_n24407_));
  NOR2_X1    g21215(.A1(new_n14102_), .A2(new_n24404_), .ZN(new_n24408_));
  AOI21_X1   g21216(.A1(new_n24408_), .A2(new_n24375_), .B(pi0660), .ZN(new_n24409_));
  INV_X1     g21217(.I(new_n24392_), .ZN(new_n24410_));
  NAND2_X1   g21218(.A1(new_n24400_), .A2(pi0609), .ZN(new_n24411_));
  XOR2_X1    g21219(.A1(new_n24411_), .A2(new_n14694_), .Z(new_n24412_));
  NAND3_X1   g21220(.A1(new_n24412_), .A2(pi0785), .A3(new_n24410_), .ZN(new_n24413_));
  AOI21_X1   g21221(.A1(new_n24407_), .A2(new_n24409_), .B(new_n24413_), .ZN(new_n24414_));
  NOR2_X1    g21222(.A1(new_n24414_), .A2(new_n24401_), .ZN(new_n24415_));
  AOI21_X1   g21223(.A1(new_n24410_), .A2(new_n13805_), .B(new_n24380_), .ZN(new_n24416_));
  INV_X1     g21224(.I(new_n24416_), .ZN(new_n24417_));
  NAND2_X1   g21225(.A1(new_n24415_), .A2(pi0618), .ZN(new_n24418_));
  XOR2_X1    g21226(.A1(new_n24418_), .A2(new_n13818_), .Z(new_n24419_));
  NOR2_X1    g21227(.A1(new_n24380_), .A2(pi1154), .ZN(new_n24420_));
  NOR2_X1    g21228(.A1(new_n16464_), .A2(new_n24420_), .ZN(new_n24421_));
  AOI21_X1   g21229(.A1(new_n24377_), .A2(new_n24421_), .B(pi0627), .ZN(new_n24422_));
  OAI21_X1   g21230(.A1(new_n24419_), .A2(new_n24417_), .B(new_n24422_), .ZN(new_n24423_));
  NOR2_X1    g21231(.A1(new_n16460_), .A2(new_n24420_), .ZN(new_n24424_));
  AOI21_X1   g21232(.A1(new_n24377_), .A2(new_n24424_), .B(pi0627), .ZN(new_n24425_));
  NAND2_X1   g21233(.A1(new_n24423_), .A2(new_n24425_), .ZN(new_n24426_));
  NAND2_X1   g21234(.A1(new_n24415_), .A2(pi1154), .ZN(new_n24427_));
  XOR2_X1    g21235(.A1(new_n24427_), .A2(new_n13818_), .Z(new_n24428_));
  NOR2_X1    g21236(.A1(new_n24428_), .A2(new_n24417_), .ZN(new_n24429_));
  AOI21_X1   g21237(.A1(new_n24426_), .A2(new_n24429_), .B(new_n13855_), .ZN(new_n24430_));
  XOR2_X1    g21238(.A1(new_n24430_), .A2(new_n18857_), .Z(new_n24431_));
  NAND2_X1   g21239(.A1(new_n24410_), .A2(new_n15437_), .ZN(new_n24432_));
  OAI21_X1   g21240(.A1(new_n24432_), .A2(new_n13918_), .B(new_n24385_), .ZN(new_n24433_));
  NAND3_X1   g21241(.A1(new_n13901_), .A2(pi0641), .A3(pi1158), .ZN(new_n24434_));
  OAI21_X1   g21242(.A1(new_n24433_), .A2(new_n24434_), .B(new_n18862_), .ZN(new_n24435_));
  AOI21_X1   g21243(.A1(new_n24380_), .A2(pi1158), .B(pi0626), .ZN(new_n24436_));
  NOR3_X1    g21244(.A1(new_n16388_), .A2(new_n24378_), .A3(new_n24436_), .ZN(new_n24437_));
  OAI21_X1   g21245(.A1(new_n24437_), .A2(pi0641), .B(new_n14140_), .ZN(new_n24438_));
  NOR2_X1    g21246(.A1(new_n24433_), .A2(new_n24438_), .ZN(new_n24439_));
  NOR2_X1    g21247(.A1(new_n24378_), .A2(new_n18869_), .ZN(new_n24440_));
  OAI21_X1   g21248(.A1(new_n24378_), .A2(new_n16476_), .B(new_n13915_), .ZN(new_n24441_));
  XNOR2_X1   g21249(.A1(new_n24441_), .A2(new_n24440_), .ZN(new_n24442_));
  NAND2_X1   g21250(.A1(new_n24385_), .A2(new_n13896_), .ZN(new_n24443_));
  NAND4_X1   g21251(.A1(new_n24442_), .A2(new_n16697_), .A3(new_n18868_), .A4(new_n24443_), .ZN(new_n24444_));
  OAI21_X1   g21252(.A1(new_n24444_), .A2(new_n24432_), .B(new_n15479_), .ZN(new_n24445_));
  AOI21_X1   g21253(.A1(new_n24435_), .A2(new_n24439_), .B(new_n24445_), .ZN(new_n24446_));
  NOR3_X1    g21254(.A1(new_n24431_), .A2(new_n24415_), .A3(new_n24446_), .ZN(new_n24447_));
  NAND2_X1   g21255(.A1(new_n24379_), .A2(new_n16372_), .ZN(new_n24448_));
  NAND2_X1   g21256(.A1(new_n24448_), .A2(new_n14010_), .ZN(new_n24449_));
  NOR2_X1    g21257(.A1(new_n24449_), .A2(pi0647), .ZN(new_n24450_));
  OAI21_X1   g21258(.A1(new_n24450_), .A2(new_n18879_), .B(new_n14010_), .ZN(new_n24451_));
  NOR2_X1    g21259(.A1(new_n24449_), .A2(pi1157), .ZN(new_n24452_));
  OAI22_X1   g21260(.A1(new_n24452_), .A2(new_n18882_), .B1(new_n14058_), .B2(new_n24394_), .ZN(new_n24453_));
  AND3_X2    g21261(.A1(new_n16418_), .A2(pi0630), .A3(pi0787), .Z(new_n24454_));
  AND4_X2    g21262(.A1(new_n24395_), .A2(new_n24453_), .A3(new_n24451_), .A4(new_n24454_), .Z(new_n24455_));
  AOI21_X1   g21263(.A1(new_n24448_), .A2(new_n13970_), .B(pi0629), .ZN(new_n24456_));
  NAND2_X1   g21264(.A1(new_n24448_), .A2(new_n13942_), .ZN(new_n24457_));
  AOI21_X1   g21265(.A1(new_n24457_), .A2(pi0629), .B(pi1156), .ZN(new_n24458_));
  OAI21_X1   g21266(.A1(new_n24380_), .A2(pi0792), .B(pi0628), .ZN(new_n24459_));
  NOR4_X1    g21267(.A1(new_n24458_), .A2(new_n24394_), .A3(new_n24456_), .A4(new_n24459_), .ZN(new_n24460_));
  OAI21_X1   g21268(.A1(new_n24447_), .A2(new_n24455_), .B(new_n24460_), .ZN(new_n24461_));
  NAND2_X1   g21269(.A1(new_n24461_), .A2(pi0644), .ZN(new_n24462_));
  XOR2_X1    g21270(.A1(new_n24462_), .A2(new_n14217_), .Z(new_n24463_));
  NAND4_X1   g21271(.A1(new_n24463_), .A2(new_n14203_), .A3(new_n24383_), .A4(new_n24396_), .ZN(new_n24464_));
  INV_X1     g21272(.I(new_n24396_), .ZN(new_n24465_));
  NAND2_X1   g21273(.A1(new_n24461_), .A2(pi0715), .ZN(new_n24466_));
  XOR2_X1    g21274(.A1(new_n24466_), .A2(new_n14205_), .Z(new_n24467_));
  NOR2_X1    g21275(.A1(new_n24467_), .A2(new_n24465_), .ZN(new_n24468_));
  AOI21_X1   g21276(.A1(new_n24464_), .A2(new_n24468_), .B(new_n14799_), .ZN(new_n24469_));
  XOR2_X1    g21277(.A1(new_n24469_), .A2(new_n14800_), .Z(new_n24470_));
  OAI21_X1   g21278(.A1(new_n5371_), .A2(new_n8642_), .B(new_n14799_), .ZN(new_n24471_));
  NOR2_X1    g21279(.A1(new_n24461_), .A2(new_n24471_), .ZN(new_n24472_));
  AOI22_X1   g21280(.A1(new_n24470_), .A2(new_n24472_), .B1(new_n5371_), .B2(new_n24374_), .ZN(new_n24473_));
  AOI21_X1   g21281(.A1(new_n24373_), .A2(new_n14204_), .B(new_n24473_), .ZN(new_n24474_));
  NAND2_X1   g21282(.A1(new_n24359_), .A2(new_n24474_), .ZN(new_n24475_));
  AOI21_X1   g21283(.A1(new_n24346_), .A2(new_n24370_), .B(new_n24475_), .ZN(po0346));
  NOR2_X1    g21284(.A1(new_n14652_), .A2(new_n17943_), .ZN(new_n24477_));
  INV_X1     g21285(.I(new_n24477_), .ZN(new_n24478_));
  NOR2_X1    g21286(.A1(new_n9992_), .A2(pi0190), .ZN(new_n24479_));
  NOR2_X1    g21287(.A1(new_n24479_), .A2(pi1153), .ZN(new_n24480_));
  NAND2_X1   g21288(.A1(new_n24478_), .A2(new_n24480_), .ZN(new_n24481_));
  INV_X1     g21289(.I(new_n24481_), .ZN(new_n24482_));
  NOR2_X1    g21290(.A1(new_n24482_), .A2(new_n13748_), .ZN(new_n24483_));
  AOI21_X1   g21291(.A1(new_n13218_), .A2(pi0699), .B(new_n24479_), .ZN(new_n24484_));
  INV_X1     g21292(.I(new_n24484_), .ZN(new_n24485_));
  AOI21_X1   g21293(.A1(new_n24478_), .A2(new_n24485_), .B(new_n13614_), .ZN(new_n24486_));
  INV_X1     g21294(.I(new_n24486_), .ZN(new_n24487_));
  NOR3_X1    g21295(.A1(new_n24487_), .A2(new_n13748_), .A3(new_n24485_), .ZN(new_n24488_));
  XNOR2_X1   g21296(.A1(new_n24488_), .A2(new_n24483_), .ZN(new_n24489_));
  NAND2_X1   g21297(.A1(new_n24489_), .A2(new_n14049_), .ZN(new_n24490_));
  NOR2_X1    g21298(.A1(new_n24490_), .A2(new_n14051_), .ZN(new_n24491_));
  INV_X1     g21299(.I(new_n24491_), .ZN(new_n24492_));
  NOR2_X1    g21300(.A1(new_n24492_), .A2(new_n14163_), .ZN(new_n24493_));
  NAND2_X1   g21301(.A1(new_n24493_), .A2(new_n18929_), .ZN(new_n24494_));
  NOR2_X1    g21302(.A1(new_n24494_), .A2(new_n14060_), .ZN(new_n24495_));
  INV_X1     g21303(.I(new_n24479_), .ZN(new_n24496_));
  NAND3_X1   g21304(.A1(new_n24495_), .A2(pi0647), .A3(pi1157), .ZN(new_n24497_));
  OR3_X2     g21305(.A1(new_n24495_), .A2(new_n14005_), .A3(pi1157), .Z(new_n24498_));
  AOI21_X1   g21306(.A1(new_n24498_), .A2(new_n24497_), .B(new_n24496_), .ZN(new_n24499_));
  INV_X1     g21307(.I(new_n24499_), .ZN(new_n24500_));
  NOR2_X1    g21308(.A1(new_n24496_), .A2(pi0647), .ZN(new_n24501_));
  AOI21_X1   g21309(.A1(new_n24495_), .A2(pi0647), .B(new_n24501_), .ZN(new_n24502_));
  AOI21_X1   g21310(.A1(new_n24502_), .A2(pi1157), .B(new_n12776_), .ZN(new_n24503_));
  AOI22_X1   g21311(.A1(new_n24500_), .A2(new_n24503_), .B1(new_n12776_), .B2(new_n24495_), .ZN(new_n24504_));
  INV_X1     g21312(.I(new_n24504_), .ZN(new_n24505_));
  NOR2_X1    g21313(.A1(new_n13105_), .A2(new_n17912_), .ZN(new_n24506_));
  INV_X1     g21314(.I(new_n24506_), .ZN(new_n24507_));
  NOR2_X1    g21315(.A1(new_n24506_), .A2(new_n24479_), .ZN(new_n24508_));
  INV_X1     g21316(.I(new_n24508_), .ZN(new_n24509_));
  NAND3_X1   g21317(.A1(new_n24509_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n24510_));
  AOI21_X1   g21318(.A1(new_n24510_), .A2(new_n16444_), .B(new_n24507_), .ZN(new_n24511_));
  NOR2_X1    g21319(.A1(new_n24511_), .A2(new_n13801_), .ZN(new_n24512_));
  NOR2_X1    g21320(.A1(new_n24479_), .A2(pi1155), .ZN(new_n24513_));
  NOR3_X1    g21321(.A1(new_n24507_), .A2(new_n16444_), .A3(new_n24513_), .ZN(new_n24514_));
  NAND4_X1   g21322(.A1(new_n24514_), .A2(new_n24509_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n24515_));
  XOR2_X1    g21323(.A1(new_n24512_), .A2(new_n24515_), .Z(new_n24516_));
  NOR2_X1    g21324(.A1(new_n24516_), .A2(new_n13817_), .ZN(new_n24517_));
  OAI21_X1   g21325(.A1(new_n24517_), .A2(pi0618), .B(new_n9992_), .ZN(new_n24518_));
  NAND2_X1   g21326(.A1(new_n24518_), .A2(pi0781), .ZN(new_n24519_));
  OAI21_X1   g21327(.A1(new_n24517_), .A2(new_n9992_), .B(pi0618), .ZN(new_n24520_));
  NOR3_X1    g21328(.A1(new_n24520_), .A2(new_n13855_), .A3(new_n24516_), .ZN(new_n24521_));
  XOR2_X1    g21329(.A1(new_n24521_), .A2(new_n24519_), .Z(new_n24522_));
  NOR2_X1    g21330(.A1(new_n24522_), .A2(new_n13868_), .ZN(new_n24523_));
  OAI21_X1   g21331(.A1(new_n24523_), .A2(pi0619), .B(new_n9992_), .ZN(new_n24524_));
  NAND2_X1   g21332(.A1(new_n24524_), .A2(pi0789), .ZN(new_n24525_));
  OAI21_X1   g21333(.A1(new_n24523_), .A2(new_n9992_), .B(pi0619), .ZN(new_n24526_));
  NOR3_X1    g21334(.A1(new_n24526_), .A2(new_n13896_), .A3(new_n24522_), .ZN(new_n24527_));
  XOR2_X1    g21335(.A1(new_n24527_), .A2(new_n24525_), .Z(new_n24528_));
  NAND2_X1   g21336(.A1(new_n24528_), .A2(new_n16372_), .ZN(new_n24529_));
  OAI21_X1   g21337(.A1(new_n16372_), .A2(new_n24479_), .B(new_n24529_), .ZN(new_n24530_));
  NOR2_X1    g21338(.A1(new_n24530_), .A2(new_n18968_), .ZN(new_n24531_));
  NAND2_X1   g21339(.A1(new_n18967_), .A2(new_n24479_), .ZN(new_n24532_));
  XOR2_X1    g21340(.A1(new_n24531_), .A2(new_n24532_), .Z(new_n24533_));
  AOI21_X1   g21341(.A1(new_n24496_), .A2(new_n14254_), .B(pi0644), .ZN(new_n24534_));
  NAND2_X1   g21342(.A1(new_n24528_), .A2(new_n13962_), .ZN(new_n24535_));
  XOR2_X1    g21343(.A1(new_n24535_), .A2(new_n18976_), .Z(new_n24536_));
  AOI22_X1   g21344(.A1(new_n24536_), .A2(new_n24479_), .B1(new_n16639_), .B2(new_n24493_), .ZN(new_n24537_));
  NOR2_X1    g21345(.A1(new_n24484_), .A2(new_n13203_), .ZN(new_n24538_));
  NAND2_X1   g21346(.A1(new_n24538_), .A2(pi0625), .ZN(new_n24539_));
  NAND3_X1   g21347(.A1(new_n24539_), .A2(pi1153), .A3(new_n24508_), .ZN(new_n24540_));
  NOR2_X1    g21348(.A1(new_n24482_), .A2(new_n14081_), .ZN(new_n24541_));
  AOI21_X1   g21349(.A1(new_n24541_), .A2(new_n24540_), .B(new_n13748_), .ZN(new_n24542_));
  NOR2_X1    g21350(.A1(new_n24509_), .A2(new_n24538_), .ZN(new_n24543_));
  INV_X1     g21351(.I(new_n24539_), .ZN(new_n24544_));
  OAI21_X1   g21352(.A1(new_n24543_), .A2(new_n24544_), .B(new_n24480_), .ZN(new_n24545_));
  NAND4_X1   g21353(.A1(new_n24545_), .A2(new_n13749_), .A3(new_n24487_), .A4(new_n24543_), .ZN(new_n24546_));
  XNOR2_X1   g21354(.A1(new_n24546_), .A2(new_n24542_), .ZN(new_n24547_));
  NAND2_X1   g21355(.A1(new_n24547_), .A2(new_n13801_), .ZN(new_n24548_));
  NOR2_X1    g21356(.A1(new_n24511_), .A2(pi0660), .ZN(new_n24551_));
  NOR2_X1    g21357(.A1(new_n24547_), .A2(new_n13766_), .ZN(new_n24552_));
  XOR2_X1    g21358(.A1(new_n24552_), .A2(new_n14090_), .Z(new_n24553_));
  NOR2_X1    g21359(.A1(new_n24489_), .A2(new_n13801_), .ZN(new_n24554_));
  NAND2_X1   g21360(.A1(new_n24553_), .A2(new_n24554_), .ZN(new_n24555_));
  OAI21_X1   g21361(.A1(new_n24555_), .A2(new_n24551_), .B(new_n24548_), .ZN(new_n24556_));
  NAND2_X1   g21362(.A1(new_n24556_), .A2(new_n13855_), .ZN(new_n24557_));
  INV_X1     g21363(.I(new_n24490_), .ZN(new_n24558_));
  NOR2_X1    g21364(.A1(new_n24556_), .A2(new_n13816_), .ZN(new_n24559_));
  XOR2_X1    g21365(.A1(new_n24559_), .A2(new_n13818_), .Z(new_n24560_));
  NAND2_X1   g21366(.A1(new_n24560_), .A2(new_n24558_), .ZN(new_n24561_));
  NAND3_X1   g21367(.A1(new_n24561_), .A2(new_n13823_), .A3(new_n24520_), .ZN(new_n24562_));
  NAND3_X1   g21368(.A1(new_n24562_), .A2(new_n13823_), .A3(new_n24518_), .ZN(new_n24563_));
  NOR2_X1    g21369(.A1(new_n24556_), .A2(new_n13817_), .ZN(new_n24564_));
  XOR2_X1    g21370(.A1(new_n24564_), .A2(new_n13818_), .Z(new_n24565_));
  NAND4_X1   g21371(.A1(new_n24563_), .A2(pi0781), .A3(new_n24558_), .A4(new_n24565_), .ZN(new_n24566_));
  NAND2_X1   g21372(.A1(new_n24566_), .A2(new_n24557_), .ZN(new_n24567_));
  NOR2_X1    g21373(.A1(new_n24567_), .A2(new_n13860_), .ZN(new_n24568_));
  XOR2_X1    g21374(.A1(new_n24568_), .A2(new_n13904_), .Z(new_n24569_));
  NOR2_X1    g21375(.A1(new_n24569_), .A2(new_n24492_), .ZN(new_n24570_));
  NAND2_X1   g21376(.A1(new_n24526_), .A2(new_n13884_), .ZN(new_n24571_));
  INV_X1     g21377(.I(new_n24567_), .ZN(new_n24572_));
  AOI21_X1   g21378(.A1(new_n24572_), .A2(new_n14143_), .B(pi0789), .ZN(new_n24573_));
  OAI21_X1   g21379(.A1(new_n24570_), .A2(new_n24571_), .B(new_n24573_), .ZN(new_n24574_));
  NOR2_X1    g21380(.A1(new_n24567_), .A2(new_n13868_), .ZN(new_n24575_));
  XOR2_X1    g21381(.A1(new_n24575_), .A2(new_n13903_), .Z(new_n24576_));
  NAND2_X1   g21382(.A1(new_n24524_), .A2(new_n19018_), .ZN(new_n24577_));
  AOI21_X1   g21383(.A1(new_n24576_), .A2(new_n24491_), .B(new_n24577_), .ZN(new_n24578_));
  AOI21_X1   g21384(.A1(new_n24574_), .A2(new_n24578_), .B(new_n24537_), .ZN(new_n24579_));
  NAND3_X1   g21385(.A1(new_n24530_), .A2(new_n18929_), .A3(new_n24493_), .ZN(new_n24580_));
  NAND2_X1   g21386(.A1(new_n24580_), .A2(new_n16569_), .ZN(new_n24581_));
  XOR2_X1    g21387(.A1(new_n24581_), .A2(new_n16572_), .Z(new_n24582_));
  AOI21_X1   g21388(.A1(new_n19022_), .A2(new_n24580_), .B(new_n24582_), .ZN(new_n24583_));
  NAND2_X1   g21389(.A1(new_n24528_), .A2(new_n13963_), .ZN(new_n24584_));
  XNOR2_X1   g21390(.A1(new_n24584_), .A2(new_n19028_), .ZN(new_n24585_));
  NOR3_X1    g21391(.A1(new_n24585_), .A2(new_n16424_), .A3(new_n24496_), .ZN(new_n24586_));
  OAI21_X1   g21392(.A1(new_n24583_), .A2(new_n16574_), .B(new_n24586_), .ZN(new_n24587_));
  NOR2_X1    g21393(.A1(new_n24530_), .A2(new_n13994_), .ZN(new_n24588_));
  XNOR2_X1   g21394(.A1(new_n24588_), .A2(new_n19033_), .ZN(new_n24589_));
  AOI22_X1   g21395(.A1(new_n24589_), .A2(new_n24479_), .B1(new_n14206_), .B2(new_n24502_), .ZN(new_n24590_));
  NOR3_X1    g21396(.A1(new_n24590_), .A2(new_n14010_), .A3(new_n24500_), .ZN(new_n24591_));
  OAI22_X1   g21397(.A1(new_n24579_), .A2(new_n24587_), .B1(new_n12776_), .B2(new_n24591_), .ZN(new_n24592_));
  NAND2_X1   g21398(.A1(new_n24592_), .A2(pi0644), .ZN(new_n24593_));
  XOR2_X1    g21399(.A1(new_n24593_), .A2(new_n14205_), .Z(new_n24594_));
  NOR2_X1    g21400(.A1(new_n24594_), .A2(new_n24504_), .ZN(new_n24595_));
  NAND2_X1   g21401(.A1(new_n24533_), .A2(pi0715), .ZN(new_n24596_));
  XOR2_X1    g21402(.A1(new_n24596_), .A2(new_n14205_), .Z(new_n24597_));
  OAI21_X1   g21403(.A1(new_n24597_), .A2(new_n24496_), .B(new_n19043_), .ZN(new_n24598_));
  OAI22_X1   g21404(.A1(new_n24595_), .A2(new_n24598_), .B1(new_n24533_), .B2(new_n24534_), .ZN(new_n24599_));
  NAND2_X1   g21405(.A1(new_n24592_), .A2(pi0715), .ZN(new_n24600_));
  XOR2_X1    g21406(.A1(new_n24600_), .A2(new_n14217_), .Z(new_n24601_));
  AOI21_X1   g21407(.A1(po1038), .A2(new_n10656_), .B(pi0832), .ZN(new_n24602_));
  NAND4_X1   g21408(.A1(new_n24599_), .A2(new_n24505_), .A3(new_n24601_), .A4(new_n24602_), .ZN(new_n24603_));
  NOR2_X1    g21409(.A1(new_n14428_), .A2(pi0190), .ZN(new_n24604_));
  INV_X1     g21410(.I(new_n24604_), .ZN(new_n24605_));
  OAI22_X1   g21411(.A1(new_n17127_), .A2(new_n10656_), .B1(new_n17912_), .B2(new_n19052_), .ZN(new_n24606_));
  OAI21_X1   g21412(.A1(pi0190), .A2(new_n14299_), .B(new_n14301_), .ZN(new_n24607_));
  NAND2_X1   g21413(.A1(new_n14299_), .A2(pi0763), .ZN(new_n24608_));
  NAND4_X1   g21414(.A1(new_n24607_), .A2(new_n17912_), .A3(new_n14362_), .A4(new_n24608_), .ZN(new_n24609_));
  NAND3_X1   g21415(.A1(new_n24609_), .A2(pi0038), .A3(pi0190), .ZN(new_n24610_));
  NAND2_X1   g21416(.A1(new_n24610_), .A2(new_n3183_), .ZN(new_n24611_));
  NAND2_X1   g21417(.A1(new_n13109_), .A2(new_n10656_), .ZN(new_n24612_));
  NAND4_X1   g21418(.A1(new_n24611_), .A2(pi0038), .A3(new_n24606_), .A4(new_n24612_), .ZN(new_n24613_));
  AOI21_X1   g21419(.A1(new_n24613_), .A2(new_n17912_), .B(new_n13107_), .ZN(new_n24614_));
  NAND2_X1   g21420(.A1(new_n24614_), .A2(new_n3289_), .ZN(new_n24615_));
  NAND2_X1   g21421(.A1(new_n3290_), .A2(new_n10656_), .ZN(new_n24616_));
  NAND3_X1   g21422(.A1(new_n24615_), .A2(new_n13776_), .A3(new_n24616_), .ZN(new_n24617_));
  NAND2_X1   g21423(.A1(new_n24605_), .A2(new_n13780_), .ZN(new_n24618_));
  NAND2_X1   g21424(.A1(new_n24617_), .A2(new_n24618_), .ZN(new_n24619_));
  NAND2_X1   g21425(.A1(new_n24619_), .A2(pi0609), .ZN(new_n24620_));
  NAND2_X1   g21426(.A1(new_n24620_), .A2(pi0785), .ZN(new_n24621_));
  NAND2_X1   g21427(.A1(new_n24615_), .A2(new_n24616_), .ZN(new_n24622_));
  NOR2_X1    g21428(.A1(new_n24605_), .A2(new_n13776_), .ZN(new_n24623_));
  AOI21_X1   g21429(.A1(new_n24622_), .A2(new_n13776_), .B(new_n24623_), .ZN(new_n24624_));
  AOI21_X1   g21430(.A1(new_n24605_), .A2(new_n14467_), .B(pi0609), .ZN(new_n24625_));
  OR2_X2     g21431(.A1(new_n24617_), .A2(new_n24625_), .Z(new_n24626_));
  NOR3_X1    g21432(.A1(new_n24626_), .A2(new_n13801_), .A3(new_n24624_), .ZN(new_n24627_));
  XNOR2_X1   g21433(.A1(new_n24627_), .A2(new_n24621_), .ZN(new_n24628_));
  NAND3_X1   g21434(.A1(new_n24628_), .A2(pi0618), .A3(pi1154), .ZN(new_n24629_));
  XOR2_X1    g21435(.A1(new_n24627_), .A2(new_n24621_), .Z(new_n24630_));
  NAND3_X1   g21436(.A1(new_n24630_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n24631_));
  NAND2_X1   g21437(.A1(new_n24629_), .A2(new_n24631_), .ZN(new_n24632_));
  NAND2_X1   g21438(.A1(new_n24632_), .A2(new_n24604_), .ZN(new_n24633_));
  NAND2_X1   g21439(.A1(new_n24633_), .A2(pi0781), .ZN(new_n24634_));
  NAND3_X1   g21440(.A1(new_n24628_), .A2(pi0618), .A3(pi1154), .ZN(new_n24635_));
  NAND3_X1   g21441(.A1(new_n24630_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n24636_));
  AOI21_X1   g21442(.A1(new_n24635_), .A2(new_n24636_), .B(new_n24605_), .ZN(new_n24637_));
  NOR2_X1    g21443(.A1(new_n24630_), .A2(new_n13855_), .ZN(new_n24638_));
  NAND3_X1   g21444(.A1(new_n24634_), .A2(new_n24637_), .A3(new_n24638_), .ZN(new_n24639_));
  NAND2_X1   g21445(.A1(new_n24637_), .A2(new_n24638_), .ZN(new_n24640_));
  NAND3_X1   g21446(.A1(new_n24640_), .A2(new_n24633_), .A3(pi0781), .ZN(new_n24641_));
  NAND2_X1   g21447(.A1(new_n24639_), .A2(new_n24641_), .ZN(new_n24642_));
  NAND3_X1   g21448(.A1(new_n24642_), .A2(pi0619), .A3(pi1159), .ZN(new_n24643_));
  INV_X1     g21449(.I(new_n24642_), .ZN(new_n24644_));
  NAND3_X1   g21450(.A1(new_n24644_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n24645_));
  AOI21_X1   g21451(.A1(new_n24645_), .A2(new_n24643_), .B(new_n24605_), .ZN(new_n24646_));
  NAND2_X1   g21452(.A1(new_n24605_), .A2(new_n13879_), .ZN(new_n24647_));
  OAI21_X1   g21453(.A1(new_n13721_), .A2(new_n17943_), .B(new_n10656_), .ZN(new_n24648_));
  NAND2_X1   g21454(.A1(new_n24648_), .A2(new_n13108_), .ZN(new_n24649_));
  NAND2_X1   g21455(.A1(new_n10656_), .A2(new_n17943_), .ZN(new_n24650_));
  NAND4_X1   g21456(.A1(new_n13634_), .A2(pi0190), .A3(new_n3290_), .A4(new_n24650_), .ZN(new_n24651_));
  NOR3_X1    g21457(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n10656_), .ZN(new_n24652_));
  NOR3_X1    g21458(.A1(new_n14422_), .A2(pi0038), .A3(new_n10656_), .ZN(new_n24653_));
  OAI21_X1   g21459(.A1(new_n24652_), .A2(new_n24653_), .B(new_n15655_), .ZN(new_n24654_));
  AOI21_X1   g21460(.A1(new_n24649_), .A2(new_n24651_), .B(new_n24654_), .ZN(new_n24655_));
  NOR2_X1    g21461(.A1(new_n24604_), .A2(new_n13613_), .ZN(new_n24656_));
  XOR2_X1    g21462(.A1(new_n24656_), .A2(new_n13615_), .Z(new_n24657_));
  NAND2_X1   g21463(.A1(new_n24657_), .A2(new_n24655_), .ZN(new_n24658_));
  NAND2_X1   g21464(.A1(new_n24658_), .A2(pi0778), .ZN(new_n24659_));
  NOR2_X1    g21465(.A1(new_n24604_), .A2(new_n13614_), .ZN(new_n24660_));
  XOR2_X1    g21466(.A1(new_n24660_), .A2(new_n13615_), .Z(new_n24661_));
  NAND3_X1   g21467(.A1(new_n24661_), .A2(pi0778), .A3(new_n24655_), .ZN(new_n24662_));
  XOR2_X1    g21468(.A1(new_n24659_), .A2(new_n24662_), .Z(new_n24663_));
  INV_X1     g21469(.I(new_n24663_), .ZN(new_n24664_));
  NAND2_X1   g21470(.A1(new_n24604_), .A2(new_n13803_), .ZN(new_n24665_));
  OAI21_X1   g21471(.A1(new_n24664_), .A2(new_n13803_), .B(new_n24665_), .ZN(new_n24666_));
  OAI21_X1   g21472(.A1(new_n24666_), .A2(new_n13879_), .B(new_n24647_), .ZN(new_n24667_));
  INV_X1     g21473(.I(new_n24614_), .ZN(new_n24668_));
  NOR2_X1    g21474(.A1(new_n10656_), .A2(new_n17912_), .ZN(new_n24669_));
  INV_X1     g21475(.I(new_n24669_), .ZN(new_n24670_));
  NAND2_X1   g21476(.A1(new_n13461_), .A2(pi0763), .ZN(new_n24671_));
  XOR2_X1    g21477(.A1(new_n24671_), .A2(new_n24670_), .Z(new_n24672_));
  NAND2_X1   g21478(.A1(new_n24672_), .A2(new_n13521_), .ZN(new_n24673_));
  NAND3_X1   g21479(.A1(new_n14270_), .A2(pi0190), .A3(pi0763), .ZN(new_n24674_));
  NAND3_X1   g21480(.A1(new_n14272_), .A2(pi0190), .A3(new_n17912_), .ZN(new_n24675_));
  AOI21_X1   g21481(.A1(new_n24674_), .A2(new_n24675_), .B(new_n13152_), .ZN(new_n24676_));
  NAND3_X1   g21482(.A1(new_n13198_), .A2(pi0190), .A3(pi0763), .ZN(new_n24677_));
  NAND3_X1   g21483(.A1(new_n13200_), .A2(new_n10656_), .A3(pi0763), .ZN(new_n24678_));
  AOI21_X1   g21484(.A1(new_n24678_), .A2(new_n24677_), .B(new_n13191_), .ZN(new_n24679_));
  OAI21_X1   g21485(.A1(new_n24676_), .A2(new_n3212_), .B(new_n24679_), .ZN(new_n24680_));
  NAND3_X1   g21486(.A1(new_n24673_), .A2(new_n3183_), .A3(new_n24680_), .ZN(new_n24681_));
  NOR2_X1    g21487(.A1(new_n14284_), .A2(new_n10656_), .ZN(new_n24682_));
  XOR2_X1    g21488(.A1(new_n24682_), .A2(new_n24669_), .Z(new_n24683_));
  NAND3_X1   g21489(.A1(new_n24681_), .A2(new_n24683_), .A3(new_n13359_), .ZN(new_n24684_));
  NAND3_X1   g21490(.A1(new_n24684_), .A2(new_n17943_), .A3(new_n3290_), .ZN(new_n24685_));
  NAND2_X1   g21491(.A1(new_n3290_), .A2(pi0190), .ZN(new_n24686_));
  NAND2_X1   g21492(.A1(new_n5504_), .A2(new_n10656_), .ZN(new_n24687_));
  NOR2_X1    g21493(.A1(new_n24507_), .A2(new_n16751_), .ZN(new_n24688_));
  AOI21_X1   g21494(.A1(new_n24687_), .A2(new_n24688_), .B(pi0038), .ZN(new_n24689_));
  NOR4_X1    g21495(.A1(new_n19135_), .A2(new_n24689_), .A3(new_n24686_), .A4(new_n24670_), .ZN(new_n24690_));
  NAND2_X1   g21496(.A1(new_n24685_), .A2(new_n24690_), .ZN(new_n24691_));
  AOI21_X1   g21497(.A1(new_n24691_), .A2(new_n24668_), .B(new_n17943_), .ZN(new_n24692_));
  NOR2_X1    g21498(.A1(new_n24622_), .A2(new_n13613_), .ZN(new_n24693_));
  XOR2_X1    g21499(.A1(new_n24693_), .A2(new_n13615_), .Z(new_n24694_));
  NAND2_X1   g21500(.A1(new_n24694_), .A2(new_n24692_), .ZN(new_n24695_));
  AOI21_X1   g21501(.A1(new_n24661_), .A2(new_n24655_), .B(pi0608), .ZN(new_n24696_));
  NAND2_X1   g21502(.A1(new_n24658_), .A2(new_n14081_), .ZN(new_n24697_));
  AOI21_X1   g21503(.A1(new_n24695_), .A2(new_n24696_), .B(new_n24697_), .ZN(new_n24698_));
  NOR2_X1    g21504(.A1(new_n24622_), .A2(new_n13614_), .ZN(new_n24699_));
  XOR2_X1    g21505(.A1(new_n24699_), .A2(new_n13615_), .Z(new_n24700_));
  NAND3_X1   g21506(.A1(new_n24700_), .A2(new_n24692_), .A3(pi0778), .ZN(new_n24701_));
  OAI22_X1   g21507(.A1(new_n24698_), .A2(new_n24701_), .B1(pi0778), .B2(new_n24692_), .ZN(new_n24702_));
  NAND3_X1   g21508(.A1(new_n24702_), .A2(pi0609), .A3(pi1155), .ZN(new_n24703_));
  INV_X1     g21509(.I(new_n24702_), .ZN(new_n24704_));
  NAND3_X1   g21510(.A1(new_n24704_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n24705_));
  AOI21_X1   g21511(.A1(new_n24705_), .A2(new_n24703_), .B(new_n24664_), .ZN(new_n24706_));
  NAND2_X1   g21512(.A1(new_n24620_), .A2(pi0660), .ZN(new_n24707_));
  NAND2_X1   g21513(.A1(new_n24626_), .A2(new_n13783_), .ZN(new_n24708_));
  INV_X1     g21514(.I(new_n24708_), .ZN(new_n24709_));
  OAI21_X1   g21515(.A1(new_n24706_), .A2(new_n24707_), .B(new_n24709_), .ZN(new_n24710_));
  AOI21_X1   g21516(.A1(new_n24704_), .A2(pi0609), .B(new_n14694_), .ZN(new_n24711_));
  NOR3_X1    g21517(.A1(new_n24702_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n24712_));
  NOR2_X1    g21518(.A1(new_n24664_), .A2(new_n13801_), .ZN(new_n24713_));
  OAI21_X1   g21519(.A1(new_n24711_), .A2(new_n24712_), .B(new_n24713_), .ZN(new_n24714_));
  INV_X1     g21520(.I(new_n24714_), .ZN(new_n24715_));
  AOI22_X1   g21521(.A1(new_n24710_), .A2(new_n24715_), .B1(new_n13801_), .B2(new_n24702_), .ZN(new_n24716_));
  AOI21_X1   g21522(.A1(new_n24716_), .A2(pi1154), .B(new_n13819_), .ZN(new_n24717_));
  INV_X1     g21523(.I(new_n24716_), .ZN(new_n24718_));
  NOR3_X1    g21524(.A1(new_n24718_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n24719_));
  OAI21_X1   g21525(.A1(new_n24719_), .A2(new_n24717_), .B(new_n24666_), .ZN(new_n24720_));
  NAND2_X1   g21526(.A1(new_n24633_), .A2(pi0627), .ZN(new_n24721_));
  INV_X1     g21527(.I(new_n24721_), .ZN(new_n24722_));
  AOI21_X1   g21528(.A1(new_n24720_), .A2(new_n24722_), .B(new_n13855_), .ZN(new_n24723_));
  NAND3_X1   g21529(.A1(new_n24718_), .A2(pi0618), .A3(pi1154), .ZN(new_n24724_));
  NAND3_X1   g21530(.A1(new_n24716_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n24725_));
  NAND2_X1   g21531(.A1(new_n24724_), .A2(new_n24725_), .ZN(new_n24726_));
  AND2_X2    g21532(.A1(new_n24726_), .A2(new_n24666_), .Z(new_n24727_));
  INV_X1     g21533(.I(new_n24637_), .ZN(new_n24728_));
  NAND3_X1   g21534(.A1(new_n24718_), .A2(new_n19177_), .A3(new_n24728_), .ZN(new_n24729_));
  NOR3_X1    g21535(.A1(new_n24727_), .A2(new_n24723_), .A3(new_n24729_), .ZN(new_n24730_));
  INV_X1     g21536(.I(new_n24723_), .ZN(new_n24731_));
  NOR2_X1    g21537(.A1(new_n24727_), .A2(new_n24729_), .ZN(new_n24732_));
  NOR2_X1    g21538(.A1(new_n24732_), .A2(new_n24731_), .ZN(new_n24733_));
  NOR2_X1    g21539(.A1(new_n24733_), .A2(new_n24730_), .ZN(new_n24734_));
  AOI21_X1   g21540(.A1(new_n24734_), .A2(pi1159), .B(new_n13904_), .ZN(new_n24735_));
  NOR4_X1    g21541(.A1(new_n24733_), .A2(pi0619), .A3(new_n13868_), .A4(new_n24730_), .ZN(new_n24736_));
  OAI21_X1   g21542(.A1(new_n24735_), .A2(new_n24736_), .B(new_n24667_), .ZN(new_n24737_));
  NAND2_X1   g21543(.A1(new_n24737_), .A2(new_n16474_), .ZN(new_n24738_));
  NAND3_X1   g21544(.A1(new_n24642_), .A2(pi0619), .A3(pi1159), .ZN(new_n24739_));
  NAND3_X1   g21545(.A1(new_n24644_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n24740_));
  AOI21_X1   g21546(.A1(new_n24740_), .A2(new_n24739_), .B(new_n24605_), .ZN(new_n24741_));
  NAND4_X1   g21547(.A1(new_n24646_), .A2(new_n24741_), .A3(pi0789), .A4(new_n24642_), .ZN(new_n24742_));
  NOR2_X1    g21548(.A1(new_n24646_), .A2(new_n13896_), .ZN(new_n24743_));
  NAND3_X1   g21549(.A1(new_n24741_), .A2(pi0789), .A3(new_n24642_), .ZN(new_n24744_));
  NAND2_X1   g21550(.A1(new_n24744_), .A2(new_n24743_), .ZN(new_n24745_));
  NAND2_X1   g21551(.A1(new_n24745_), .A2(new_n24742_), .ZN(new_n24746_));
  NAND3_X1   g21552(.A1(new_n24746_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n24747_));
  INV_X1     g21553(.I(new_n24746_), .ZN(new_n24748_));
  NAND3_X1   g21554(.A1(new_n24748_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n24749_));
  AOI21_X1   g21555(.A1(new_n24749_), .A2(new_n24747_), .B(new_n24605_), .ZN(new_n24750_));
  NOR2_X1    g21556(.A1(new_n24667_), .A2(new_n13918_), .ZN(new_n24751_));
  AOI21_X1   g21557(.A1(new_n13918_), .A2(new_n24604_), .B(new_n24751_), .ZN(new_n24752_));
  NOR2_X1    g21558(.A1(new_n24752_), .A2(new_n14162_), .ZN(new_n24753_));
  OAI21_X1   g21559(.A1(new_n24750_), .A2(new_n24753_), .B(new_n19204_), .ZN(new_n24754_));
  NOR2_X1    g21560(.A1(new_n24734_), .A2(pi0789), .ZN(new_n24755_));
  NOR2_X1    g21561(.A1(new_n24746_), .A2(new_n19208_), .ZN(new_n24756_));
  XOR2_X1    g21562(.A1(new_n24756_), .A2(new_n19028_), .Z(new_n24757_));
  NOR4_X1    g21563(.A1(new_n24757_), .A2(new_n15479_), .A3(new_n24605_), .A4(new_n24755_), .ZN(new_n24758_));
  AOI22_X1   g21564(.A1(new_n24738_), .A2(new_n24646_), .B1(new_n24758_), .B2(new_n24754_), .ZN(new_n24759_));
  AOI21_X1   g21565(.A1(new_n24734_), .A2(pi0619), .B(new_n13904_), .ZN(new_n24760_));
  NOR4_X1    g21566(.A1(new_n24733_), .A2(new_n13860_), .A3(pi1159), .A4(new_n24730_), .ZN(new_n24761_));
  OAI21_X1   g21567(.A1(new_n24760_), .A2(new_n24761_), .B(new_n24667_), .ZN(new_n24762_));
  NOR2_X1    g21568(.A1(new_n24741_), .A2(pi0648), .ZN(new_n24763_));
  NAND2_X1   g21569(.A1(new_n24762_), .A2(new_n24763_), .ZN(new_n24764_));
  NOR2_X1    g21570(.A1(new_n24604_), .A2(new_n16372_), .ZN(new_n24765_));
  INV_X1     g21571(.I(new_n24765_), .ZN(new_n24766_));
  NAND3_X1   g21572(.A1(new_n24745_), .A2(new_n16372_), .A3(new_n24742_), .ZN(new_n24767_));
  AOI21_X1   g21573(.A1(new_n24767_), .A2(new_n24766_), .B(new_n13993_), .ZN(new_n24768_));
  NOR2_X1    g21574(.A1(new_n24604_), .A2(new_n13994_), .ZN(new_n24769_));
  OR2_X2     g21575(.A1(new_n24768_), .A2(new_n24769_), .Z(new_n24770_));
  NAND2_X1   g21576(.A1(new_n24752_), .A2(new_n13966_), .ZN(new_n24771_));
  OAI21_X1   g21577(.A1(new_n13966_), .A2(new_n24604_), .B(new_n24771_), .ZN(new_n24772_));
  NAND2_X1   g21578(.A1(new_n24772_), .A2(new_n12777_), .ZN(new_n24773_));
  NOR2_X1    g21579(.A1(new_n24604_), .A2(new_n13942_), .ZN(new_n24774_));
  AOI21_X1   g21580(.A1(new_n24772_), .A2(new_n13942_), .B(new_n24774_), .ZN(new_n24775_));
  NOR2_X1    g21581(.A1(new_n24775_), .A2(pi1156), .ZN(new_n24776_));
  NOR2_X1    g21582(.A1(new_n24604_), .A2(pi0628), .ZN(new_n24777_));
  AOI21_X1   g21583(.A1(new_n24772_), .A2(pi0628), .B(new_n24777_), .ZN(new_n24778_));
  NOR2_X1    g21584(.A1(new_n24778_), .A2(new_n13969_), .ZN(new_n24779_));
  OAI21_X1   g21585(.A1(new_n24776_), .A2(new_n24779_), .B(pi0792), .ZN(new_n24780_));
  NAND2_X1   g21586(.A1(new_n24780_), .A2(new_n24773_), .ZN(new_n24781_));
  NAND2_X1   g21587(.A1(new_n24781_), .A2(new_n14005_), .ZN(new_n24782_));
  NAND2_X1   g21588(.A1(new_n24605_), .A2(pi0647), .ZN(new_n24783_));
  AOI21_X1   g21589(.A1(new_n24782_), .A2(new_n24783_), .B(new_n14012_), .ZN(new_n24784_));
  NOR2_X1    g21590(.A1(new_n24604_), .A2(pi0647), .ZN(new_n24785_));
  AOI21_X1   g21591(.A1(new_n24781_), .A2(pi0647), .B(new_n24785_), .ZN(new_n24786_));
  NAND2_X1   g21592(.A1(new_n24786_), .A2(new_n14206_), .ZN(new_n24787_));
  OR2_X2     g21593(.A1(new_n24784_), .A2(new_n24787_), .Z(new_n24788_));
  NAND2_X1   g21594(.A1(new_n24784_), .A2(new_n24787_), .ZN(new_n24789_));
  AOI21_X1   g21595(.A1(new_n24788_), .A2(new_n24789_), .B(new_n12776_), .ZN(new_n24790_));
  NOR2_X1    g21596(.A1(new_n24790_), .A2(new_n24770_), .ZN(new_n24791_));
  OAI22_X1   g21597(.A1(new_n24759_), .A2(new_n24764_), .B1(new_n16891_), .B2(new_n24791_), .ZN(new_n24792_));
  AOI21_X1   g21598(.A1(new_n24748_), .A2(new_n16372_), .B(new_n24765_), .ZN(new_n24793_));
  NOR2_X1    g21599(.A1(new_n24775_), .A2(new_n15270_), .ZN(new_n24794_));
  NAND2_X1   g21600(.A1(new_n24778_), .A2(new_n13990_), .ZN(new_n24795_));
  XNOR2_X1   g21601(.A1(new_n24794_), .A2(new_n24795_), .ZN(new_n24796_));
  NAND2_X1   g21602(.A1(new_n24796_), .A2(pi0792), .ZN(new_n24797_));
  AOI21_X1   g21603(.A1(new_n24793_), .A2(new_n24797_), .B(new_n16875_), .ZN(new_n24798_));
  NAND2_X1   g21604(.A1(new_n24781_), .A2(new_n12776_), .ZN(new_n24799_));
  AOI21_X1   g21605(.A1(new_n24782_), .A2(new_n24783_), .B(pi1157), .ZN(new_n24800_));
  NOR2_X1    g21606(.A1(new_n24786_), .A2(new_n14006_), .ZN(new_n24801_));
  OAI21_X1   g21607(.A1(new_n24801_), .A2(new_n24800_), .B(pi0787), .ZN(new_n24802_));
  NAND2_X1   g21608(.A1(new_n24802_), .A2(new_n24799_), .ZN(new_n24803_));
  INV_X1     g21609(.I(new_n24803_), .ZN(new_n24804_));
  OAI21_X1   g21610(.A1(new_n24768_), .A2(new_n24769_), .B(new_n14211_), .ZN(new_n24805_));
  NOR2_X1    g21611(.A1(new_n24604_), .A2(new_n14211_), .ZN(new_n24806_));
  INV_X1     g21612(.I(new_n24806_), .ZN(new_n24807_));
  NOR2_X1    g21613(.A1(new_n14243_), .A2(pi0644), .ZN(new_n24808_));
  AOI21_X1   g21614(.A1(new_n24805_), .A2(new_n24807_), .B(new_n24808_), .ZN(new_n24809_));
  AOI21_X1   g21615(.A1(new_n24809_), .A2(pi0715), .B(pi0644), .ZN(new_n24810_));
  AOI21_X1   g21616(.A1(new_n24770_), .A2(new_n14211_), .B(new_n24806_), .ZN(new_n24811_));
  AOI21_X1   g21617(.A1(new_n24604_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n24812_));
  NOR2_X1    g21618(.A1(new_n24812_), .A2(pi0644), .ZN(new_n24813_));
  NOR2_X1    g21619(.A1(new_n24811_), .A2(new_n24813_), .ZN(new_n24814_));
  AOI21_X1   g21620(.A1(new_n24814_), .A2(pi0715), .B(new_n24803_), .ZN(new_n24815_));
  OAI22_X1   g21621(.A1(new_n24815_), .A2(new_n14204_), .B1(new_n24810_), .B2(new_n24804_), .ZN(new_n24816_));
  AOI22_X1   g21622(.A1(new_n24792_), .A2(new_n24798_), .B1(new_n24816_), .B2(new_n19269_), .ZN(new_n24817_));
  NOR3_X1    g21623(.A1(new_n24811_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n24818_));
  NOR3_X1    g21624(.A1(new_n24814_), .A2(pi0644), .A3(new_n12775_), .ZN(new_n24819_));
  NOR2_X1    g21625(.A1(new_n24592_), .A2(pi0790), .ZN(new_n24820_));
  NOR4_X1    g21626(.A1(new_n24811_), .A2(new_n14799_), .A3(new_n24808_), .A4(new_n24820_), .ZN(new_n24821_));
  OAI21_X1   g21627(.A1(new_n24819_), .A2(new_n24818_), .B(new_n24821_), .ZN(new_n24822_));
  OAI21_X1   g21628(.A1(new_n24817_), .A2(new_n24822_), .B(new_n24603_), .ZN(po0347));
  NOR2_X1    g21629(.A1(new_n14652_), .A2(new_n17987_), .ZN(new_n24824_));
  INV_X1     g21630(.I(new_n24824_), .ZN(new_n24825_));
  NOR2_X1    g21631(.A1(new_n9992_), .A2(pi0191), .ZN(new_n24826_));
  NOR2_X1    g21632(.A1(new_n24826_), .A2(pi1153), .ZN(new_n24827_));
  NAND2_X1   g21633(.A1(new_n24825_), .A2(new_n24827_), .ZN(new_n24828_));
  INV_X1     g21634(.I(new_n24828_), .ZN(new_n24829_));
  NOR2_X1    g21635(.A1(new_n24829_), .A2(new_n13748_), .ZN(new_n24830_));
  AOI21_X1   g21636(.A1(new_n13218_), .A2(pi0729), .B(new_n24826_), .ZN(new_n24831_));
  INV_X1     g21637(.I(new_n24831_), .ZN(new_n24832_));
  AOI21_X1   g21638(.A1(new_n24825_), .A2(new_n24832_), .B(new_n13614_), .ZN(new_n24833_));
  INV_X1     g21639(.I(new_n24833_), .ZN(new_n24834_));
  NOR3_X1    g21640(.A1(new_n24834_), .A2(new_n13748_), .A3(new_n24832_), .ZN(new_n24835_));
  XNOR2_X1   g21641(.A1(new_n24835_), .A2(new_n24830_), .ZN(new_n24836_));
  NAND2_X1   g21642(.A1(new_n24836_), .A2(new_n14049_), .ZN(new_n24837_));
  NOR2_X1    g21643(.A1(new_n24837_), .A2(new_n14051_), .ZN(new_n24838_));
  INV_X1     g21644(.I(new_n24838_), .ZN(new_n24839_));
  NOR2_X1    g21645(.A1(new_n24839_), .A2(new_n14163_), .ZN(new_n24840_));
  NAND2_X1   g21646(.A1(new_n24840_), .A2(new_n18929_), .ZN(new_n24841_));
  NOR2_X1    g21647(.A1(new_n24841_), .A2(new_n14060_), .ZN(new_n24842_));
  INV_X1     g21648(.I(new_n24826_), .ZN(new_n24843_));
  NAND3_X1   g21649(.A1(new_n24842_), .A2(pi0647), .A3(pi1157), .ZN(new_n24844_));
  OR3_X2     g21650(.A1(new_n24842_), .A2(new_n14005_), .A3(pi1157), .Z(new_n24845_));
  AOI21_X1   g21651(.A1(new_n24845_), .A2(new_n24844_), .B(new_n24843_), .ZN(new_n24846_));
  INV_X1     g21652(.I(new_n24846_), .ZN(new_n24847_));
  NOR2_X1    g21653(.A1(new_n24843_), .A2(pi0647), .ZN(new_n24848_));
  AOI21_X1   g21654(.A1(new_n24842_), .A2(pi0647), .B(new_n24848_), .ZN(new_n24849_));
  AOI21_X1   g21655(.A1(new_n24849_), .A2(pi1157), .B(new_n12776_), .ZN(new_n24850_));
  AOI22_X1   g21656(.A1(new_n24847_), .A2(new_n24850_), .B1(new_n12776_), .B2(new_n24842_), .ZN(new_n24851_));
  INV_X1     g21657(.I(new_n24851_), .ZN(new_n24852_));
  NOR2_X1    g21658(.A1(new_n13105_), .A2(new_n17956_), .ZN(new_n24853_));
  INV_X1     g21659(.I(new_n24853_), .ZN(new_n24854_));
  NOR2_X1    g21660(.A1(new_n24853_), .A2(new_n24826_), .ZN(new_n24855_));
  INV_X1     g21661(.I(new_n24855_), .ZN(new_n24856_));
  NAND3_X1   g21662(.A1(new_n24856_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n24857_));
  AOI21_X1   g21663(.A1(new_n24857_), .A2(new_n16444_), .B(new_n24854_), .ZN(new_n24858_));
  NOR2_X1    g21664(.A1(new_n24858_), .A2(new_n13801_), .ZN(new_n24859_));
  NOR2_X1    g21665(.A1(new_n24826_), .A2(pi1155), .ZN(new_n24860_));
  NOR3_X1    g21666(.A1(new_n24854_), .A2(new_n16444_), .A3(new_n24860_), .ZN(new_n24861_));
  NAND4_X1   g21667(.A1(new_n24861_), .A2(new_n24856_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n24862_));
  XOR2_X1    g21668(.A1(new_n24859_), .A2(new_n24862_), .Z(new_n24863_));
  NOR2_X1    g21669(.A1(new_n24863_), .A2(new_n13817_), .ZN(new_n24864_));
  OAI21_X1   g21670(.A1(new_n24864_), .A2(pi0618), .B(new_n9992_), .ZN(new_n24865_));
  NAND2_X1   g21671(.A1(new_n24865_), .A2(pi0781), .ZN(new_n24866_));
  OAI21_X1   g21672(.A1(new_n24864_), .A2(new_n9992_), .B(pi0618), .ZN(new_n24867_));
  NOR3_X1    g21673(.A1(new_n24867_), .A2(new_n13855_), .A3(new_n24863_), .ZN(new_n24868_));
  XOR2_X1    g21674(.A1(new_n24868_), .A2(new_n24866_), .Z(new_n24869_));
  NOR2_X1    g21675(.A1(new_n24869_), .A2(new_n13868_), .ZN(new_n24870_));
  OAI21_X1   g21676(.A1(new_n24870_), .A2(pi0619), .B(new_n9992_), .ZN(new_n24871_));
  NAND2_X1   g21677(.A1(new_n24871_), .A2(pi0789), .ZN(new_n24872_));
  OAI21_X1   g21678(.A1(new_n24870_), .A2(new_n9992_), .B(pi0619), .ZN(new_n24873_));
  NOR3_X1    g21679(.A1(new_n24873_), .A2(new_n13896_), .A3(new_n24869_), .ZN(new_n24874_));
  XOR2_X1    g21680(.A1(new_n24874_), .A2(new_n24872_), .Z(new_n24875_));
  NAND2_X1   g21681(.A1(new_n24875_), .A2(new_n16372_), .ZN(new_n24876_));
  OAI21_X1   g21682(.A1(new_n16372_), .A2(new_n24826_), .B(new_n24876_), .ZN(new_n24877_));
  NOR2_X1    g21683(.A1(new_n24877_), .A2(new_n18968_), .ZN(new_n24878_));
  NAND2_X1   g21684(.A1(new_n18967_), .A2(new_n24826_), .ZN(new_n24879_));
  XOR2_X1    g21685(.A1(new_n24878_), .A2(new_n24879_), .Z(new_n24880_));
  AOI21_X1   g21686(.A1(new_n24843_), .A2(new_n14254_), .B(pi0644), .ZN(new_n24881_));
  NAND2_X1   g21687(.A1(new_n24875_), .A2(new_n13962_), .ZN(new_n24882_));
  XOR2_X1    g21688(.A1(new_n24882_), .A2(new_n18976_), .Z(new_n24883_));
  AOI22_X1   g21689(.A1(new_n24883_), .A2(new_n24826_), .B1(new_n16639_), .B2(new_n24840_), .ZN(new_n24884_));
  NOR2_X1    g21690(.A1(new_n24831_), .A2(new_n13203_), .ZN(new_n24885_));
  NAND2_X1   g21691(.A1(new_n24885_), .A2(pi0625), .ZN(new_n24886_));
  NAND3_X1   g21692(.A1(new_n24886_), .A2(pi1153), .A3(new_n24855_), .ZN(new_n24887_));
  NOR2_X1    g21693(.A1(new_n24829_), .A2(new_n14081_), .ZN(new_n24888_));
  AOI21_X1   g21694(.A1(new_n24888_), .A2(new_n24887_), .B(new_n13748_), .ZN(new_n24889_));
  NOR2_X1    g21695(.A1(new_n24856_), .A2(new_n24885_), .ZN(new_n24890_));
  INV_X1     g21696(.I(new_n24886_), .ZN(new_n24891_));
  OAI21_X1   g21697(.A1(new_n24890_), .A2(new_n24891_), .B(new_n24827_), .ZN(new_n24892_));
  NAND4_X1   g21698(.A1(new_n24892_), .A2(new_n13749_), .A3(new_n24834_), .A4(new_n24890_), .ZN(new_n24893_));
  XNOR2_X1   g21699(.A1(new_n24893_), .A2(new_n24889_), .ZN(new_n24894_));
  NAND2_X1   g21700(.A1(new_n24894_), .A2(new_n13801_), .ZN(new_n24895_));
  NOR2_X1    g21701(.A1(new_n24858_), .A2(pi0660), .ZN(new_n24898_));
  NOR2_X1    g21702(.A1(new_n24894_), .A2(new_n13766_), .ZN(new_n24899_));
  XOR2_X1    g21703(.A1(new_n24899_), .A2(new_n14090_), .Z(new_n24900_));
  NOR2_X1    g21704(.A1(new_n24836_), .A2(new_n13801_), .ZN(new_n24901_));
  NAND2_X1   g21705(.A1(new_n24900_), .A2(new_n24901_), .ZN(new_n24902_));
  OAI21_X1   g21706(.A1(new_n24902_), .A2(new_n24898_), .B(new_n24895_), .ZN(new_n24903_));
  NAND2_X1   g21707(.A1(new_n24903_), .A2(new_n13855_), .ZN(new_n24904_));
  INV_X1     g21708(.I(new_n24837_), .ZN(new_n24905_));
  NOR2_X1    g21709(.A1(new_n24903_), .A2(new_n13816_), .ZN(new_n24906_));
  XOR2_X1    g21710(.A1(new_n24906_), .A2(new_n13818_), .Z(new_n24907_));
  NAND2_X1   g21711(.A1(new_n24907_), .A2(new_n24905_), .ZN(new_n24908_));
  NAND3_X1   g21712(.A1(new_n24908_), .A2(new_n13823_), .A3(new_n24867_), .ZN(new_n24909_));
  NAND3_X1   g21713(.A1(new_n24909_), .A2(new_n13823_), .A3(new_n24865_), .ZN(new_n24910_));
  NOR2_X1    g21714(.A1(new_n24903_), .A2(new_n13817_), .ZN(new_n24911_));
  XOR2_X1    g21715(.A1(new_n24911_), .A2(new_n13818_), .Z(new_n24912_));
  NAND4_X1   g21716(.A1(new_n24910_), .A2(pi0781), .A3(new_n24905_), .A4(new_n24912_), .ZN(new_n24913_));
  NAND2_X1   g21717(.A1(new_n24913_), .A2(new_n24904_), .ZN(new_n24914_));
  NOR2_X1    g21718(.A1(new_n24914_), .A2(new_n13860_), .ZN(new_n24915_));
  XOR2_X1    g21719(.A1(new_n24915_), .A2(new_n13904_), .Z(new_n24916_));
  NOR2_X1    g21720(.A1(new_n24916_), .A2(new_n24839_), .ZN(new_n24917_));
  NAND2_X1   g21721(.A1(new_n24873_), .A2(new_n13884_), .ZN(new_n24918_));
  INV_X1     g21722(.I(new_n24914_), .ZN(new_n24919_));
  AOI21_X1   g21723(.A1(new_n24919_), .A2(new_n14143_), .B(pi0789), .ZN(new_n24920_));
  OAI21_X1   g21724(.A1(new_n24917_), .A2(new_n24918_), .B(new_n24920_), .ZN(new_n24921_));
  NOR2_X1    g21725(.A1(new_n24914_), .A2(new_n13868_), .ZN(new_n24922_));
  XOR2_X1    g21726(.A1(new_n24922_), .A2(new_n13903_), .Z(new_n24923_));
  NAND2_X1   g21727(.A1(new_n24871_), .A2(new_n19018_), .ZN(new_n24924_));
  AOI21_X1   g21728(.A1(new_n24923_), .A2(new_n24838_), .B(new_n24924_), .ZN(new_n24925_));
  AOI21_X1   g21729(.A1(new_n24921_), .A2(new_n24925_), .B(new_n24884_), .ZN(new_n24926_));
  NAND3_X1   g21730(.A1(new_n24877_), .A2(new_n18929_), .A3(new_n24840_), .ZN(new_n24927_));
  NAND2_X1   g21731(.A1(new_n24927_), .A2(new_n16569_), .ZN(new_n24928_));
  XOR2_X1    g21732(.A1(new_n24928_), .A2(new_n16572_), .Z(new_n24929_));
  AOI21_X1   g21733(.A1(new_n19022_), .A2(new_n24927_), .B(new_n24929_), .ZN(new_n24930_));
  NAND2_X1   g21734(.A1(new_n24875_), .A2(new_n13963_), .ZN(new_n24931_));
  XNOR2_X1   g21735(.A1(new_n24931_), .A2(new_n19028_), .ZN(new_n24932_));
  NOR3_X1    g21736(.A1(new_n24932_), .A2(new_n16424_), .A3(new_n24843_), .ZN(new_n24933_));
  OAI21_X1   g21737(.A1(new_n24930_), .A2(new_n16574_), .B(new_n24933_), .ZN(new_n24934_));
  NOR2_X1    g21738(.A1(new_n24877_), .A2(new_n13994_), .ZN(new_n24935_));
  XNOR2_X1   g21739(.A1(new_n24935_), .A2(new_n19033_), .ZN(new_n24936_));
  AOI22_X1   g21740(.A1(new_n24936_), .A2(new_n24826_), .B1(new_n14206_), .B2(new_n24849_), .ZN(new_n24937_));
  NOR3_X1    g21741(.A1(new_n24937_), .A2(new_n14010_), .A3(new_n24847_), .ZN(new_n24938_));
  OAI22_X1   g21742(.A1(new_n24926_), .A2(new_n24934_), .B1(new_n12776_), .B2(new_n24938_), .ZN(new_n24939_));
  NAND2_X1   g21743(.A1(new_n24939_), .A2(pi0644), .ZN(new_n24940_));
  XOR2_X1    g21744(.A1(new_n24940_), .A2(new_n14205_), .Z(new_n24941_));
  NOR2_X1    g21745(.A1(new_n24941_), .A2(new_n24851_), .ZN(new_n24942_));
  NAND2_X1   g21746(.A1(new_n24880_), .A2(pi0715), .ZN(new_n24943_));
  XOR2_X1    g21747(.A1(new_n24943_), .A2(new_n14205_), .Z(new_n24944_));
  OAI21_X1   g21748(.A1(new_n24944_), .A2(new_n24843_), .B(new_n19043_), .ZN(new_n24945_));
  OAI22_X1   g21749(.A1(new_n24942_), .A2(new_n24945_), .B1(new_n24880_), .B2(new_n24881_), .ZN(new_n24946_));
  NAND2_X1   g21750(.A1(new_n24939_), .A2(pi0715), .ZN(new_n24947_));
  XOR2_X1    g21751(.A1(new_n24947_), .A2(new_n14217_), .Z(new_n24948_));
  AOI21_X1   g21752(.A1(po1038), .A2(new_n12167_), .B(pi0832), .ZN(new_n24949_));
  NAND4_X1   g21753(.A1(new_n24946_), .A2(new_n24852_), .A3(new_n24948_), .A4(new_n24949_), .ZN(new_n24950_));
  NOR2_X1    g21754(.A1(new_n14428_), .A2(pi0191), .ZN(new_n24951_));
  INV_X1     g21755(.I(new_n24951_), .ZN(new_n24952_));
  OAI22_X1   g21756(.A1(new_n17127_), .A2(new_n12167_), .B1(new_n17956_), .B2(new_n19052_), .ZN(new_n24953_));
  OAI21_X1   g21757(.A1(pi0191), .A2(new_n14299_), .B(new_n14301_), .ZN(new_n24954_));
  NAND2_X1   g21758(.A1(new_n14299_), .A2(pi0746), .ZN(new_n24955_));
  NAND4_X1   g21759(.A1(new_n24954_), .A2(new_n17956_), .A3(new_n14362_), .A4(new_n24955_), .ZN(new_n24956_));
  NAND3_X1   g21760(.A1(new_n24956_), .A2(pi0038), .A3(pi0191), .ZN(new_n24957_));
  NAND2_X1   g21761(.A1(new_n24957_), .A2(new_n3183_), .ZN(new_n24958_));
  NAND2_X1   g21762(.A1(new_n13109_), .A2(new_n12167_), .ZN(new_n24959_));
  NAND4_X1   g21763(.A1(new_n24958_), .A2(pi0038), .A3(new_n24953_), .A4(new_n24959_), .ZN(new_n24960_));
  AOI21_X1   g21764(.A1(new_n24960_), .A2(new_n17956_), .B(new_n13107_), .ZN(new_n24961_));
  NAND2_X1   g21765(.A1(new_n24961_), .A2(new_n3289_), .ZN(new_n24962_));
  NAND2_X1   g21766(.A1(new_n3290_), .A2(new_n12167_), .ZN(new_n24963_));
  NAND3_X1   g21767(.A1(new_n24962_), .A2(new_n13776_), .A3(new_n24963_), .ZN(new_n24964_));
  NAND2_X1   g21768(.A1(new_n24952_), .A2(new_n13780_), .ZN(new_n24965_));
  NAND2_X1   g21769(.A1(new_n24964_), .A2(new_n24965_), .ZN(new_n24966_));
  NAND2_X1   g21770(.A1(new_n24966_), .A2(pi0609), .ZN(new_n24967_));
  NAND2_X1   g21771(.A1(new_n24967_), .A2(pi0785), .ZN(new_n24968_));
  NAND2_X1   g21772(.A1(new_n24962_), .A2(new_n24963_), .ZN(new_n24969_));
  NOR2_X1    g21773(.A1(new_n24952_), .A2(new_n13776_), .ZN(new_n24970_));
  AOI21_X1   g21774(.A1(new_n24969_), .A2(new_n13776_), .B(new_n24970_), .ZN(new_n24971_));
  AOI21_X1   g21775(.A1(new_n24952_), .A2(new_n14467_), .B(pi0609), .ZN(new_n24972_));
  OR2_X2     g21776(.A1(new_n24964_), .A2(new_n24972_), .Z(new_n24973_));
  NOR3_X1    g21777(.A1(new_n24973_), .A2(new_n13801_), .A3(new_n24971_), .ZN(new_n24974_));
  XNOR2_X1   g21778(.A1(new_n24974_), .A2(new_n24968_), .ZN(new_n24975_));
  NAND3_X1   g21779(.A1(new_n24975_), .A2(pi0618), .A3(pi1154), .ZN(new_n24976_));
  XOR2_X1    g21780(.A1(new_n24974_), .A2(new_n24968_), .Z(new_n24977_));
  NAND3_X1   g21781(.A1(new_n24977_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n24978_));
  NAND2_X1   g21782(.A1(new_n24976_), .A2(new_n24978_), .ZN(new_n24979_));
  NAND2_X1   g21783(.A1(new_n24979_), .A2(new_n24951_), .ZN(new_n24980_));
  NAND2_X1   g21784(.A1(new_n24980_), .A2(pi0781), .ZN(new_n24981_));
  NAND3_X1   g21785(.A1(new_n24975_), .A2(pi0618), .A3(pi1154), .ZN(new_n24982_));
  NAND3_X1   g21786(.A1(new_n24977_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n24983_));
  AOI21_X1   g21787(.A1(new_n24982_), .A2(new_n24983_), .B(new_n24952_), .ZN(new_n24984_));
  NOR2_X1    g21788(.A1(new_n24977_), .A2(new_n13855_), .ZN(new_n24985_));
  NAND3_X1   g21789(.A1(new_n24981_), .A2(new_n24984_), .A3(new_n24985_), .ZN(new_n24986_));
  NAND2_X1   g21790(.A1(new_n24984_), .A2(new_n24985_), .ZN(new_n24987_));
  NAND3_X1   g21791(.A1(new_n24987_), .A2(new_n24980_), .A3(pi0781), .ZN(new_n24988_));
  NAND2_X1   g21792(.A1(new_n24986_), .A2(new_n24988_), .ZN(new_n24989_));
  NAND3_X1   g21793(.A1(new_n24989_), .A2(pi0619), .A3(pi1159), .ZN(new_n24990_));
  INV_X1     g21794(.I(new_n24989_), .ZN(new_n24991_));
  NAND3_X1   g21795(.A1(new_n24991_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n24992_));
  AOI21_X1   g21796(.A1(new_n24992_), .A2(new_n24990_), .B(new_n24952_), .ZN(new_n24993_));
  NAND2_X1   g21797(.A1(new_n24952_), .A2(new_n13879_), .ZN(new_n24994_));
  OAI21_X1   g21798(.A1(new_n13721_), .A2(new_n17987_), .B(new_n12167_), .ZN(new_n24995_));
  NAND2_X1   g21799(.A1(new_n24995_), .A2(new_n13108_), .ZN(new_n24996_));
  NAND2_X1   g21800(.A1(new_n12167_), .A2(new_n17987_), .ZN(new_n24997_));
  NAND4_X1   g21801(.A1(new_n13634_), .A2(pi0191), .A3(new_n3290_), .A4(new_n24997_), .ZN(new_n24998_));
  NOR3_X1    g21802(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n12167_), .ZN(new_n24999_));
  NOR3_X1    g21803(.A1(new_n14422_), .A2(pi0038), .A3(new_n12167_), .ZN(new_n25000_));
  OAI21_X1   g21804(.A1(new_n24999_), .A2(new_n25000_), .B(new_n15655_), .ZN(new_n25001_));
  AOI21_X1   g21805(.A1(new_n24996_), .A2(new_n24998_), .B(new_n25001_), .ZN(new_n25002_));
  NOR2_X1    g21806(.A1(new_n24951_), .A2(new_n13613_), .ZN(new_n25003_));
  XOR2_X1    g21807(.A1(new_n25003_), .A2(new_n13615_), .Z(new_n25004_));
  NAND2_X1   g21808(.A1(new_n25004_), .A2(new_n25002_), .ZN(new_n25005_));
  NAND2_X1   g21809(.A1(new_n25005_), .A2(pi0778), .ZN(new_n25006_));
  NOR2_X1    g21810(.A1(new_n24951_), .A2(new_n13614_), .ZN(new_n25007_));
  XOR2_X1    g21811(.A1(new_n25007_), .A2(new_n13615_), .Z(new_n25008_));
  NAND3_X1   g21812(.A1(new_n25008_), .A2(pi0778), .A3(new_n25002_), .ZN(new_n25009_));
  XOR2_X1    g21813(.A1(new_n25006_), .A2(new_n25009_), .Z(new_n25010_));
  INV_X1     g21814(.I(new_n25010_), .ZN(new_n25011_));
  NAND2_X1   g21815(.A1(new_n24951_), .A2(new_n13803_), .ZN(new_n25012_));
  OAI21_X1   g21816(.A1(new_n25011_), .A2(new_n13803_), .B(new_n25012_), .ZN(new_n25013_));
  OAI21_X1   g21817(.A1(new_n25013_), .A2(new_n13879_), .B(new_n24994_), .ZN(new_n25014_));
  INV_X1     g21818(.I(new_n24961_), .ZN(new_n25015_));
  NOR2_X1    g21819(.A1(new_n12167_), .A2(new_n17956_), .ZN(new_n25016_));
  INV_X1     g21820(.I(new_n25016_), .ZN(new_n25017_));
  NAND2_X1   g21821(.A1(new_n13461_), .A2(pi0746), .ZN(new_n25018_));
  XOR2_X1    g21822(.A1(new_n25018_), .A2(new_n25017_), .Z(new_n25019_));
  NAND2_X1   g21823(.A1(new_n25019_), .A2(new_n13521_), .ZN(new_n25020_));
  NAND3_X1   g21824(.A1(new_n14270_), .A2(pi0191), .A3(pi0746), .ZN(new_n25021_));
  NAND3_X1   g21825(.A1(new_n14272_), .A2(pi0191), .A3(new_n17956_), .ZN(new_n25022_));
  AOI21_X1   g21826(.A1(new_n25021_), .A2(new_n25022_), .B(new_n13152_), .ZN(new_n25023_));
  NAND3_X1   g21827(.A1(new_n13198_), .A2(pi0191), .A3(pi0746), .ZN(new_n25024_));
  NAND3_X1   g21828(.A1(new_n13200_), .A2(new_n12167_), .A3(pi0746), .ZN(new_n25025_));
  AOI21_X1   g21829(.A1(new_n25025_), .A2(new_n25024_), .B(new_n13191_), .ZN(new_n25026_));
  OAI21_X1   g21830(.A1(new_n25023_), .A2(new_n3212_), .B(new_n25026_), .ZN(new_n25027_));
  NAND3_X1   g21831(.A1(new_n25020_), .A2(new_n3183_), .A3(new_n25027_), .ZN(new_n25028_));
  NOR2_X1    g21832(.A1(new_n14284_), .A2(new_n12167_), .ZN(new_n25029_));
  XOR2_X1    g21833(.A1(new_n25029_), .A2(new_n25016_), .Z(new_n25030_));
  NAND3_X1   g21834(.A1(new_n25028_), .A2(new_n25030_), .A3(new_n13359_), .ZN(new_n25031_));
  NAND3_X1   g21835(.A1(new_n25031_), .A2(new_n17987_), .A3(new_n3290_), .ZN(new_n25032_));
  NAND2_X1   g21836(.A1(new_n3290_), .A2(pi0191), .ZN(new_n25033_));
  NAND2_X1   g21837(.A1(new_n5504_), .A2(new_n12167_), .ZN(new_n25034_));
  NOR2_X1    g21838(.A1(new_n24854_), .A2(new_n16751_), .ZN(new_n25035_));
  AOI21_X1   g21839(.A1(new_n25034_), .A2(new_n25035_), .B(pi0038), .ZN(new_n25036_));
  NOR4_X1    g21840(.A1(new_n19135_), .A2(new_n25036_), .A3(new_n25033_), .A4(new_n25017_), .ZN(new_n25037_));
  NAND2_X1   g21841(.A1(new_n25032_), .A2(new_n25037_), .ZN(new_n25038_));
  AOI21_X1   g21842(.A1(new_n25038_), .A2(new_n25015_), .B(new_n17987_), .ZN(new_n25039_));
  NOR2_X1    g21843(.A1(new_n24969_), .A2(new_n13613_), .ZN(new_n25040_));
  XOR2_X1    g21844(.A1(new_n25040_), .A2(new_n13615_), .Z(new_n25041_));
  NAND2_X1   g21845(.A1(new_n25041_), .A2(new_n25039_), .ZN(new_n25042_));
  AOI21_X1   g21846(.A1(new_n25008_), .A2(new_n25002_), .B(pi0608), .ZN(new_n25043_));
  NAND2_X1   g21847(.A1(new_n25005_), .A2(new_n14081_), .ZN(new_n25044_));
  AOI21_X1   g21848(.A1(new_n25042_), .A2(new_n25043_), .B(new_n25044_), .ZN(new_n25045_));
  NOR2_X1    g21849(.A1(new_n24969_), .A2(new_n13614_), .ZN(new_n25046_));
  XOR2_X1    g21850(.A1(new_n25046_), .A2(new_n13615_), .Z(new_n25047_));
  NAND3_X1   g21851(.A1(new_n25047_), .A2(new_n25039_), .A3(pi0778), .ZN(new_n25048_));
  OAI22_X1   g21852(.A1(new_n25045_), .A2(new_n25048_), .B1(pi0778), .B2(new_n25039_), .ZN(new_n25049_));
  NAND3_X1   g21853(.A1(new_n25049_), .A2(pi0609), .A3(pi1155), .ZN(new_n25050_));
  INV_X1     g21854(.I(new_n25049_), .ZN(new_n25051_));
  NAND3_X1   g21855(.A1(new_n25051_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n25052_));
  AOI21_X1   g21856(.A1(new_n25052_), .A2(new_n25050_), .B(new_n25011_), .ZN(new_n25053_));
  NAND2_X1   g21857(.A1(new_n24967_), .A2(pi0660), .ZN(new_n25054_));
  NAND2_X1   g21858(.A1(new_n24973_), .A2(new_n13783_), .ZN(new_n25055_));
  INV_X1     g21859(.I(new_n25055_), .ZN(new_n25056_));
  OAI21_X1   g21860(.A1(new_n25053_), .A2(new_n25054_), .B(new_n25056_), .ZN(new_n25057_));
  AOI21_X1   g21861(.A1(new_n25051_), .A2(pi0609), .B(new_n14694_), .ZN(new_n25058_));
  NOR3_X1    g21862(.A1(new_n25049_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n25059_));
  NOR2_X1    g21863(.A1(new_n25011_), .A2(new_n13801_), .ZN(new_n25060_));
  OAI21_X1   g21864(.A1(new_n25058_), .A2(new_n25059_), .B(new_n25060_), .ZN(new_n25061_));
  INV_X1     g21865(.I(new_n25061_), .ZN(new_n25062_));
  AOI22_X1   g21866(.A1(new_n25057_), .A2(new_n25062_), .B1(new_n13801_), .B2(new_n25049_), .ZN(new_n25063_));
  AOI21_X1   g21867(.A1(new_n25063_), .A2(pi1154), .B(new_n13819_), .ZN(new_n25064_));
  INV_X1     g21868(.I(new_n25063_), .ZN(new_n25065_));
  NOR3_X1    g21869(.A1(new_n25065_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n25066_));
  OAI21_X1   g21870(.A1(new_n25066_), .A2(new_n25064_), .B(new_n25013_), .ZN(new_n25067_));
  NAND2_X1   g21871(.A1(new_n24980_), .A2(pi0627), .ZN(new_n25068_));
  INV_X1     g21872(.I(new_n25068_), .ZN(new_n25069_));
  AOI21_X1   g21873(.A1(new_n25067_), .A2(new_n25069_), .B(new_n13855_), .ZN(new_n25070_));
  NAND3_X1   g21874(.A1(new_n25065_), .A2(pi0618), .A3(pi1154), .ZN(new_n25071_));
  NAND3_X1   g21875(.A1(new_n25063_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n25072_));
  NAND2_X1   g21876(.A1(new_n25071_), .A2(new_n25072_), .ZN(new_n25073_));
  AND2_X2    g21877(.A1(new_n25073_), .A2(new_n25013_), .Z(new_n25074_));
  INV_X1     g21878(.I(new_n24984_), .ZN(new_n25075_));
  NAND3_X1   g21879(.A1(new_n25065_), .A2(new_n19177_), .A3(new_n25075_), .ZN(new_n25076_));
  NOR3_X1    g21880(.A1(new_n25074_), .A2(new_n25070_), .A3(new_n25076_), .ZN(new_n25077_));
  INV_X1     g21881(.I(new_n25070_), .ZN(new_n25078_));
  NOR2_X1    g21882(.A1(new_n25074_), .A2(new_n25076_), .ZN(new_n25079_));
  NOR2_X1    g21883(.A1(new_n25079_), .A2(new_n25078_), .ZN(new_n25080_));
  NOR2_X1    g21884(.A1(new_n25080_), .A2(new_n25077_), .ZN(new_n25081_));
  AOI21_X1   g21885(.A1(new_n25081_), .A2(pi1159), .B(new_n13904_), .ZN(new_n25082_));
  NOR4_X1    g21886(.A1(new_n25080_), .A2(pi0619), .A3(new_n13868_), .A4(new_n25077_), .ZN(new_n25083_));
  OAI21_X1   g21887(.A1(new_n25082_), .A2(new_n25083_), .B(new_n25014_), .ZN(new_n25084_));
  NAND2_X1   g21888(.A1(new_n25084_), .A2(new_n16474_), .ZN(new_n25085_));
  NAND3_X1   g21889(.A1(new_n24989_), .A2(pi0619), .A3(pi1159), .ZN(new_n25086_));
  NAND3_X1   g21890(.A1(new_n24991_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n25087_));
  AOI21_X1   g21891(.A1(new_n25087_), .A2(new_n25086_), .B(new_n24952_), .ZN(new_n25088_));
  NAND4_X1   g21892(.A1(new_n24993_), .A2(new_n25088_), .A3(pi0789), .A4(new_n24989_), .ZN(new_n25089_));
  NOR2_X1    g21893(.A1(new_n24993_), .A2(new_n13896_), .ZN(new_n25090_));
  NAND3_X1   g21894(.A1(new_n25088_), .A2(pi0789), .A3(new_n24989_), .ZN(new_n25091_));
  NAND2_X1   g21895(.A1(new_n25091_), .A2(new_n25090_), .ZN(new_n25092_));
  NAND2_X1   g21896(.A1(new_n25092_), .A2(new_n25089_), .ZN(new_n25093_));
  NAND3_X1   g21897(.A1(new_n25093_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n25094_));
  INV_X1     g21898(.I(new_n25093_), .ZN(new_n25095_));
  NAND3_X1   g21899(.A1(new_n25095_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n25096_));
  AOI21_X1   g21900(.A1(new_n25096_), .A2(new_n25094_), .B(new_n24952_), .ZN(new_n25097_));
  NOR2_X1    g21901(.A1(new_n25014_), .A2(new_n13918_), .ZN(new_n25098_));
  AOI21_X1   g21902(.A1(new_n13918_), .A2(new_n24951_), .B(new_n25098_), .ZN(new_n25099_));
  NOR2_X1    g21903(.A1(new_n25099_), .A2(new_n14162_), .ZN(new_n25100_));
  OAI21_X1   g21904(.A1(new_n25097_), .A2(new_n25100_), .B(new_n19204_), .ZN(new_n25101_));
  NOR2_X1    g21905(.A1(new_n25081_), .A2(pi0789), .ZN(new_n25102_));
  NOR2_X1    g21906(.A1(new_n25093_), .A2(new_n19208_), .ZN(new_n25103_));
  XOR2_X1    g21907(.A1(new_n25103_), .A2(new_n19028_), .Z(new_n25104_));
  NOR4_X1    g21908(.A1(new_n25104_), .A2(new_n15479_), .A3(new_n24952_), .A4(new_n25102_), .ZN(new_n25105_));
  AOI22_X1   g21909(.A1(new_n25085_), .A2(new_n24993_), .B1(new_n25105_), .B2(new_n25101_), .ZN(new_n25106_));
  AOI21_X1   g21910(.A1(new_n25081_), .A2(pi0619), .B(new_n13904_), .ZN(new_n25107_));
  NOR4_X1    g21911(.A1(new_n25080_), .A2(new_n13860_), .A3(pi1159), .A4(new_n25077_), .ZN(new_n25108_));
  OAI21_X1   g21912(.A1(new_n25107_), .A2(new_n25108_), .B(new_n25014_), .ZN(new_n25109_));
  NOR2_X1    g21913(.A1(new_n25088_), .A2(pi0648), .ZN(new_n25110_));
  NAND2_X1   g21914(.A1(new_n25109_), .A2(new_n25110_), .ZN(new_n25111_));
  NOR2_X1    g21915(.A1(new_n24951_), .A2(new_n16372_), .ZN(new_n25112_));
  INV_X1     g21916(.I(new_n25112_), .ZN(new_n25113_));
  NAND3_X1   g21917(.A1(new_n25092_), .A2(new_n16372_), .A3(new_n25089_), .ZN(new_n25114_));
  AOI21_X1   g21918(.A1(new_n25114_), .A2(new_n25113_), .B(new_n13993_), .ZN(new_n25115_));
  NOR2_X1    g21919(.A1(new_n24951_), .A2(new_n13994_), .ZN(new_n25116_));
  OR2_X2     g21920(.A1(new_n25115_), .A2(new_n25116_), .Z(new_n25117_));
  NAND2_X1   g21921(.A1(new_n25099_), .A2(new_n13966_), .ZN(new_n25118_));
  OAI21_X1   g21922(.A1(new_n13966_), .A2(new_n24951_), .B(new_n25118_), .ZN(new_n25119_));
  NAND2_X1   g21923(.A1(new_n25119_), .A2(new_n12777_), .ZN(new_n25120_));
  NOR2_X1    g21924(.A1(new_n24951_), .A2(new_n13942_), .ZN(new_n25121_));
  AOI21_X1   g21925(.A1(new_n25119_), .A2(new_n13942_), .B(new_n25121_), .ZN(new_n25122_));
  NOR2_X1    g21926(.A1(new_n25122_), .A2(pi1156), .ZN(new_n25123_));
  NOR2_X1    g21927(.A1(new_n24951_), .A2(pi0628), .ZN(new_n25124_));
  AOI21_X1   g21928(.A1(new_n25119_), .A2(pi0628), .B(new_n25124_), .ZN(new_n25125_));
  NOR2_X1    g21929(.A1(new_n25125_), .A2(new_n13969_), .ZN(new_n25126_));
  OAI21_X1   g21930(.A1(new_n25123_), .A2(new_n25126_), .B(pi0792), .ZN(new_n25127_));
  NAND2_X1   g21931(.A1(new_n25127_), .A2(new_n25120_), .ZN(new_n25128_));
  NAND2_X1   g21932(.A1(new_n25128_), .A2(new_n14005_), .ZN(new_n25129_));
  NAND2_X1   g21933(.A1(new_n24952_), .A2(pi0647), .ZN(new_n25130_));
  AOI21_X1   g21934(.A1(new_n25129_), .A2(new_n25130_), .B(new_n14012_), .ZN(new_n25131_));
  NOR2_X1    g21935(.A1(new_n24951_), .A2(pi0647), .ZN(new_n25132_));
  AOI21_X1   g21936(.A1(new_n25128_), .A2(pi0647), .B(new_n25132_), .ZN(new_n25133_));
  NAND2_X1   g21937(.A1(new_n25133_), .A2(new_n14206_), .ZN(new_n25134_));
  OR2_X2     g21938(.A1(new_n25131_), .A2(new_n25134_), .Z(new_n25135_));
  NAND2_X1   g21939(.A1(new_n25131_), .A2(new_n25134_), .ZN(new_n25136_));
  AOI21_X1   g21940(.A1(new_n25135_), .A2(new_n25136_), .B(new_n12776_), .ZN(new_n25137_));
  NOR2_X1    g21941(.A1(new_n25137_), .A2(new_n25117_), .ZN(new_n25138_));
  OAI22_X1   g21942(.A1(new_n25106_), .A2(new_n25111_), .B1(new_n16891_), .B2(new_n25138_), .ZN(new_n25139_));
  AOI21_X1   g21943(.A1(new_n25095_), .A2(new_n16372_), .B(new_n25112_), .ZN(new_n25140_));
  NOR2_X1    g21944(.A1(new_n25122_), .A2(new_n15270_), .ZN(new_n25141_));
  NAND2_X1   g21945(.A1(new_n25125_), .A2(new_n13990_), .ZN(new_n25142_));
  XNOR2_X1   g21946(.A1(new_n25141_), .A2(new_n25142_), .ZN(new_n25143_));
  NAND2_X1   g21947(.A1(new_n25143_), .A2(pi0792), .ZN(new_n25144_));
  AOI21_X1   g21948(.A1(new_n25140_), .A2(new_n25144_), .B(new_n16875_), .ZN(new_n25145_));
  NAND2_X1   g21949(.A1(new_n25128_), .A2(new_n12776_), .ZN(new_n25146_));
  AOI21_X1   g21950(.A1(new_n25129_), .A2(new_n25130_), .B(pi1157), .ZN(new_n25147_));
  NOR2_X1    g21951(.A1(new_n25133_), .A2(new_n14006_), .ZN(new_n25148_));
  OAI21_X1   g21952(.A1(new_n25148_), .A2(new_n25147_), .B(pi0787), .ZN(new_n25149_));
  NAND2_X1   g21953(.A1(new_n25149_), .A2(new_n25146_), .ZN(new_n25150_));
  INV_X1     g21954(.I(new_n25150_), .ZN(new_n25151_));
  OAI21_X1   g21955(.A1(new_n25115_), .A2(new_n25116_), .B(new_n14211_), .ZN(new_n25152_));
  NOR2_X1    g21956(.A1(new_n24951_), .A2(new_n14211_), .ZN(new_n25153_));
  INV_X1     g21957(.I(new_n25153_), .ZN(new_n25154_));
  NOR2_X1    g21958(.A1(new_n14243_), .A2(pi0644), .ZN(new_n25155_));
  AOI21_X1   g21959(.A1(new_n25152_), .A2(new_n25154_), .B(new_n25155_), .ZN(new_n25156_));
  AOI21_X1   g21960(.A1(new_n25156_), .A2(pi0715), .B(pi0644), .ZN(new_n25157_));
  AOI21_X1   g21961(.A1(new_n25117_), .A2(new_n14211_), .B(new_n25153_), .ZN(new_n25158_));
  AOI21_X1   g21962(.A1(new_n24951_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n25159_));
  NOR2_X1    g21963(.A1(new_n25159_), .A2(pi0644), .ZN(new_n25160_));
  NOR2_X1    g21964(.A1(new_n25158_), .A2(new_n25160_), .ZN(new_n25161_));
  AOI21_X1   g21965(.A1(new_n25161_), .A2(pi0715), .B(new_n25150_), .ZN(new_n25162_));
  OAI22_X1   g21966(.A1(new_n25162_), .A2(new_n14204_), .B1(new_n25157_), .B2(new_n25151_), .ZN(new_n25163_));
  AOI22_X1   g21967(.A1(new_n25139_), .A2(new_n25145_), .B1(new_n25163_), .B2(new_n19269_), .ZN(new_n25164_));
  NOR3_X1    g21968(.A1(new_n25158_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n25165_));
  NOR3_X1    g21969(.A1(new_n25161_), .A2(pi0644), .A3(new_n12775_), .ZN(new_n25166_));
  NOR2_X1    g21970(.A1(new_n24939_), .A2(pi0790), .ZN(new_n25167_));
  NOR4_X1    g21971(.A1(new_n25158_), .A2(new_n14799_), .A3(new_n25155_), .A4(new_n25167_), .ZN(new_n25168_));
  OAI21_X1   g21972(.A1(new_n25166_), .A2(new_n25165_), .B(new_n25168_), .ZN(new_n25169_));
  OAI21_X1   g21973(.A1(new_n25164_), .A2(new_n25169_), .B(new_n24950_), .ZN(po0348));
  NOR2_X1    g21974(.A1(new_n14652_), .A2(new_n18082_), .ZN(new_n25171_));
  INV_X1     g21975(.I(new_n25171_), .ZN(new_n25172_));
  NOR2_X1    g21976(.A1(new_n9992_), .A2(pi0192), .ZN(new_n25173_));
  NOR2_X1    g21977(.A1(new_n25173_), .A2(pi1153), .ZN(new_n25174_));
  NAND2_X1   g21978(.A1(new_n25172_), .A2(new_n25174_), .ZN(new_n25175_));
  INV_X1     g21979(.I(new_n25175_), .ZN(new_n25176_));
  NOR2_X1    g21980(.A1(new_n25176_), .A2(new_n13748_), .ZN(new_n25177_));
  AOI21_X1   g21981(.A1(new_n13218_), .A2(pi0691), .B(new_n25173_), .ZN(new_n25178_));
  INV_X1     g21982(.I(new_n25178_), .ZN(new_n25179_));
  AOI21_X1   g21983(.A1(new_n25172_), .A2(new_n25179_), .B(new_n13614_), .ZN(new_n25180_));
  INV_X1     g21984(.I(new_n25180_), .ZN(new_n25181_));
  NOR3_X1    g21985(.A1(new_n25181_), .A2(new_n13748_), .A3(new_n25179_), .ZN(new_n25182_));
  XNOR2_X1   g21986(.A1(new_n25182_), .A2(new_n25177_), .ZN(new_n25183_));
  NAND2_X1   g21987(.A1(new_n25183_), .A2(new_n14049_), .ZN(new_n25184_));
  NOR2_X1    g21988(.A1(new_n25184_), .A2(new_n14051_), .ZN(new_n25185_));
  INV_X1     g21989(.I(new_n25185_), .ZN(new_n25186_));
  NOR2_X1    g21990(.A1(new_n25186_), .A2(new_n14163_), .ZN(new_n25187_));
  NAND2_X1   g21991(.A1(new_n25187_), .A2(new_n18929_), .ZN(new_n25188_));
  NOR2_X1    g21992(.A1(new_n25188_), .A2(new_n14060_), .ZN(new_n25189_));
  INV_X1     g21993(.I(new_n25173_), .ZN(new_n25190_));
  NAND3_X1   g21994(.A1(new_n25189_), .A2(pi0647), .A3(pi1157), .ZN(new_n25191_));
  OR3_X2     g21995(.A1(new_n25189_), .A2(new_n14005_), .A3(pi1157), .Z(new_n25192_));
  AOI21_X1   g21996(.A1(new_n25192_), .A2(new_n25191_), .B(new_n25190_), .ZN(new_n25193_));
  INV_X1     g21997(.I(new_n25193_), .ZN(new_n25194_));
  NOR2_X1    g21998(.A1(new_n25190_), .A2(pi0647), .ZN(new_n25195_));
  AOI21_X1   g21999(.A1(new_n25189_), .A2(pi0647), .B(new_n25195_), .ZN(new_n25196_));
  AOI21_X1   g22000(.A1(new_n25196_), .A2(pi1157), .B(new_n12776_), .ZN(new_n25197_));
  AOI22_X1   g22001(.A1(new_n25194_), .A2(new_n25197_), .B1(new_n12776_), .B2(new_n25189_), .ZN(new_n25198_));
  INV_X1     g22002(.I(new_n25198_), .ZN(new_n25199_));
  NOR2_X1    g22003(.A1(new_n13105_), .A2(new_n18051_), .ZN(new_n25200_));
  INV_X1     g22004(.I(new_n25200_), .ZN(new_n25201_));
  NOR2_X1    g22005(.A1(new_n25200_), .A2(new_n25173_), .ZN(new_n25202_));
  INV_X1     g22006(.I(new_n25202_), .ZN(new_n25203_));
  NAND3_X1   g22007(.A1(new_n25203_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n25204_));
  AOI21_X1   g22008(.A1(new_n25204_), .A2(new_n16444_), .B(new_n25201_), .ZN(new_n25205_));
  NOR2_X1    g22009(.A1(new_n25205_), .A2(new_n13801_), .ZN(new_n25206_));
  NOR2_X1    g22010(.A1(new_n25173_), .A2(pi1155), .ZN(new_n25207_));
  NOR3_X1    g22011(.A1(new_n25201_), .A2(new_n16444_), .A3(new_n25207_), .ZN(new_n25208_));
  NAND4_X1   g22012(.A1(new_n25208_), .A2(new_n25203_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n25209_));
  XOR2_X1    g22013(.A1(new_n25206_), .A2(new_n25209_), .Z(new_n25210_));
  NOR2_X1    g22014(.A1(new_n25210_), .A2(new_n13817_), .ZN(new_n25211_));
  OAI21_X1   g22015(.A1(new_n25211_), .A2(pi0618), .B(new_n9992_), .ZN(new_n25212_));
  NAND2_X1   g22016(.A1(new_n25212_), .A2(pi0781), .ZN(new_n25213_));
  OAI21_X1   g22017(.A1(new_n25211_), .A2(new_n9992_), .B(pi0618), .ZN(new_n25214_));
  NOR3_X1    g22018(.A1(new_n25214_), .A2(new_n13855_), .A3(new_n25210_), .ZN(new_n25215_));
  XOR2_X1    g22019(.A1(new_n25215_), .A2(new_n25213_), .Z(new_n25216_));
  NOR2_X1    g22020(.A1(new_n25216_), .A2(new_n13868_), .ZN(new_n25217_));
  OAI21_X1   g22021(.A1(new_n25217_), .A2(pi0619), .B(new_n9992_), .ZN(new_n25218_));
  NAND2_X1   g22022(.A1(new_n25218_), .A2(pi0789), .ZN(new_n25219_));
  OAI21_X1   g22023(.A1(new_n25217_), .A2(new_n9992_), .B(pi0619), .ZN(new_n25220_));
  NOR3_X1    g22024(.A1(new_n25220_), .A2(new_n13896_), .A3(new_n25216_), .ZN(new_n25221_));
  XOR2_X1    g22025(.A1(new_n25221_), .A2(new_n25219_), .Z(new_n25222_));
  NAND2_X1   g22026(.A1(new_n25222_), .A2(new_n16372_), .ZN(new_n25223_));
  OAI21_X1   g22027(.A1(new_n16372_), .A2(new_n25173_), .B(new_n25223_), .ZN(new_n25224_));
  NOR2_X1    g22028(.A1(new_n25224_), .A2(new_n18968_), .ZN(new_n25225_));
  NAND2_X1   g22029(.A1(new_n18967_), .A2(new_n25173_), .ZN(new_n25226_));
  XOR2_X1    g22030(.A1(new_n25225_), .A2(new_n25226_), .Z(new_n25227_));
  AOI21_X1   g22031(.A1(new_n25190_), .A2(new_n14254_), .B(pi0644), .ZN(new_n25228_));
  NAND2_X1   g22032(.A1(new_n25222_), .A2(new_n13962_), .ZN(new_n25229_));
  XOR2_X1    g22033(.A1(new_n25229_), .A2(new_n18976_), .Z(new_n25230_));
  AOI22_X1   g22034(.A1(new_n25230_), .A2(new_n25173_), .B1(new_n16639_), .B2(new_n25187_), .ZN(new_n25231_));
  NOR2_X1    g22035(.A1(new_n25178_), .A2(new_n13203_), .ZN(new_n25232_));
  NAND2_X1   g22036(.A1(new_n25232_), .A2(pi0625), .ZN(new_n25233_));
  NAND3_X1   g22037(.A1(new_n25233_), .A2(pi1153), .A3(new_n25202_), .ZN(new_n25234_));
  NOR2_X1    g22038(.A1(new_n25176_), .A2(new_n14081_), .ZN(new_n25235_));
  AOI21_X1   g22039(.A1(new_n25235_), .A2(new_n25234_), .B(new_n13748_), .ZN(new_n25236_));
  NOR2_X1    g22040(.A1(new_n25203_), .A2(new_n25232_), .ZN(new_n25237_));
  INV_X1     g22041(.I(new_n25233_), .ZN(new_n25238_));
  OAI21_X1   g22042(.A1(new_n25237_), .A2(new_n25238_), .B(new_n25174_), .ZN(new_n25239_));
  NAND4_X1   g22043(.A1(new_n25239_), .A2(new_n13749_), .A3(new_n25181_), .A4(new_n25237_), .ZN(new_n25240_));
  XNOR2_X1   g22044(.A1(new_n25240_), .A2(new_n25236_), .ZN(new_n25241_));
  NAND2_X1   g22045(.A1(new_n25241_), .A2(new_n13801_), .ZN(new_n25242_));
  NOR2_X1    g22046(.A1(new_n25205_), .A2(pi0660), .ZN(new_n25245_));
  NOR2_X1    g22047(.A1(new_n25241_), .A2(new_n13766_), .ZN(new_n25246_));
  XOR2_X1    g22048(.A1(new_n25246_), .A2(new_n14090_), .Z(new_n25247_));
  NOR2_X1    g22049(.A1(new_n25183_), .A2(new_n13801_), .ZN(new_n25248_));
  NAND2_X1   g22050(.A1(new_n25247_), .A2(new_n25248_), .ZN(new_n25249_));
  OAI21_X1   g22051(.A1(new_n25249_), .A2(new_n25245_), .B(new_n25242_), .ZN(new_n25250_));
  NAND2_X1   g22052(.A1(new_n25250_), .A2(new_n13855_), .ZN(new_n25251_));
  INV_X1     g22053(.I(new_n25184_), .ZN(new_n25252_));
  NOR2_X1    g22054(.A1(new_n25250_), .A2(new_n13816_), .ZN(new_n25253_));
  XOR2_X1    g22055(.A1(new_n25253_), .A2(new_n13818_), .Z(new_n25254_));
  NAND2_X1   g22056(.A1(new_n25254_), .A2(new_n25252_), .ZN(new_n25255_));
  NAND3_X1   g22057(.A1(new_n25255_), .A2(new_n13823_), .A3(new_n25214_), .ZN(new_n25256_));
  NAND3_X1   g22058(.A1(new_n25256_), .A2(new_n13823_), .A3(new_n25212_), .ZN(new_n25257_));
  NOR2_X1    g22059(.A1(new_n25250_), .A2(new_n13817_), .ZN(new_n25258_));
  XOR2_X1    g22060(.A1(new_n25258_), .A2(new_n13818_), .Z(new_n25259_));
  NAND4_X1   g22061(.A1(new_n25257_), .A2(pi0781), .A3(new_n25252_), .A4(new_n25259_), .ZN(new_n25260_));
  NAND2_X1   g22062(.A1(new_n25260_), .A2(new_n25251_), .ZN(new_n25261_));
  NOR2_X1    g22063(.A1(new_n25261_), .A2(new_n13860_), .ZN(new_n25262_));
  XOR2_X1    g22064(.A1(new_n25262_), .A2(new_n13904_), .Z(new_n25263_));
  NOR2_X1    g22065(.A1(new_n25263_), .A2(new_n25186_), .ZN(new_n25264_));
  NAND2_X1   g22066(.A1(new_n25220_), .A2(new_n13884_), .ZN(new_n25265_));
  INV_X1     g22067(.I(new_n25261_), .ZN(new_n25266_));
  AOI21_X1   g22068(.A1(new_n25266_), .A2(new_n14143_), .B(pi0789), .ZN(new_n25267_));
  OAI21_X1   g22069(.A1(new_n25264_), .A2(new_n25265_), .B(new_n25267_), .ZN(new_n25268_));
  NOR2_X1    g22070(.A1(new_n25261_), .A2(new_n13868_), .ZN(new_n25269_));
  XOR2_X1    g22071(.A1(new_n25269_), .A2(new_n13903_), .Z(new_n25270_));
  NAND2_X1   g22072(.A1(new_n25218_), .A2(new_n19018_), .ZN(new_n25271_));
  AOI21_X1   g22073(.A1(new_n25270_), .A2(new_n25185_), .B(new_n25271_), .ZN(new_n25272_));
  AOI21_X1   g22074(.A1(new_n25268_), .A2(new_n25272_), .B(new_n25231_), .ZN(new_n25273_));
  NAND3_X1   g22075(.A1(new_n25224_), .A2(new_n18929_), .A3(new_n25187_), .ZN(new_n25274_));
  NAND2_X1   g22076(.A1(new_n25274_), .A2(new_n16569_), .ZN(new_n25275_));
  XOR2_X1    g22077(.A1(new_n25275_), .A2(new_n16572_), .Z(new_n25276_));
  AOI21_X1   g22078(.A1(new_n19022_), .A2(new_n25274_), .B(new_n25276_), .ZN(new_n25277_));
  NAND2_X1   g22079(.A1(new_n25222_), .A2(new_n13963_), .ZN(new_n25278_));
  XNOR2_X1   g22080(.A1(new_n25278_), .A2(new_n19028_), .ZN(new_n25279_));
  NOR3_X1    g22081(.A1(new_n25279_), .A2(new_n16424_), .A3(new_n25190_), .ZN(new_n25280_));
  OAI21_X1   g22082(.A1(new_n25277_), .A2(new_n16574_), .B(new_n25280_), .ZN(new_n25281_));
  NOR2_X1    g22083(.A1(new_n25224_), .A2(new_n13994_), .ZN(new_n25282_));
  XNOR2_X1   g22084(.A1(new_n25282_), .A2(new_n19033_), .ZN(new_n25283_));
  AOI22_X1   g22085(.A1(new_n25283_), .A2(new_n25173_), .B1(new_n14206_), .B2(new_n25196_), .ZN(new_n25284_));
  NOR3_X1    g22086(.A1(new_n25284_), .A2(new_n14010_), .A3(new_n25194_), .ZN(new_n25285_));
  OAI22_X1   g22087(.A1(new_n25273_), .A2(new_n25281_), .B1(new_n12776_), .B2(new_n25285_), .ZN(new_n25286_));
  NAND2_X1   g22088(.A1(new_n25286_), .A2(pi0644), .ZN(new_n25287_));
  XOR2_X1    g22089(.A1(new_n25287_), .A2(new_n14205_), .Z(new_n25288_));
  NOR2_X1    g22090(.A1(new_n25288_), .A2(new_n25198_), .ZN(new_n25289_));
  NAND2_X1   g22091(.A1(new_n25227_), .A2(pi0715), .ZN(new_n25290_));
  XOR2_X1    g22092(.A1(new_n25290_), .A2(new_n14205_), .Z(new_n25291_));
  OAI21_X1   g22093(.A1(new_n25291_), .A2(new_n25190_), .B(new_n19043_), .ZN(new_n25292_));
  OAI22_X1   g22094(.A1(new_n25289_), .A2(new_n25292_), .B1(new_n25227_), .B2(new_n25228_), .ZN(new_n25293_));
  NAND2_X1   g22095(.A1(new_n25286_), .A2(pi0715), .ZN(new_n25294_));
  XOR2_X1    g22096(.A1(new_n25294_), .A2(new_n14217_), .Z(new_n25295_));
  AOI21_X1   g22097(.A1(po1038), .A2(new_n12450_), .B(pi0832), .ZN(new_n25296_));
  NAND4_X1   g22098(.A1(new_n25293_), .A2(new_n25199_), .A3(new_n25295_), .A4(new_n25296_), .ZN(new_n25297_));
  NOR2_X1    g22099(.A1(new_n14428_), .A2(pi0192), .ZN(new_n25298_));
  INV_X1     g22100(.I(new_n25298_), .ZN(new_n25299_));
  OAI22_X1   g22101(.A1(new_n17127_), .A2(new_n12450_), .B1(new_n18051_), .B2(new_n19052_), .ZN(new_n25300_));
  OAI21_X1   g22102(.A1(pi0192), .A2(new_n14299_), .B(new_n14301_), .ZN(new_n25301_));
  NAND2_X1   g22103(.A1(new_n14299_), .A2(pi0764), .ZN(new_n25302_));
  NAND4_X1   g22104(.A1(new_n25301_), .A2(new_n18051_), .A3(new_n14362_), .A4(new_n25302_), .ZN(new_n25303_));
  NAND3_X1   g22105(.A1(new_n25303_), .A2(pi0038), .A3(pi0192), .ZN(new_n25304_));
  NAND2_X1   g22106(.A1(new_n25304_), .A2(new_n3183_), .ZN(new_n25305_));
  NAND2_X1   g22107(.A1(new_n13109_), .A2(new_n12450_), .ZN(new_n25306_));
  NAND4_X1   g22108(.A1(new_n25305_), .A2(pi0038), .A3(new_n25300_), .A4(new_n25306_), .ZN(new_n25307_));
  AOI21_X1   g22109(.A1(new_n25307_), .A2(new_n18051_), .B(new_n13107_), .ZN(new_n25308_));
  NAND2_X1   g22110(.A1(new_n25308_), .A2(new_n3289_), .ZN(new_n25309_));
  NAND2_X1   g22111(.A1(new_n3290_), .A2(new_n12450_), .ZN(new_n25310_));
  NAND3_X1   g22112(.A1(new_n25309_), .A2(new_n13776_), .A3(new_n25310_), .ZN(new_n25311_));
  NAND2_X1   g22113(.A1(new_n25299_), .A2(new_n13780_), .ZN(new_n25312_));
  NAND2_X1   g22114(.A1(new_n25311_), .A2(new_n25312_), .ZN(new_n25313_));
  NAND2_X1   g22115(.A1(new_n25313_), .A2(pi0609), .ZN(new_n25314_));
  NAND2_X1   g22116(.A1(new_n25314_), .A2(pi0785), .ZN(new_n25315_));
  NAND2_X1   g22117(.A1(new_n25309_), .A2(new_n25310_), .ZN(new_n25316_));
  NOR2_X1    g22118(.A1(new_n25299_), .A2(new_n13776_), .ZN(new_n25317_));
  AOI21_X1   g22119(.A1(new_n25316_), .A2(new_n13776_), .B(new_n25317_), .ZN(new_n25318_));
  AOI21_X1   g22120(.A1(new_n25299_), .A2(new_n14467_), .B(pi0609), .ZN(new_n25319_));
  OR2_X2     g22121(.A1(new_n25311_), .A2(new_n25319_), .Z(new_n25320_));
  NOR3_X1    g22122(.A1(new_n25320_), .A2(new_n13801_), .A3(new_n25318_), .ZN(new_n25321_));
  XNOR2_X1   g22123(.A1(new_n25321_), .A2(new_n25315_), .ZN(new_n25322_));
  NAND3_X1   g22124(.A1(new_n25322_), .A2(pi0618), .A3(pi1154), .ZN(new_n25323_));
  XOR2_X1    g22125(.A1(new_n25321_), .A2(new_n25315_), .Z(new_n25324_));
  NAND3_X1   g22126(.A1(new_n25324_), .A2(pi0618), .A3(new_n13819_), .ZN(new_n25325_));
  NAND2_X1   g22127(.A1(new_n25323_), .A2(new_n25325_), .ZN(new_n25326_));
  NAND2_X1   g22128(.A1(new_n25326_), .A2(new_n25298_), .ZN(new_n25327_));
  NAND2_X1   g22129(.A1(new_n25327_), .A2(pi0781), .ZN(new_n25328_));
  NAND3_X1   g22130(.A1(new_n25322_), .A2(pi0618), .A3(pi1154), .ZN(new_n25329_));
  NAND3_X1   g22131(.A1(new_n25324_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n25330_));
  AOI21_X1   g22132(.A1(new_n25329_), .A2(new_n25330_), .B(new_n25299_), .ZN(new_n25331_));
  NOR2_X1    g22133(.A1(new_n25324_), .A2(new_n13855_), .ZN(new_n25332_));
  NAND3_X1   g22134(.A1(new_n25328_), .A2(new_n25331_), .A3(new_n25332_), .ZN(new_n25333_));
  NAND2_X1   g22135(.A1(new_n25331_), .A2(new_n25332_), .ZN(new_n25334_));
  NAND3_X1   g22136(.A1(new_n25334_), .A2(new_n25327_), .A3(pi0781), .ZN(new_n25335_));
  NAND2_X1   g22137(.A1(new_n25333_), .A2(new_n25335_), .ZN(new_n25336_));
  NAND3_X1   g22138(.A1(new_n25336_), .A2(pi0619), .A3(pi1159), .ZN(new_n25337_));
  INV_X1     g22139(.I(new_n25336_), .ZN(new_n25338_));
  NAND3_X1   g22140(.A1(new_n25338_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n25339_));
  AOI21_X1   g22141(.A1(new_n25339_), .A2(new_n25337_), .B(new_n25299_), .ZN(new_n25340_));
  NAND2_X1   g22142(.A1(new_n25299_), .A2(new_n13879_), .ZN(new_n25341_));
  OAI21_X1   g22143(.A1(new_n13721_), .A2(new_n18082_), .B(new_n12450_), .ZN(new_n25342_));
  NAND2_X1   g22144(.A1(new_n25342_), .A2(new_n13108_), .ZN(new_n25343_));
  NAND2_X1   g22145(.A1(new_n12450_), .A2(new_n18082_), .ZN(new_n25344_));
  NAND4_X1   g22146(.A1(new_n13634_), .A2(pi0192), .A3(new_n3290_), .A4(new_n25344_), .ZN(new_n25345_));
  NOR3_X1    g22147(.A1(new_n14424_), .A2(new_n3259_), .A3(new_n12450_), .ZN(new_n25346_));
  NOR3_X1    g22148(.A1(new_n14422_), .A2(pi0038), .A3(new_n12450_), .ZN(new_n25347_));
  OAI21_X1   g22149(.A1(new_n25346_), .A2(new_n25347_), .B(new_n15655_), .ZN(new_n25348_));
  AOI21_X1   g22150(.A1(new_n25343_), .A2(new_n25345_), .B(new_n25348_), .ZN(new_n25349_));
  NOR2_X1    g22151(.A1(new_n25298_), .A2(new_n13613_), .ZN(new_n25350_));
  XOR2_X1    g22152(.A1(new_n25350_), .A2(new_n13615_), .Z(new_n25351_));
  NAND2_X1   g22153(.A1(new_n25351_), .A2(new_n25349_), .ZN(new_n25352_));
  NAND2_X1   g22154(.A1(new_n25352_), .A2(pi0778), .ZN(new_n25353_));
  NOR2_X1    g22155(.A1(new_n25298_), .A2(new_n13614_), .ZN(new_n25354_));
  XOR2_X1    g22156(.A1(new_n25354_), .A2(new_n13615_), .Z(new_n25355_));
  NAND3_X1   g22157(.A1(new_n25355_), .A2(pi0778), .A3(new_n25349_), .ZN(new_n25356_));
  XOR2_X1    g22158(.A1(new_n25353_), .A2(new_n25356_), .Z(new_n25357_));
  INV_X1     g22159(.I(new_n25357_), .ZN(new_n25358_));
  NAND2_X1   g22160(.A1(new_n25298_), .A2(new_n13803_), .ZN(new_n25359_));
  OAI21_X1   g22161(.A1(new_n25358_), .A2(new_n13803_), .B(new_n25359_), .ZN(new_n25360_));
  OAI21_X1   g22162(.A1(new_n25360_), .A2(new_n13879_), .B(new_n25341_), .ZN(new_n25361_));
  INV_X1     g22163(.I(new_n25308_), .ZN(new_n25362_));
  NOR2_X1    g22164(.A1(new_n12450_), .A2(new_n18051_), .ZN(new_n25363_));
  INV_X1     g22165(.I(new_n25363_), .ZN(new_n25364_));
  NAND2_X1   g22166(.A1(new_n13461_), .A2(pi0764), .ZN(new_n25365_));
  XOR2_X1    g22167(.A1(new_n25365_), .A2(new_n25364_), .Z(new_n25366_));
  NAND2_X1   g22168(.A1(new_n25366_), .A2(new_n13521_), .ZN(new_n25367_));
  NAND3_X1   g22169(.A1(new_n14270_), .A2(pi0192), .A3(pi0764), .ZN(new_n25368_));
  NAND3_X1   g22170(.A1(new_n14272_), .A2(pi0192), .A3(new_n18051_), .ZN(new_n25369_));
  AOI21_X1   g22171(.A1(new_n25368_), .A2(new_n25369_), .B(new_n13152_), .ZN(new_n25370_));
  NAND3_X1   g22172(.A1(new_n13198_), .A2(pi0192), .A3(pi0764), .ZN(new_n25371_));
  NAND3_X1   g22173(.A1(new_n13200_), .A2(new_n12450_), .A3(pi0764), .ZN(new_n25372_));
  AOI21_X1   g22174(.A1(new_n25372_), .A2(new_n25371_), .B(new_n13191_), .ZN(new_n25373_));
  OAI21_X1   g22175(.A1(new_n25370_), .A2(new_n3212_), .B(new_n25373_), .ZN(new_n25374_));
  NAND3_X1   g22176(.A1(new_n25367_), .A2(new_n3183_), .A3(new_n25374_), .ZN(new_n25375_));
  NOR2_X1    g22177(.A1(new_n14284_), .A2(new_n12450_), .ZN(new_n25376_));
  XOR2_X1    g22178(.A1(new_n25376_), .A2(new_n25363_), .Z(new_n25377_));
  NAND3_X1   g22179(.A1(new_n25375_), .A2(new_n25377_), .A3(new_n13359_), .ZN(new_n25378_));
  NAND3_X1   g22180(.A1(new_n25378_), .A2(new_n18082_), .A3(new_n3290_), .ZN(new_n25379_));
  NAND2_X1   g22181(.A1(new_n3290_), .A2(pi0192), .ZN(new_n25380_));
  NAND2_X1   g22182(.A1(new_n5504_), .A2(new_n12450_), .ZN(new_n25381_));
  NOR2_X1    g22183(.A1(new_n25201_), .A2(new_n16751_), .ZN(new_n25382_));
  AOI21_X1   g22184(.A1(new_n25381_), .A2(new_n25382_), .B(pi0038), .ZN(new_n25383_));
  NOR4_X1    g22185(.A1(new_n19135_), .A2(new_n25383_), .A3(new_n25380_), .A4(new_n25364_), .ZN(new_n25384_));
  NAND2_X1   g22186(.A1(new_n25379_), .A2(new_n25384_), .ZN(new_n25385_));
  AOI21_X1   g22187(.A1(new_n25385_), .A2(new_n25362_), .B(new_n18082_), .ZN(new_n25386_));
  NOR2_X1    g22188(.A1(new_n25316_), .A2(new_n13613_), .ZN(new_n25387_));
  XOR2_X1    g22189(.A1(new_n25387_), .A2(new_n13615_), .Z(new_n25388_));
  NAND2_X1   g22190(.A1(new_n25388_), .A2(new_n25386_), .ZN(new_n25389_));
  AOI21_X1   g22191(.A1(new_n25355_), .A2(new_n25349_), .B(pi0608), .ZN(new_n25390_));
  NAND2_X1   g22192(.A1(new_n25352_), .A2(new_n14081_), .ZN(new_n25391_));
  AOI21_X1   g22193(.A1(new_n25389_), .A2(new_n25390_), .B(new_n25391_), .ZN(new_n25392_));
  NOR2_X1    g22194(.A1(new_n25316_), .A2(new_n13614_), .ZN(new_n25393_));
  XOR2_X1    g22195(.A1(new_n25393_), .A2(new_n13615_), .Z(new_n25394_));
  NAND3_X1   g22196(.A1(new_n25394_), .A2(new_n25386_), .A3(pi0778), .ZN(new_n25395_));
  OAI22_X1   g22197(.A1(new_n25392_), .A2(new_n25395_), .B1(pi0778), .B2(new_n25386_), .ZN(new_n25396_));
  NAND3_X1   g22198(.A1(new_n25396_), .A2(pi0609), .A3(pi1155), .ZN(new_n25397_));
  INV_X1     g22199(.I(new_n25396_), .ZN(new_n25398_));
  NAND3_X1   g22200(.A1(new_n25398_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n25399_));
  AOI21_X1   g22201(.A1(new_n25399_), .A2(new_n25397_), .B(new_n25358_), .ZN(new_n25400_));
  NAND2_X1   g22202(.A1(new_n25314_), .A2(pi0660), .ZN(new_n25401_));
  NAND2_X1   g22203(.A1(new_n25320_), .A2(new_n13783_), .ZN(new_n25402_));
  INV_X1     g22204(.I(new_n25402_), .ZN(new_n25403_));
  OAI21_X1   g22205(.A1(new_n25400_), .A2(new_n25401_), .B(new_n25403_), .ZN(new_n25404_));
  AOI21_X1   g22206(.A1(new_n25398_), .A2(pi0609), .B(new_n14694_), .ZN(new_n25405_));
  NOR3_X1    g22207(.A1(new_n25396_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n25406_));
  NOR2_X1    g22208(.A1(new_n25358_), .A2(new_n13801_), .ZN(new_n25407_));
  OAI21_X1   g22209(.A1(new_n25405_), .A2(new_n25406_), .B(new_n25407_), .ZN(new_n25408_));
  INV_X1     g22210(.I(new_n25408_), .ZN(new_n25409_));
  AOI22_X1   g22211(.A1(new_n25404_), .A2(new_n25409_), .B1(new_n13801_), .B2(new_n25396_), .ZN(new_n25410_));
  AOI21_X1   g22212(.A1(new_n25410_), .A2(pi1154), .B(new_n13819_), .ZN(new_n25411_));
  INV_X1     g22213(.I(new_n25410_), .ZN(new_n25412_));
  NOR3_X1    g22214(.A1(new_n25412_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n25413_));
  OAI21_X1   g22215(.A1(new_n25413_), .A2(new_n25411_), .B(new_n25360_), .ZN(new_n25414_));
  NAND2_X1   g22216(.A1(new_n25327_), .A2(pi0627), .ZN(new_n25415_));
  INV_X1     g22217(.I(new_n25415_), .ZN(new_n25416_));
  AOI21_X1   g22218(.A1(new_n25414_), .A2(new_n25416_), .B(new_n13855_), .ZN(new_n25417_));
  NAND3_X1   g22219(.A1(new_n25412_), .A2(pi0618), .A3(pi1154), .ZN(new_n25418_));
  NAND3_X1   g22220(.A1(new_n25410_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n25419_));
  NAND2_X1   g22221(.A1(new_n25418_), .A2(new_n25419_), .ZN(new_n25420_));
  AND2_X2    g22222(.A1(new_n25420_), .A2(new_n25360_), .Z(new_n25421_));
  INV_X1     g22223(.I(new_n25331_), .ZN(new_n25422_));
  NAND3_X1   g22224(.A1(new_n25412_), .A2(new_n19177_), .A3(new_n25422_), .ZN(new_n25423_));
  NOR3_X1    g22225(.A1(new_n25421_), .A2(new_n25417_), .A3(new_n25423_), .ZN(new_n25424_));
  INV_X1     g22226(.I(new_n25417_), .ZN(new_n25425_));
  NOR2_X1    g22227(.A1(new_n25421_), .A2(new_n25423_), .ZN(new_n25426_));
  NOR2_X1    g22228(.A1(new_n25426_), .A2(new_n25425_), .ZN(new_n25427_));
  NOR2_X1    g22229(.A1(new_n25427_), .A2(new_n25424_), .ZN(new_n25428_));
  AOI21_X1   g22230(.A1(new_n25428_), .A2(pi1159), .B(new_n13904_), .ZN(new_n25429_));
  NOR4_X1    g22231(.A1(new_n25427_), .A2(pi0619), .A3(new_n13868_), .A4(new_n25424_), .ZN(new_n25430_));
  OAI21_X1   g22232(.A1(new_n25429_), .A2(new_n25430_), .B(new_n25361_), .ZN(new_n25431_));
  NAND2_X1   g22233(.A1(new_n25431_), .A2(new_n16474_), .ZN(new_n25432_));
  NAND3_X1   g22234(.A1(new_n25336_), .A2(pi0619), .A3(pi1159), .ZN(new_n25433_));
  NAND3_X1   g22235(.A1(new_n25338_), .A2(pi1159), .A3(new_n13904_), .ZN(new_n25434_));
  AOI21_X1   g22236(.A1(new_n25434_), .A2(new_n25433_), .B(new_n25299_), .ZN(new_n25435_));
  NAND4_X1   g22237(.A1(new_n25340_), .A2(new_n25435_), .A3(pi0789), .A4(new_n25336_), .ZN(new_n25436_));
  NOR2_X1    g22238(.A1(new_n25340_), .A2(new_n13896_), .ZN(new_n25437_));
  NAND3_X1   g22239(.A1(new_n25435_), .A2(pi0789), .A3(new_n25336_), .ZN(new_n25438_));
  NAND2_X1   g22240(.A1(new_n25438_), .A2(new_n25437_), .ZN(new_n25439_));
  NAND2_X1   g22241(.A1(new_n25439_), .A2(new_n25436_), .ZN(new_n25440_));
  NAND3_X1   g22242(.A1(new_n25440_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n25441_));
  INV_X1     g22243(.I(new_n25440_), .ZN(new_n25442_));
  NAND3_X1   g22244(.A1(new_n25442_), .A2(new_n13962_), .A3(new_n18976_), .ZN(new_n25443_));
  AOI21_X1   g22245(.A1(new_n25443_), .A2(new_n25441_), .B(new_n25299_), .ZN(new_n25444_));
  NOR2_X1    g22246(.A1(new_n25361_), .A2(new_n13918_), .ZN(new_n25445_));
  AOI21_X1   g22247(.A1(new_n13918_), .A2(new_n25298_), .B(new_n25445_), .ZN(new_n25446_));
  NOR2_X1    g22248(.A1(new_n25446_), .A2(new_n14162_), .ZN(new_n25447_));
  OAI21_X1   g22249(.A1(new_n25444_), .A2(new_n25447_), .B(new_n19204_), .ZN(new_n25448_));
  NOR2_X1    g22250(.A1(new_n25428_), .A2(pi0789), .ZN(new_n25449_));
  NOR2_X1    g22251(.A1(new_n25440_), .A2(new_n19208_), .ZN(new_n25450_));
  XOR2_X1    g22252(.A1(new_n25450_), .A2(new_n19028_), .Z(new_n25451_));
  NOR4_X1    g22253(.A1(new_n25451_), .A2(new_n15479_), .A3(new_n25299_), .A4(new_n25449_), .ZN(new_n25452_));
  AOI22_X1   g22254(.A1(new_n25432_), .A2(new_n25340_), .B1(new_n25452_), .B2(new_n25448_), .ZN(new_n25453_));
  AOI21_X1   g22255(.A1(new_n25428_), .A2(pi0619), .B(new_n13904_), .ZN(new_n25454_));
  NOR4_X1    g22256(.A1(new_n25427_), .A2(new_n13860_), .A3(pi1159), .A4(new_n25424_), .ZN(new_n25455_));
  OAI21_X1   g22257(.A1(new_n25454_), .A2(new_n25455_), .B(new_n25361_), .ZN(new_n25456_));
  NOR2_X1    g22258(.A1(new_n25435_), .A2(pi0648), .ZN(new_n25457_));
  NAND2_X1   g22259(.A1(new_n25456_), .A2(new_n25457_), .ZN(new_n25458_));
  NOR2_X1    g22260(.A1(new_n25298_), .A2(new_n16372_), .ZN(new_n25459_));
  INV_X1     g22261(.I(new_n25459_), .ZN(new_n25460_));
  NAND3_X1   g22262(.A1(new_n25439_), .A2(new_n16372_), .A3(new_n25436_), .ZN(new_n25461_));
  AOI21_X1   g22263(.A1(new_n25461_), .A2(new_n25460_), .B(new_n13993_), .ZN(new_n25462_));
  NOR2_X1    g22264(.A1(new_n25298_), .A2(new_n13994_), .ZN(new_n25463_));
  OR2_X2     g22265(.A1(new_n25462_), .A2(new_n25463_), .Z(new_n25464_));
  NAND2_X1   g22266(.A1(new_n25446_), .A2(new_n13966_), .ZN(new_n25465_));
  OAI21_X1   g22267(.A1(new_n13966_), .A2(new_n25298_), .B(new_n25465_), .ZN(new_n25466_));
  NAND2_X1   g22268(.A1(new_n25466_), .A2(new_n12777_), .ZN(new_n25467_));
  NOR2_X1    g22269(.A1(new_n25298_), .A2(new_n13942_), .ZN(new_n25468_));
  AOI21_X1   g22270(.A1(new_n25466_), .A2(new_n13942_), .B(new_n25468_), .ZN(new_n25469_));
  NOR2_X1    g22271(.A1(new_n25469_), .A2(pi1156), .ZN(new_n25470_));
  NOR2_X1    g22272(.A1(new_n25298_), .A2(pi0628), .ZN(new_n25471_));
  AOI21_X1   g22273(.A1(new_n25466_), .A2(pi0628), .B(new_n25471_), .ZN(new_n25472_));
  NOR2_X1    g22274(.A1(new_n25472_), .A2(new_n13969_), .ZN(new_n25473_));
  OAI21_X1   g22275(.A1(new_n25470_), .A2(new_n25473_), .B(pi0792), .ZN(new_n25474_));
  NAND2_X1   g22276(.A1(new_n25474_), .A2(new_n25467_), .ZN(new_n25475_));
  NAND2_X1   g22277(.A1(new_n25475_), .A2(new_n14005_), .ZN(new_n25476_));
  NAND2_X1   g22278(.A1(new_n25299_), .A2(pi0647), .ZN(new_n25477_));
  AOI21_X1   g22279(.A1(new_n25476_), .A2(new_n25477_), .B(new_n14012_), .ZN(new_n25478_));
  NOR2_X1    g22280(.A1(new_n25298_), .A2(pi0647), .ZN(new_n25479_));
  AOI21_X1   g22281(.A1(new_n25475_), .A2(pi0647), .B(new_n25479_), .ZN(new_n25480_));
  NAND2_X1   g22282(.A1(new_n25480_), .A2(new_n14206_), .ZN(new_n25481_));
  OR2_X2     g22283(.A1(new_n25478_), .A2(new_n25481_), .Z(new_n25482_));
  NAND2_X1   g22284(.A1(new_n25478_), .A2(new_n25481_), .ZN(new_n25483_));
  AOI21_X1   g22285(.A1(new_n25482_), .A2(new_n25483_), .B(new_n12776_), .ZN(new_n25484_));
  NOR2_X1    g22286(.A1(new_n25484_), .A2(new_n25464_), .ZN(new_n25485_));
  OAI22_X1   g22287(.A1(new_n25453_), .A2(new_n25458_), .B1(new_n16891_), .B2(new_n25485_), .ZN(new_n25486_));
  AOI21_X1   g22288(.A1(new_n25442_), .A2(new_n16372_), .B(new_n25459_), .ZN(new_n25487_));
  NOR2_X1    g22289(.A1(new_n25469_), .A2(new_n15270_), .ZN(new_n25488_));
  NAND2_X1   g22290(.A1(new_n25472_), .A2(new_n13990_), .ZN(new_n25489_));
  XNOR2_X1   g22291(.A1(new_n25488_), .A2(new_n25489_), .ZN(new_n25490_));
  NAND2_X1   g22292(.A1(new_n25490_), .A2(pi0792), .ZN(new_n25491_));
  AOI21_X1   g22293(.A1(new_n25487_), .A2(new_n25491_), .B(new_n16875_), .ZN(new_n25492_));
  NAND2_X1   g22294(.A1(new_n25475_), .A2(new_n12776_), .ZN(new_n25493_));
  AOI21_X1   g22295(.A1(new_n25476_), .A2(new_n25477_), .B(pi1157), .ZN(new_n25494_));
  NOR2_X1    g22296(.A1(new_n25480_), .A2(new_n14006_), .ZN(new_n25495_));
  OAI21_X1   g22297(.A1(new_n25495_), .A2(new_n25494_), .B(pi0787), .ZN(new_n25496_));
  NAND2_X1   g22298(.A1(new_n25496_), .A2(new_n25493_), .ZN(new_n25497_));
  INV_X1     g22299(.I(new_n25497_), .ZN(new_n25498_));
  OAI21_X1   g22300(.A1(new_n25462_), .A2(new_n25463_), .B(new_n14211_), .ZN(new_n25499_));
  NOR2_X1    g22301(.A1(new_n25298_), .A2(new_n14211_), .ZN(new_n25500_));
  INV_X1     g22302(.I(new_n25500_), .ZN(new_n25501_));
  NOR2_X1    g22303(.A1(new_n14243_), .A2(pi0644), .ZN(new_n25502_));
  AOI21_X1   g22304(.A1(new_n25499_), .A2(new_n25501_), .B(new_n25502_), .ZN(new_n25503_));
  AOI21_X1   g22305(.A1(new_n25503_), .A2(pi0715), .B(pi0644), .ZN(new_n25504_));
  AOI21_X1   g22306(.A1(new_n25464_), .A2(new_n14211_), .B(new_n25500_), .ZN(new_n25505_));
  AOI21_X1   g22307(.A1(new_n25298_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n25506_));
  NOR2_X1    g22308(.A1(new_n25506_), .A2(pi0644), .ZN(new_n25507_));
  NOR2_X1    g22309(.A1(new_n25505_), .A2(new_n25507_), .ZN(new_n25508_));
  AOI21_X1   g22310(.A1(new_n25508_), .A2(pi0715), .B(new_n25497_), .ZN(new_n25509_));
  OAI22_X1   g22311(.A1(new_n25509_), .A2(new_n14204_), .B1(new_n25504_), .B2(new_n25498_), .ZN(new_n25510_));
  AOI22_X1   g22312(.A1(new_n25486_), .A2(new_n25492_), .B1(new_n25510_), .B2(new_n19269_), .ZN(new_n25511_));
  NOR3_X1    g22313(.A1(new_n25505_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n25512_));
  NOR3_X1    g22314(.A1(new_n25508_), .A2(pi0644), .A3(new_n12775_), .ZN(new_n25513_));
  NOR2_X1    g22315(.A1(new_n25286_), .A2(pi0790), .ZN(new_n25514_));
  NOR4_X1    g22316(.A1(new_n25505_), .A2(new_n14799_), .A3(new_n25502_), .A4(new_n25514_), .ZN(new_n25515_));
  OAI21_X1   g22317(.A1(new_n25513_), .A2(new_n25512_), .B(new_n25515_), .ZN(new_n25516_));
  OAI21_X1   g22318(.A1(new_n25511_), .A2(new_n25516_), .B(new_n25297_), .ZN(po0349));
  NAND2_X1   g22319(.A1(new_n13627_), .A2(new_n7342_), .ZN(new_n25518_));
  INV_X1     g22320(.I(new_n25518_), .ZN(new_n25519_));
  NOR2_X1    g22321(.A1(new_n25519_), .A2(new_n13966_), .ZN(new_n25520_));
  NOR2_X1    g22322(.A1(new_n25518_), .A2(new_n13919_), .ZN(new_n25521_));
  NOR2_X1    g22323(.A1(new_n25519_), .A2(new_n13880_), .ZN(new_n25522_));
  OAI21_X1   g22324(.A1(new_n13721_), .A2(new_n18129_), .B(new_n7342_), .ZN(new_n25523_));
  NAND2_X1   g22325(.A1(new_n16715_), .A2(new_n7342_), .ZN(new_n25524_));
  NAND4_X1   g22326(.A1(new_n15655_), .A2(new_n13108_), .A3(new_n25523_), .A4(new_n25524_), .ZN(new_n25525_));
  NAND2_X1   g22327(.A1(new_n25525_), .A2(new_n14424_), .ZN(new_n25526_));
  NAND2_X1   g22328(.A1(new_n25526_), .A2(pi0193), .ZN(new_n25527_));
  OAI21_X1   g22329(.A1(new_n25527_), .A2(new_n25518_), .B(new_n18129_), .ZN(new_n25528_));
  NAND2_X1   g22330(.A1(new_n25528_), .A2(new_n3289_), .ZN(new_n25529_));
  NAND2_X1   g22331(.A1(new_n25529_), .A2(pi0625), .ZN(new_n25530_));
  XOR2_X1    g22332(.A1(new_n25530_), .A2(new_n13620_), .Z(new_n25531_));
  NAND2_X1   g22333(.A1(new_n25531_), .A2(new_n25519_), .ZN(new_n25532_));
  NAND2_X1   g22334(.A1(new_n25532_), .A2(pi0778), .ZN(new_n25533_));
  NAND2_X1   g22335(.A1(new_n25529_), .A2(pi1153), .ZN(new_n25534_));
  XOR2_X1    g22336(.A1(new_n25534_), .A2(new_n13620_), .Z(new_n25535_));
  NAND2_X1   g22337(.A1(new_n25535_), .A2(new_n25519_), .ZN(new_n25536_));
  NOR3_X1    g22338(.A1(new_n25536_), .A2(new_n13748_), .A3(new_n25529_), .ZN(new_n25537_));
  XNOR2_X1   g22339(.A1(new_n25537_), .A2(new_n25533_), .ZN(new_n25538_));
  INV_X1     g22340(.I(new_n25538_), .ZN(new_n25539_));
  NAND2_X1   g22341(.A1(new_n25519_), .A2(new_n13803_), .ZN(new_n25540_));
  OAI21_X1   g22342(.A1(new_n25539_), .A2(new_n13803_), .B(new_n25540_), .ZN(new_n25541_));
  INV_X1     g22343(.I(new_n25541_), .ZN(new_n25542_));
  AOI21_X1   g22344(.A1(new_n25542_), .A2(new_n13880_), .B(new_n25522_), .ZN(new_n25543_));
  AOI21_X1   g22345(.A1(new_n25543_), .A2(new_n13919_), .B(new_n25521_), .ZN(new_n25544_));
  AOI21_X1   g22346(.A1(new_n25544_), .A2(new_n13966_), .B(new_n25520_), .ZN(new_n25545_));
  INV_X1     g22347(.I(new_n25545_), .ZN(new_n25546_));
  NAND3_X1   g22348(.A1(new_n25546_), .A2(pi0628), .A3(pi1156), .ZN(new_n25547_));
  NAND3_X1   g22349(.A1(new_n25545_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n25548_));
  AOI21_X1   g22350(.A1(new_n25547_), .A2(new_n25548_), .B(new_n25518_), .ZN(new_n25549_));
  NAND3_X1   g22351(.A1(new_n25546_), .A2(pi0628), .A3(pi1156), .ZN(new_n25550_));
  NAND3_X1   g22352(.A1(new_n25545_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n25551_));
  AOI21_X1   g22353(.A1(new_n25550_), .A2(new_n25551_), .B(new_n25518_), .ZN(new_n25552_));
  NAND4_X1   g22354(.A1(new_n25552_), .A2(new_n25549_), .A3(pi0792), .A4(new_n25546_), .ZN(new_n25553_));
  NOR2_X1    g22355(.A1(new_n25549_), .A2(new_n12777_), .ZN(new_n25554_));
  NAND3_X1   g22356(.A1(new_n25552_), .A2(pi0792), .A3(new_n25546_), .ZN(new_n25555_));
  NAND2_X1   g22357(.A1(new_n25555_), .A2(new_n25554_), .ZN(new_n25556_));
  NAND2_X1   g22358(.A1(new_n25556_), .A2(new_n25553_), .ZN(new_n25557_));
  NAND2_X1   g22359(.A1(new_n25519_), .A2(new_n14005_), .ZN(new_n25558_));
  NAND2_X1   g22360(.A1(new_n25558_), .A2(pi1157), .ZN(new_n25559_));
  AOI21_X1   g22361(.A1(new_n25557_), .A2(pi0647), .B(new_n25559_), .ZN(new_n25560_));
  AOI21_X1   g22362(.A1(new_n25556_), .A2(new_n25553_), .B(pi0647), .ZN(new_n25561_));
  NOR2_X1    g22363(.A1(new_n25518_), .A2(new_n14005_), .ZN(new_n25562_));
  NOR3_X1    g22364(.A1(new_n25561_), .A2(pi1157), .A3(new_n25562_), .ZN(new_n25563_));
  OAI21_X1   g22365(.A1(new_n25563_), .A2(new_n25560_), .B(pi0787), .ZN(new_n25564_));
  OAI21_X1   g22366(.A1(pi0787), .A2(new_n25557_), .B(new_n25564_), .ZN(new_n25565_));
  NOR2_X1    g22367(.A1(new_n25519_), .A2(new_n16372_), .ZN(new_n25566_));
  INV_X1     g22368(.I(new_n25566_), .ZN(new_n25567_));
  AOI21_X1   g22369(.A1(new_n7342_), .A2(new_n18095_), .B(pi0038), .ZN(new_n25568_));
  NAND2_X1   g22370(.A1(new_n13097_), .A2(new_n25568_), .ZN(new_n25569_));
  OAI22_X1   g22371(.A1(new_n7342_), .A2(new_n13107_), .B1(new_n13109_), .B2(new_n18095_), .ZN(new_n25570_));
  NAND2_X1   g22372(.A1(new_n25570_), .A2(pi0038), .ZN(new_n25571_));
  NAND2_X1   g22373(.A1(new_n25569_), .A2(new_n25571_), .ZN(new_n25572_));
  NAND2_X1   g22374(.A1(new_n3290_), .A2(new_n7342_), .ZN(new_n25573_));
  OAI21_X1   g22375(.A1(new_n25572_), .A2(new_n3290_), .B(new_n25573_), .ZN(new_n25574_));
  INV_X1     g22376(.I(new_n25574_), .ZN(new_n25575_));
  NAND2_X1   g22377(.A1(new_n25575_), .A2(new_n13776_), .ZN(new_n25576_));
  OAI21_X1   g22378(.A1(new_n15147_), .A2(new_n25519_), .B(new_n25576_), .ZN(new_n25577_));
  NAND2_X1   g22379(.A1(new_n25577_), .A2(pi0609), .ZN(new_n25578_));
  NAND2_X1   g22380(.A1(new_n25578_), .A2(pi0785), .ZN(new_n25579_));
  AOI21_X1   g22381(.A1(new_n25518_), .A2(new_n14467_), .B(pi0609), .ZN(new_n25580_));
  NOR2_X1    g22382(.A1(new_n25576_), .A2(new_n25580_), .ZN(new_n25581_));
  NAND2_X1   g22383(.A1(new_n25574_), .A2(new_n13776_), .ZN(new_n25582_));
  OAI21_X1   g22384(.A1(new_n13776_), .A2(new_n25518_), .B(new_n25582_), .ZN(new_n25583_));
  NAND3_X1   g22385(.A1(new_n25581_), .A2(new_n25583_), .A3(pi0785), .ZN(new_n25584_));
  XNOR2_X1   g22386(.A1(new_n25579_), .A2(new_n25584_), .ZN(new_n25585_));
  NAND2_X1   g22387(.A1(new_n25585_), .A2(pi0618), .ZN(new_n25586_));
  XOR2_X1    g22388(.A1(new_n25586_), .A2(new_n13819_), .Z(new_n25587_));
  NAND2_X1   g22389(.A1(new_n25587_), .A2(new_n25519_), .ZN(new_n25588_));
  NAND2_X1   g22390(.A1(new_n25588_), .A2(pi0781), .ZN(new_n25589_));
  NAND2_X1   g22391(.A1(new_n25585_), .A2(pi1154), .ZN(new_n25590_));
  XOR2_X1    g22392(.A1(new_n25590_), .A2(new_n13819_), .Z(new_n25591_));
  NAND2_X1   g22393(.A1(new_n25591_), .A2(new_n25519_), .ZN(new_n25592_));
  NOR3_X1    g22394(.A1(new_n25592_), .A2(new_n13855_), .A3(new_n25585_), .ZN(new_n25593_));
  XNOR2_X1   g22395(.A1(new_n25593_), .A2(new_n25589_), .ZN(new_n25594_));
  NOR2_X1    g22396(.A1(new_n25594_), .A2(new_n13860_), .ZN(new_n25595_));
  NOR2_X1    g22397(.A1(new_n25595_), .A2(new_n13904_), .ZN(new_n25596_));
  INV_X1     g22398(.I(new_n25596_), .ZN(new_n25597_));
  NAND2_X1   g22399(.A1(new_n25595_), .A2(new_n13904_), .ZN(new_n25598_));
  AOI21_X1   g22400(.A1(new_n25597_), .A2(new_n25598_), .B(new_n25518_), .ZN(new_n25599_));
  NAND3_X1   g22401(.A1(new_n25594_), .A2(pi0619), .A3(pi1159), .ZN(new_n25600_));
  NOR2_X1    g22402(.A1(new_n25594_), .A2(new_n13868_), .ZN(new_n25601_));
  NAND2_X1   g22403(.A1(new_n25601_), .A2(new_n13904_), .ZN(new_n25602_));
  AOI21_X1   g22404(.A1(new_n25602_), .A2(new_n25600_), .B(new_n25518_), .ZN(new_n25603_));
  NAND4_X1   g22405(.A1(new_n25599_), .A2(new_n25603_), .A3(pi0789), .A4(new_n25594_), .ZN(new_n25604_));
  INV_X1     g22406(.I(new_n25598_), .ZN(new_n25605_));
  OAI21_X1   g22407(.A1(new_n25605_), .A2(new_n25596_), .B(new_n25519_), .ZN(new_n25606_));
  NAND3_X1   g22408(.A1(new_n25603_), .A2(pi0789), .A3(new_n25594_), .ZN(new_n25607_));
  NAND3_X1   g22409(.A1(new_n25607_), .A2(pi0789), .A3(new_n25606_), .ZN(new_n25608_));
  NAND3_X1   g22410(.A1(new_n25608_), .A2(new_n25604_), .A3(new_n16372_), .ZN(new_n25609_));
  AOI21_X1   g22411(.A1(new_n25609_), .A2(new_n25567_), .B(new_n13993_), .ZN(new_n25610_));
  NOR2_X1    g22412(.A1(new_n25519_), .A2(new_n13994_), .ZN(new_n25611_));
  OAI21_X1   g22413(.A1(new_n25610_), .A2(new_n25611_), .B(new_n14211_), .ZN(new_n25612_));
  INV_X1     g22414(.I(new_n25612_), .ZN(new_n25613_));
  NOR2_X1    g22415(.A1(new_n25519_), .A2(new_n14211_), .ZN(new_n25614_));
  NOR2_X1    g22416(.A1(new_n14243_), .A2(pi0644), .ZN(new_n25615_));
  INV_X1     g22417(.I(new_n25615_), .ZN(new_n25616_));
  OAI21_X1   g22418(.A1(new_n25613_), .A2(new_n25614_), .B(new_n25616_), .ZN(new_n25617_));
  OAI21_X1   g22419(.A1(new_n25617_), .A2(new_n14200_), .B(new_n14204_), .ZN(new_n25618_));
  NAND2_X1   g22420(.A1(new_n25618_), .A2(new_n25565_), .ZN(new_n25619_));
  NOR2_X1    g22421(.A1(new_n25613_), .A2(new_n25614_), .ZN(new_n25620_));
  AOI21_X1   g22422(.A1(new_n25519_), .A2(new_n14204_), .B(new_n14255_), .ZN(new_n25621_));
  NOR2_X1    g22423(.A1(new_n25621_), .A2(pi0644), .ZN(new_n25622_));
  NOR3_X1    g22424(.A1(new_n25620_), .A2(new_n14200_), .A3(new_n25622_), .ZN(new_n25623_));
  OAI21_X1   g22425(.A1(new_n25623_), .A2(new_n25565_), .B(pi0644), .ZN(new_n25624_));
  AOI21_X1   g22426(.A1(new_n25624_), .A2(new_n25619_), .B(new_n12775_), .ZN(new_n25625_));
  INV_X1     g22427(.I(new_n25614_), .ZN(new_n25626_));
  AOI21_X1   g22428(.A1(new_n25612_), .A2(new_n25626_), .B(new_n25622_), .ZN(new_n25627_));
  NAND3_X1   g22429(.A1(new_n25627_), .A2(pi0644), .A3(pi0790), .ZN(new_n25628_));
  OR3_X2     g22430(.A1(new_n25627_), .A2(new_n12775_), .A3(new_n19379_), .Z(new_n25629_));
  AOI21_X1   g22431(.A1(new_n25629_), .A2(new_n25628_), .B(new_n25617_), .ZN(new_n25630_));
  NAND2_X1   g22432(.A1(new_n25557_), .A2(pi0647), .ZN(new_n25631_));
  OR2_X2     g22433(.A1(new_n25561_), .A2(new_n25562_), .Z(new_n25632_));
  NAND4_X1   g22434(.A1(new_n25631_), .A2(new_n14010_), .A3(pi1157), .A4(new_n25558_), .ZN(new_n25634_));
  NAND2_X1   g22435(.A1(new_n25560_), .A2(new_n14010_), .ZN(new_n25635_));
  NAND3_X1   g22436(.A1(new_n25635_), .A2(new_n25632_), .A3(new_n14011_), .ZN(new_n25636_));
  AOI21_X1   g22437(.A1(new_n25636_), .A2(new_n25634_), .B(new_n12776_), .ZN(new_n25637_));
  NOR3_X1    g22438(.A1(new_n25637_), .A2(new_n25610_), .A3(new_n25611_), .ZN(new_n25638_));
  NOR2_X1    g22439(.A1(new_n25638_), .A2(new_n16867_), .ZN(new_n25639_));
  NOR3_X1    g22440(.A1(new_n25625_), .A2(new_n25639_), .A3(new_n25630_), .ZN(new_n25640_));
  NOR2_X1    g22441(.A1(new_n7342_), .A2(new_n18095_), .ZN(new_n25641_));
  INV_X1     g22442(.I(new_n25641_), .ZN(new_n25642_));
  NOR2_X1    g22443(.A1(new_n14284_), .A2(new_n7342_), .ZN(new_n25643_));
  XOR2_X1    g22444(.A1(new_n25643_), .A2(new_n25642_), .Z(new_n25644_));
  NAND2_X1   g22445(.A1(new_n13461_), .A2(pi0739), .ZN(new_n25645_));
  XOR2_X1    g22446(.A1(new_n25645_), .A2(new_n25641_), .Z(new_n25646_));
  NOR2_X1    g22447(.A1(new_n25646_), .A2(new_n14262_), .ZN(new_n25647_));
  NOR2_X1    g22448(.A1(new_n13198_), .A2(new_n18095_), .ZN(new_n25648_));
  XOR2_X1    g22449(.A1(new_n25648_), .A2(new_n25641_), .Z(new_n25649_));
  AOI21_X1   g22450(.A1(new_n25649_), .A2(new_n13190_), .B(new_n3262_), .ZN(new_n25650_));
  AOI21_X1   g22451(.A1(new_n14272_), .A2(pi0193), .B(new_n25642_), .ZN(new_n25651_));
  NOR3_X1    g22452(.A1(new_n14270_), .A2(new_n7342_), .A3(pi0739), .ZN(new_n25652_));
  OAI21_X1   g22453(.A1(new_n25651_), .A2(new_n25652_), .B(new_n14269_), .ZN(new_n25653_));
  OAI21_X1   g22454(.A1(new_n25653_), .A2(new_n25650_), .B(new_n3183_), .ZN(new_n25654_));
  OAI21_X1   g22455(.A1(new_n25647_), .A2(new_n25654_), .B(new_n13359_), .ZN(new_n25655_));
  NOR2_X1    g22456(.A1(new_n3289_), .A2(pi0690), .ZN(new_n25656_));
  OAI21_X1   g22457(.A1(new_n25655_), .A2(new_n25644_), .B(new_n25656_), .ZN(new_n25657_));
  NAND2_X1   g22458(.A1(new_n5504_), .A2(new_n7342_), .ZN(new_n25658_));
  NOR2_X1    g22459(.A1(new_n13105_), .A2(new_n18095_), .ZN(new_n25659_));
  INV_X1     g22460(.I(new_n25659_), .ZN(new_n25660_));
  NOR2_X1    g22461(.A1(new_n25660_), .A2(new_n16751_), .ZN(new_n25661_));
  AOI21_X1   g22462(.A1(new_n25658_), .A2(new_n25661_), .B(pi0038), .ZN(new_n25662_));
  NOR4_X1    g22463(.A1(new_n19135_), .A2(new_n25662_), .A3(new_n3289_), .A4(new_n25642_), .ZN(new_n25663_));
  NAND2_X1   g22464(.A1(new_n25657_), .A2(new_n25663_), .ZN(new_n25664_));
  AOI22_X1   g22465(.A1(new_n25664_), .A2(new_n18129_), .B1(new_n25569_), .B2(new_n25571_), .ZN(new_n25665_));
  INV_X1     g22466(.I(new_n25665_), .ZN(new_n25666_));
  NAND3_X1   g22467(.A1(new_n25665_), .A2(pi0625), .A3(pi1153), .ZN(new_n25667_));
  OR3_X2     g22468(.A1(new_n25665_), .A2(new_n13613_), .A3(new_n13615_), .Z(new_n25668_));
  NAND2_X1   g22469(.A1(new_n25668_), .A2(new_n25667_), .ZN(new_n25669_));
  NAND2_X1   g22470(.A1(new_n25669_), .A2(new_n25574_), .ZN(new_n25670_));
  NAND3_X1   g22471(.A1(new_n25670_), .A2(new_n14081_), .A3(new_n25536_), .ZN(new_n25671_));
  NOR2_X1    g22472(.A1(new_n25665_), .A2(new_n13614_), .ZN(new_n25672_));
  XOR2_X1    g22473(.A1(new_n25672_), .A2(new_n13615_), .Z(new_n25673_));
  AOI21_X1   g22474(.A1(new_n25673_), .A2(new_n25574_), .B(pi0608), .ZN(new_n25674_));
  NAND2_X1   g22475(.A1(new_n25671_), .A2(new_n25674_), .ZN(new_n25675_));
  NOR2_X1    g22476(.A1(new_n25532_), .A2(new_n13748_), .ZN(new_n25676_));
  AOI22_X1   g22477(.A1(new_n25675_), .A2(new_n25676_), .B1(new_n13748_), .B2(new_n25666_), .ZN(new_n25677_));
  AOI21_X1   g22478(.A1(new_n25677_), .A2(pi1155), .B(new_n14694_), .ZN(new_n25678_));
  INV_X1     g22479(.I(new_n25678_), .ZN(new_n25679_));
  NAND3_X1   g22480(.A1(new_n25677_), .A2(pi1155), .A3(new_n14694_), .ZN(new_n25680_));
  AOI21_X1   g22481(.A1(new_n25679_), .A2(new_n25680_), .B(new_n25539_), .ZN(new_n25681_));
  NAND2_X1   g22482(.A1(new_n25578_), .A2(pi0660), .ZN(new_n25682_));
  NOR2_X1    g22483(.A1(new_n25581_), .A2(pi0660), .ZN(new_n25683_));
  OAI21_X1   g22484(.A1(new_n25681_), .A2(new_n25682_), .B(new_n25683_), .ZN(new_n25684_));
  INV_X1     g22485(.I(new_n25684_), .ZN(new_n25685_));
  INV_X1     g22486(.I(new_n25677_), .ZN(new_n25686_));
  NAND3_X1   g22487(.A1(new_n25686_), .A2(pi0609), .A3(pi1155), .ZN(new_n25687_));
  NAND3_X1   g22488(.A1(new_n25677_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n25688_));
  NAND2_X1   g22489(.A1(new_n25687_), .A2(new_n25688_), .ZN(new_n25689_));
  NOR2_X1    g22490(.A1(new_n25539_), .A2(new_n13801_), .ZN(new_n25690_));
  NAND2_X1   g22491(.A1(new_n25689_), .A2(new_n25690_), .ZN(new_n25691_));
  OAI22_X1   g22492(.A1(new_n25685_), .A2(new_n25691_), .B1(pi0785), .B2(new_n25677_), .ZN(new_n25692_));
  NAND3_X1   g22493(.A1(new_n25692_), .A2(pi0618), .A3(pi1154), .ZN(new_n25693_));
  INV_X1     g22494(.I(new_n25691_), .ZN(new_n25694_));
  AOI22_X1   g22495(.A1(new_n25694_), .A2(new_n25684_), .B1(new_n13801_), .B2(new_n25686_), .ZN(new_n25695_));
  NAND3_X1   g22496(.A1(new_n25695_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n25696_));
  AOI21_X1   g22497(.A1(new_n25693_), .A2(new_n25696_), .B(new_n25542_), .ZN(new_n25697_));
  NAND2_X1   g22498(.A1(new_n25588_), .A2(pi0627), .ZN(new_n25698_));
  OAI21_X1   g22499(.A1(new_n25697_), .A2(new_n25698_), .B(pi0781), .ZN(new_n25699_));
  NAND3_X1   g22500(.A1(new_n25692_), .A2(pi0618), .A3(pi1154), .ZN(new_n25700_));
  NAND3_X1   g22501(.A1(new_n25695_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n25701_));
  NAND2_X1   g22502(.A1(new_n25700_), .A2(new_n25701_), .ZN(new_n25702_));
  NAND3_X1   g22503(.A1(new_n25692_), .A2(new_n19177_), .A3(new_n25592_), .ZN(new_n25703_));
  AOI21_X1   g22504(.A1(new_n25702_), .A2(new_n25541_), .B(new_n25703_), .ZN(new_n25704_));
  NAND2_X1   g22505(.A1(new_n25699_), .A2(new_n25704_), .ZN(new_n25705_));
  AOI21_X1   g22506(.A1(new_n25695_), .A2(pi1154), .B(new_n13819_), .ZN(new_n25706_));
  NOR3_X1    g22507(.A1(new_n25692_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n25707_));
  OAI21_X1   g22508(.A1(new_n25707_), .A2(new_n25706_), .B(new_n25541_), .ZN(new_n25708_));
  INV_X1     g22509(.I(new_n25698_), .ZN(new_n25709_));
  AOI21_X1   g22510(.A1(new_n25708_), .A2(new_n25709_), .B(new_n13855_), .ZN(new_n25710_));
  AOI21_X1   g22511(.A1(new_n25695_), .A2(pi0618), .B(new_n13819_), .ZN(new_n25711_));
  NOR3_X1    g22512(.A1(new_n25692_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n25712_));
  OAI21_X1   g22513(.A1(new_n25712_), .A2(new_n25711_), .B(new_n25541_), .ZN(new_n25713_));
  INV_X1     g22514(.I(new_n25703_), .ZN(new_n25714_));
  NAND2_X1   g22515(.A1(new_n25713_), .A2(new_n25714_), .ZN(new_n25715_));
  NAND2_X1   g22516(.A1(new_n25710_), .A2(new_n25715_), .ZN(new_n25716_));
  NAND2_X1   g22517(.A1(new_n25716_), .A2(new_n25705_), .ZN(new_n25717_));
  NAND3_X1   g22518(.A1(new_n25717_), .A2(pi0619), .A3(pi1159), .ZN(new_n25718_));
  NAND4_X1   g22519(.A1(new_n25716_), .A2(new_n25705_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n25719_));
  AOI21_X1   g22520(.A1(new_n25718_), .A2(new_n25719_), .B(new_n25543_), .ZN(new_n25720_));
  OAI21_X1   g22521(.A1(new_n25720_), .A2(new_n20003_), .B(new_n25599_), .ZN(new_n25721_));
  NAND2_X1   g22522(.A1(new_n25717_), .A2(new_n13896_), .ZN(new_n25722_));
  NAND2_X1   g22523(.A1(new_n25608_), .A2(new_n25604_), .ZN(new_n25723_));
  NAND3_X1   g22524(.A1(new_n25723_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n25724_));
  NAND4_X1   g22525(.A1(new_n25608_), .A2(new_n25604_), .A3(new_n13901_), .A4(new_n13962_), .ZN(new_n25725_));
  AOI21_X1   g22526(.A1(new_n25724_), .A2(new_n25725_), .B(new_n25518_), .ZN(new_n25726_));
  NOR2_X1    g22527(.A1(new_n25544_), .A2(new_n14162_), .ZN(new_n25727_));
  OAI21_X1   g22528(.A1(new_n25726_), .A2(new_n25727_), .B(new_n19204_), .ZN(new_n25728_));
  NOR2_X1    g22529(.A1(new_n25723_), .A2(new_n19208_), .ZN(new_n25729_));
  XNOR2_X1   g22530(.A1(new_n25729_), .A2(new_n19028_), .ZN(new_n25730_));
  NOR2_X1    g22531(.A1(new_n25518_), .A2(new_n15479_), .ZN(new_n25731_));
  NAND4_X1   g22532(.A1(new_n25722_), .A2(new_n25728_), .A3(new_n25730_), .A4(new_n25731_), .ZN(new_n25732_));
  NOR2_X1    g22533(.A1(new_n25710_), .A2(new_n25715_), .ZN(new_n25733_));
  NOR2_X1    g22534(.A1(new_n25699_), .A2(new_n25704_), .ZN(new_n25734_));
  NOR3_X1    g22535(.A1(new_n25733_), .A2(new_n25734_), .A3(new_n13860_), .ZN(new_n25735_));
  NOR2_X1    g22536(.A1(new_n25735_), .A2(new_n13904_), .ZN(new_n25736_));
  NOR4_X1    g22537(.A1(new_n25733_), .A2(new_n25734_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n25737_));
  NOR2_X1    g22538(.A1(new_n25736_), .A2(new_n25737_), .ZN(new_n25738_));
  NOR3_X1    g22539(.A1(new_n25603_), .A2(pi0648), .A3(new_n16419_), .ZN(new_n25739_));
  OAI21_X1   g22540(.A1(new_n25738_), .A2(new_n25543_), .B(new_n25739_), .ZN(new_n25740_));
  AOI21_X1   g22541(.A1(new_n25721_), .A2(new_n25732_), .B(new_n25740_), .ZN(new_n25741_));
  NOR2_X1    g22542(.A1(new_n25549_), .A2(new_n13976_), .ZN(new_n25742_));
  NOR2_X1    g22543(.A1(new_n25552_), .A2(pi0629), .ZN(new_n25743_));
  NOR2_X1    g22544(.A1(new_n25743_), .A2(new_n25742_), .ZN(new_n25744_));
  AOI21_X1   g22545(.A1(new_n25609_), .A2(new_n25567_), .B(new_n16874_), .ZN(new_n25745_));
  NOR2_X1    g22546(.A1(new_n14652_), .A2(new_n18129_), .ZN(new_n25746_));
  INV_X1     g22547(.I(new_n25746_), .ZN(new_n25747_));
  NOR2_X1    g22548(.A1(new_n9992_), .A2(pi0193), .ZN(new_n25748_));
  NOR2_X1    g22549(.A1(new_n25748_), .A2(pi1153), .ZN(new_n25749_));
  NAND2_X1   g22550(.A1(new_n25747_), .A2(new_n25749_), .ZN(new_n25750_));
  INV_X1     g22551(.I(new_n25750_), .ZN(new_n25751_));
  NOR2_X1    g22552(.A1(new_n25751_), .A2(new_n13748_), .ZN(new_n25752_));
  AOI21_X1   g22553(.A1(new_n13218_), .A2(pi0690), .B(new_n25748_), .ZN(new_n25753_));
  INV_X1     g22554(.I(new_n25753_), .ZN(new_n25754_));
  AOI21_X1   g22555(.A1(new_n25747_), .A2(new_n25754_), .B(new_n13614_), .ZN(new_n25755_));
  INV_X1     g22556(.I(new_n25755_), .ZN(new_n25756_));
  NOR3_X1    g22557(.A1(new_n25756_), .A2(new_n13748_), .A3(new_n25754_), .ZN(new_n25757_));
  XNOR2_X1   g22558(.A1(new_n25757_), .A2(new_n25752_), .ZN(new_n25758_));
  NAND2_X1   g22559(.A1(new_n25758_), .A2(new_n14049_), .ZN(new_n25759_));
  NOR2_X1    g22560(.A1(new_n25759_), .A2(new_n14051_), .ZN(new_n25760_));
  INV_X1     g22561(.I(new_n25760_), .ZN(new_n25761_));
  NOR4_X1    g22562(.A1(new_n25761_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n25762_));
  NOR2_X1    g22563(.A1(new_n25762_), .A2(new_n14005_), .ZN(new_n25763_));
  XOR2_X1    g22564(.A1(new_n25763_), .A2(new_n14007_), .Z(new_n25764_));
  NAND2_X1   g22565(.A1(new_n25764_), .A2(new_n25748_), .ZN(new_n25765_));
  INV_X1     g22566(.I(new_n25748_), .ZN(new_n25766_));
  NOR2_X1    g22567(.A1(new_n25766_), .A2(pi0647), .ZN(new_n25767_));
  AOI21_X1   g22568(.A1(new_n25762_), .A2(pi0647), .B(new_n25767_), .ZN(new_n25768_));
  AOI21_X1   g22569(.A1(new_n25768_), .A2(pi1157), .B(new_n12776_), .ZN(new_n25769_));
  AOI22_X1   g22570(.A1(new_n25765_), .A2(new_n25769_), .B1(new_n12776_), .B2(new_n25762_), .ZN(new_n25770_));
  NOR2_X1    g22571(.A1(new_n25761_), .A2(new_n14163_), .ZN(new_n25771_));
  NOR2_X1    g22572(.A1(new_n25659_), .A2(new_n25748_), .ZN(new_n25772_));
  INV_X1     g22573(.I(new_n25772_), .ZN(new_n25773_));
  NAND3_X1   g22574(.A1(new_n25773_), .A2(pi1155), .A3(new_n18184_), .ZN(new_n25774_));
  AOI21_X1   g22575(.A1(new_n25774_), .A2(new_n16444_), .B(new_n25660_), .ZN(new_n25775_));
  NOR2_X1    g22576(.A1(new_n25775_), .A2(new_n13801_), .ZN(new_n25776_));
  NOR2_X1    g22577(.A1(new_n25748_), .A2(pi1155), .ZN(new_n25777_));
  NOR3_X1    g22578(.A1(new_n25660_), .A2(new_n16444_), .A3(new_n25777_), .ZN(new_n25778_));
  NAND4_X1   g22579(.A1(new_n25778_), .A2(new_n25773_), .A3(pi0785), .A4(new_n18184_), .ZN(new_n25779_));
  XOR2_X1    g22580(.A1(new_n25776_), .A2(new_n25779_), .Z(new_n25780_));
  NOR2_X1    g22581(.A1(new_n25780_), .A2(new_n13817_), .ZN(new_n25781_));
  OAI21_X1   g22582(.A1(new_n25781_), .A2(pi0618), .B(new_n9992_), .ZN(new_n25782_));
  NAND2_X1   g22583(.A1(new_n25782_), .A2(pi0781), .ZN(new_n25783_));
  OAI21_X1   g22584(.A1(new_n25781_), .A2(new_n9992_), .B(pi0618), .ZN(new_n25784_));
  NOR3_X1    g22585(.A1(new_n25784_), .A2(new_n13855_), .A3(new_n25780_), .ZN(new_n25785_));
  XOR2_X1    g22586(.A1(new_n25785_), .A2(new_n25783_), .Z(new_n25786_));
  NOR2_X1    g22587(.A1(new_n25786_), .A2(new_n13868_), .ZN(new_n25787_));
  OAI21_X1   g22588(.A1(new_n25787_), .A2(pi0619), .B(new_n9992_), .ZN(new_n25788_));
  NAND2_X1   g22589(.A1(new_n25788_), .A2(pi0789), .ZN(new_n25789_));
  OAI21_X1   g22590(.A1(new_n25787_), .A2(new_n9992_), .B(pi0619), .ZN(new_n25790_));
  NOR3_X1    g22591(.A1(new_n25790_), .A2(new_n13896_), .A3(new_n25786_), .ZN(new_n25791_));
  XOR2_X1    g22592(.A1(new_n25791_), .A2(new_n25789_), .Z(new_n25792_));
  NAND2_X1   g22593(.A1(new_n25792_), .A2(new_n13962_), .ZN(new_n25793_));
  XOR2_X1    g22594(.A1(new_n25793_), .A2(new_n18976_), .Z(new_n25794_));
  AOI22_X1   g22595(.A1(new_n25794_), .A2(new_n25748_), .B1(new_n16639_), .B2(new_n25771_), .ZN(new_n25795_));
  NOR2_X1    g22596(.A1(new_n25753_), .A2(new_n13203_), .ZN(new_n25796_));
  NAND2_X1   g22597(.A1(new_n25796_), .A2(pi0625), .ZN(new_n25797_));
  NAND3_X1   g22598(.A1(new_n25797_), .A2(pi1153), .A3(new_n25772_), .ZN(new_n25798_));
  NOR2_X1    g22599(.A1(new_n25751_), .A2(new_n14081_), .ZN(new_n25799_));
  AOI21_X1   g22600(.A1(new_n25799_), .A2(new_n25798_), .B(new_n13748_), .ZN(new_n25800_));
  NOR2_X1    g22601(.A1(new_n25773_), .A2(new_n25796_), .ZN(new_n25801_));
  INV_X1     g22602(.I(new_n25797_), .ZN(new_n25802_));
  OAI21_X1   g22603(.A1(new_n25801_), .A2(new_n25802_), .B(new_n25749_), .ZN(new_n25803_));
  NAND4_X1   g22604(.A1(new_n25803_), .A2(new_n13749_), .A3(new_n25756_), .A4(new_n25801_), .ZN(new_n25804_));
  XNOR2_X1   g22605(.A1(new_n25804_), .A2(new_n25800_), .ZN(new_n25805_));
  NAND2_X1   g22606(.A1(new_n25805_), .A2(new_n13801_), .ZN(new_n25806_));
  NOR2_X1    g22607(.A1(new_n25775_), .A2(pi0660), .ZN(new_n25810_));
  NOR2_X1    g22608(.A1(new_n25805_), .A2(new_n13766_), .ZN(new_n25811_));
  XOR2_X1    g22609(.A1(new_n25811_), .A2(new_n14090_), .Z(new_n25812_));
  NOR2_X1    g22610(.A1(new_n25758_), .A2(new_n13801_), .ZN(new_n25813_));
  NAND2_X1   g22611(.A1(new_n25812_), .A2(new_n25813_), .ZN(new_n25814_));
  OAI21_X1   g22612(.A1(new_n25814_), .A2(new_n25810_), .B(new_n25806_), .ZN(new_n25815_));
  NAND2_X1   g22613(.A1(new_n25815_), .A2(new_n13855_), .ZN(new_n25816_));
  INV_X1     g22614(.I(new_n25759_), .ZN(new_n25817_));
  NOR2_X1    g22615(.A1(new_n25815_), .A2(new_n13816_), .ZN(new_n25818_));
  XOR2_X1    g22616(.A1(new_n25818_), .A2(new_n13818_), .Z(new_n25819_));
  NAND2_X1   g22617(.A1(new_n25819_), .A2(new_n25817_), .ZN(new_n25820_));
  NAND3_X1   g22618(.A1(new_n25820_), .A2(new_n13823_), .A3(new_n25784_), .ZN(new_n25821_));
  NAND3_X1   g22619(.A1(new_n25821_), .A2(new_n13823_), .A3(new_n25782_), .ZN(new_n25822_));
  NOR2_X1    g22620(.A1(new_n25815_), .A2(new_n13817_), .ZN(new_n25823_));
  XOR2_X1    g22621(.A1(new_n25823_), .A2(new_n13818_), .Z(new_n25824_));
  NAND4_X1   g22622(.A1(new_n25822_), .A2(pi0781), .A3(new_n25817_), .A4(new_n25824_), .ZN(new_n25825_));
  NAND2_X1   g22623(.A1(new_n25825_), .A2(new_n25816_), .ZN(new_n25826_));
  NOR2_X1    g22624(.A1(new_n25826_), .A2(new_n13860_), .ZN(new_n25827_));
  XOR2_X1    g22625(.A1(new_n25827_), .A2(new_n13904_), .Z(new_n25828_));
  NOR2_X1    g22626(.A1(new_n25828_), .A2(new_n25761_), .ZN(new_n25829_));
  NAND2_X1   g22627(.A1(new_n25790_), .A2(new_n13884_), .ZN(new_n25830_));
  INV_X1     g22628(.I(new_n25826_), .ZN(new_n25831_));
  AOI21_X1   g22629(.A1(new_n25831_), .A2(new_n14143_), .B(pi0789), .ZN(new_n25832_));
  OAI21_X1   g22630(.A1(new_n25829_), .A2(new_n25830_), .B(new_n25832_), .ZN(new_n25833_));
  NOR2_X1    g22631(.A1(new_n25826_), .A2(new_n13868_), .ZN(new_n25834_));
  XOR2_X1    g22632(.A1(new_n25834_), .A2(new_n13903_), .Z(new_n25835_));
  NAND2_X1   g22633(.A1(new_n25788_), .A2(new_n19018_), .ZN(new_n25836_));
  AOI21_X1   g22634(.A1(new_n25835_), .A2(new_n25760_), .B(new_n25836_), .ZN(new_n25837_));
  AOI21_X1   g22635(.A1(new_n25833_), .A2(new_n25837_), .B(new_n25795_), .ZN(new_n25838_));
  NAND2_X1   g22636(.A1(new_n25792_), .A2(new_n16372_), .ZN(new_n25839_));
  OAI21_X1   g22637(.A1(new_n16372_), .A2(new_n25748_), .B(new_n25839_), .ZN(new_n25840_));
  NAND3_X1   g22638(.A1(new_n25840_), .A2(new_n18929_), .A3(new_n25771_), .ZN(new_n25841_));
  NAND2_X1   g22639(.A1(new_n25841_), .A2(new_n16569_), .ZN(new_n25842_));
  XOR2_X1    g22640(.A1(new_n25842_), .A2(new_n16572_), .Z(new_n25843_));
  AOI21_X1   g22641(.A1(new_n19022_), .A2(new_n25841_), .B(new_n25843_), .ZN(new_n25844_));
  NAND2_X1   g22642(.A1(new_n25792_), .A2(new_n13963_), .ZN(new_n25845_));
  XNOR2_X1   g22643(.A1(new_n25845_), .A2(new_n19028_), .ZN(new_n25846_));
  NOR3_X1    g22644(.A1(new_n25846_), .A2(new_n16424_), .A3(new_n25766_), .ZN(new_n25847_));
  OAI21_X1   g22645(.A1(new_n25844_), .A2(new_n16574_), .B(new_n25847_), .ZN(new_n25848_));
  NOR2_X1    g22646(.A1(new_n25840_), .A2(new_n13994_), .ZN(new_n25849_));
  XNOR2_X1   g22647(.A1(new_n25849_), .A2(new_n19033_), .ZN(new_n25850_));
  AOI22_X1   g22648(.A1(new_n25850_), .A2(new_n25748_), .B1(new_n14206_), .B2(new_n25768_), .ZN(new_n25851_));
  NOR3_X1    g22649(.A1(new_n25851_), .A2(new_n14010_), .A3(new_n25765_), .ZN(new_n25852_));
  OAI22_X1   g22650(.A1(new_n25838_), .A2(new_n25848_), .B1(new_n12776_), .B2(new_n25852_), .ZN(new_n25853_));
  NAND2_X1   g22651(.A1(new_n25853_), .A2(pi0644), .ZN(new_n25854_));
  XOR2_X1    g22652(.A1(new_n25854_), .A2(new_n14205_), .Z(new_n25855_));
  NOR2_X1    g22653(.A1(new_n25855_), .A2(new_n25770_), .ZN(new_n25856_));
  NOR2_X1    g22654(.A1(new_n25840_), .A2(new_n18968_), .ZN(new_n25857_));
  NAND2_X1   g22655(.A1(new_n18967_), .A2(new_n25748_), .ZN(new_n25858_));
  XOR2_X1    g22656(.A1(new_n25857_), .A2(new_n25858_), .Z(new_n25859_));
  NAND2_X1   g22657(.A1(new_n25859_), .A2(pi0715), .ZN(new_n25860_));
  XOR2_X1    g22658(.A1(new_n25860_), .A2(new_n14205_), .Z(new_n25861_));
  OAI21_X1   g22659(.A1(new_n25861_), .A2(new_n25766_), .B(new_n14203_), .ZN(new_n25862_));
  NAND2_X1   g22660(.A1(new_n25859_), .A2(pi0644), .ZN(new_n25863_));
  XOR2_X1    g22661(.A1(new_n25863_), .A2(new_n14217_), .Z(new_n25864_));
  AOI21_X1   g22662(.A1(new_n25864_), .A2(new_n25748_), .B(pi1160), .ZN(new_n25865_));
  OAI21_X1   g22663(.A1(new_n25856_), .A2(new_n25862_), .B(new_n25865_), .ZN(new_n25866_));
  NAND2_X1   g22664(.A1(new_n25853_), .A2(pi0715), .ZN(new_n25867_));
  XOR2_X1    g22665(.A1(new_n25867_), .A2(new_n14205_), .Z(new_n25868_));
  NOR2_X1    g22666(.A1(new_n25868_), .A2(new_n25770_), .ZN(new_n25869_));
  AOI21_X1   g22667(.A1(new_n25866_), .A2(new_n25869_), .B(new_n14799_), .ZN(new_n25870_));
  XOR2_X1    g22668(.A1(new_n25870_), .A2(new_n14800_), .Z(new_n25871_));
  OAI21_X1   g22669(.A1(new_n7240_), .A2(pi0193), .B(new_n14799_), .ZN(new_n25872_));
  NOR2_X1    g22670(.A1(new_n25853_), .A2(new_n25872_), .ZN(new_n25873_));
  AOI21_X1   g22671(.A1(new_n25871_), .A2(new_n25873_), .B(po1038), .ZN(new_n25874_));
  NOR3_X1    g22672(.A1(new_n25745_), .A2(new_n25744_), .A3(new_n25874_), .ZN(new_n25875_));
  OAI21_X1   g22673(.A1(new_n25741_), .A2(pi0792), .B(new_n25875_), .ZN(new_n25876_));
  NOR2_X1    g22674(.A1(new_n25876_), .A2(new_n25640_), .ZN(po0350));
  XOR2_X1    g22675(.A1(new_n22960_), .A2(new_n12528_), .Z(new_n25878_));
  NAND2_X1   g22676(.A1(new_n25878_), .A2(new_n13624_), .ZN(new_n25879_));
  NAND2_X1   g22677(.A1(new_n19323_), .A2(pi0194), .ZN(new_n25880_));
  NAND2_X1   g22678(.A1(new_n19329_), .A2(new_n12522_), .ZN(new_n25881_));
  NAND2_X1   g22679(.A1(new_n25880_), .A2(new_n25881_), .ZN(new_n25882_));
  NAND2_X1   g22680(.A1(new_n25882_), .A2(pi0748), .ZN(new_n25883_));
  OAI21_X1   g22681(.A1(new_n25879_), .A2(pi0748), .B(new_n25883_), .ZN(new_n25884_));
  NOR2_X1    g22682(.A1(new_n3289_), .A2(pi0194), .ZN(new_n25885_));
  AOI21_X1   g22683(.A1(new_n25884_), .A2(new_n3289_), .B(new_n25885_), .ZN(new_n25886_));
  NOR2_X1    g22684(.A1(new_n18025_), .A2(new_n18000_), .ZN(new_n25887_));
  AOI21_X1   g22685(.A1(new_n15607_), .A2(new_n25887_), .B(pi0194), .ZN(new_n25888_));
  NOR2_X1    g22686(.A1(new_n12522_), .A2(new_n18000_), .ZN(new_n25889_));
  NOR2_X1    g22687(.A1(new_n19395_), .A2(new_n15630_), .ZN(new_n25890_));
  OAI21_X1   g22688(.A1(new_n15615_), .A2(new_n25889_), .B(new_n25890_), .ZN(new_n25891_));
  OAI21_X1   g22689(.A1(new_n25891_), .A2(new_n25888_), .B(new_n15595_), .ZN(new_n25892_));
  NAND2_X1   g22690(.A1(new_n25892_), .A2(pi0194), .ZN(new_n25893_));
  NAND2_X1   g22691(.A1(new_n25893_), .A2(new_n3289_), .ZN(new_n25894_));
  NAND3_X1   g22692(.A1(new_n25882_), .A2(pi0730), .A3(pi0748), .ZN(new_n25895_));
  NAND4_X1   g22693(.A1(new_n25880_), .A2(new_n25881_), .A3(new_n18025_), .A4(pi0748), .ZN(new_n25896_));
  NAND2_X1   g22694(.A1(new_n25895_), .A2(new_n25896_), .ZN(new_n25897_));
  NOR2_X1    g22695(.A1(new_n3290_), .A2(new_n12522_), .ZN(new_n25898_));
  NAND4_X1   g22696(.A1(new_n25897_), .A2(new_n13624_), .A3(new_n25878_), .A4(new_n25898_), .ZN(new_n25899_));
  INV_X1     g22697(.I(new_n25899_), .ZN(new_n25900_));
  NAND2_X1   g22698(.A1(new_n25894_), .A2(new_n25900_), .ZN(new_n25901_));
  AOI21_X1   g22699(.A1(new_n25892_), .A2(pi0194), .B(new_n3290_), .ZN(new_n25902_));
  NAND2_X1   g22700(.A1(new_n25902_), .A2(new_n25899_), .ZN(new_n25903_));
  NAND3_X1   g22701(.A1(new_n25901_), .A2(new_n25903_), .A3(pi1153), .ZN(new_n25904_));
  NAND2_X1   g22702(.A1(new_n25904_), .A2(new_n13615_), .ZN(new_n25905_));
  XOR2_X1    g22703(.A1(new_n25902_), .A2(new_n25899_), .Z(new_n25906_));
  NAND3_X1   g22704(.A1(new_n25906_), .A2(pi1153), .A3(new_n13620_), .ZN(new_n25907_));
  AOI21_X1   g22705(.A1(new_n25905_), .A2(new_n25907_), .B(new_n25886_), .ZN(new_n25908_));
  NOR2_X1    g22706(.A1(new_n14428_), .A2(pi0194), .ZN(new_n25909_));
  NOR2_X1    g22707(.A1(new_n19287_), .A2(new_n3290_), .ZN(new_n25910_));
  OAI21_X1   g22708(.A1(new_n25879_), .A2(pi0730), .B(new_n25910_), .ZN(new_n25911_));
  NAND2_X1   g22709(.A1(pi0194), .A2(pi0730), .ZN(new_n25912_));
  NAND2_X1   g22710(.A1(new_n25911_), .A2(new_n25912_), .ZN(new_n25913_));
  INV_X1     g22711(.I(new_n25913_), .ZN(new_n25914_));
  AOI21_X1   g22712(.A1(new_n25914_), .A2(pi0625), .B(new_n13620_), .ZN(new_n25915_));
  NOR3_X1    g22713(.A1(new_n25913_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n25916_));
  OAI21_X1   g22714(.A1(new_n25915_), .A2(new_n25916_), .B(new_n25909_), .ZN(new_n25917_));
  NAND2_X1   g22715(.A1(new_n25917_), .A2(pi0608), .ZN(new_n25918_));
  OAI21_X1   g22716(.A1(new_n25908_), .A2(new_n25918_), .B(pi0778), .ZN(new_n25919_));
  INV_X1     g22717(.I(new_n25886_), .ZN(new_n25920_));
  NAND3_X1   g22718(.A1(new_n25901_), .A2(new_n25903_), .A3(pi0625), .ZN(new_n25921_));
  NAND2_X1   g22719(.A1(new_n25921_), .A2(new_n13615_), .ZN(new_n25922_));
  NAND3_X1   g22720(.A1(new_n25906_), .A2(pi0625), .A3(new_n13620_), .ZN(new_n25923_));
  NAND2_X1   g22721(.A1(new_n25922_), .A2(new_n25923_), .ZN(new_n25924_));
  AOI21_X1   g22722(.A1(new_n25914_), .A2(pi1153), .B(new_n13620_), .ZN(new_n25925_));
  NOR3_X1    g22723(.A1(new_n25913_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n25926_));
  OAI21_X1   g22724(.A1(new_n25925_), .A2(new_n25926_), .B(new_n25909_), .ZN(new_n25927_));
  NOR2_X1    g22725(.A1(new_n25906_), .A2(new_n13750_), .ZN(new_n25928_));
  NAND2_X1   g22726(.A1(new_n25928_), .A2(new_n25927_), .ZN(new_n25929_));
  AOI21_X1   g22727(.A1(new_n25924_), .A2(new_n25920_), .B(new_n25929_), .ZN(new_n25930_));
  NAND2_X1   g22728(.A1(new_n25919_), .A2(new_n25930_), .ZN(new_n25931_));
  AOI21_X1   g22729(.A1(new_n25906_), .A2(pi1153), .B(new_n13620_), .ZN(new_n25932_));
  NOR2_X1    g22730(.A1(new_n25904_), .A2(new_n13615_), .ZN(new_n25933_));
  OAI21_X1   g22731(.A1(new_n25933_), .A2(new_n25932_), .B(new_n25920_), .ZN(new_n25934_));
  INV_X1     g22732(.I(new_n25918_), .ZN(new_n25935_));
  AOI21_X1   g22733(.A1(new_n25934_), .A2(new_n25935_), .B(new_n13748_), .ZN(new_n25936_));
  AOI21_X1   g22734(.A1(new_n25906_), .A2(pi0625), .B(new_n13620_), .ZN(new_n25937_));
  NOR2_X1    g22735(.A1(new_n25921_), .A2(new_n13615_), .ZN(new_n25938_));
  OAI21_X1   g22736(.A1(new_n25938_), .A2(new_n25937_), .B(new_n25920_), .ZN(new_n25939_));
  NAND3_X1   g22737(.A1(new_n25939_), .A2(new_n25927_), .A3(new_n25928_), .ZN(new_n25940_));
  NAND2_X1   g22738(.A1(new_n25936_), .A2(new_n25940_), .ZN(new_n25941_));
  NAND2_X1   g22739(.A1(new_n25941_), .A2(new_n25931_), .ZN(new_n25942_));
  NAND2_X1   g22740(.A1(new_n25917_), .A2(pi0778), .ZN(new_n25943_));
  NOR3_X1    g22741(.A1(new_n25927_), .A2(new_n13748_), .A3(new_n25914_), .ZN(new_n25944_));
  NAND2_X1   g22742(.A1(new_n25944_), .A2(new_n25943_), .ZN(new_n25945_));
  NOR2_X1    g22743(.A1(new_n25944_), .A2(new_n25943_), .ZN(new_n25946_));
  INV_X1     g22744(.I(new_n25946_), .ZN(new_n25947_));
  NAND2_X1   g22745(.A1(new_n25947_), .A2(new_n25945_), .ZN(new_n25948_));
  NAND2_X1   g22746(.A1(new_n25886_), .A2(new_n13776_), .ZN(new_n25949_));
  NOR2_X1    g22747(.A1(new_n25909_), .A2(new_n15147_), .ZN(new_n25951_));
  OAI21_X1   g22748(.A1(new_n25948_), .A2(new_n13785_), .B(new_n13766_), .ZN(new_n25952_));
  AOI21_X1   g22749(.A1(new_n25947_), .A2(new_n25945_), .B(new_n13766_), .ZN(new_n25953_));
  INV_X1     g22750(.I(new_n25909_), .ZN(new_n25954_));
  AOI21_X1   g22751(.A1(new_n25954_), .A2(new_n14467_), .B(pi0609), .ZN(new_n25955_));
  NOR2_X1    g22752(.A1(new_n25949_), .A2(new_n25955_), .ZN(new_n25956_));
  NOR2_X1    g22753(.A1(new_n25956_), .A2(new_n14465_), .ZN(new_n25957_));
  INV_X1     g22754(.I(new_n25957_), .ZN(new_n25958_));
  OAI21_X1   g22755(.A1(new_n25953_), .A2(new_n25958_), .B(new_n13766_), .ZN(new_n25959_));
  NAND4_X1   g22756(.A1(new_n25942_), .A2(pi0785), .A3(new_n25959_), .A4(new_n25952_), .ZN(new_n25960_));
  NAND2_X1   g22757(.A1(new_n25942_), .A2(new_n25952_), .ZN(new_n25961_));
  NAND3_X1   g22758(.A1(new_n25942_), .A2(pi0785), .A3(new_n25959_), .ZN(new_n25962_));
  NAND3_X1   g22759(.A1(new_n25962_), .A2(new_n25961_), .A3(pi0785), .ZN(new_n25963_));
  NAND2_X1   g22760(.A1(new_n25963_), .A2(new_n25960_), .ZN(new_n25964_));
  AOI21_X1   g22761(.A1(new_n25886_), .A2(new_n13776_), .B(new_n25951_), .ZN(new_n25965_));
  OAI21_X1   g22762(.A1(new_n25965_), .A2(new_n13766_), .B(pi0785), .ZN(new_n25966_));
  NAND2_X1   g22763(.A1(new_n25909_), .A2(new_n13775_), .ZN(new_n25967_));
  OAI21_X1   g22764(.A1(new_n25886_), .A2(new_n13775_), .B(new_n25967_), .ZN(new_n25968_));
  NAND3_X1   g22765(.A1(new_n25956_), .A2(pi0785), .A3(new_n25968_), .ZN(new_n25969_));
  XOR2_X1    g22766(.A1(new_n25969_), .A2(new_n25966_), .Z(new_n25970_));
  NAND3_X1   g22767(.A1(new_n25970_), .A2(pi0618), .A3(pi1154), .ZN(new_n25971_));
  NOR3_X1    g22768(.A1(new_n25970_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n25972_));
  INV_X1     g22769(.I(new_n25972_), .ZN(new_n25973_));
  AOI21_X1   g22770(.A1(new_n25973_), .A2(new_n25971_), .B(new_n25954_), .ZN(new_n25974_));
  AOI21_X1   g22771(.A1(new_n25947_), .A2(new_n25945_), .B(new_n13803_), .ZN(new_n25975_));
  NOR2_X1    g22772(.A1(new_n25954_), .A2(new_n13805_), .ZN(new_n25976_));
  NOR2_X1    g22773(.A1(new_n25975_), .A2(new_n25976_), .ZN(new_n25977_));
  OAI21_X1   g22774(.A1(new_n25977_), .A2(pi0618), .B(new_n13824_), .ZN(new_n25978_));
  OAI21_X1   g22775(.A1(new_n25978_), .A2(new_n25974_), .B(new_n13816_), .ZN(new_n25979_));
  NAND3_X1   g22776(.A1(new_n25970_), .A2(pi0618), .A3(pi1154), .ZN(new_n25980_));
  XNOR2_X1   g22777(.A1(new_n25969_), .A2(new_n25966_), .ZN(new_n25981_));
  NAND3_X1   g22778(.A1(new_n25981_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n25982_));
  AOI21_X1   g22779(.A1(new_n25982_), .A2(new_n25980_), .B(new_n25954_), .ZN(new_n25983_));
  INV_X1     g22780(.I(new_n25945_), .ZN(new_n25984_));
  OAI21_X1   g22781(.A1(new_n25984_), .A2(new_n25946_), .B(new_n13805_), .ZN(new_n25985_));
  INV_X1     g22782(.I(new_n25976_), .ZN(new_n25986_));
  AOI21_X1   g22783(.A1(new_n25985_), .A2(new_n25986_), .B(new_n13816_), .ZN(new_n25987_));
  NOR3_X1    g22784(.A1(new_n25987_), .A2(new_n25983_), .A3(new_n13837_), .ZN(new_n25988_));
  NOR2_X1    g22785(.A1(new_n25988_), .A2(pi0618), .ZN(new_n25989_));
  INV_X1     g22786(.I(new_n25989_), .ZN(new_n25990_));
  NAND4_X1   g22787(.A1(new_n25964_), .A2(pi0781), .A3(new_n25979_), .A4(new_n25990_), .ZN(new_n25991_));
  INV_X1     g22788(.I(new_n25960_), .ZN(new_n25992_));
  NOR2_X1    g22789(.A1(new_n25936_), .A2(new_n25940_), .ZN(new_n25993_));
  NOR2_X1    g22790(.A1(new_n25919_), .A2(new_n25930_), .ZN(new_n25994_));
  NOR2_X1    g22791(.A1(new_n25993_), .A2(new_n25994_), .ZN(new_n25995_));
  NOR2_X1    g22792(.A1(new_n25984_), .A2(new_n25946_), .ZN(new_n25996_));
  AOI21_X1   g22793(.A1(new_n25996_), .A2(new_n13784_), .B(pi0609), .ZN(new_n25997_));
  OAI21_X1   g22794(.A1(new_n25995_), .A2(new_n25997_), .B(pi0785), .ZN(new_n25998_));
  OAI21_X1   g22795(.A1(new_n25984_), .A2(new_n25946_), .B(pi0609), .ZN(new_n25999_));
  AOI21_X1   g22796(.A1(new_n25999_), .A2(new_n25957_), .B(pi0609), .ZN(new_n26000_));
  NOR3_X1    g22797(.A1(new_n25995_), .A2(new_n13801_), .A3(new_n26000_), .ZN(new_n26001_));
  NOR2_X1    g22798(.A1(new_n26001_), .A2(new_n25998_), .ZN(new_n26002_));
  OAI21_X1   g22799(.A1(new_n26002_), .A2(new_n25992_), .B(new_n25979_), .ZN(new_n26003_));
  AOI21_X1   g22800(.A1(new_n25981_), .A2(pi1154), .B(new_n13819_), .ZN(new_n26004_));
  NOR3_X1    g22801(.A1(new_n25970_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n26005_));
  OAI21_X1   g22802(.A1(new_n26004_), .A2(new_n26005_), .B(new_n25909_), .ZN(new_n26006_));
  OAI21_X1   g22803(.A1(new_n25975_), .A2(new_n25976_), .B(pi0618), .ZN(new_n26007_));
  NAND3_X1   g22804(.A1(new_n26007_), .A2(new_n26006_), .A3(new_n13836_), .ZN(new_n26008_));
  AOI21_X1   g22805(.A1(new_n26008_), .A2(new_n13816_), .B(new_n13855_), .ZN(new_n26009_));
  OAI21_X1   g22806(.A1(new_n26002_), .A2(new_n25992_), .B(new_n26009_), .ZN(new_n26010_));
  NAND3_X1   g22807(.A1(new_n26010_), .A2(new_n26003_), .A3(pi0781), .ZN(new_n26011_));
  NAND2_X1   g22808(.A1(new_n26011_), .A2(new_n25991_), .ZN(new_n26012_));
  NAND4_X1   g22809(.A1(new_n25974_), .A2(new_n25983_), .A3(pi0781), .A4(new_n25970_), .ZN(new_n26013_));
  INV_X1     g22810(.I(new_n25971_), .ZN(new_n26014_));
  OAI21_X1   g22811(.A1(new_n26014_), .A2(new_n25972_), .B(new_n25909_), .ZN(new_n26015_));
  NAND3_X1   g22812(.A1(new_n25983_), .A2(pi0781), .A3(new_n25970_), .ZN(new_n26016_));
  NAND3_X1   g22813(.A1(new_n26016_), .A2(pi0781), .A3(new_n26015_), .ZN(new_n26017_));
  NAND2_X1   g22814(.A1(new_n26017_), .A2(new_n26013_), .ZN(new_n26018_));
  NAND3_X1   g22815(.A1(new_n26018_), .A2(pi0619), .A3(pi1159), .ZN(new_n26019_));
  NAND4_X1   g22816(.A1(new_n26017_), .A2(pi0619), .A3(new_n26013_), .A4(new_n13868_), .ZN(new_n26020_));
  AOI21_X1   g22817(.A1(new_n26019_), .A2(new_n26020_), .B(new_n25954_), .ZN(new_n26021_));
  NAND2_X1   g22818(.A1(new_n25985_), .A2(new_n25986_), .ZN(new_n26022_));
  NOR2_X1    g22819(.A1(new_n25909_), .A2(new_n13880_), .ZN(new_n26023_));
  INV_X1     g22820(.I(new_n26023_), .ZN(new_n26024_));
  OAI21_X1   g22821(.A1(new_n26022_), .A2(new_n13879_), .B(new_n26024_), .ZN(new_n26025_));
  OAI21_X1   g22822(.A1(new_n26025_), .A2(pi0619), .B(new_n13885_), .ZN(new_n26026_));
  OAI21_X1   g22823(.A1(new_n26021_), .A2(new_n26026_), .B(new_n13860_), .ZN(new_n26027_));
  NAND3_X1   g22824(.A1(new_n26018_), .A2(pi0619), .A3(pi1159), .ZN(new_n26028_));
  NAND4_X1   g22825(.A1(new_n26017_), .A2(new_n13860_), .A3(new_n26013_), .A4(pi1159), .ZN(new_n26029_));
  AOI21_X1   g22826(.A1(new_n26028_), .A2(new_n26029_), .B(new_n25954_), .ZN(new_n26030_));
  OAI21_X1   g22827(.A1(new_n26025_), .A2(new_n13860_), .B(new_n13892_), .ZN(new_n26031_));
  OAI21_X1   g22828(.A1(new_n26030_), .A2(new_n26031_), .B(new_n13860_), .ZN(new_n26032_));
  NAND4_X1   g22829(.A1(new_n26027_), .A2(new_n26032_), .A3(pi0789), .A4(new_n26012_), .ZN(new_n26033_));
  INV_X1     g22830(.I(new_n26033_), .ZN(new_n26034_));
  AOI21_X1   g22831(.A1(pi0781), .A2(new_n26003_), .B(new_n26010_), .ZN(new_n26035_));
  AOI21_X1   g22832(.A1(new_n26022_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n26036_));
  AOI21_X1   g22833(.A1(new_n26036_), .A2(new_n26015_), .B(pi0618), .ZN(new_n26037_));
  AOI21_X1   g22834(.A1(new_n25963_), .A2(new_n25960_), .B(new_n26037_), .ZN(new_n26038_));
  OAI21_X1   g22835(.A1(new_n25988_), .A2(pi0618), .B(pi0781), .ZN(new_n26039_));
  AOI21_X1   g22836(.A1(new_n25963_), .A2(new_n25960_), .B(new_n26039_), .ZN(new_n26040_));
  NOR3_X1    g22837(.A1(new_n26040_), .A2(new_n26038_), .A3(new_n13855_), .ZN(new_n26041_));
  NOR2_X1    g22838(.A1(new_n26035_), .A2(new_n26041_), .ZN(new_n26042_));
  NOR4_X1    g22839(.A1(new_n26015_), .A2(new_n26006_), .A3(new_n13855_), .A4(new_n25981_), .ZN(new_n26043_));
  NOR3_X1    g22840(.A1(new_n26006_), .A2(new_n13855_), .A3(new_n25981_), .ZN(new_n26044_));
  NOR3_X1    g22841(.A1(new_n26044_), .A2(new_n13855_), .A3(new_n25974_), .ZN(new_n26045_));
  NOR2_X1    g22842(.A1(new_n26045_), .A2(new_n26043_), .ZN(new_n26046_));
  AOI21_X1   g22843(.A1(new_n26046_), .A2(pi0619), .B(new_n13904_), .ZN(new_n26047_));
  INV_X1     g22844(.I(new_n26020_), .ZN(new_n26048_));
  OAI21_X1   g22845(.A1(new_n26047_), .A2(new_n26048_), .B(new_n25909_), .ZN(new_n26049_));
  INV_X1     g22846(.I(new_n26026_), .ZN(new_n26050_));
  AOI21_X1   g22847(.A1(new_n26049_), .A2(new_n26050_), .B(pi0619), .ZN(new_n26051_));
  OAI21_X1   g22848(.A1(new_n26051_), .A2(new_n26042_), .B(pi0789), .ZN(new_n26052_));
  AOI21_X1   g22849(.A1(new_n26046_), .A2(pi1159), .B(new_n13904_), .ZN(new_n26053_));
  INV_X1     g22850(.I(new_n26029_), .ZN(new_n26054_));
  OAI21_X1   g22851(.A1(new_n26053_), .A2(new_n26054_), .B(new_n25909_), .ZN(new_n26055_));
  INV_X1     g22852(.I(new_n26031_), .ZN(new_n26056_));
  AOI21_X1   g22853(.A1(new_n26055_), .A2(new_n26056_), .B(pi0619), .ZN(new_n26057_));
  OAI21_X1   g22854(.A1(new_n26035_), .A2(new_n26041_), .B(pi0789), .ZN(new_n26058_));
  NOR2_X1    g22855(.A1(new_n26057_), .A2(new_n26058_), .ZN(new_n26059_));
  NOR2_X1    g22856(.A1(new_n26052_), .A2(new_n26059_), .ZN(new_n26060_));
  NOR2_X1    g22857(.A1(new_n26060_), .A2(new_n26034_), .ZN(new_n26061_));
  NAND4_X1   g22858(.A1(new_n26021_), .A2(new_n26030_), .A3(pi0789), .A4(new_n26018_), .ZN(new_n26062_));
  NOR2_X1    g22859(.A1(new_n26046_), .A2(new_n13896_), .ZN(new_n26063_));
  NAND2_X1   g22860(.A1(new_n26030_), .A2(new_n26063_), .ZN(new_n26064_));
  NAND3_X1   g22861(.A1(new_n26064_), .A2(pi0789), .A3(new_n26049_), .ZN(new_n26065_));
  AOI21_X1   g22862(.A1(new_n25977_), .A2(new_n13880_), .B(new_n26023_), .ZN(new_n26066_));
  NOR2_X1    g22863(.A1(new_n25954_), .A2(new_n13919_), .ZN(new_n26067_));
  AOI21_X1   g22864(.A1(new_n26066_), .A2(new_n13919_), .B(new_n26067_), .ZN(new_n26068_));
  NOR2_X1    g22865(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n26069_));
  INV_X1     g22866(.I(new_n26069_), .ZN(new_n26070_));
  AOI21_X1   g22867(.A1(new_n26065_), .A2(new_n26062_), .B(new_n26070_), .ZN(new_n26071_));
  INV_X1     g22868(.I(new_n26067_), .ZN(new_n26072_));
  OAI21_X1   g22869(.A1(new_n26025_), .A2(new_n13918_), .B(new_n26072_), .ZN(new_n26073_));
  NOR3_X1    g22870(.A1(new_n26061_), .A2(new_n13901_), .A3(new_n13937_), .ZN(new_n26077_));
  AOI21_X1   g22871(.A1(new_n26027_), .A2(new_n26012_), .B(new_n13896_), .ZN(new_n26078_));
  AOI21_X1   g22872(.A1(new_n26011_), .A2(new_n25991_), .B(new_n13896_), .ZN(new_n26079_));
  NAND2_X1   g22873(.A1(new_n26032_), .A2(new_n26079_), .ZN(new_n26080_));
  NAND2_X1   g22874(.A1(new_n26078_), .A2(new_n26080_), .ZN(new_n26081_));
  INV_X1     g22875(.I(new_n26062_), .ZN(new_n26082_));
  NAND2_X1   g22876(.A1(new_n26049_), .A2(pi0789), .ZN(new_n26083_));
  NOR3_X1    g22877(.A1(new_n26055_), .A2(new_n13896_), .A3(new_n26046_), .ZN(new_n26084_));
  NOR2_X1    g22878(.A1(new_n26084_), .A2(new_n26083_), .ZN(new_n26085_));
  OAI21_X1   g22879(.A1(new_n26085_), .A2(new_n26082_), .B(new_n26069_), .ZN(new_n26086_));
  AOI22_X1   g22880(.A1(new_n26086_), .A2(new_n13901_), .B1(new_n26081_), .B2(new_n26033_), .ZN(new_n26087_));
  AOI21_X1   g22881(.A1(new_n26081_), .A2(new_n26033_), .B(new_n15258_), .ZN(new_n26088_));
  NOR3_X1    g22882(.A1(new_n26087_), .A2(new_n13937_), .A3(new_n26088_), .ZN(new_n26089_));
  NOR2_X1    g22883(.A1(new_n26089_), .A2(new_n26077_), .ZN(new_n26090_));
  NOR2_X1    g22884(.A1(new_n25909_), .A2(new_n16372_), .ZN(new_n26091_));
  NOR3_X1    g22885(.A1(new_n26085_), .A2(new_n26082_), .A3(new_n14142_), .ZN(new_n26092_));
  NOR2_X1    g22886(.A1(new_n26092_), .A2(new_n26091_), .ZN(new_n26093_));
  NOR2_X1    g22887(.A1(new_n25909_), .A2(new_n13966_), .ZN(new_n26094_));
  INV_X1     g22888(.I(new_n26094_), .ZN(new_n26095_));
  OAI21_X1   g22889(.A1(new_n26073_), .A2(new_n13965_), .B(new_n26095_), .ZN(new_n26096_));
  NAND3_X1   g22890(.A1(new_n26096_), .A2(pi0628), .A3(pi1156), .ZN(new_n26097_));
  AOI21_X1   g22891(.A1(new_n26068_), .A2(new_n13966_), .B(new_n26094_), .ZN(new_n26098_));
  NAND3_X1   g22892(.A1(new_n26098_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n26099_));
  AOI21_X1   g22893(.A1(new_n26099_), .A2(new_n26097_), .B(new_n25954_), .ZN(new_n26100_));
  NOR2_X1    g22894(.A1(new_n26100_), .A2(new_n15270_), .ZN(new_n26101_));
  INV_X1     g22895(.I(new_n26101_), .ZN(new_n26102_));
  INV_X1     g22896(.I(new_n26091_), .ZN(new_n26104_));
  NAND3_X1   g22897(.A1(new_n26065_), .A2(new_n16372_), .A3(new_n26062_), .ZN(new_n26105_));
  NAND2_X1   g22898(.A1(new_n26105_), .A2(new_n26104_), .ZN(new_n26106_));
  NAND3_X1   g22899(.A1(new_n26096_), .A2(pi0628), .A3(pi1156), .ZN(new_n26108_));
  NAND3_X1   g22900(.A1(new_n26098_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n26109_));
  AOI21_X1   g22901(.A1(new_n26109_), .A2(new_n26108_), .B(new_n25954_), .ZN(new_n26110_));
  NOR3_X1    g22902(.A1(new_n26090_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n26112_));
  NAND2_X1   g22903(.A1(new_n26081_), .A2(new_n26033_), .ZN(new_n26113_));
  NAND3_X1   g22904(.A1(new_n26113_), .A2(pi0626), .A3(pi0788), .ZN(new_n26114_));
  OAI22_X1   g22905(.A1(new_n26060_), .A2(new_n26034_), .B1(new_n26071_), .B2(pi0626), .ZN(new_n26115_));
  OAI21_X1   g22906(.A1(new_n26060_), .A2(new_n26034_), .B(new_n14577_), .ZN(new_n26116_));
  NAND3_X1   g22907(.A1(new_n26115_), .A2(new_n26116_), .A3(pi0788), .ZN(new_n26117_));
  AOI21_X1   g22908(.A1(new_n26106_), .A2(new_n26101_), .B(pi0628), .ZN(new_n26118_));
  AOI21_X1   g22909(.A1(new_n26117_), .A2(new_n26114_), .B(new_n26118_), .ZN(new_n26119_));
  AOI21_X1   g22910(.A1(new_n26117_), .A2(new_n26114_), .B(new_n15296_), .ZN(new_n26120_));
  NOR3_X1    g22911(.A1(new_n26119_), .A2(new_n26120_), .A3(new_n12777_), .ZN(new_n26121_));
  NOR2_X1    g22912(.A1(new_n26121_), .A2(new_n26112_), .ZN(new_n26122_));
  NOR2_X1    g22913(.A1(new_n26100_), .A2(new_n12777_), .ZN(new_n26123_));
  NAND3_X1   g22914(.A1(new_n26110_), .A2(pi0792), .A3(new_n26096_), .ZN(new_n26124_));
  XOR2_X1    g22915(.A1(new_n26124_), .A2(new_n26123_), .Z(new_n26125_));
  AOI21_X1   g22916(.A1(new_n26125_), .A2(pi0647), .B(new_n14008_), .ZN(new_n26126_));
  NAND4_X1   g22917(.A1(new_n26100_), .A2(new_n26110_), .A3(pi0792), .A4(new_n26096_), .ZN(new_n26127_));
  NAND2_X1   g22918(.A1(new_n26124_), .A2(new_n26123_), .ZN(new_n26128_));
  NAND2_X1   g22919(.A1(new_n26128_), .A2(new_n26127_), .ZN(new_n26129_));
  NOR3_X1    g22920(.A1(new_n26129_), .A2(new_n14005_), .A3(pi1157), .ZN(new_n26130_));
  OAI21_X1   g22921(.A1(new_n26126_), .A2(new_n26130_), .B(new_n25909_), .ZN(new_n26131_));
  AOI21_X1   g22922(.A1(new_n26105_), .A2(new_n26104_), .B(new_n13993_), .ZN(new_n26132_));
  NOR2_X1    g22923(.A1(new_n25909_), .A2(new_n13994_), .ZN(new_n26133_));
  NOR2_X1    g22924(.A1(new_n26132_), .A2(new_n26133_), .ZN(new_n26134_));
  AOI21_X1   g22925(.A1(new_n26134_), .A2(new_n14005_), .B(new_n14012_), .ZN(new_n26135_));
  AOI21_X1   g22926(.A1(new_n26135_), .A2(new_n26131_), .B(pi0647), .ZN(new_n26136_));
  NAND3_X1   g22927(.A1(new_n26129_), .A2(pi0647), .A3(pi1157), .ZN(new_n26137_));
  NAND4_X1   g22928(.A1(new_n26128_), .A2(new_n26127_), .A3(new_n14005_), .A4(pi1157), .ZN(new_n26138_));
  AOI21_X1   g22929(.A1(new_n26137_), .A2(new_n26138_), .B(new_n25954_), .ZN(new_n26139_));
  NOR3_X1    g22930(.A1(new_n26132_), .A2(new_n14005_), .A3(new_n26133_), .ZN(new_n26140_));
  NOR3_X1    g22931(.A1(new_n26139_), .A2(new_n26140_), .A3(new_n16329_), .ZN(new_n26141_));
  NOR2_X1    g22932(.A1(new_n26141_), .A2(pi0647), .ZN(new_n26142_));
  NOR4_X1    g22933(.A1(new_n26122_), .A2(new_n12776_), .A3(new_n26136_), .A4(new_n26142_), .ZN(new_n26143_));
  NAND2_X1   g22934(.A1(new_n26117_), .A2(new_n26114_), .ZN(new_n26144_));
  NAND3_X1   g22935(.A1(new_n26144_), .A2(pi0628), .A3(pi0792), .ZN(new_n26145_));
  OAI21_X1   g22936(.A1(new_n26093_), .A2(new_n26102_), .B(new_n13942_), .ZN(new_n26146_));
  OAI21_X1   g22937(.A1(new_n26089_), .A2(new_n26077_), .B(new_n26146_), .ZN(new_n26147_));
  OAI21_X1   g22938(.A1(new_n26089_), .A2(new_n26077_), .B(new_n14606_), .ZN(new_n26148_));
  NAND3_X1   g22939(.A1(new_n26147_), .A2(new_n26148_), .A3(pi0792), .ZN(new_n26149_));
  AOI21_X1   g22940(.A1(new_n26149_), .A2(new_n26145_), .B(new_n26136_), .ZN(new_n26150_));
  OAI21_X1   g22941(.A1(new_n26141_), .A2(pi0647), .B(pi0787), .ZN(new_n26151_));
  AOI21_X1   g22942(.A1(new_n26149_), .A2(new_n26145_), .B(new_n26151_), .ZN(new_n26152_));
  NOR3_X1    g22943(.A1(new_n26150_), .A2(new_n26152_), .A3(new_n12776_), .ZN(new_n26153_));
  OAI21_X1   g22944(.A1(new_n26153_), .A2(new_n26143_), .B(new_n12775_), .ZN(new_n26154_));
  NOR2_X1    g22945(.A1(new_n9992_), .A2(pi0194), .ZN(new_n26155_));
  NOR2_X1    g22946(.A1(new_n14652_), .A2(new_n18025_), .ZN(new_n26156_));
  AOI21_X1   g22947(.A1(new_n13218_), .A2(pi0730), .B(new_n26155_), .ZN(new_n26157_));
  INV_X1     g22948(.I(new_n26157_), .ZN(new_n26158_));
  NAND3_X1   g22949(.A1(new_n26158_), .A2(new_n26156_), .A3(new_n26155_), .ZN(new_n26159_));
  NOR3_X1    g22950(.A1(new_n26156_), .A2(new_n13614_), .A3(new_n26157_), .ZN(new_n26160_));
  XNOR2_X1   g22951(.A1(new_n26159_), .A2(new_n26160_), .ZN(new_n26161_));
  NAND2_X1   g22952(.A1(new_n26161_), .A2(pi0778), .ZN(new_n26162_));
  NAND2_X1   g22953(.A1(new_n26158_), .A2(new_n13748_), .ZN(new_n26163_));
  NAND2_X1   g22954(.A1(new_n26162_), .A2(new_n26163_), .ZN(new_n26164_));
  INV_X1     g22955(.I(new_n26164_), .ZN(new_n26165_));
  NOR2_X1    g22956(.A1(new_n26165_), .A2(new_n14048_), .ZN(new_n26166_));
  INV_X1     g22957(.I(new_n26166_), .ZN(new_n26167_));
  NOR2_X1    g22958(.A1(new_n26167_), .A2(new_n14051_), .ZN(new_n26168_));
  INV_X1     g22959(.I(new_n26168_), .ZN(new_n26169_));
  NOR2_X1    g22960(.A1(new_n26169_), .A2(new_n14163_), .ZN(new_n26170_));
  AOI21_X1   g22961(.A1(new_n13104_), .A2(pi0748), .B(new_n26155_), .ZN(new_n26171_));
  NOR2_X1    g22962(.A1(new_n14096_), .A2(new_n26171_), .ZN(new_n26172_));
  AOI21_X1   g22963(.A1(new_n26172_), .A2(new_n14094_), .B(pi1155), .ZN(new_n26173_));
  NOR2_X1    g22964(.A1(new_n26173_), .A2(new_n13801_), .ZN(new_n26174_));
  AOI21_X1   g22965(.A1(new_n26171_), .A2(pi1155), .B(new_n9992_), .ZN(new_n26175_));
  NOR2_X1    g22966(.A1(new_n26175_), .A2(new_n14102_), .ZN(new_n26176_));
  NAND3_X1   g22967(.A1(new_n26176_), .A2(new_n26172_), .A3(pi0785), .ZN(new_n26177_));
  XOR2_X1    g22968(.A1(new_n26174_), .A2(new_n26177_), .Z(new_n26178_));
  NOR2_X1    g22969(.A1(new_n26178_), .A2(new_n13817_), .ZN(new_n26179_));
  OAI21_X1   g22970(.A1(new_n26179_), .A2(pi0618), .B(new_n9992_), .ZN(new_n26180_));
  NAND2_X1   g22971(.A1(new_n26180_), .A2(pi0781), .ZN(new_n26181_));
  OAI21_X1   g22972(.A1(new_n26179_), .A2(new_n9992_), .B(pi0618), .ZN(new_n26182_));
  NOR3_X1    g22973(.A1(new_n26182_), .A2(new_n13855_), .A3(new_n26178_), .ZN(new_n26183_));
  XOR2_X1    g22974(.A1(new_n26183_), .A2(new_n26181_), .Z(new_n26184_));
  NAND2_X1   g22975(.A1(new_n26184_), .A2(pi0619), .ZN(new_n26185_));
  XOR2_X1    g22976(.A1(new_n26185_), .A2(new_n13904_), .Z(new_n26186_));
  NAND2_X1   g22977(.A1(new_n26186_), .A2(new_n26155_), .ZN(new_n26187_));
  NAND2_X1   g22978(.A1(new_n26187_), .A2(pi0789), .ZN(new_n26188_));
  NAND2_X1   g22979(.A1(new_n26184_), .A2(pi1159), .ZN(new_n26189_));
  XOR2_X1    g22980(.A1(new_n26189_), .A2(new_n13904_), .Z(new_n26190_));
  NAND2_X1   g22981(.A1(new_n26190_), .A2(new_n26155_), .ZN(new_n26191_));
  NOR3_X1    g22982(.A1(new_n26191_), .A2(new_n13896_), .A3(new_n26184_), .ZN(new_n26192_));
  XOR2_X1    g22983(.A1(new_n26192_), .A2(new_n26188_), .Z(new_n26193_));
  NAND2_X1   g22984(.A1(new_n26193_), .A2(new_n13962_), .ZN(new_n26194_));
  XOR2_X1    g22985(.A1(new_n26194_), .A2(new_n18976_), .Z(new_n26195_));
  AOI22_X1   g22986(.A1(new_n26195_), .A2(new_n26155_), .B1(new_n16639_), .B2(new_n26170_), .ZN(new_n26196_));
  NOR2_X1    g22987(.A1(new_n26157_), .A2(new_n13203_), .ZN(new_n26197_));
  INV_X1     g22988(.I(new_n26197_), .ZN(new_n26198_));
  NOR2_X1    g22989(.A1(new_n26198_), .A2(new_n13613_), .ZN(new_n26199_));
  NOR2_X1    g22990(.A1(new_n26155_), .A2(pi1153), .ZN(new_n26200_));
  INV_X1     g22991(.I(new_n26200_), .ZN(new_n26201_));
  OAI21_X1   g22992(.A1(new_n26156_), .A2(new_n26201_), .B(pi0608), .ZN(new_n26202_));
  NOR2_X1    g22993(.A1(new_n26171_), .A2(pi1153), .ZN(new_n26203_));
  NAND2_X1   g22994(.A1(new_n26202_), .A2(new_n26203_), .ZN(new_n26204_));
  AOI21_X1   g22995(.A1(new_n26204_), .A2(new_n26199_), .B(new_n13748_), .ZN(new_n26205_));
  NOR2_X1    g22996(.A1(new_n26157_), .A2(new_n14082_), .ZN(new_n26206_));
  NAND2_X1   g22997(.A1(new_n26156_), .A2(new_n26200_), .ZN(new_n26207_));
  OAI22_X1   g22998(.A1(new_n26198_), .A2(new_n13613_), .B1(new_n26207_), .B2(new_n26206_), .ZN(new_n26208_));
  NAND4_X1   g22999(.A1(new_n26208_), .A2(pi0778), .A3(new_n26171_), .A4(new_n26198_), .ZN(new_n26209_));
  XNOR2_X1   g23000(.A1(new_n26209_), .A2(new_n26205_), .ZN(new_n26210_));
  NAND2_X1   g23001(.A1(new_n26210_), .A2(new_n13801_), .ZN(new_n26211_));
  NOR2_X1    g23002(.A1(new_n26210_), .A2(new_n13778_), .ZN(new_n26212_));
  XOR2_X1    g23003(.A1(new_n26212_), .A2(new_n14694_), .Z(new_n26213_));
  NOR2_X1    g23004(.A1(new_n26213_), .A2(new_n26165_), .ZN(new_n26214_));
  NOR3_X1    g23005(.A1(new_n26214_), .A2(new_n13783_), .A3(new_n26173_), .ZN(new_n26215_));
  NOR3_X1    g23006(.A1(new_n26215_), .A2(pi0660), .A3(new_n26176_), .ZN(new_n26216_));
  NOR2_X1    g23007(.A1(new_n26210_), .A2(new_n13766_), .ZN(new_n26217_));
  XOR2_X1    g23008(.A1(new_n26217_), .A2(new_n14090_), .Z(new_n26218_));
  NAND3_X1   g23009(.A1(new_n26218_), .A2(pi0785), .A3(new_n26164_), .ZN(new_n26219_));
  OAI21_X1   g23010(.A1(new_n26216_), .A2(new_n26219_), .B(new_n26211_), .ZN(new_n26220_));
  NAND2_X1   g23011(.A1(new_n26220_), .A2(new_n13855_), .ZN(new_n26221_));
  NOR2_X1    g23012(.A1(new_n26220_), .A2(new_n13816_), .ZN(new_n26222_));
  XOR2_X1    g23013(.A1(new_n26222_), .A2(new_n13818_), .Z(new_n26223_));
  NAND2_X1   g23014(.A1(new_n26223_), .A2(new_n26166_), .ZN(new_n26224_));
  NAND3_X1   g23015(.A1(new_n26224_), .A2(new_n13823_), .A3(new_n26182_), .ZN(new_n26225_));
  AND3_X2    g23016(.A1(new_n26225_), .A2(new_n13823_), .A3(new_n26180_), .Z(new_n26226_));
  NOR2_X1    g23017(.A1(new_n26220_), .A2(new_n13817_), .ZN(new_n26227_));
  XOR2_X1    g23018(.A1(new_n26227_), .A2(new_n13819_), .Z(new_n26228_));
  NOR3_X1    g23019(.A1(new_n26228_), .A2(new_n13855_), .A3(new_n26167_), .ZN(new_n26229_));
  INV_X1     g23020(.I(new_n26229_), .ZN(new_n26230_));
  OAI21_X1   g23021(.A1(new_n26226_), .A2(new_n26230_), .B(new_n26221_), .ZN(new_n26231_));
  NOR2_X1    g23022(.A1(new_n26231_), .A2(new_n13860_), .ZN(new_n26232_));
  XOR2_X1    g23023(.A1(new_n26232_), .A2(new_n13904_), .Z(new_n26233_));
  NOR2_X1    g23024(.A1(new_n26233_), .A2(new_n26169_), .ZN(new_n26234_));
  NAND2_X1   g23025(.A1(new_n26191_), .A2(new_n13884_), .ZN(new_n26235_));
  INV_X1     g23026(.I(new_n26231_), .ZN(new_n26236_));
  AOI21_X1   g23027(.A1(new_n26236_), .A2(new_n14143_), .B(pi0789), .ZN(new_n26237_));
  OAI21_X1   g23028(.A1(new_n26234_), .A2(new_n26235_), .B(new_n26237_), .ZN(new_n26238_));
  NOR2_X1    g23029(.A1(new_n26231_), .A2(new_n13868_), .ZN(new_n26239_));
  XOR2_X1    g23030(.A1(new_n26239_), .A2(new_n13903_), .Z(new_n26240_));
  NAND2_X1   g23031(.A1(new_n26187_), .A2(new_n19018_), .ZN(new_n26241_));
  AOI21_X1   g23032(.A1(new_n26240_), .A2(new_n26168_), .B(new_n26241_), .ZN(new_n26242_));
  AOI21_X1   g23033(.A1(new_n26238_), .A2(new_n26242_), .B(new_n26196_), .ZN(new_n26243_));
  NAND2_X1   g23034(.A1(new_n26193_), .A2(new_n16372_), .ZN(new_n26244_));
  OAI21_X1   g23035(.A1(new_n16372_), .A2(new_n26155_), .B(new_n26244_), .ZN(new_n26245_));
  NAND3_X1   g23036(.A1(new_n26245_), .A2(new_n18929_), .A3(new_n26170_), .ZN(new_n26246_));
  NAND2_X1   g23037(.A1(new_n26246_), .A2(new_n16569_), .ZN(new_n26247_));
  XOR2_X1    g23038(.A1(new_n26247_), .A2(new_n16572_), .Z(new_n26248_));
  AOI21_X1   g23039(.A1(new_n19022_), .A2(new_n26246_), .B(new_n26248_), .ZN(new_n26249_));
  INV_X1     g23040(.I(new_n26155_), .ZN(new_n26250_));
  NAND2_X1   g23041(.A1(new_n26193_), .A2(new_n13963_), .ZN(new_n26251_));
  XNOR2_X1   g23042(.A1(new_n26251_), .A2(new_n19028_), .ZN(new_n26252_));
  NOR3_X1    g23043(.A1(new_n26252_), .A2(new_n16424_), .A3(new_n26250_), .ZN(new_n26253_));
  OAI21_X1   g23044(.A1(new_n26249_), .A2(new_n16574_), .B(new_n26253_), .ZN(new_n26254_));
  NOR4_X1    g23045(.A1(new_n26169_), .A2(new_n14060_), .A3(new_n14163_), .A4(new_n18928_), .ZN(new_n26255_));
  NOR2_X1    g23046(.A1(new_n26255_), .A2(new_n14005_), .ZN(new_n26256_));
  XOR2_X1    g23047(.A1(new_n26256_), .A2(new_n14007_), .Z(new_n26257_));
  NAND2_X1   g23048(.A1(new_n26257_), .A2(new_n26155_), .ZN(new_n26258_));
  NOR2_X1    g23049(.A1(new_n26250_), .A2(pi0647), .ZN(new_n26259_));
  AOI21_X1   g23050(.A1(new_n26255_), .A2(pi0647), .B(new_n26259_), .ZN(new_n26260_));
  NOR2_X1    g23051(.A1(new_n26245_), .A2(new_n13994_), .ZN(new_n26261_));
  XNOR2_X1   g23052(.A1(new_n26261_), .A2(new_n19033_), .ZN(new_n26262_));
  AOI22_X1   g23053(.A1(new_n26262_), .A2(new_n26155_), .B1(new_n14206_), .B2(new_n26260_), .ZN(new_n26263_));
  NOR3_X1    g23054(.A1(new_n26263_), .A2(new_n14010_), .A3(new_n26258_), .ZN(new_n26264_));
  OAI22_X1   g23055(.A1(new_n26243_), .A2(new_n26254_), .B1(new_n12776_), .B2(new_n26264_), .ZN(new_n26265_));
  AOI21_X1   g23056(.A1(new_n26260_), .A2(pi1157), .B(new_n12776_), .ZN(new_n26266_));
  AOI22_X1   g23057(.A1(new_n26258_), .A2(new_n26266_), .B1(new_n12776_), .B2(new_n26255_), .ZN(new_n26267_));
  NAND2_X1   g23058(.A1(new_n26265_), .A2(pi0644), .ZN(new_n26268_));
  XOR2_X1    g23059(.A1(new_n26268_), .A2(new_n14205_), .Z(new_n26269_));
  NOR2_X1    g23060(.A1(new_n26269_), .A2(new_n26267_), .ZN(new_n26270_));
  NOR2_X1    g23061(.A1(new_n26245_), .A2(new_n18968_), .ZN(new_n26271_));
  NAND2_X1   g23062(.A1(new_n18967_), .A2(new_n26155_), .ZN(new_n26272_));
  XOR2_X1    g23063(.A1(new_n26271_), .A2(new_n26272_), .Z(new_n26273_));
  NAND2_X1   g23064(.A1(new_n26273_), .A2(pi0715), .ZN(new_n26274_));
  XOR2_X1    g23065(.A1(new_n26274_), .A2(new_n14205_), .Z(new_n26275_));
  OAI21_X1   g23066(.A1(new_n26275_), .A2(new_n26250_), .B(new_n14203_), .ZN(new_n26276_));
  NAND2_X1   g23067(.A1(new_n26273_), .A2(pi0644), .ZN(new_n26277_));
  XOR2_X1    g23068(.A1(new_n26277_), .A2(new_n14217_), .Z(new_n26278_));
  AOI21_X1   g23069(.A1(new_n26278_), .A2(new_n26155_), .B(pi1160), .ZN(new_n26279_));
  OAI21_X1   g23070(.A1(new_n26270_), .A2(new_n26276_), .B(new_n26279_), .ZN(new_n26280_));
  NAND2_X1   g23071(.A1(new_n26265_), .A2(pi0715), .ZN(new_n26281_));
  XOR2_X1    g23072(.A1(new_n26281_), .A2(new_n14205_), .Z(new_n26282_));
  NOR2_X1    g23073(.A1(new_n26282_), .A2(new_n26267_), .ZN(new_n26283_));
  AOI21_X1   g23074(.A1(new_n26280_), .A2(new_n26283_), .B(new_n14799_), .ZN(new_n26284_));
  XOR2_X1    g23075(.A1(new_n26284_), .A2(new_n14801_), .Z(new_n26285_));
  NOR2_X1    g23076(.A1(new_n7240_), .A2(pi0194), .ZN(new_n26286_));
  NOR4_X1    g23077(.A1(new_n26285_), .A2(pi0832), .A3(new_n26265_), .A4(new_n26286_), .ZN(new_n26287_));
  AOI21_X1   g23078(.A1(new_n26154_), .A2(new_n7240_), .B(new_n26287_), .ZN(new_n26288_));
  NOR3_X1    g23079(.A1(new_n26153_), .A2(new_n26143_), .A3(new_n14200_), .ZN(new_n26289_));
  NOR2_X1    g23080(.A1(new_n26289_), .A2(new_n14217_), .ZN(new_n26290_));
  NOR4_X1    g23081(.A1(new_n26153_), .A2(new_n26143_), .A3(pi0644), .A4(new_n14200_), .ZN(new_n26291_));
  NOR2_X1    g23082(.A1(new_n26290_), .A2(new_n26291_), .ZN(new_n26292_));
  OAI21_X1   g23083(.A1(new_n12776_), .A2(new_n26150_), .B(new_n26152_), .ZN(new_n26293_));
  INV_X1     g23084(.I(new_n26136_), .ZN(new_n26294_));
  OAI21_X1   g23085(.A1(new_n26112_), .A2(new_n26121_), .B(new_n26294_), .ZN(new_n26295_));
  NAND2_X1   g23086(.A1(new_n26137_), .A2(new_n26138_), .ZN(new_n26296_));
  NAND2_X1   g23087(.A1(new_n26296_), .A2(new_n25909_), .ZN(new_n26297_));
  NOR2_X1    g23088(.A1(new_n26140_), .A2(new_n16329_), .ZN(new_n26298_));
  NAND2_X1   g23089(.A1(new_n26298_), .A2(new_n26297_), .ZN(new_n26299_));
  AOI21_X1   g23090(.A1(new_n26299_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n26300_));
  OAI21_X1   g23091(.A1(new_n26112_), .A2(new_n26121_), .B(new_n26300_), .ZN(new_n26301_));
  NAND3_X1   g23092(.A1(new_n26301_), .A2(new_n26295_), .A3(pi0787), .ZN(new_n26302_));
  NOR4_X1    g23093(.A1(new_n26297_), .A2(new_n26131_), .A3(new_n12776_), .A4(new_n26125_), .ZN(new_n26303_));
  NAND3_X1   g23094(.A1(new_n26139_), .A2(pi0787), .A3(new_n26129_), .ZN(new_n26304_));
  AND3_X2    g23095(.A1(new_n26304_), .A2(pi0787), .A3(new_n26131_), .Z(new_n26305_));
  NOR2_X1    g23096(.A1(new_n26305_), .A2(new_n26303_), .ZN(new_n26306_));
  INV_X1     g23097(.I(new_n14815_), .ZN(new_n26307_));
  NOR2_X1    g23098(.A1(new_n25954_), .A2(new_n14211_), .ZN(new_n26308_));
  AOI21_X1   g23099(.A1(new_n26134_), .A2(new_n14211_), .B(new_n26308_), .ZN(new_n26309_));
  OAI21_X1   g23100(.A1(new_n25954_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n26310_));
  AOI21_X1   g23101(.A1(new_n26309_), .A2(new_n26310_), .B(new_n26307_), .ZN(new_n26311_));
  OAI21_X1   g23102(.A1(new_n26306_), .A2(new_n14204_), .B(new_n26311_), .ZN(new_n26312_));
  AOI22_X1   g23103(.A1(new_n26302_), .A2(new_n26293_), .B1(new_n14204_), .B2(new_n26312_), .ZN(new_n26313_));
  AOI21_X1   g23104(.A1(new_n25954_), .A2(new_n14254_), .B(pi0644), .ZN(new_n26314_));
  NOR3_X1    g23105(.A1(new_n26306_), .A2(new_n26309_), .A3(new_n26314_), .ZN(new_n26315_));
  OAI21_X1   g23106(.A1(new_n26313_), .A2(pi0790), .B(new_n26315_), .ZN(new_n26316_));
  NOR3_X1    g23107(.A1(new_n26292_), .A2(new_n26316_), .A3(new_n26288_), .ZN(po0351));
  NOR2_X1    g23108(.A1(pi0171), .A2(pi0299), .ZN(new_n26318_));
  OAI21_X1   g23109(.A1(new_n6448_), .A2(new_n26318_), .B(pi0232), .ZN(new_n26319_));
  NAND2_X1   g23110(.A1(new_n9281_), .A2(pi0192), .ZN(new_n26320_));
  XOR2_X1    g23111(.A1(new_n26320_), .A2(new_n12449_), .Z(new_n26321_));
  NAND2_X1   g23112(.A1(new_n12737_), .A2(new_n26321_), .ZN(new_n26322_));
  XNOR2_X1   g23113(.A1(new_n26322_), .A2(new_n26319_), .ZN(new_n26323_));
  NOR2_X1    g23114(.A1(new_n12456_), .A2(new_n3098_), .ZN(new_n26324_));
  AOI21_X1   g23115(.A1(new_n7855_), .A2(new_n26324_), .B(pi0171), .ZN(new_n26325_));
  OAI21_X1   g23116(.A1(new_n12745_), .A2(new_n26325_), .B(new_n5551_), .ZN(new_n26326_));
  NOR3_X1    g23117(.A1(new_n12686_), .A2(new_n12450_), .A3(new_n12749_), .ZN(new_n26327_));
  AOI21_X1   g23118(.A1(new_n26327_), .A2(new_n26326_), .B(pi0192), .ZN(new_n26328_));
  NAND2_X1   g23119(.A1(new_n12753_), .A2(pi0192), .ZN(new_n26329_));
  NAND2_X1   g23120(.A1(new_n12695_), .A2(new_n12450_), .ZN(new_n26330_));
  AOI21_X1   g23121(.A1(new_n26330_), .A2(new_n26329_), .B(new_n5551_), .ZN(new_n26331_));
  NOR2_X1    g23122(.A1(new_n12757_), .A2(new_n3989_), .ZN(new_n26332_));
  OAI21_X1   g23123(.A1(new_n26331_), .A2(new_n7605_), .B(new_n26332_), .ZN(new_n26333_));
  AOI21_X1   g23124(.A1(new_n26333_), .A2(new_n3417_), .B(new_n12752_), .ZN(new_n26334_));
  OAI21_X1   g23125(.A1(new_n26334_), .A2(new_n12761_), .B(new_n12762_), .ZN(new_n26335_));
  NOR3_X1    g23126(.A1(new_n26328_), .A2(new_n12678_), .A3(new_n26335_), .ZN(new_n26336_));
  NAND2_X1   g23127(.A1(new_n12723_), .A2(new_n7954_), .ZN(new_n26337_));
  NOR2_X1    g23128(.A1(new_n26337_), .A2(new_n7957_), .ZN(new_n26338_));
  NAND2_X1   g23129(.A1(new_n26338_), .A2(new_n3225_), .ZN(new_n26339_));
  AOI21_X1   g23130(.A1(new_n7956_), .A2(new_n10754_), .B(new_n26339_), .ZN(new_n26340_));
  AOI22_X1   g23131(.A1(new_n8346_), .A2(pi0195), .B1(new_n12723_), .B2(new_n7954_), .ZN(new_n26341_));
  NOR3_X1    g23132(.A1(new_n26341_), .A2(new_n3183_), .A3(new_n7957_), .ZN(new_n26342_));
  OAI21_X1   g23133(.A1(new_n12672_), .A2(new_n26342_), .B(new_n12442_), .ZN(new_n26343_));
  NOR2_X1    g23134(.A1(new_n12712_), .A2(new_n26343_), .ZN(new_n26344_));
  OAI21_X1   g23135(.A1(new_n26336_), .A2(new_n26340_), .B(new_n26344_), .ZN(new_n26345_));
  AOI21_X1   g23136(.A1(new_n26345_), .A2(new_n3183_), .B(new_n26323_), .ZN(po0352));
  NOR2_X1    g23137(.A1(new_n10694_), .A2(new_n6448_), .ZN(new_n26347_));
  OAI21_X1   g23138(.A1(new_n5689_), .A2(new_n4150_), .B(new_n9241_), .ZN(new_n26348_));
  OAI21_X1   g23139(.A1(new_n26347_), .A2(new_n26348_), .B(pi0232), .ZN(new_n26349_));
  NAND2_X1   g23140(.A1(new_n10297_), .A2(pi0232), .ZN(new_n26350_));
  NOR3_X1    g23141(.A1(new_n9283_), .A2(new_n12664_), .A3(new_n26350_), .ZN(new_n26351_));
  XOR2_X1    g23142(.A1(new_n26351_), .A2(new_n26349_), .Z(new_n26352_));
  NOR2_X1    g23143(.A1(new_n26352_), .A2(new_n3098_), .ZN(new_n26353_));
  OAI21_X1   g23144(.A1(new_n9281_), .A2(pi0299), .B(pi0039), .ZN(new_n26354_));
  NOR2_X1    g23145(.A1(new_n26353_), .A2(new_n26354_), .ZN(new_n26355_));
  XOR2_X1    g23146(.A1(new_n26355_), .A2(new_n3262_), .Z(new_n26356_));
  AOI21_X1   g23147(.A1(new_n12673_), .A2(new_n8648_), .B(new_n12520_), .ZN(new_n26357_));
  AOI21_X1   g23148(.A1(new_n26356_), .A2(new_n26357_), .B(new_n8345_), .ZN(new_n26358_));
  NOR2_X1    g23149(.A1(new_n8345_), .A2(new_n12522_), .ZN(new_n26359_));
  XOR2_X1    g23150(.A1(new_n26358_), .A2(new_n26359_), .Z(new_n26360_));
  NAND2_X1   g23151(.A1(new_n26352_), .A2(pi0039), .ZN(new_n26361_));
  XOR2_X1    g23152(.A1(new_n26361_), .A2(new_n4368_), .Z(new_n26362_));
  OAI21_X1   g23153(.A1(new_n12673_), .A2(new_n6494_), .B(new_n3098_), .ZN(new_n26363_));
  NAND4_X1   g23154(.A1(new_n26360_), .A2(pi0170), .A3(new_n26362_), .A4(new_n26363_), .ZN(new_n26364_));
  AOI21_X1   g23155(.A1(new_n12700_), .A2(pi0232), .B(new_n12694_), .ZN(new_n26365_));
  AOI21_X1   g23156(.A1(new_n4150_), .A2(new_n7613_), .B(new_n12704_), .ZN(new_n26366_));
  NOR2_X1    g23157(.A1(new_n7604_), .A2(new_n3183_), .ZN(new_n26367_));
  OAI21_X1   g23158(.A1(new_n26366_), .A2(new_n7440_), .B(new_n26367_), .ZN(new_n26368_));
  NOR2_X1    g23159(.A1(new_n26365_), .A2(new_n26368_), .ZN(new_n26369_));
  OAI21_X1   g23160(.A1(new_n26369_), .A2(pi0232), .B(new_n12702_), .ZN(new_n26370_));
  NAND3_X1   g23161(.A1(new_n26370_), .A2(new_n3259_), .A3(pi0194), .ZN(new_n26371_));
  INV_X1     g23162(.I(new_n26371_), .ZN(new_n26372_));
  INV_X1     g23163(.I(new_n26369_), .ZN(new_n26373_));
  AOI21_X1   g23164(.A1(new_n3259_), .A2(new_n12522_), .B(new_n26373_), .ZN(new_n26374_));
  INV_X1     g23165(.I(new_n12678_), .ZN(new_n26375_));
  OAI21_X1   g23166(.A1(new_n26371_), .A2(new_n12749_), .B(new_n5551_), .ZN(new_n26376_));
  AOI21_X1   g23167(.A1(new_n26375_), .A2(new_n26374_), .B(new_n26376_), .ZN(new_n26377_));
  NOR3_X1    g23168(.A1(new_n7776_), .A2(new_n7855_), .A3(new_n12520_), .ZN(new_n26378_));
  NOR3_X1    g23169(.A1(new_n7775_), .A2(new_n7854_), .A3(new_n12520_), .ZN(new_n26379_));
  NOR2_X1    g23170(.A1(new_n3462_), .A2(new_n3098_), .ZN(new_n26380_));
  OAI21_X1   g23171(.A1(new_n26378_), .A2(new_n26379_), .B(new_n26380_), .ZN(new_n26381_));
  OAI22_X1   g23172(.A1(new_n26377_), .A2(new_n26381_), .B1(new_n26372_), .B2(new_n26374_), .ZN(new_n26382_));
  NAND4_X1   g23173(.A1(new_n26382_), .A2(new_n12687_), .A3(new_n12713_), .A4(new_n12715_), .ZN(new_n26383_));
  AOI21_X1   g23174(.A1(new_n26383_), .A2(new_n3225_), .B(new_n10754_), .ZN(new_n26384_));
  NOR2_X1    g23175(.A1(new_n26384_), .A2(new_n7957_), .ZN(new_n26385_));
  XNOR2_X1   g23176(.A1(new_n26385_), .A2(new_n26338_), .ZN(new_n26386_));
  NOR2_X1    g23177(.A1(new_n26384_), .A2(new_n26337_), .ZN(new_n26387_));
  NOR3_X1    g23178(.A1(new_n26337_), .A2(new_n7956_), .A3(pi0196), .ZN(new_n26388_));
  XNOR2_X1   g23179(.A1(new_n26387_), .A2(new_n26388_), .ZN(new_n26389_));
  AOI21_X1   g23180(.A1(new_n26386_), .A2(new_n26389_), .B(new_n26364_), .ZN(po0353));
  NOR2_X1    g23181(.A1(new_n5800_), .A2(pi0767), .ZN(new_n26391_));
  NOR2_X1    g23182(.A1(new_n14298_), .A2(new_n26391_), .ZN(new_n26392_));
  XOR2_X1    g23183(.A1(new_n26392_), .A2(new_n13094_), .Z(new_n26393_));
  NAND2_X1   g23184(.A1(new_n26393_), .A2(pi0197), .ZN(new_n26394_));
  NAND3_X1   g23185(.A1(new_n17057_), .A2(pi0197), .A3(pi0767), .ZN(new_n26395_));
  NAND3_X1   g23186(.A1(new_n17058_), .A2(pi0197), .A3(new_n16517_), .ZN(new_n26396_));
  NAND2_X1   g23187(.A1(new_n26396_), .A2(new_n26395_), .ZN(new_n26397_));
  AOI21_X1   g23188(.A1(new_n26397_), .A2(new_n17042_), .B(pi0039), .ZN(new_n26398_));
  NOR2_X1    g23189(.A1(new_n5665_), .A2(new_n3098_), .ZN(new_n26399_));
  XOR2_X1    g23190(.A1(new_n17157_), .A2(new_n26399_), .Z(new_n26400_));
  OAI21_X1   g23191(.A1(new_n16973_), .A2(new_n16517_), .B(new_n5665_), .ZN(new_n26401_));
  NOR2_X1    g23192(.A1(new_n16981_), .A2(new_n3259_), .ZN(new_n26402_));
  NAND4_X1   g23193(.A1(new_n26400_), .A2(new_n16971_), .A3(new_n26401_), .A4(new_n26402_), .ZN(new_n26403_));
  OAI21_X1   g23194(.A1(new_n26398_), .A2(new_n26403_), .B(new_n26394_), .ZN(new_n26404_));
  AOI21_X1   g23195(.A1(new_n26404_), .A2(new_n16970_), .B(new_n16550_), .ZN(new_n26405_));
  NOR3_X1    g23196(.A1(new_n17125_), .A2(new_n5665_), .A3(new_n3098_), .ZN(new_n26406_));
  NOR3_X1    g23197(.A1(new_n17076_), .A2(new_n3098_), .A3(new_n26399_), .ZN(new_n26407_));
  OAI21_X1   g23198(.A1(new_n26406_), .A2(new_n26407_), .B(new_n17133_), .ZN(new_n26408_));
  OAI21_X1   g23199(.A1(pi0197), .A2(new_n16971_), .B(new_n17087_), .ZN(new_n26409_));
  NOR2_X1    g23200(.A1(pi0039), .A2(pi0197), .ZN(new_n26410_));
  NOR3_X1    g23201(.A1(new_n26410_), .A2(new_n3259_), .A3(pi0767), .ZN(new_n26411_));
  OAI21_X1   g23202(.A1(new_n13109_), .A2(new_n26391_), .B(new_n26411_), .ZN(new_n26412_));
  AOI21_X1   g23203(.A1(new_n26394_), .A2(new_n3259_), .B(new_n26412_), .ZN(new_n26413_));
  NAND4_X1   g23204(.A1(new_n26408_), .A2(new_n14366_), .A3(new_n26409_), .A4(new_n26413_), .ZN(new_n26414_));
  NAND2_X1   g23205(.A1(new_n26414_), .A2(new_n5665_), .ZN(new_n26415_));
  OR3_X2     g23206(.A1(new_n17176_), .A2(new_n16517_), .A3(new_n5800_), .Z(new_n26416_));
  NAND4_X1   g23207(.A1(new_n13624_), .A2(pi0197), .A3(pi0698), .A4(new_n13108_), .ZN(new_n26417_));
  AOI21_X1   g23208(.A1(new_n3259_), .A2(new_n26416_), .B(new_n26417_), .ZN(new_n26418_));
  NAND2_X1   g23209(.A1(new_n26415_), .A2(new_n26418_), .ZN(new_n26419_));
  OAI21_X1   g23210(.A1(new_n26405_), .A2(new_n26419_), .B(new_n8297_), .ZN(new_n26420_));
  AOI21_X1   g23211(.A1(new_n26405_), .A2(new_n26419_), .B(new_n26420_), .ZN(new_n26421_));
  XOR2_X1    g23212(.A1(new_n26421_), .A2(new_n17184_), .Z(new_n26422_));
  AOI21_X1   g23213(.A1(new_n16550_), .A2(new_n16968_), .B(new_n26391_), .ZN(new_n26423_));
  NOR2_X1    g23214(.A1(new_n26423_), .A2(new_n14799_), .ZN(new_n26424_));
  XOR2_X1    g23215(.A1(new_n26424_), .A2(new_n16913_), .Z(new_n26425_));
  OAI21_X1   g23216(.A1(new_n26422_), .A2(new_n26425_), .B(pi0197), .ZN(po0354));
  NAND2_X1   g23217(.A1(new_n13417_), .A2(pi0198), .ZN(new_n26427_));
  NAND2_X1   g23218(.A1(new_n26427_), .A2(new_n5398_), .ZN(new_n26428_));
  XOR2_X1    g23219(.A1(new_n26428_), .A2(new_n12981_), .Z(new_n26429_));
  INV_X1     g23220(.I(new_n26429_), .ZN(new_n26430_));
  NAND3_X1   g23221(.A1(new_n12922_), .A2(pi0198), .A3(new_n5383_), .ZN(new_n26431_));
  NAND3_X1   g23222(.A1(new_n12930_), .A2(pi0198), .A3(new_n5796_), .ZN(new_n26432_));
  AOI21_X1   g23223(.A1(new_n26432_), .A2(new_n26431_), .B(new_n12862_), .ZN(new_n26433_));
  NOR2_X1    g23224(.A1(new_n13334_), .A2(new_n3072_), .ZN(new_n26434_));
  NOR2_X1    g23225(.A1(new_n12784_), .A2(new_n3072_), .ZN(new_n26435_));
  OAI21_X1   g23226(.A1(po1101), .A2(new_n26435_), .B(new_n26434_), .ZN(new_n26436_));
  NOR2_X1    g23227(.A1(new_n26436_), .A2(new_n3090_), .ZN(new_n26437_));
  OAI21_X1   g23228(.A1(new_n26437_), .A2(new_n26433_), .B(new_n5398_), .ZN(new_n26438_));
  NAND2_X1   g23229(.A1(new_n26438_), .A2(new_n3098_), .ZN(new_n26439_));
  INV_X1     g23230(.I(new_n26435_), .ZN(new_n26440_));
  NOR2_X1    g23231(.A1(new_n12949_), .A2(new_n3072_), .ZN(new_n26441_));
  NAND2_X1   g23232(.A1(new_n26441_), .A2(po1101), .ZN(new_n26442_));
  OAI21_X1   g23233(.A1(po1101), .A2(new_n26440_), .B(new_n26442_), .ZN(new_n26443_));
  AOI21_X1   g23234(.A1(new_n26440_), .A2(new_n3091_), .B(pi0223), .ZN(new_n26444_));
  NAND4_X1   g23235(.A1(new_n26430_), .A2(new_n26439_), .A3(new_n26443_), .A4(new_n26444_), .ZN(new_n26445_));
  NOR3_X1    g23236(.A1(new_n3290_), .A2(pi0038), .A3(new_n3183_), .ZN(new_n26446_));
  AND2_X2    g23237(.A1(new_n26445_), .A2(new_n26446_), .Z(new_n26447_));
  NAND2_X1   g23238(.A1(new_n26427_), .A2(new_n5454_), .ZN(new_n26448_));
  XOR2_X1    g23239(.A1(new_n26448_), .A2(new_n13516_), .Z(new_n26449_));
  INV_X1     g23240(.I(new_n26449_), .ZN(new_n26450_));
  NOR2_X1    g23241(.A1(new_n26436_), .A2(new_n3111_), .ZN(new_n26451_));
  OAI21_X1   g23242(.A1(new_n26451_), .A2(new_n26433_), .B(new_n5454_), .ZN(new_n26452_));
  NAND2_X1   g23243(.A1(new_n26452_), .A2(new_n3098_), .ZN(new_n26453_));
  NOR2_X1    g23244(.A1(new_n26435_), .A2(new_n3313_), .ZN(new_n26454_));
  NOR3_X1    g23245(.A1(new_n26454_), .A2(new_n3072_), .A3(pi0215), .ZN(new_n26455_));
  AND4_X2    g23246(.A1(new_n26443_), .A2(new_n26450_), .A3(new_n26453_), .A4(new_n26455_), .Z(new_n26456_));
  NOR2_X1    g23247(.A1(new_n26447_), .A2(new_n26456_), .ZN(new_n26457_));
  NOR2_X1    g23248(.A1(new_n26457_), .A2(new_n13994_), .ZN(new_n26458_));
  INV_X1     g23249(.I(new_n26458_), .ZN(new_n26459_));
  INV_X1     g23250(.I(new_n26457_), .ZN(new_n26460_));
  NOR2_X1    g23251(.A1(new_n26460_), .A2(new_n16372_), .ZN(new_n26461_));
  INV_X1     g23252(.I(new_n26461_), .ZN(new_n26462_));
  INV_X1     g23253(.I(pi0633), .ZN(new_n26463_));
  NOR2_X1    g23254(.A1(new_n3072_), .A2(new_n26463_), .ZN(new_n26464_));
  NAND3_X1   g23255(.A1(new_n12794_), .A2(new_n13203_), .A3(new_n26464_), .ZN(new_n26465_));
  INV_X1     g23256(.I(new_n26464_), .ZN(new_n26466_));
  NAND3_X1   g23257(.A1(new_n12794_), .A2(new_n13103_), .A3(new_n26466_), .ZN(new_n26467_));
  NAND2_X1   g23258(.A1(new_n26465_), .A2(new_n26467_), .ZN(new_n26468_));
  NOR2_X1    g23259(.A1(new_n26468_), .A2(new_n3259_), .ZN(new_n26469_));
  XOR2_X1    g23260(.A1(new_n26469_), .A2(new_n3262_), .Z(new_n26470_));
  AOI21_X1   g23261(.A1(new_n26470_), .A2(pi0198), .B(new_n3290_), .ZN(new_n26471_));
  INV_X1     g23262(.I(new_n26471_), .ZN(new_n26472_));
  NOR2_X1    g23263(.A1(new_n12818_), .A2(new_n3072_), .ZN(new_n26473_));
  AOI21_X1   g23264(.A1(pi0633), .A2(new_n13423_), .B(new_n26473_), .ZN(new_n26474_));
  NOR2_X1    g23265(.A1(new_n26474_), .A2(new_n5794_), .ZN(new_n26475_));
  NOR2_X1    g23266(.A1(new_n26475_), .A2(new_n5636_), .ZN(new_n26476_));
  NOR3_X1    g23267(.A1(new_n12809_), .A2(new_n13102_), .A3(new_n26466_), .ZN(new_n26477_));
  NOR3_X1    g23268(.A1(new_n12809_), .A2(new_n13230_), .A3(new_n26464_), .ZN(new_n26478_));
  NOR2_X1    g23269(.A1(new_n26477_), .A2(new_n26478_), .ZN(new_n26479_));
  NOR2_X1    g23270(.A1(new_n13336_), .A2(pi0603), .ZN(new_n26480_));
  NAND2_X1   g23271(.A1(new_n26474_), .A2(new_n5373_), .ZN(new_n26482_));
  AOI21_X1   g23272(.A1(new_n13336_), .A2(new_n26475_), .B(new_n26482_), .ZN(new_n26483_));
  NAND3_X1   g23273(.A1(new_n26483_), .A2(new_n5378_), .A3(new_n26473_), .ZN(new_n26484_));
  XOR2_X1    g23274(.A1(new_n26484_), .A2(new_n26476_), .Z(new_n26485_));
  INV_X1     g23275(.I(new_n26479_), .ZN(new_n26486_));
  XOR2_X1    g23276(.A1(new_n26475_), .A2(new_n13282_), .Z(new_n26487_));
  NAND2_X1   g23277(.A1(new_n26487_), .A2(new_n26486_), .ZN(new_n26488_));
  NAND2_X1   g23278(.A1(new_n26488_), .A2(new_n5378_), .ZN(new_n26489_));
  NOR2_X1    g23279(.A1(new_n5382_), .A2(new_n5379_), .ZN(new_n26490_));
  NAND4_X1   g23280(.A1(new_n26486_), .A2(pi0603), .A3(new_n5381_), .A4(new_n26435_), .ZN(new_n26491_));
  AOI21_X1   g23281(.A1(new_n5379_), .A2(new_n26491_), .B(new_n26488_), .ZN(new_n26492_));
  NAND4_X1   g23282(.A1(new_n26492_), .A2(new_n5794_), .A3(new_n5378_), .A4(new_n26441_), .ZN(new_n26493_));
  XNOR2_X1   g23283(.A1(new_n26493_), .A2(new_n26489_), .ZN(new_n26494_));
  NAND2_X1   g23284(.A1(new_n26494_), .A2(new_n5454_), .ZN(new_n26495_));
  XOR2_X1    g23285(.A1(new_n26495_), .A2(new_n13516_), .Z(new_n26496_));
  OAI21_X1   g23286(.A1(new_n26496_), .A2(new_n26485_), .B(new_n3111_), .ZN(new_n26497_));
  NOR2_X1    g23287(.A1(new_n26479_), .A2(new_n5794_), .ZN(new_n26498_));
  AOI21_X1   g23288(.A1(new_n5794_), .A2(new_n26440_), .B(new_n26498_), .ZN(new_n26499_));
  NOR2_X1    g23289(.A1(new_n26499_), .A2(new_n3313_), .ZN(new_n26500_));
  AOI21_X1   g23290(.A1(new_n26497_), .A2(new_n26500_), .B(new_n5827_), .ZN(new_n26501_));
  NOR4_X1    g23291(.A1(new_n12862_), .A2(new_n26463_), .A3(new_n12809_), .A4(new_n13102_), .ZN(new_n26502_));
  NOR2_X1    g23292(.A1(new_n12862_), .A2(new_n3072_), .ZN(new_n26503_));
  OAI21_X1   g23293(.A1(new_n26502_), .A2(new_n26503_), .B(new_n5378_), .ZN(new_n26504_));
  NOR2_X1    g23294(.A1(new_n12922_), .A2(new_n13364_), .ZN(new_n26505_));
  NOR3_X1    g23295(.A1(new_n26433_), .A2(pi0633), .A3(new_n26505_), .ZN(new_n26506_));
  NOR3_X1    g23296(.A1(new_n26506_), .A2(new_n13388_), .A3(new_n14306_), .ZN(new_n26507_));
  XOR2_X1    g23297(.A1(new_n26507_), .A2(new_n26504_), .Z(new_n26508_));
  INV_X1     g23298(.I(new_n26508_), .ZN(new_n26509_));
  NOR3_X1    g23299(.A1(new_n26434_), .A2(pi0603), .A3(new_n26502_), .ZN(new_n26510_));
  NOR3_X1    g23300(.A1(new_n26510_), .A2(new_n5386_), .A3(new_n26486_), .ZN(new_n26511_));
  NOR2_X1    g23301(.A1(new_n26511_), .A2(new_n5636_), .ZN(new_n26512_));
  OAI21_X1   g23302(.A1(new_n26440_), .A2(pi0603), .B(new_n13336_), .ZN(new_n26513_));
  INV_X1     g23303(.I(new_n26499_), .ZN(new_n26514_));
  NAND3_X1   g23304(.A1(new_n26511_), .A2(new_n13336_), .A3(new_n26514_), .ZN(new_n26515_));
  XOR2_X1    g23305(.A1(new_n26515_), .A2(new_n26513_), .Z(new_n26516_));
  NAND3_X1   g23306(.A1(new_n26516_), .A2(new_n5378_), .A3(new_n26434_), .ZN(new_n26517_));
  XOR2_X1    g23307(.A1(new_n26517_), .A2(new_n26512_), .Z(new_n26518_));
  NAND2_X1   g23308(.A1(new_n26518_), .A2(pi0215), .ZN(new_n26519_));
  XOR2_X1    g23309(.A1(new_n26519_), .A2(new_n13309_), .Z(new_n26520_));
  NAND2_X1   g23310(.A1(new_n26520_), .A2(new_n26509_), .ZN(new_n26521_));
  OR2_X2     g23311(.A1(new_n13177_), .A2(new_n13175_), .Z(new_n26522_));
  NOR2_X1    g23312(.A1(new_n26522_), .A2(pi0198), .ZN(new_n26523_));
  AOI21_X1   g23313(.A1(pi0198), .A2(new_n14979_), .B(new_n26523_), .ZN(new_n26524_));
  NOR2_X1    g23314(.A1(new_n5794_), .A2(new_n26463_), .ZN(new_n26525_));
  NAND2_X1   g23315(.A1(new_n26524_), .A2(new_n26525_), .ZN(new_n26526_));
  NOR2_X1    g23316(.A1(new_n14336_), .A2(new_n3072_), .ZN(new_n26527_));
  NAND2_X1   g23317(.A1(new_n26527_), .A2(new_n26525_), .ZN(new_n26528_));
  XNOR2_X1   g23318(.A1(new_n26526_), .A2(new_n26528_), .ZN(new_n26529_));
  NAND2_X1   g23319(.A1(new_n26529_), .A2(pi0299), .ZN(new_n26530_));
  XOR2_X1    g23320(.A1(new_n26530_), .A2(new_n5827_), .Z(new_n26531_));
  NOR3_X1    g23321(.A1(new_n13160_), .A2(new_n3072_), .A3(new_n13039_), .ZN(new_n26532_));
  NOR2_X1    g23322(.A1(new_n13119_), .A2(new_n3072_), .ZN(new_n26533_));
  INV_X1     g23323(.I(new_n26533_), .ZN(new_n26534_));
  NOR3_X1    g23324(.A1(new_n13166_), .A2(new_n3072_), .A3(new_n13142_), .ZN(new_n26535_));
  AOI21_X1   g23325(.A1(new_n26534_), .A2(new_n26535_), .B(new_n26463_), .ZN(new_n26536_));
  OAI21_X1   g23326(.A1(new_n26534_), .A2(new_n26535_), .B(new_n26536_), .ZN(new_n26537_));
  INV_X1     g23327(.I(new_n26537_), .ZN(new_n26538_));
  OAI22_X1   g23328(.A1(new_n26538_), .A2(new_n26532_), .B1(pi0603), .B2(new_n14972_), .ZN(new_n26539_));
  OR2_X2     g23329(.A1(new_n26539_), .A2(new_n3259_), .Z(new_n26540_));
  OAI22_X1   g23330(.A1(new_n26501_), .A2(new_n26521_), .B1(new_n26531_), .B2(new_n26540_), .ZN(new_n26541_));
  NAND2_X1   g23331(.A1(new_n26514_), .A2(new_n3091_), .ZN(new_n26542_));
  NAND2_X1   g23332(.A1(new_n26518_), .A2(pi0223), .ZN(new_n26543_));
  XOR2_X1    g23333(.A1(new_n26543_), .A2(new_n13466_), .Z(new_n26544_));
  NOR2_X1    g23334(.A1(new_n26508_), .A2(new_n3098_), .ZN(new_n26545_));
  AOI22_X1   g23335(.A1(new_n26544_), .A2(new_n26545_), .B1(new_n3090_), .B2(new_n26542_), .ZN(new_n26546_));
  NAND2_X1   g23336(.A1(new_n26494_), .A2(new_n5398_), .ZN(new_n26547_));
  XOR2_X1    g23337(.A1(new_n26547_), .A2(new_n12981_), .Z(new_n26548_));
  NOR2_X1    g23338(.A1(new_n3290_), .A2(new_n3072_), .ZN(new_n26549_));
  INV_X1     g23339(.I(new_n26549_), .ZN(new_n26550_));
  NOR4_X1    g23340(.A1(new_n26546_), .A2(new_n26548_), .A3(new_n26485_), .A4(new_n26550_), .ZN(new_n26551_));
  NAND3_X1   g23341(.A1(new_n26541_), .A2(new_n26472_), .A3(new_n26551_), .ZN(new_n26552_));
  INV_X1     g23342(.I(new_n26552_), .ZN(new_n26553_));
  AOI21_X1   g23343(.A1(new_n26541_), .A2(new_n26551_), .B(new_n26472_), .ZN(new_n26554_));
  NOR2_X1    g23344(.A1(new_n13776_), .A2(new_n13766_), .ZN(new_n26555_));
  INV_X1     g23345(.I(new_n26555_), .ZN(new_n26556_));
  NOR3_X1    g23346(.A1(new_n26553_), .A2(new_n26554_), .A3(new_n26556_), .ZN(new_n26557_));
  NOR2_X1    g23347(.A1(new_n26457_), .A2(new_n26556_), .ZN(new_n26558_));
  INV_X1     g23348(.I(new_n26558_), .ZN(new_n26559_));
  NOR2_X1    g23349(.A1(new_n26557_), .A2(new_n26559_), .ZN(new_n26560_));
  NOR4_X1    g23350(.A1(new_n26553_), .A2(new_n26460_), .A3(new_n26554_), .A4(new_n26556_), .ZN(new_n26561_));
  NOR3_X1    g23351(.A1(new_n26560_), .A2(pi1155), .A3(new_n26561_), .ZN(new_n26562_));
  INV_X1     g23352(.I(new_n26554_), .ZN(new_n26563_));
  AOI21_X1   g23353(.A1(new_n26563_), .A2(new_n26552_), .B(new_n13775_), .ZN(new_n26564_));
  NOR2_X1    g23354(.A1(new_n26457_), .A2(new_n13776_), .ZN(new_n26565_));
  OAI21_X1   g23355(.A1(new_n26564_), .A2(new_n26565_), .B(pi0785), .ZN(new_n26566_));
  NOR4_X1    g23356(.A1(new_n26566_), .A2(new_n26560_), .A3(new_n13778_), .A4(new_n26561_), .ZN(new_n26567_));
  OAI21_X1   g23357(.A1(new_n13801_), .A2(new_n26562_), .B(new_n26567_), .ZN(new_n26568_));
  NOR2_X1    g23358(.A1(new_n26562_), .A2(new_n13801_), .ZN(new_n26569_));
  NOR2_X1    g23359(.A1(new_n26560_), .A2(new_n26561_), .ZN(new_n26570_));
  OAI21_X1   g23360(.A1(new_n26553_), .A2(new_n26554_), .B(new_n13776_), .ZN(new_n26571_));
  INV_X1     g23361(.I(new_n26565_), .ZN(new_n26572_));
  AOI21_X1   g23362(.A1(new_n26571_), .A2(new_n26572_), .B(new_n13801_), .ZN(new_n26573_));
  NAND3_X1   g23363(.A1(new_n26570_), .A2(pi1155), .A3(new_n26573_), .ZN(new_n26574_));
  NAND2_X1   g23364(.A1(new_n26569_), .A2(new_n26574_), .ZN(new_n26575_));
  NAND2_X1   g23365(.A1(new_n26575_), .A2(new_n26568_), .ZN(new_n26576_));
  NAND3_X1   g23366(.A1(new_n26576_), .A2(pi0618), .A3(pi1154), .ZN(new_n26577_));
  INV_X1     g23367(.I(new_n26570_), .ZN(new_n26578_));
  NOR4_X1    g23368(.A1(new_n26578_), .A2(pi0785), .A3(new_n13778_), .A4(new_n26566_), .ZN(new_n26579_));
  NOR3_X1    g23369(.A1(new_n26567_), .A2(new_n13801_), .A3(new_n26562_), .ZN(new_n26580_));
  NOR2_X1    g23370(.A1(new_n26579_), .A2(new_n26580_), .ZN(new_n26581_));
  NAND3_X1   g23371(.A1(new_n26581_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n26582_));
  AOI21_X1   g23372(.A1(new_n26577_), .A2(new_n26582_), .B(new_n26457_), .ZN(new_n26583_));
  NAND3_X1   g23373(.A1(new_n26576_), .A2(pi0618), .A3(pi1154), .ZN(new_n26584_));
  NAND3_X1   g23374(.A1(new_n26581_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n26585_));
  AOI21_X1   g23375(.A1(new_n26584_), .A2(new_n26585_), .B(new_n26457_), .ZN(new_n26586_));
  NAND4_X1   g23376(.A1(new_n26583_), .A2(new_n26586_), .A3(pi0781), .A4(new_n26576_), .ZN(new_n26587_));
  AOI21_X1   g23377(.A1(new_n26581_), .A2(pi0618), .B(new_n13819_), .ZN(new_n26588_));
  NOR3_X1    g23378(.A1(new_n26576_), .A2(new_n13816_), .A3(new_n13818_), .ZN(new_n26589_));
  OAI21_X1   g23379(.A1(new_n26589_), .A2(new_n26588_), .B(new_n26460_), .ZN(new_n26590_));
  NOR2_X1    g23380(.A1(new_n26581_), .A2(new_n13855_), .ZN(new_n26591_));
  NAND2_X1   g23381(.A1(new_n26586_), .A2(new_n26591_), .ZN(new_n26592_));
  NAND3_X1   g23382(.A1(new_n26592_), .A2(pi0781), .A3(new_n26590_), .ZN(new_n26593_));
  NAND2_X1   g23383(.A1(new_n26593_), .A2(new_n26587_), .ZN(new_n26594_));
  NAND3_X1   g23384(.A1(new_n26594_), .A2(pi0619), .A3(pi1159), .ZN(new_n26595_));
  AOI21_X1   g23385(.A1(new_n26581_), .A2(pi1154), .B(new_n13819_), .ZN(new_n26596_));
  NOR3_X1    g23386(.A1(new_n26576_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n26597_));
  OAI21_X1   g23387(.A1(new_n26597_), .A2(new_n26596_), .B(new_n26460_), .ZN(new_n26598_));
  NOR4_X1    g23388(.A1(new_n26598_), .A2(new_n26590_), .A3(new_n13855_), .A4(new_n26581_), .ZN(new_n26599_));
  NAND2_X1   g23389(.A1(new_n26590_), .A2(pi0781), .ZN(new_n26600_));
  NOR3_X1    g23390(.A1(new_n26598_), .A2(new_n13855_), .A3(new_n26581_), .ZN(new_n26601_));
  NOR2_X1    g23391(.A1(new_n26601_), .A2(new_n26600_), .ZN(new_n26602_));
  NOR2_X1    g23392(.A1(new_n26602_), .A2(new_n26599_), .ZN(new_n26603_));
  NAND3_X1   g23393(.A1(new_n26603_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n26604_));
  AOI21_X1   g23394(.A1(new_n26604_), .A2(new_n26595_), .B(new_n26457_), .ZN(new_n26605_));
  NAND3_X1   g23395(.A1(new_n26594_), .A2(pi0619), .A3(pi1159), .ZN(new_n26606_));
  NAND4_X1   g23396(.A1(new_n26593_), .A2(new_n13860_), .A3(pi1159), .A4(new_n26587_), .ZN(new_n26607_));
  AOI21_X1   g23397(.A1(new_n26606_), .A2(new_n26607_), .B(new_n26457_), .ZN(new_n26608_));
  NAND4_X1   g23398(.A1(new_n26605_), .A2(new_n26608_), .A3(pi0789), .A4(new_n26594_), .ZN(new_n26609_));
  AOI21_X1   g23399(.A1(new_n26603_), .A2(pi0619), .B(new_n13904_), .ZN(new_n26610_));
  NOR3_X1    g23400(.A1(new_n26594_), .A2(new_n13860_), .A3(pi1159), .ZN(new_n26611_));
  OAI21_X1   g23401(.A1(new_n26610_), .A2(new_n26611_), .B(new_n26460_), .ZN(new_n26612_));
  NOR2_X1    g23402(.A1(new_n26603_), .A2(new_n13896_), .ZN(new_n26613_));
  NAND2_X1   g23403(.A1(new_n26608_), .A2(new_n26613_), .ZN(new_n26614_));
  NAND3_X1   g23404(.A1(new_n26614_), .A2(pi0789), .A3(new_n26612_), .ZN(new_n26615_));
  NAND3_X1   g23405(.A1(new_n26615_), .A2(new_n16372_), .A3(new_n26609_), .ZN(new_n26616_));
  NAND3_X1   g23406(.A1(new_n26616_), .A2(new_n13994_), .A3(new_n26462_), .ZN(new_n26617_));
  NAND3_X1   g23407(.A1(new_n26617_), .A2(new_n16867_), .A3(new_n26459_), .ZN(new_n26618_));
  NOR2_X1    g23408(.A1(new_n26457_), .A2(pi0647), .ZN(new_n26619_));
  NOR2_X1    g23409(.A1(new_n26457_), .A2(new_n13880_), .ZN(new_n26620_));
  INV_X1     g23410(.I(new_n26620_), .ZN(new_n26621_));
  NOR2_X1    g23411(.A1(new_n26460_), .A2(new_n13805_), .ZN(new_n26622_));
  INV_X1     g23412(.I(new_n26622_), .ZN(new_n26623_));
  INV_X1     g23413(.I(pi0634), .ZN(new_n26624_));
  NOR2_X1    g23414(.A1(new_n3072_), .A2(new_n26624_), .ZN(new_n26625_));
  INV_X1     g23415(.I(new_n26625_), .ZN(new_n26626_));
  NAND3_X1   g23416(.A1(new_n12794_), .A2(new_n13205_), .A3(new_n26626_), .ZN(new_n26627_));
  NAND3_X1   g23417(.A1(new_n12794_), .A2(new_n13206_), .A3(new_n26625_), .ZN(new_n26628_));
  NAND3_X1   g23418(.A1(new_n26628_), .A2(new_n26627_), .A3(pi0038), .ZN(new_n26629_));
  XOR2_X1    g23419(.A1(new_n26629_), .A2(new_n4368_), .Z(new_n26630_));
  AOI21_X1   g23420(.A1(new_n26630_), .A2(pi0198), .B(new_n3290_), .ZN(new_n26631_));
  AOI21_X1   g23421(.A1(pi0634), .A2(new_n13246_), .B(new_n26435_), .ZN(new_n26632_));
  INV_X1     g23422(.I(new_n26632_), .ZN(new_n26633_));
  NOR2_X1    g23423(.A1(new_n26633_), .A2(new_n5386_), .ZN(new_n26634_));
  NOR3_X1    g23424(.A1(new_n13258_), .A2(new_n12862_), .A3(new_n26626_), .ZN(new_n26635_));
  NOR3_X1    g23425(.A1(new_n13246_), .A2(new_n12862_), .A3(new_n26625_), .ZN(new_n26636_));
  NOR2_X1    g23426(.A1(new_n26635_), .A2(new_n26636_), .ZN(new_n26637_));
  INV_X1     g23427(.I(new_n26637_), .ZN(new_n26638_));
  AOI21_X1   g23428(.A1(new_n26638_), .A2(new_n5386_), .B(new_n26634_), .ZN(new_n26639_));
  NAND2_X1   g23429(.A1(new_n13234_), .A2(new_n5383_), .ZN(new_n26640_));
  NAND2_X1   g23430(.A1(new_n26639_), .A2(new_n13234_), .ZN(new_n26641_));
  XOR2_X1    g23431(.A1(new_n26641_), .A2(new_n26640_), .Z(new_n26642_));
  AOI22_X1   g23432(.A1(new_n26642_), .A2(new_n26632_), .B1(new_n5378_), .B2(new_n26639_), .ZN(new_n26643_));
  NAND2_X1   g23433(.A1(new_n26433_), .A2(new_n5375_), .ZN(new_n26644_));
  NOR4_X1    g23434(.A1(new_n26643_), .A2(new_n3072_), .A3(new_n13334_), .A4(new_n26644_), .ZN(new_n26645_));
  NOR2_X1    g23435(.A1(new_n26632_), .A2(new_n5373_), .ZN(new_n26646_));
  AOI21_X1   g23436(.A1(new_n26637_), .A2(new_n5373_), .B(new_n26646_), .ZN(new_n26647_));
  NAND2_X1   g23437(.A1(new_n26647_), .A2(new_n13234_), .ZN(new_n26648_));
  XNOR2_X1   g23438(.A1(new_n26648_), .A2(new_n26640_), .ZN(new_n26649_));
  OAI21_X1   g23439(.A1(new_n26649_), .A2(new_n26637_), .B(new_n26644_), .ZN(new_n26650_));
  NAND3_X1   g23440(.A1(new_n26650_), .A2(new_n5378_), .A3(new_n26638_), .ZN(new_n26651_));
  NAND2_X1   g23441(.A1(new_n26651_), .A2(pi0215), .ZN(new_n26652_));
  XOR2_X1    g23442(.A1(new_n26652_), .A2(new_n13309_), .Z(new_n26653_));
  AOI21_X1   g23443(.A1(new_n26653_), .A2(new_n26645_), .B(pi0299), .ZN(new_n26654_));
  NOR4_X1    g23444(.A1(new_n12949_), .A2(new_n3072_), .A3(new_n5375_), .A4(new_n5796_), .ZN(new_n26655_));
  NOR3_X1    g23445(.A1(new_n26441_), .A2(pi0680), .A3(new_n5796_), .ZN(new_n26656_));
  NOR2_X1    g23446(.A1(new_n26656_), .A2(new_n26655_), .ZN(new_n26657_));
  NAND2_X1   g23447(.A1(new_n13242_), .A2(pi0634), .ZN(new_n26658_));
  OAI21_X1   g23448(.A1(new_n3072_), .A2(new_n12818_), .B(new_n26658_), .ZN(new_n26659_));
  INV_X1     g23449(.I(new_n26659_), .ZN(new_n26660_));
  AOI21_X1   g23450(.A1(new_n26660_), .A2(new_n5386_), .B(new_n26634_), .ZN(new_n26661_));
  NAND2_X1   g23451(.A1(new_n26661_), .A2(new_n13234_), .ZN(new_n26662_));
  XNOR2_X1   g23452(.A1(new_n26662_), .A2(new_n26640_), .ZN(new_n26663_));
  OAI22_X1   g23453(.A1(new_n26663_), .A2(new_n26633_), .B1(new_n26440_), .B2(new_n26657_), .ZN(new_n26664_));
  NOR2_X1    g23454(.A1(new_n26661_), .A2(new_n5636_), .ZN(new_n26665_));
  NAND2_X1   g23455(.A1(new_n26664_), .A2(new_n26665_), .ZN(new_n26666_));
  NAND2_X1   g23456(.A1(new_n26666_), .A2(new_n5454_), .ZN(new_n26667_));
  XOR2_X1    g23457(.A1(new_n26667_), .A2(new_n14371_), .Z(new_n26668_));
  INV_X1     g23458(.I(new_n26646_), .ZN(new_n26669_));
  OAI21_X1   g23459(.A1(new_n26660_), .A2(new_n5386_), .B(new_n26669_), .ZN(new_n26670_));
  NOR2_X1    g23460(.A1(new_n26670_), .A2(new_n13296_), .ZN(new_n26671_));
  XNOR2_X1   g23461(.A1(new_n26671_), .A2(new_n26640_), .ZN(new_n26672_));
  AOI22_X1   g23462(.A1(new_n26672_), .A2(new_n26660_), .B1(pi0198), .B2(new_n13671_), .ZN(new_n26673_));
  NOR3_X1    g23463(.A1(new_n26673_), .A2(new_n5636_), .A3(new_n26659_), .ZN(new_n26674_));
  NOR3_X1    g23464(.A1(new_n26435_), .A2(pi0634), .A3(pi0680), .ZN(new_n26675_));
  NOR2_X1    g23465(.A1(new_n26675_), .A2(new_n13258_), .ZN(new_n26676_));
  NAND2_X1   g23466(.A1(new_n26676_), .A2(new_n3312_), .ZN(new_n26677_));
  NAND4_X1   g23467(.A1(new_n26668_), .A2(new_n3111_), .A3(new_n26674_), .A4(new_n26677_), .ZN(new_n26678_));
  NOR2_X1    g23468(.A1(new_n26678_), .A2(new_n26654_), .ZN(new_n26679_));
  NAND2_X1   g23469(.A1(new_n26651_), .A2(pi0223), .ZN(new_n26680_));
  XOR2_X1    g23470(.A1(new_n26680_), .A2(new_n13466_), .Z(new_n26681_));
  NAND2_X1   g23471(.A1(new_n26681_), .A2(new_n26645_), .ZN(new_n26682_));
  NAND2_X1   g23472(.A1(new_n26682_), .A2(new_n3098_), .ZN(new_n26683_));
  NOR2_X1    g23473(.A1(new_n26679_), .A2(new_n26683_), .ZN(new_n26684_));
  NOR2_X1    g23474(.A1(new_n26624_), .A2(new_n5375_), .ZN(new_n26685_));
  NAND2_X1   g23475(.A1(new_n13141_), .A2(new_n3072_), .ZN(new_n26686_));
  OAI21_X1   g23476(.A1(new_n3072_), .A2(new_n13155_), .B(new_n26686_), .ZN(new_n26687_));
  NAND2_X1   g23477(.A1(new_n26687_), .A2(new_n26685_), .ZN(new_n26688_));
  INV_X1     g23478(.I(new_n26685_), .ZN(new_n26689_));
  OAI21_X1   g23479(.A1(new_n14336_), .A2(new_n3072_), .B(new_n26689_), .ZN(new_n26690_));
  NAND3_X1   g23480(.A1(new_n26688_), .A2(pi0299), .A3(new_n26690_), .ZN(new_n26691_));
  XOR2_X1    g23481(.A1(new_n26691_), .A2(new_n11324_), .Z(new_n26692_));
  AOI21_X1   g23482(.A1(new_n13125_), .A2(new_n3072_), .B(new_n26689_), .ZN(new_n26693_));
  NOR2_X1    g23483(.A1(new_n13120_), .A2(new_n13124_), .ZN(new_n26694_));
  NOR4_X1    g23484(.A1(new_n26694_), .A2(new_n26693_), .A3(new_n3072_), .A4(new_n26532_), .ZN(new_n26695_));
  AND3_X2    g23485(.A1(new_n26692_), .A2(pi0038), .A3(new_n26695_), .Z(new_n26696_));
  NAND2_X1   g23486(.A1(new_n26666_), .A2(new_n5398_), .ZN(new_n26697_));
  XOR2_X1    g23487(.A1(new_n26697_), .A2(new_n12982_), .Z(new_n26698_));
  NAND2_X1   g23488(.A1(new_n26698_), .A2(new_n26674_), .ZN(new_n26699_));
  NAND4_X1   g23489(.A1(new_n26676_), .A2(pi0198), .A3(new_n3091_), .A4(new_n3289_), .ZN(new_n26700_));
  AOI21_X1   g23490(.A1(new_n26699_), .A2(new_n3090_), .B(new_n26700_), .ZN(new_n26701_));
  OAI21_X1   g23491(.A1(new_n26696_), .A2(pi0039), .B(new_n26701_), .ZN(new_n26702_));
  NOR2_X1    g23492(.A1(new_n26702_), .A2(new_n26684_), .ZN(new_n26703_));
  XOR2_X1    g23493(.A1(new_n26703_), .A2(new_n26631_), .Z(new_n26704_));
  AND3_X2    g23494(.A1(new_n26704_), .A2(pi0625), .A3(pi1153), .Z(new_n26705_));
  NOR3_X1    g23495(.A1(new_n26704_), .A2(new_n13613_), .A3(new_n13615_), .ZN(new_n26706_));
  OAI21_X1   g23496(.A1(new_n26705_), .A2(new_n26706_), .B(new_n26460_), .ZN(new_n26707_));
  NAND2_X1   g23497(.A1(new_n26707_), .A2(pi0778), .ZN(new_n26708_));
  NOR2_X1    g23498(.A1(new_n26704_), .A2(new_n13614_), .ZN(new_n26709_));
  XOR2_X1    g23499(.A1(new_n26709_), .A2(new_n13615_), .Z(new_n26710_));
  NAND4_X1   g23500(.A1(new_n26710_), .A2(pi0778), .A3(new_n26460_), .A4(new_n26704_), .ZN(new_n26711_));
  INV_X1     g23501(.I(new_n26711_), .ZN(new_n26712_));
  NAND2_X1   g23502(.A1(new_n26712_), .A2(new_n26708_), .ZN(new_n26713_));
  NAND3_X1   g23503(.A1(new_n26711_), .A2(pi0778), .A3(new_n26707_), .ZN(new_n26714_));
  NAND3_X1   g23504(.A1(new_n26713_), .A2(new_n13805_), .A3(new_n26714_), .ZN(new_n26715_));
  NAND3_X1   g23505(.A1(new_n26715_), .A2(new_n13880_), .A3(new_n26623_), .ZN(new_n26716_));
  NAND2_X1   g23506(.A1(new_n26716_), .A2(new_n26621_), .ZN(new_n26717_));
  NAND3_X1   g23507(.A1(new_n26717_), .A2(new_n15395_), .A3(new_n26460_), .ZN(new_n26718_));
  INV_X1     g23508(.I(new_n26717_), .ZN(new_n26719_));
  NAND3_X1   g23509(.A1(new_n26719_), .A2(new_n15395_), .A3(new_n26457_), .ZN(new_n26720_));
  NAND2_X1   g23510(.A1(new_n26720_), .A2(new_n26718_), .ZN(new_n26721_));
  NAND3_X1   g23511(.A1(new_n26721_), .A2(pi0628), .A3(pi1156), .ZN(new_n26722_));
  NAND4_X1   g23512(.A1(new_n26720_), .A2(pi0628), .A3(new_n13969_), .A4(new_n26718_), .ZN(new_n26723_));
  AOI21_X1   g23513(.A1(new_n26722_), .A2(new_n26723_), .B(new_n26457_), .ZN(new_n26724_));
  NOR2_X1    g23514(.A1(new_n26460_), .A2(pi0628), .ZN(new_n26725_));
  AOI21_X1   g23515(.A1(new_n26721_), .A2(pi0628), .B(new_n26725_), .ZN(new_n26726_));
  OAI21_X1   g23516(.A1(new_n26726_), .A2(new_n13969_), .B(pi0792), .ZN(new_n26727_));
  OAI22_X1   g23517(.A1(new_n26727_), .A2(new_n26724_), .B1(pi0792), .B2(new_n26721_), .ZN(new_n26728_));
  AOI21_X1   g23518(.A1(new_n26728_), .A2(pi0647), .B(new_n26619_), .ZN(new_n26729_));
  AOI21_X1   g23519(.A1(new_n26729_), .A2(new_n14206_), .B(pi0787), .ZN(new_n26730_));
  NAND3_X1   g23520(.A1(new_n26728_), .A2(pi0647), .A3(pi1157), .ZN(new_n26731_));
  INV_X1     g23521(.I(new_n26728_), .ZN(new_n26732_));
  NAND3_X1   g23522(.A1(new_n26732_), .A2(pi0647), .A3(new_n14006_), .ZN(new_n26733_));
  AOI21_X1   g23523(.A1(new_n26733_), .A2(new_n26731_), .B(new_n26457_), .ZN(new_n26734_));
  NAND2_X1   g23524(.A1(new_n26734_), .A2(pi0630), .ZN(new_n26735_));
  AOI21_X1   g23525(.A1(new_n26618_), .A2(new_n26730_), .B(new_n26735_), .ZN(new_n26736_));
  NOR2_X1    g23526(.A1(new_n26553_), .A2(new_n26554_), .ZN(new_n26737_));
  INV_X1     g23527(.I(new_n26737_), .ZN(new_n26738_));
  NOR3_X1    g23528(.A1(new_n26468_), .A2(pi0634), .A3(new_n13213_), .ZN(new_n26739_));
  OAI21_X1   g23529(.A1(new_n26739_), .A2(new_n14291_), .B(pi0038), .ZN(new_n26740_));
  XOR2_X1    g23530(.A1(new_n26740_), .A2(new_n4368_), .Z(new_n26741_));
  AOI21_X1   g23531(.A1(new_n26741_), .A2(pi0198), .B(new_n3290_), .ZN(new_n26742_));
  NOR2_X1    g23532(.A1(new_n26506_), .A2(new_n13388_), .ZN(new_n26743_));
  INV_X1     g23533(.I(new_n26647_), .ZN(new_n26744_));
  NOR2_X1    g23534(.A1(new_n26480_), .A2(new_n5386_), .ZN(new_n26745_));
  NOR2_X1    g23535(.A1(new_n13316_), .A2(pi0634), .ZN(new_n26746_));
  AOI21_X1   g23536(.A1(new_n26746_), .A2(new_n26479_), .B(new_n13124_), .ZN(new_n26747_));
  NOR2_X1    g23537(.A1(new_n26747_), .A2(new_n5794_), .ZN(new_n26748_));
  AOI22_X1   g23538(.A1(new_n26748_), .A2(new_n13365_), .B1(new_n26486_), .B2(new_n26745_), .ZN(new_n26749_));
  AOI21_X1   g23539(.A1(new_n26749_), .A2(new_n26744_), .B(new_n13282_), .ZN(new_n26750_));
  INV_X1     g23540(.I(new_n26503_), .ZN(new_n26751_));
  NOR3_X1    g23541(.A1(new_n26751_), .A2(new_n26624_), .A3(new_n26502_), .ZN(new_n26754_));
  AOI21_X1   g23542(.A1(new_n26749_), .A2(new_n26754_), .B(pi0603), .ZN(new_n26755_));
  NOR3_X1    g23543(.A1(new_n26750_), .A2(new_n26755_), .A3(new_n13365_), .ZN(new_n26756_));
  NOR2_X1    g23544(.A1(new_n26754_), .A2(new_n5636_), .ZN(new_n26757_));
  NAND2_X1   g23545(.A1(new_n5378_), .A2(pi0603), .ZN(new_n26758_));
  XOR2_X1    g23546(.A1(new_n26757_), .A2(new_n26758_), .Z(new_n26759_));
  OAI22_X1   g23547(.A1(new_n26756_), .A2(new_n13296_), .B1(new_n26637_), .B2(new_n26759_), .ZN(new_n26760_));
  NAND3_X1   g23548(.A1(new_n26760_), .A2(pi0680), .A3(new_n26743_), .ZN(new_n26761_));
  INV_X1     g23549(.I(new_n26761_), .ZN(new_n26762_));
  NOR2_X1    g23550(.A1(new_n26754_), .A2(new_n5794_), .ZN(new_n26763_));
  XOR2_X1    g23551(.A1(new_n26763_), .A2(new_n13282_), .Z(new_n26764_));
  NAND2_X1   g23552(.A1(new_n26764_), .A2(new_n26747_), .ZN(new_n26765_));
  NOR2_X1    g23553(.A1(new_n26765_), .A2(new_n5636_), .ZN(new_n26766_));
  NOR2_X1    g23554(.A1(new_n26766_), .A2(pi0603), .ZN(new_n26767_));
  NOR2_X1    g23555(.A1(new_n26632_), .A2(pi0603), .ZN(new_n26768_));
  NOR2_X1    g23556(.A1(new_n26748_), .A2(new_n26768_), .ZN(new_n26769_));
  AOI21_X1   g23557(.A1(new_n26769_), .A2(new_n13365_), .B(new_n13296_), .ZN(new_n26770_));
  NOR3_X1    g23558(.A1(new_n26770_), .A2(new_n13336_), .A3(new_n26768_), .ZN(new_n26771_));
  OAI22_X1   g23559(.A1(new_n26767_), .A2(new_n26639_), .B1(new_n26765_), .B2(new_n26771_), .ZN(new_n26772_));
  NAND3_X1   g23560(.A1(new_n26772_), .A2(pi0680), .A3(new_n26516_), .ZN(new_n26773_));
  NAND2_X1   g23561(.A1(new_n26773_), .A2(pi0223), .ZN(new_n26774_));
  XOR2_X1    g23562(.A1(new_n26774_), .A2(new_n13466_), .Z(new_n26775_));
  NOR3_X1    g23563(.A1(new_n26474_), .A2(new_n5794_), .A3(new_n5636_), .ZN(new_n26776_));
  OAI21_X1   g23564(.A1(new_n26776_), .A2(new_n13203_), .B(new_n26660_), .ZN(new_n26777_));
  OAI21_X1   g23565(.A1(new_n26624_), .A2(new_n13233_), .B(new_n26474_), .ZN(new_n26778_));
  NAND2_X1   g23566(.A1(new_n26778_), .A2(new_n5386_), .ZN(new_n26779_));
  AOI22_X1   g23567(.A1(new_n26779_), .A2(new_n5383_), .B1(new_n5373_), .B2(new_n26749_), .ZN(new_n26780_));
  NOR2_X1    g23568(.A1(new_n26780_), .A2(new_n13296_), .ZN(new_n26781_));
  OAI21_X1   g23569(.A1(new_n26781_), .A2(new_n26670_), .B(pi0603), .ZN(new_n26782_));
  NAND2_X1   g23570(.A1(new_n26483_), .A2(pi0680), .ZN(new_n26783_));
  AOI21_X1   g23571(.A1(new_n26782_), .A2(new_n26777_), .B(new_n26783_), .ZN(new_n26784_));
  INV_X1     g23572(.I(new_n26747_), .ZN(new_n26785_));
  NAND2_X1   g23573(.A1(new_n26778_), .A2(pi0603), .ZN(new_n26786_));
  XOR2_X1    g23574(.A1(new_n26786_), .A2(new_n13282_), .Z(new_n26787_));
  OAI21_X1   g23575(.A1(new_n26787_), .A2(new_n26785_), .B(new_n12845_), .ZN(new_n26788_));
  NOR2_X1    g23576(.A1(new_n26661_), .A2(new_n5794_), .ZN(new_n26789_));
  AOI21_X1   g23577(.A1(new_n26788_), .A2(new_n26789_), .B(new_n5375_), .ZN(new_n26790_));
  NOR4_X1    g23578(.A1(new_n26747_), .A2(new_n26768_), .A3(new_n5794_), .A4(new_n5379_), .ZN(new_n26791_));
  NOR2_X1    g23579(.A1(new_n26791_), .A2(new_n5382_), .ZN(new_n26792_));
  NOR2_X1    g23580(.A1(new_n12845_), .A2(new_n5382_), .ZN(new_n26793_));
  XOR2_X1    g23581(.A1(new_n26792_), .A2(new_n26793_), .Z(new_n26794_));
  NAND4_X1   g23582(.A1(new_n26492_), .A2(pi0680), .A3(new_n26769_), .A4(new_n26794_), .ZN(new_n26795_));
  XOR2_X1    g23583(.A1(new_n26790_), .A2(new_n26795_), .Z(new_n26796_));
  NAND2_X1   g23584(.A1(new_n26796_), .A2(new_n5454_), .ZN(new_n26797_));
  XOR2_X1    g23585(.A1(new_n26797_), .A2(new_n14371_), .Z(new_n26798_));
  AOI21_X1   g23586(.A1(new_n26798_), .A2(new_n26784_), .B(pi0215), .ZN(new_n26799_));
  NAND3_X1   g23587(.A1(new_n26499_), .A2(new_n26624_), .A3(new_n13324_), .ZN(new_n26800_));
  NAND3_X1   g23588(.A1(new_n26800_), .A2(new_n13258_), .A3(new_n26440_), .ZN(new_n26801_));
  NOR3_X1    g23589(.A1(new_n26799_), .A2(new_n3313_), .A3(new_n26801_), .ZN(new_n26802_));
  NOR2_X1    g23590(.A1(new_n26802_), .A2(new_n5827_), .ZN(new_n26803_));
  NAND2_X1   g23591(.A1(new_n26773_), .A2(pi0215), .ZN(new_n26804_));
  XOR2_X1    g23592(.A1(new_n26804_), .A2(new_n5456_), .Z(new_n26805_));
  NOR4_X1    g23593(.A1(new_n26803_), .A2(new_n3098_), .A3(new_n26761_), .A4(new_n26805_), .ZN(new_n26806_));
  AOI21_X1   g23594(.A1(new_n26762_), .A2(new_n26775_), .B(new_n26806_), .ZN(new_n26807_));
  NAND2_X1   g23595(.A1(new_n26796_), .A2(new_n5398_), .ZN(new_n26808_));
  XOR2_X1    g23596(.A1(new_n26808_), .A2(new_n12982_), .Z(new_n26809_));
  AND2_X2    g23597(.A1(new_n26809_), .A2(new_n26784_), .Z(new_n26810_));
  NOR3_X1    g23598(.A1(new_n26801_), .A2(new_n3259_), .A3(new_n3092_), .ZN(new_n26811_));
  OAI21_X1   g23599(.A1(new_n26810_), .A2(pi0223), .B(new_n26811_), .ZN(new_n26812_));
  OAI21_X1   g23600(.A1(new_n26807_), .A2(new_n26812_), .B(new_n3183_), .ZN(new_n26813_));
  OAI21_X1   g23601(.A1(new_n13176_), .A2(new_n13168_), .B(pi0634), .ZN(new_n26814_));
  NOR2_X1    g23602(.A1(new_n26694_), .A2(new_n26626_), .ZN(new_n26815_));
  NAND2_X1   g23603(.A1(new_n26815_), .A2(new_n26532_), .ZN(new_n26816_));
  XNOR2_X1   g23604(.A1(new_n26816_), .A2(new_n26814_), .ZN(new_n26817_));
  NAND2_X1   g23605(.A1(new_n26537_), .A2(new_n5794_), .ZN(new_n26818_));
  NAND2_X1   g23606(.A1(new_n26624_), .A2(new_n13124_), .ZN(new_n26819_));
  NAND4_X1   g23607(.A1(new_n13121_), .A2(pi0680), .A3(new_n26464_), .A4(new_n26819_), .ZN(new_n26820_));
  AOI21_X1   g23608(.A1(new_n26695_), .A2(new_n5794_), .B(new_n26820_), .ZN(new_n26821_));
  AOI21_X1   g23609(.A1(new_n26818_), .A2(new_n26821_), .B(pi0633), .ZN(new_n26822_));
  OAI21_X1   g23610(.A1(new_n26822_), .A2(new_n26817_), .B(new_n3098_), .ZN(new_n26823_));
  OR2_X2     g23611(.A1(new_n26529_), .A2(new_n26685_), .Z(new_n26824_));
  NOR3_X1    g23612(.A1(new_n26539_), .A2(new_n3098_), .A3(new_n5375_), .ZN(new_n26825_));
  NAND3_X1   g23613(.A1(new_n26824_), .A2(new_n26823_), .A3(new_n26825_), .ZN(new_n26826_));
  NAND2_X1   g23614(.A1(new_n26826_), .A2(new_n26689_), .ZN(new_n26827_));
  NAND2_X1   g23615(.A1(new_n13141_), .A2(pi0633), .ZN(new_n26828_));
  XOR2_X1    g23616(.A1(new_n26828_), .A2(new_n26464_), .Z(new_n26829_));
  OR3_X2     g23617(.A1(new_n26829_), .A2(new_n13124_), .A3(new_n26524_), .Z(new_n26830_));
  NAND2_X1   g23618(.A1(new_n26830_), .A2(pi0603), .ZN(new_n26831_));
  NAND2_X1   g23619(.A1(new_n13155_), .A2(new_n3072_), .ZN(new_n26833_));
  NAND3_X1   g23620(.A1(new_n26687_), .A2(new_n13192_), .A3(new_n26833_), .ZN(new_n26834_));
  XOR2_X1    g23621(.A1(new_n26831_), .A2(new_n26834_), .Z(new_n26835_));
  NAND4_X1   g23622(.A1(new_n26813_), .A2(new_n26549_), .A3(new_n26827_), .A4(new_n26835_), .ZN(new_n26836_));
  XOR2_X1    g23623(.A1(new_n26836_), .A2(new_n26742_), .Z(new_n26837_));
  NAND2_X1   g23624(.A1(new_n26837_), .A2(pi0625), .ZN(new_n26838_));
  XOR2_X1    g23625(.A1(new_n26838_), .A2(new_n13620_), .Z(new_n26839_));
  NAND2_X1   g23626(.A1(new_n26710_), .A2(new_n26460_), .ZN(new_n26840_));
  NAND2_X1   g23627(.A1(new_n26840_), .A2(new_n14081_), .ZN(new_n26841_));
  AOI21_X1   g23628(.A1(new_n26839_), .A2(new_n26738_), .B(new_n26841_), .ZN(new_n26842_));
  NAND2_X1   g23629(.A1(new_n26707_), .A2(new_n14081_), .ZN(new_n26843_));
  NAND2_X1   g23630(.A1(new_n26837_), .A2(pi1153), .ZN(new_n26844_));
  XOR2_X1    g23631(.A1(new_n26844_), .A2(new_n13615_), .Z(new_n26845_));
  NOR3_X1    g23632(.A1(new_n26845_), .A2(new_n13748_), .A3(new_n26737_), .ZN(new_n26846_));
  OAI21_X1   g23633(.A1(new_n26842_), .A2(new_n26843_), .B(new_n26846_), .ZN(new_n26847_));
  NAND2_X1   g23634(.A1(new_n26837_), .A2(new_n13748_), .ZN(new_n26848_));
  NAND2_X1   g23635(.A1(new_n26847_), .A2(new_n26848_), .ZN(new_n26849_));
  AND2_X2    g23636(.A1(new_n26713_), .A2(new_n26714_), .Z(new_n26850_));
  NOR2_X1    g23637(.A1(new_n13783_), .A2(new_n13778_), .ZN(new_n26851_));
  AOI21_X1   g23638(.A1(new_n26850_), .A2(new_n26851_), .B(pi0609), .ZN(new_n26852_));
  INV_X1     g23639(.I(new_n26852_), .ZN(new_n26853_));
  AOI21_X1   g23640(.A1(new_n26849_), .A2(new_n26853_), .B(new_n13801_), .ZN(new_n26854_));
  AOI21_X1   g23641(.A1(new_n13783_), .A2(new_n13778_), .B(pi0609), .ZN(new_n26855_));
  NOR2_X1    g23642(.A1(new_n26855_), .A2(new_n13801_), .ZN(new_n26856_));
  NAND2_X1   g23643(.A1(new_n26849_), .A2(new_n26856_), .ZN(new_n26857_));
  NOR2_X1    g23644(.A1(new_n26854_), .A2(new_n26857_), .ZN(new_n26858_));
  INV_X1     g23645(.I(new_n26858_), .ZN(new_n26859_));
  NAND2_X1   g23646(.A1(new_n26854_), .A2(new_n26857_), .ZN(new_n26860_));
  AOI21_X1   g23647(.A1(new_n26850_), .A2(new_n13805_), .B(new_n26622_), .ZN(new_n26861_));
  NAND2_X1   g23648(.A1(new_n26861_), .A2(new_n13816_), .ZN(new_n26862_));
  NAND2_X1   g23649(.A1(new_n26862_), .A2(new_n13824_), .ZN(new_n26863_));
  OAI21_X1   g23650(.A1(new_n26863_), .A2(new_n26583_), .B(new_n13816_), .ZN(new_n26864_));
  INV_X1     g23651(.I(new_n26864_), .ZN(new_n26865_));
  AOI21_X1   g23652(.A1(new_n26859_), .A2(new_n26860_), .B(new_n26865_), .ZN(new_n26866_));
  AOI21_X1   g23653(.A1(new_n26598_), .A2(new_n13836_), .B(pi0618), .ZN(new_n26867_));
  NOR2_X1    g23654(.A1(new_n26867_), .A2(new_n13855_), .ZN(new_n26868_));
  INV_X1     g23655(.I(new_n26868_), .ZN(new_n26869_));
  AOI21_X1   g23656(.A1(new_n26859_), .A2(new_n26860_), .B(new_n26869_), .ZN(new_n26870_));
  OAI21_X1   g23657(.A1(new_n13855_), .A2(new_n26866_), .B(new_n26870_), .ZN(new_n26871_));
  INV_X1     g23658(.I(new_n26860_), .ZN(new_n26872_));
  OAI21_X1   g23659(.A1(new_n26872_), .A2(new_n26858_), .B(new_n26864_), .ZN(new_n26873_));
  OAI21_X1   g23660(.A1(new_n26872_), .A2(new_n26858_), .B(new_n26868_), .ZN(new_n26874_));
  NAND3_X1   g23661(.A1(new_n26873_), .A2(new_n26874_), .A3(pi0781), .ZN(new_n26875_));
  NAND2_X1   g23662(.A1(new_n26871_), .A2(new_n26875_), .ZN(new_n26876_));
  AOI21_X1   g23663(.A1(new_n26876_), .A2(new_n13896_), .B(new_n15479_), .ZN(new_n26877_));
  AOI21_X1   g23664(.A1(pi0781), .A2(new_n26873_), .B(new_n26874_), .ZN(new_n26878_));
  NOR3_X1    g23665(.A1(new_n26866_), .A2(new_n26870_), .A3(new_n13855_), .ZN(new_n26879_));
  NOR2_X1    g23666(.A1(new_n26878_), .A2(new_n26879_), .ZN(new_n26880_));
  AOI21_X1   g23667(.A1(new_n26603_), .A2(pi1159), .B(new_n13904_), .ZN(new_n26881_));
  INV_X1     g23668(.I(new_n26607_), .ZN(new_n26882_));
  OAI21_X1   g23669(.A1(new_n26881_), .A2(new_n26882_), .B(new_n26460_), .ZN(new_n26883_));
  AOI21_X1   g23670(.A1(new_n26883_), .A2(new_n13892_), .B(pi0619), .ZN(new_n26884_));
  OAI21_X1   g23671(.A1(new_n26880_), .A2(new_n26884_), .B(new_n13896_), .ZN(new_n26885_));
  AOI21_X1   g23672(.A1(new_n26717_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n26886_));
  AOI21_X1   g23673(.A1(new_n26612_), .A2(new_n26886_), .B(pi0619), .ZN(new_n26887_));
  NOR3_X1    g23674(.A1(new_n26880_), .A2(new_n12777_), .A3(new_n26887_), .ZN(new_n26888_));
  OAI21_X1   g23675(.A1(new_n26877_), .A2(new_n26885_), .B(new_n26888_), .ZN(new_n26889_));
  NOR4_X1    g23676(.A1(new_n26612_), .A2(new_n26883_), .A3(new_n13896_), .A4(new_n26603_), .ZN(new_n26890_));
  NAND2_X1   g23677(.A1(new_n26612_), .A2(pi0789), .ZN(new_n26891_));
  NOR3_X1    g23678(.A1(new_n26883_), .A2(new_n13896_), .A3(new_n26603_), .ZN(new_n26892_));
  NOR2_X1    g23679(.A1(new_n26892_), .A2(new_n26891_), .ZN(new_n26893_));
  NOR2_X1    g23680(.A1(new_n26893_), .A2(new_n26890_), .ZN(new_n26894_));
  AOI21_X1   g23681(.A1(new_n26894_), .A2(new_n13963_), .B(new_n19028_), .ZN(new_n26895_));
  NAND2_X1   g23682(.A1(new_n26615_), .A2(new_n26609_), .ZN(new_n26896_));
  NOR3_X1    g23683(.A1(new_n26896_), .A2(pi0626), .A3(new_n19208_), .ZN(new_n26897_));
  OAI21_X1   g23684(.A1(new_n26895_), .A2(new_n26897_), .B(new_n26460_), .ZN(new_n26898_));
  NOR2_X1    g23685(.A1(new_n26717_), .A2(new_n14162_), .ZN(new_n26899_));
  XOR2_X1    g23686(.A1(new_n26899_), .A2(new_n16828_), .Z(new_n26900_));
  AOI21_X1   g23687(.A1(new_n26900_), .A2(new_n26460_), .B(pi0788), .ZN(new_n26901_));
  NAND2_X1   g23688(.A1(new_n26898_), .A2(new_n26901_), .ZN(new_n26902_));
  AOI21_X1   g23689(.A1(new_n26894_), .A2(new_n13962_), .B(new_n18976_), .ZN(new_n26903_));
  NOR3_X1    g23690(.A1(new_n26896_), .A2(new_n18974_), .A3(new_n18975_), .ZN(new_n26904_));
  NOR2_X1    g23691(.A1(new_n26903_), .A2(new_n26904_), .ZN(new_n26905_));
  OR2_X2     g23692(.A1(new_n26726_), .A2(new_n19489_), .Z(new_n26906_));
  NAND2_X1   g23693(.A1(new_n26724_), .A2(pi0629), .ZN(new_n26907_));
  AOI21_X1   g23694(.A1(new_n26907_), .A2(new_n26906_), .B(new_n16875_), .ZN(new_n26908_));
  NAND4_X1   g23695(.A1(new_n26894_), .A2(new_n16372_), .A3(new_n26460_), .A4(new_n26908_), .ZN(new_n26909_));
  NOR2_X1    g23696(.A1(new_n26905_), .A2(new_n26909_), .ZN(new_n26910_));
  NAND2_X1   g23697(.A1(new_n26616_), .A2(new_n26462_), .ZN(new_n26911_));
  NAND2_X1   g23698(.A1(new_n26911_), .A2(new_n26908_), .ZN(new_n26912_));
  OAI21_X1   g23699(.A1(new_n26912_), .A2(new_n16424_), .B(new_n16419_), .ZN(new_n26913_));
  AOI21_X1   g23700(.A1(new_n26902_), .A2(new_n26910_), .B(new_n26913_), .ZN(new_n26914_));
  AOI21_X1   g23701(.A1(new_n26914_), .A2(new_n26889_), .B(new_n26736_), .ZN(new_n26915_));
  AOI21_X1   g23702(.A1(new_n26894_), .A2(new_n16372_), .B(new_n26461_), .ZN(new_n26916_));
  AOI21_X1   g23703(.A1(new_n26916_), .A2(new_n13994_), .B(new_n26458_), .ZN(new_n26917_));
  NOR2_X1    g23704(.A1(new_n26460_), .A2(new_n14211_), .ZN(new_n26918_));
  AOI21_X1   g23705(.A1(new_n26917_), .A2(new_n14211_), .B(new_n26918_), .ZN(new_n26919_));
  AOI21_X1   g23706(.A1(new_n26919_), .A2(pi0715), .B(new_n14217_), .ZN(new_n26920_));
  INV_X1     g23707(.I(new_n26918_), .ZN(new_n26921_));
  NAND3_X1   g23708(.A1(new_n26617_), .A2(new_n14211_), .A3(new_n26459_), .ZN(new_n26922_));
  AND4_X2    g23709(.A1(new_n14204_), .A2(new_n26922_), .A3(pi0715), .A4(new_n26921_), .Z(new_n26923_));
  OAI21_X1   g23710(.A1(new_n26920_), .A2(new_n26923_), .B(new_n26460_), .ZN(new_n26924_));
  NAND2_X1   g23711(.A1(new_n26729_), .A2(pi1157), .ZN(new_n26925_));
  NAND2_X1   g23712(.A1(new_n26925_), .A2(pi0787), .ZN(new_n26926_));
  OAI22_X1   g23713(.A1(new_n26926_), .A2(new_n26734_), .B1(pi0787), .B2(new_n26732_), .ZN(new_n26927_));
  AOI21_X1   g23714(.A1(new_n26927_), .A2(pi0644), .B(new_n15386_), .ZN(new_n26928_));
  AOI21_X1   g23715(.A1(new_n26924_), .A2(new_n26928_), .B(new_n26915_), .ZN(new_n26929_));
  OAI21_X1   g23716(.A1(new_n26929_), .A2(new_n14204_), .B(pi0790), .ZN(new_n26930_));
  NAND3_X1   g23717(.A1(new_n26922_), .A2(pi0644), .A3(new_n26921_), .ZN(new_n26931_));
  XOR2_X1    g23718(.A1(new_n26931_), .A2(new_n14205_), .Z(new_n26932_));
  AOI21_X1   g23719(.A1(new_n26927_), .A2(new_n14204_), .B(new_n19370_), .ZN(new_n26933_));
  OAI21_X1   g23720(.A1(new_n26932_), .A2(new_n26457_), .B(new_n26933_), .ZN(new_n26934_));
  NAND2_X1   g23721(.A1(new_n26915_), .A2(pi0790), .ZN(new_n26935_));
  AOI21_X1   g23722(.A1(new_n26934_), .A2(new_n14204_), .B(new_n26935_), .ZN(new_n26936_));
  AND2_X2    g23723(.A1(new_n26618_), .A2(new_n26730_), .Z(new_n26937_));
  OAI21_X1   g23724(.A1(new_n26880_), .A2(pi0789), .B(new_n14143_), .ZN(new_n26938_));
  INV_X1     g23725(.I(new_n26884_), .ZN(new_n26939_));
  AOI21_X1   g23726(.A1(new_n26876_), .A2(new_n26939_), .B(pi0789), .ZN(new_n26940_));
  NOR2_X1    g23727(.A1(new_n26887_), .A2(new_n12777_), .ZN(new_n26941_));
  NAND2_X1   g23728(.A1(new_n26876_), .A2(new_n26941_), .ZN(new_n26942_));
  AOI21_X1   g23729(.A1(new_n26938_), .A2(new_n26940_), .B(new_n26942_), .ZN(new_n26943_));
  NAND3_X1   g23730(.A1(new_n26896_), .A2(pi0626), .A3(new_n13963_), .ZN(new_n26944_));
  NAND3_X1   g23731(.A1(new_n26894_), .A2(new_n13901_), .A3(new_n13963_), .ZN(new_n26945_));
  NAND2_X1   g23732(.A1(new_n26945_), .A2(new_n26944_), .ZN(new_n26946_));
  INV_X1     g23733(.I(new_n26901_), .ZN(new_n26947_));
  AOI21_X1   g23734(.A1(new_n26946_), .A2(new_n26460_), .B(new_n26947_), .ZN(new_n26948_));
  INV_X1     g23735(.I(new_n26908_), .ZN(new_n26949_));
  NOR4_X1    g23736(.A1(new_n26949_), .A2(new_n26896_), .A3(new_n14142_), .A4(new_n26457_), .ZN(new_n26950_));
  OAI21_X1   g23737(.A1(new_n26904_), .A2(new_n26903_), .B(new_n26950_), .ZN(new_n26951_));
  AOI21_X1   g23738(.A1(new_n26462_), .A2(new_n26616_), .B(new_n26949_), .ZN(new_n26952_));
  AOI21_X1   g23739(.A1(new_n26952_), .A2(new_n16423_), .B(new_n16574_), .ZN(new_n26953_));
  OAI21_X1   g23740(.A1(new_n26948_), .A2(new_n26951_), .B(new_n26953_), .ZN(new_n26954_));
  OAI22_X1   g23741(.A1(new_n26954_), .A2(new_n26943_), .B1(new_n26937_), .B2(new_n26735_), .ZN(new_n26955_));
  NOR3_X1    g23742(.A1(new_n26955_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n26958_));
  NOR2_X1    g23743(.A1(new_n26958_), .A2(po1038), .ZN(new_n26959_));
  OAI21_X1   g23744(.A1(new_n26930_), .A2(new_n26936_), .B(new_n26959_), .ZN(new_n26960_));
  NAND2_X1   g23745(.A1(new_n26960_), .A2(new_n12658_), .ZN(po0355));
  NOR2_X1    g23746(.A1(new_n7240_), .A2(new_n8549_), .ZN(new_n26962_));
  INV_X1     g23747(.I(new_n26962_), .ZN(new_n26963_));
  INV_X1     g23748(.I(pi0617), .ZN(new_n26964_));
  NAND3_X1   g23749(.A1(new_n19325_), .A2(new_n19326_), .A3(pi0199), .ZN(new_n26965_));
  NOR2_X1    g23750(.A1(new_n3259_), .A2(new_n8549_), .ZN(new_n26966_));
  NAND2_X1   g23751(.A1(new_n26965_), .A2(new_n26966_), .ZN(new_n26967_));
  NAND3_X1   g23752(.A1(new_n14362_), .A2(new_n3259_), .A3(pi0199), .ZN(new_n26968_));
  OAI21_X1   g23753(.A1(new_n15561_), .A2(new_n15559_), .B(new_n15555_), .ZN(new_n26969_));
  AOI21_X1   g23754(.A1(new_n26967_), .A2(new_n26968_), .B(new_n26969_), .ZN(new_n26970_));
  OAI21_X1   g23755(.A1(new_n26970_), .A2(pi0199), .B(new_n19321_), .ZN(new_n26971_));
  NOR3_X1    g23756(.A1(new_n26971_), .A2(new_n26964_), .A3(new_n3290_), .ZN(new_n26972_));
  NOR3_X1    g23757(.A1(new_n14362_), .A2(new_n3259_), .A3(new_n8549_), .ZN(new_n26973_));
  NOR2_X1    g23758(.A1(new_n26965_), .A2(new_n26966_), .ZN(new_n26974_));
  AOI21_X1   g23759(.A1(new_n16113_), .A2(new_n16112_), .B(new_n19328_), .ZN(new_n26975_));
  OAI21_X1   g23760(.A1(new_n26973_), .A2(new_n26974_), .B(new_n26975_), .ZN(new_n26976_));
  AOI21_X1   g23761(.A1(new_n26976_), .A2(new_n8549_), .B(new_n19641_), .ZN(new_n26977_));
  NOR3_X1    g23762(.A1(new_n26977_), .A2(new_n26964_), .A3(new_n3289_), .ZN(new_n26978_));
  NOR2_X1    g23763(.A1(new_n8549_), .A2(new_n26964_), .ZN(new_n26979_));
  OAI21_X1   g23764(.A1(new_n26972_), .A2(new_n26978_), .B(new_n26979_), .ZN(new_n26980_));
  AOI21_X1   g23765(.A1(new_n26980_), .A2(new_n8549_), .B(new_n13627_), .ZN(new_n26981_));
  NOR2_X1    g23766(.A1(new_n26981_), .A2(new_n13613_), .ZN(new_n26982_));
  INV_X1     g23767(.I(pi0637), .ZN(new_n26983_));
  NOR2_X1    g23768(.A1(new_n13613_), .A2(new_n26983_), .ZN(new_n26984_));
  XOR2_X1    g23769(.A1(new_n26982_), .A2(new_n26984_), .Z(new_n26985_));
  NOR2_X1    g23770(.A1(new_n3183_), .A2(new_n8549_), .ZN(new_n26986_));
  XOR2_X1    g23771(.A1(new_n13717_), .A2(new_n26986_), .Z(new_n26987_));
  NOR2_X1    g23772(.A1(new_n16149_), .A2(new_n8549_), .ZN(new_n26988_));
  NOR2_X1    g23773(.A1(new_n26988_), .A2(pi0038), .ZN(new_n26989_));
  OAI21_X1   g23774(.A1(new_n26987_), .A2(new_n13686_), .B(new_n26989_), .ZN(new_n26990_));
  INV_X1     g23775(.I(new_n13197_), .ZN(new_n26991_));
  NAND3_X1   g23776(.A1(new_n13165_), .A2(pi0039), .A3(pi0199), .ZN(new_n26992_));
  OR3_X2     g23777(.A1(new_n13165_), .A2(new_n8549_), .A3(new_n26986_), .Z(new_n26993_));
  AOI21_X1   g23778(.A1(new_n26993_), .A2(new_n26992_), .B(new_n26991_), .ZN(new_n26994_));
  AOI21_X1   g23779(.A1(new_n26990_), .A2(new_n26994_), .B(new_n26983_), .ZN(new_n26995_));
  NAND2_X1   g23780(.A1(new_n3289_), .A2(pi0637), .ZN(new_n26996_));
  XOR2_X1    g23781(.A1(new_n26995_), .A2(new_n26996_), .Z(new_n26997_));
  NOR2_X1    g23782(.A1(new_n26997_), .A2(new_n8549_), .ZN(new_n26998_));
  NOR2_X1    g23783(.A1(new_n14428_), .A2(new_n8549_), .ZN(new_n26999_));
  OAI21_X1   g23784(.A1(pi0199), .A2(pi1153), .B(pi0625), .ZN(new_n27000_));
  OAI22_X1   g23785(.A1(new_n26999_), .A2(pi0637), .B1(new_n13627_), .B2(new_n27000_), .ZN(new_n27001_));
  NAND2_X1   g23786(.A1(new_n26998_), .A2(new_n27001_), .ZN(new_n27002_));
  NAND2_X1   g23787(.A1(new_n27002_), .A2(new_n14081_), .ZN(new_n27003_));
  NAND3_X1   g23788(.A1(new_n26977_), .A2(pi0617), .A3(new_n3289_), .ZN(new_n27004_));
  NAND3_X1   g23789(.A1(new_n26971_), .A2(pi0617), .A3(new_n3290_), .ZN(new_n27005_));
  INV_X1     g23790(.I(new_n26979_), .ZN(new_n27006_));
  AOI21_X1   g23791(.A1(new_n27005_), .A2(new_n27004_), .B(new_n27006_), .ZN(new_n27007_));
  OAI21_X1   g23792(.A1(new_n27007_), .A2(pi0199), .B(new_n14428_), .ZN(new_n27008_));
  NAND2_X1   g23793(.A1(new_n27008_), .A2(new_n13613_), .ZN(new_n27009_));
  NAND2_X1   g23794(.A1(new_n15585_), .A2(new_n15578_), .ZN(new_n27010_));
  NAND3_X1   g23795(.A1(new_n27010_), .A2(new_n3259_), .A3(pi0199), .ZN(new_n27011_));
  NAND2_X1   g23796(.A1(new_n26964_), .A2(pi0199), .ZN(new_n27012_));
  OAI21_X1   g23797(.A1(new_n15588_), .A2(new_n27012_), .B(new_n3290_), .ZN(new_n27013_));
  NAND3_X1   g23798(.A1(new_n19390_), .A2(new_n27011_), .A3(new_n27013_), .ZN(new_n27014_));
  AOI21_X1   g23799(.A1(new_n15607_), .A2(pi0199), .B(new_n26964_), .ZN(new_n27015_));
  NOR4_X1    g23800(.A1(new_n27015_), .A2(new_n15628_), .A3(pi0199), .A4(new_n3290_), .ZN(new_n27016_));
  NAND2_X1   g23801(.A1(new_n27014_), .A2(new_n27016_), .ZN(new_n27017_));
  NOR2_X1    g23802(.A1(new_n27017_), .A2(new_n13614_), .ZN(new_n27018_));
  NAND4_X1   g23803(.A1(new_n26985_), .A2(new_n27003_), .A3(new_n27009_), .A4(new_n27018_), .ZN(new_n27019_));
  NAND2_X1   g23804(.A1(new_n27008_), .A2(pi0637), .ZN(new_n27020_));
  XOR2_X1    g23805(.A1(new_n27020_), .A2(new_n26984_), .Z(new_n27021_));
  NAND2_X1   g23806(.A1(new_n27008_), .A2(new_n26983_), .ZN(new_n27022_));
  OAI21_X1   g23807(.A1(new_n27017_), .A2(new_n26983_), .B(new_n27022_), .ZN(new_n27023_));
  NOR4_X1    g23808(.A1(new_n26982_), .A2(new_n13748_), .A3(pi1153), .A4(new_n27017_), .ZN(new_n27024_));
  NAND3_X1   g23809(.A1(new_n27003_), .A2(new_n27024_), .A3(new_n27023_), .ZN(new_n27025_));
  NOR2_X1    g23810(.A1(new_n27025_), .A2(new_n27021_), .ZN(new_n27026_));
  INV_X1     g23811(.I(new_n27026_), .ZN(new_n27027_));
  AOI21_X1   g23812(.A1(pi0778), .A2(new_n27019_), .B(new_n27027_), .ZN(new_n27028_));
  NAND2_X1   g23813(.A1(new_n27019_), .A2(pi0778), .ZN(new_n27029_));
  NOR2_X1    g23814(.A1(new_n27029_), .A2(new_n27026_), .ZN(new_n27030_));
  NOR2_X1    g23815(.A1(new_n27028_), .A2(new_n27030_), .ZN(new_n27031_));
  NAND2_X1   g23816(.A1(new_n26999_), .A2(new_n13775_), .ZN(new_n27032_));
  INV_X1     g23817(.I(new_n27032_), .ZN(new_n27033_));
  AOI21_X1   g23818(.A1(new_n26981_), .A2(new_n13776_), .B(new_n27033_), .ZN(new_n27034_));
  AOI21_X1   g23819(.A1(new_n27034_), .A2(pi0609), .B(new_n14694_), .ZN(new_n27035_));
  OAI21_X1   g23820(.A1(new_n27008_), .A2(new_n13775_), .B(new_n27032_), .ZN(new_n27036_));
  NOR3_X1    g23821(.A1(new_n27036_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n27037_));
  OAI21_X1   g23822(.A1(new_n27035_), .A2(new_n27037_), .B(new_n26999_), .ZN(new_n27038_));
  NOR2_X1    g23823(.A1(new_n26999_), .A2(pi0637), .ZN(new_n27039_));
  NOR3_X1    g23824(.A1(new_n26998_), .A2(new_n13748_), .A3(new_n27039_), .ZN(new_n27040_));
  MUX2_X1    g23825(.I0(new_n27040_), .I1(pi0778), .S(new_n27002_), .Z(new_n27041_));
  AOI21_X1   g23826(.A1(new_n27041_), .A2(new_n13766_), .B(new_n13785_), .ZN(new_n27042_));
  AOI21_X1   g23827(.A1(new_n27042_), .A2(new_n27038_), .B(pi0609), .ZN(new_n27043_));
  OAI21_X1   g23828(.A1(new_n27031_), .A2(new_n27043_), .B(pi0785), .ZN(new_n27044_));
  AOI21_X1   g23829(.A1(new_n27034_), .A2(pi1155), .B(new_n14694_), .ZN(new_n27045_));
  NOR3_X1    g23830(.A1(new_n27036_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n27046_));
  OAI21_X1   g23831(.A1(new_n27045_), .A2(new_n27046_), .B(new_n26999_), .ZN(new_n27047_));
  AOI21_X1   g23832(.A1(new_n27041_), .A2(pi0609), .B(new_n14465_), .ZN(new_n27048_));
  AOI21_X1   g23833(.A1(new_n27048_), .A2(new_n27047_), .B(pi0609), .ZN(new_n27049_));
  NOR3_X1    g23834(.A1(new_n27031_), .A2(new_n13801_), .A3(new_n27049_), .ZN(new_n27050_));
  XOR2_X1    g23835(.A1(new_n27050_), .A2(new_n27044_), .Z(new_n27051_));
  NOR4_X1    g23836(.A1(new_n27038_), .A2(new_n27047_), .A3(new_n13801_), .A4(new_n27034_), .ZN(new_n27052_));
  NAND2_X1   g23837(.A1(new_n27038_), .A2(pi0785), .ZN(new_n27053_));
  NOR3_X1    g23838(.A1(new_n27047_), .A2(new_n13801_), .A3(new_n27034_), .ZN(new_n27054_));
  NOR2_X1    g23839(.A1(new_n27054_), .A2(new_n27053_), .ZN(new_n27055_));
  NOR2_X1    g23840(.A1(new_n27055_), .A2(new_n27052_), .ZN(new_n27056_));
  AOI21_X1   g23841(.A1(new_n27056_), .A2(pi0618), .B(new_n13819_), .ZN(new_n27057_));
  INV_X1     g23842(.I(new_n26999_), .ZN(new_n27058_));
  NAND3_X1   g23843(.A1(new_n27036_), .A2(pi0609), .A3(pi1155), .ZN(new_n27059_));
  INV_X1     g23844(.I(new_n27037_), .ZN(new_n27060_));
  AOI21_X1   g23845(.A1(new_n27060_), .A2(new_n27059_), .B(new_n27058_), .ZN(new_n27061_));
  NAND3_X1   g23846(.A1(new_n27036_), .A2(pi0609), .A3(pi1155), .ZN(new_n27062_));
  NAND3_X1   g23847(.A1(new_n27034_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n27063_));
  AOI21_X1   g23848(.A1(new_n27063_), .A2(new_n27062_), .B(new_n27058_), .ZN(new_n27064_));
  NAND4_X1   g23849(.A1(new_n27061_), .A2(new_n27064_), .A3(pi0785), .A4(new_n27036_), .ZN(new_n27065_));
  NOR2_X1    g23850(.A1(new_n27034_), .A2(new_n13801_), .ZN(new_n27066_));
  NAND2_X1   g23851(.A1(new_n27064_), .A2(new_n27066_), .ZN(new_n27067_));
  NAND3_X1   g23852(.A1(new_n27067_), .A2(pi0785), .A3(new_n27038_), .ZN(new_n27068_));
  NAND2_X1   g23853(.A1(new_n27068_), .A2(new_n27065_), .ZN(new_n27069_));
  NOR3_X1    g23854(.A1(new_n27069_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n27070_));
  OAI21_X1   g23855(.A1(new_n27057_), .A2(new_n27070_), .B(new_n26999_), .ZN(new_n27071_));
  NOR2_X1    g23856(.A1(new_n27041_), .A2(new_n13803_), .ZN(new_n27072_));
  AOI21_X1   g23857(.A1(new_n13803_), .A2(new_n26999_), .B(new_n27072_), .ZN(new_n27073_));
  AOI21_X1   g23858(.A1(new_n27073_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n27074_));
  AOI21_X1   g23859(.A1(new_n27071_), .A2(new_n27074_), .B(pi0618), .ZN(new_n27075_));
  OAI21_X1   g23860(.A1(new_n27051_), .A2(new_n27075_), .B(pi0781), .ZN(new_n27076_));
  AOI21_X1   g23861(.A1(new_n27056_), .A2(pi1154), .B(new_n13819_), .ZN(new_n27077_));
  NAND4_X1   g23862(.A1(new_n27068_), .A2(new_n27065_), .A3(new_n13816_), .A4(pi1154), .ZN(new_n27078_));
  INV_X1     g23863(.I(new_n27078_), .ZN(new_n27079_));
  OAI21_X1   g23864(.A1(new_n27077_), .A2(new_n27079_), .B(new_n26999_), .ZN(new_n27080_));
  AOI21_X1   g23865(.A1(new_n27073_), .A2(pi0618), .B(new_n13837_), .ZN(new_n27081_));
  AOI21_X1   g23866(.A1(new_n27080_), .A2(new_n27081_), .B(pi0618), .ZN(new_n27082_));
  NOR3_X1    g23867(.A1(new_n27051_), .A2(new_n13855_), .A3(new_n27082_), .ZN(new_n27083_));
  NAND2_X1   g23868(.A1(new_n27083_), .A2(new_n27076_), .ZN(new_n27084_));
  XNOR2_X1   g23869(.A1(new_n27050_), .A2(new_n27044_), .ZN(new_n27085_));
  INV_X1     g23870(.I(new_n27075_), .ZN(new_n27086_));
  AOI21_X1   g23871(.A1(new_n27085_), .A2(new_n27086_), .B(new_n13855_), .ZN(new_n27087_));
  INV_X1     g23872(.I(new_n27082_), .ZN(new_n27088_));
  NAND3_X1   g23873(.A1(new_n27085_), .A2(pi0781), .A3(new_n27088_), .ZN(new_n27089_));
  NAND2_X1   g23874(.A1(new_n27087_), .A2(new_n27089_), .ZN(new_n27090_));
  NAND2_X1   g23875(.A1(new_n27090_), .A2(new_n27084_), .ZN(new_n27091_));
  NAND3_X1   g23876(.A1(new_n27069_), .A2(pi0618), .A3(pi1154), .ZN(new_n27092_));
  NAND3_X1   g23877(.A1(new_n27056_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n27093_));
  AOI21_X1   g23878(.A1(new_n27093_), .A2(new_n27092_), .B(new_n27058_), .ZN(new_n27094_));
  NAND3_X1   g23879(.A1(new_n27069_), .A2(pi0618), .A3(pi1154), .ZN(new_n27095_));
  AOI21_X1   g23880(.A1(new_n27095_), .A2(new_n27078_), .B(new_n27058_), .ZN(new_n27096_));
  NAND4_X1   g23881(.A1(new_n27094_), .A2(new_n27096_), .A3(pi0781), .A4(new_n27069_), .ZN(new_n27097_));
  NOR2_X1    g23882(.A1(new_n27056_), .A2(new_n13855_), .ZN(new_n27098_));
  NAND2_X1   g23883(.A1(new_n27096_), .A2(new_n27098_), .ZN(new_n27099_));
  NAND3_X1   g23884(.A1(new_n27099_), .A2(pi0781), .A3(new_n27071_), .ZN(new_n27100_));
  NAND2_X1   g23885(.A1(new_n27100_), .A2(new_n27097_), .ZN(new_n27101_));
  NAND3_X1   g23886(.A1(new_n27101_), .A2(pi0619), .A3(pi1159), .ZN(new_n27102_));
  NAND4_X1   g23887(.A1(new_n27100_), .A2(pi0619), .A3(new_n13868_), .A4(new_n27097_), .ZN(new_n27103_));
  AOI21_X1   g23888(.A1(new_n27102_), .A2(new_n27103_), .B(new_n27058_), .ZN(new_n27104_));
  NOR2_X1    g23889(.A1(new_n26999_), .A2(new_n13880_), .ZN(new_n27105_));
  AOI21_X1   g23890(.A1(new_n27073_), .A2(new_n13880_), .B(new_n27105_), .ZN(new_n27106_));
  INV_X1     g23891(.I(new_n27106_), .ZN(new_n27107_));
  AOI21_X1   g23892(.A1(new_n27107_), .A2(new_n13860_), .B(new_n14538_), .ZN(new_n27108_));
  INV_X1     g23893(.I(new_n27108_), .ZN(new_n27109_));
  OAI21_X1   g23894(.A1(new_n27104_), .A2(new_n27109_), .B(new_n13860_), .ZN(new_n27110_));
  NAND3_X1   g23895(.A1(new_n27101_), .A2(pi0619), .A3(pi1159), .ZN(new_n27111_));
  NAND4_X1   g23896(.A1(new_n27100_), .A2(new_n13860_), .A3(pi1159), .A4(new_n27097_), .ZN(new_n27112_));
  AOI21_X1   g23897(.A1(new_n27111_), .A2(new_n27112_), .B(new_n27058_), .ZN(new_n27113_));
  AOI21_X1   g23898(.A1(new_n27107_), .A2(pi0619), .B(new_n15217_), .ZN(new_n27114_));
  INV_X1     g23899(.I(new_n27114_), .ZN(new_n27115_));
  OAI21_X1   g23900(.A1(new_n27113_), .A2(new_n27115_), .B(new_n13860_), .ZN(new_n27116_));
  NAND4_X1   g23901(.A1(new_n27110_), .A2(new_n27116_), .A3(pi0789), .A4(new_n27091_), .ZN(new_n27117_));
  AOI21_X1   g23902(.A1(new_n27110_), .A2(new_n27091_), .B(new_n13896_), .ZN(new_n27118_));
  AOI21_X1   g23903(.A1(new_n27090_), .A2(new_n27084_), .B(new_n13896_), .ZN(new_n27119_));
  NAND2_X1   g23904(.A1(new_n27116_), .A2(new_n27119_), .ZN(new_n27120_));
  NAND2_X1   g23905(.A1(new_n27118_), .A2(new_n27120_), .ZN(new_n27121_));
  NAND2_X1   g23906(.A1(new_n27121_), .A2(new_n27117_), .ZN(new_n27122_));
  NAND4_X1   g23907(.A1(new_n27104_), .A2(new_n27113_), .A3(pi0789), .A4(new_n27101_), .ZN(new_n27123_));
  NOR4_X1    g23908(.A1(new_n27071_), .A2(new_n27080_), .A3(new_n13855_), .A4(new_n27056_), .ZN(new_n27124_));
  NAND2_X1   g23909(.A1(new_n27071_), .A2(pi0781), .ZN(new_n27125_));
  NOR3_X1    g23910(.A1(new_n27080_), .A2(new_n13855_), .A3(new_n27056_), .ZN(new_n27126_));
  NOR2_X1    g23911(.A1(new_n27126_), .A2(new_n27125_), .ZN(new_n27127_));
  NOR2_X1    g23912(.A1(new_n27127_), .A2(new_n27124_), .ZN(new_n27128_));
  AOI21_X1   g23913(.A1(new_n27128_), .A2(pi0619), .B(new_n13904_), .ZN(new_n27129_));
  INV_X1     g23914(.I(new_n27103_), .ZN(new_n27130_));
  OAI21_X1   g23915(.A1(new_n27129_), .A2(new_n27130_), .B(new_n26999_), .ZN(new_n27131_));
  NOR2_X1    g23916(.A1(new_n27128_), .A2(new_n13896_), .ZN(new_n27132_));
  NAND2_X1   g23917(.A1(new_n27113_), .A2(new_n27132_), .ZN(new_n27133_));
  NAND3_X1   g23918(.A1(new_n27133_), .A2(pi0789), .A3(new_n27131_), .ZN(new_n27134_));
  NOR2_X1    g23919(.A1(new_n27058_), .A2(new_n13919_), .ZN(new_n27135_));
  AOI21_X1   g23920(.A1(new_n27106_), .A2(new_n13919_), .B(new_n27135_), .ZN(new_n27136_));
  NOR2_X1    g23921(.A1(new_n13901_), .A2(new_n13922_), .ZN(new_n27137_));
  INV_X1     g23922(.I(new_n27137_), .ZN(new_n27138_));
  AOI21_X1   g23923(.A1(new_n27134_), .A2(new_n27123_), .B(new_n27138_), .ZN(new_n27139_));
  NAND3_X1   g23924(.A1(new_n27122_), .A2(pi0626), .A3(pi0788), .ZN(new_n27143_));
  INV_X1     g23925(.I(new_n27117_), .ZN(new_n27144_));
  NOR2_X1    g23926(.A1(new_n27087_), .A2(new_n27089_), .ZN(new_n27145_));
  NOR2_X1    g23927(.A1(new_n27083_), .A2(new_n27076_), .ZN(new_n27146_));
  NOR2_X1    g23928(.A1(new_n27145_), .A2(new_n27146_), .ZN(new_n27147_));
  AOI21_X1   g23929(.A1(new_n27131_), .A2(new_n27108_), .B(pi0619), .ZN(new_n27148_));
  OAI21_X1   g23930(.A1(new_n27148_), .A2(new_n27147_), .B(pi0789), .ZN(new_n27149_));
  AOI21_X1   g23931(.A1(new_n27128_), .A2(pi1159), .B(new_n13904_), .ZN(new_n27150_));
  INV_X1     g23932(.I(new_n27112_), .ZN(new_n27151_));
  OAI21_X1   g23933(.A1(new_n27150_), .A2(new_n27151_), .B(new_n26999_), .ZN(new_n27152_));
  AOI21_X1   g23934(.A1(new_n27152_), .A2(new_n27114_), .B(pi0619), .ZN(new_n27153_));
  OAI21_X1   g23935(.A1(new_n27145_), .A2(new_n27146_), .B(pi0789), .ZN(new_n27154_));
  NOR2_X1    g23936(.A1(new_n27153_), .A2(new_n27154_), .ZN(new_n27155_));
  NOR2_X1    g23937(.A1(new_n27149_), .A2(new_n27155_), .ZN(new_n27156_));
  OAI22_X1   g23938(.A1(new_n27156_), .A2(new_n27144_), .B1(new_n27139_), .B2(pi0626), .ZN(new_n27157_));
  OAI21_X1   g23939(.A1(new_n27156_), .A2(new_n27144_), .B(new_n14577_), .ZN(new_n27158_));
  NAND3_X1   g23940(.A1(new_n27157_), .A2(new_n27158_), .A3(pi0788), .ZN(new_n27159_));
  NAND2_X1   g23941(.A1(new_n27159_), .A2(new_n27143_), .ZN(new_n27160_));
  INV_X1     g23942(.I(new_n27123_), .ZN(new_n27161_));
  NAND2_X1   g23943(.A1(new_n27131_), .A2(pi0789), .ZN(new_n27162_));
  NOR3_X1    g23944(.A1(new_n27152_), .A2(new_n13896_), .A3(new_n27128_), .ZN(new_n27163_));
  NOR2_X1    g23945(.A1(new_n27163_), .A2(new_n27162_), .ZN(new_n27164_));
  OAI21_X1   g23946(.A1(new_n27164_), .A2(new_n27161_), .B(new_n16372_), .ZN(new_n27165_));
  NOR2_X1    g23947(.A1(new_n26999_), .A2(new_n16372_), .ZN(new_n27166_));
  INV_X1     g23948(.I(new_n27166_), .ZN(new_n27167_));
  NAND2_X1   g23949(.A1(new_n27165_), .A2(new_n27167_), .ZN(new_n27168_));
  NOR2_X1    g23950(.A1(new_n26999_), .A2(new_n13966_), .ZN(new_n27169_));
  INV_X1     g23951(.I(new_n27169_), .ZN(new_n27170_));
  NAND2_X1   g23952(.A1(new_n27136_), .A2(new_n13966_), .ZN(new_n27171_));
  NAND2_X1   g23953(.A1(new_n27171_), .A2(new_n27170_), .ZN(new_n27172_));
  NAND3_X1   g23954(.A1(new_n27172_), .A2(pi0628), .A3(pi1156), .ZN(new_n27173_));
  NAND4_X1   g23955(.A1(new_n27171_), .A2(pi0628), .A3(new_n13969_), .A4(new_n27170_), .ZN(new_n27174_));
  AOI21_X1   g23956(.A1(new_n27173_), .A2(new_n27174_), .B(new_n27058_), .ZN(new_n27175_));
  NOR2_X1    g23957(.A1(new_n27175_), .A2(new_n15270_), .ZN(new_n27176_));
  INV_X1     g23958(.I(new_n27176_), .ZN(new_n27177_));
  NAND2_X1   g23959(.A1(new_n27134_), .A2(new_n27123_), .ZN(new_n27179_));
  AOI21_X1   g23960(.A1(new_n27179_), .A2(new_n16372_), .B(new_n27166_), .ZN(new_n27180_));
  NAND3_X1   g23961(.A1(new_n27172_), .A2(pi0628), .A3(pi1156), .ZN(new_n27182_));
  NAND4_X1   g23962(.A1(new_n27171_), .A2(new_n13942_), .A3(pi1156), .A4(new_n27170_), .ZN(new_n27183_));
  AOI21_X1   g23963(.A1(new_n27182_), .A2(new_n27183_), .B(new_n27058_), .ZN(new_n27184_));
  NAND3_X1   g23964(.A1(new_n27160_), .A2(pi0628), .A3(pi0792), .ZN(new_n27186_));
  NOR2_X1    g23965(.A1(new_n27156_), .A2(new_n27144_), .ZN(new_n27187_));
  NOR3_X1    g23966(.A1(new_n27187_), .A2(new_n13901_), .A3(new_n13937_), .ZN(new_n27188_));
  OAI21_X1   g23967(.A1(new_n27164_), .A2(new_n27161_), .B(new_n27137_), .ZN(new_n27189_));
  AOI22_X1   g23968(.A1(new_n27189_), .A2(new_n13901_), .B1(new_n27121_), .B2(new_n27117_), .ZN(new_n27190_));
  AOI21_X1   g23969(.A1(new_n27121_), .A2(new_n27117_), .B(new_n15258_), .ZN(new_n27191_));
  NOR3_X1    g23970(.A1(new_n27190_), .A2(new_n13937_), .A3(new_n27191_), .ZN(new_n27192_));
  OAI21_X1   g23971(.A1(new_n27168_), .A2(new_n27177_), .B(new_n13942_), .ZN(new_n27193_));
  OAI21_X1   g23972(.A1(new_n27192_), .A2(new_n27188_), .B(new_n27193_), .ZN(new_n27194_));
  OAI21_X1   g23973(.A1(new_n27192_), .A2(new_n27188_), .B(new_n14606_), .ZN(new_n27195_));
  NAND3_X1   g23974(.A1(new_n27194_), .A2(new_n27195_), .A3(pi0792), .ZN(new_n27196_));
  NAND2_X1   g23975(.A1(new_n27196_), .A2(new_n27186_), .ZN(new_n27197_));
  NOR2_X1    g23976(.A1(new_n26999_), .A2(new_n13994_), .ZN(new_n27198_));
  AOI21_X1   g23977(.A1(new_n27168_), .A2(new_n13994_), .B(new_n27198_), .ZN(new_n27199_));
  INV_X1     g23978(.I(new_n27199_), .ZN(new_n27200_));
  NAND4_X1   g23979(.A1(new_n27175_), .A2(new_n27184_), .A3(pi0792), .A4(new_n27172_), .ZN(new_n27201_));
  NOR2_X1    g23980(.A1(new_n27175_), .A2(new_n12777_), .ZN(new_n27202_));
  NAND3_X1   g23981(.A1(new_n27184_), .A2(pi0792), .A3(new_n27172_), .ZN(new_n27203_));
  NAND2_X1   g23982(.A1(new_n27203_), .A2(new_n27202_), .ZN(new_n27204_));
  NAND2_X1   g23983(.A1(new_n27204_), .A2(new_n27201_), .ZN(new_n27205_));
  INV_X1     g23984(.I(new_n27205_), .ZN(new_n27206_));
  AOI21_X1   g23985(.A1(new_n27206_), .A2(pi0647), .B(new_n14008_), .ZN(new_n27207_));
  NOR3_X1    g23986(.A1(new_n27205_), .A2(new_n14005_), .A3(pi1157), .ZN(new_n27208_));
  OAI21_X1   g23987(.A1(new_n27207_), .A2(new_n27208_), .B(new_n26999_), .ZN(new_n27209_));
  NAND2_X1   g23988(.A1(new_n27209_), .A2(new_n14011_), .ZN(new_n27210_));
  OAI21_X1   g23989(.A1(new_n27200_), .A2(new_n27210_), .B(new_n14005_), .ZN(new_n27211_));
  NAND3_X1   g23990(.A1(new_n27205_), .A2(pi0647), .A3(pi1157), .ZN(new_n27212_));
  NAND3_X1   g23991(.A1(new_n27206_), .A2(pi1157), .A3(new_n14008_), .ZN(new_n27213_));
  NAND2_X1   g23992(.A1(new_n27213_), .A2(new_n27212_), .ZN(new_n27214_));
  AOI21_X1   g23993(.A1(new_n27214_), .A2(new_n26999_), .B(new_n16329_), .ZN(new_n27215_));
  OAI21_X1   g23994(.A1(new_n27199_), .A2(new_n14005_), .B(new_n27215_), .ZN(new_n27216_));
  NAND2_X1   g23995(.A1(new_n27216_), .A2(new_n14005_), .ZN(new_n27217_));
  NAND4_X1   g23996(.A1(new_n27197_), .A2(pi0787), .A3(new_n27211_), .A4(new_n27217_), .ZN(new_n27218_));
  NOR2_X1    g23997(.A1(new_n27192_), .A2(new_n27188_), .ZN(new_n27219_));
  NOR3_X1    g23998(.A1(new_n27219_), .A2(new_n13942_), .A3(new_n12777_), .ZN(new_n27220_));
  AOI21_X1   g23999(.A1(new_n27180_), .A2(new_n27176_), .B(pi0628), .ZN(new_n27221_));
  AOI21_X1   g24000(.A1(new_n27159_), .A2(new_n27143_), .B(new_n27221_), .ZN(new_n27222_));
  AOI21_X1   g24001(.A1(new_n27159_), .A2(new_n27143_), .B(new_n15296_), .ZN(new_n27223_));
  NOR3_X1    g24002(.A1(new_n27222_), .A2(new_n27223_), .A3(new_n12777_), .ZN(new_n27224_));
  OAI21_X1   g24003(.A1(new_n27224_), .A2(new_n27220_), .B(new_n27211_), .ZN(new_n27225_));
  AOI21_X1   g24004(.A1(new_n27216_), .A2(new_n14005_), .B(new_n12776_), .ZN(new_n27226_));
  OAI21_X1   g24005(.A1(new_n27224_), .A2(new_n27220_), .B(new_n27226_), .ZN(new_n27227_));
  NAND3_X1   g24006(.A1(new_n27225_), .A2(new_n27227_), .A3(pi0787), .ZN(new_n27228_));
  NAND2_X1   g24007(.A1(new_n26999_), .A2(new_n14210_), .ZN(new_n27229_));
  NAND2_X1   g24008(.A1(new_n27199_), .A2(new_n14211_), .ZN(new_n27230_));
  NAND2_X1   g24009(.A1(new_n27230_), .A2(new_n27229_), .ZN(new_n27231_));
  NAND4_X1   g24010(.A1(new_n27214_), .A2(pi0787), .A3(new_n26999_), .A4(new_n27205_), .ZN(new_n27232_));
  AOI21_X1   g24011(.A1(pi0787), .A2(new_n27209_), .B(new_n27232_), .ZN(new_n27233_));
  NAND2_X1   g24012(.A1(new_n27209_), .A2(pi0787), .ZN(new_n27234_));
  INV_X1     g24013(.I(new_n27232_), .ZN(new_n27235_));
  NOR2_X1    g24014(.A1(new_n27235_), .A2(new_n27234_), .ZN(new_n27236_));
  OAI21_X1   g24015(.A1(new_n27236_), .A2(new_n27233_), .B(pi0644), .ZN(new_n27237_));
  NOR2_X1    g24016(.A1(new_n14204_), .A2(pi0715), .ZN(new_n27238_));
  NAND3_X1   g24017(.A1(new_n27237_), .A2(new_n27231_), .A3(new_n27238_), .ZN(new_n27239_));
  AOI22_X1   g24018(.A1(new_n27228_), .A2(new_n27218_), .B1(new_n14204_), .B2(new_n27239_), .ZN(new_n27240_));
  INV_X1     g24019(.I(new_n27231_), .ZN(new_n27241_));
  NAND2_X1   g24020(.A1(pi0644), .A2(pi0715), .ZN(new_n27244_));
  OAI21_X1   g24021(.A1(new_n27241_), .A2(new_n27244_), .B(new_n14204_), .ZN(new_n27245_));
  NAND2_X1   g24022(.A1(new_n27245_), .A2(pi0790), .ZN(new_n27246_));
  AOI21_X1   g24023(.A1(new_n27228_), .A2(new_n27218_), .B(new_n27246_), .ZN(new_n27247_));
  NOR3_X1    g24024(.A1(new_n27240_), .A2(new_n27247_), .A3(new_n12775_), .ZN(new_n27248_));
  NAND2_X1   g24025(.A1(new_n27228_), .A2(new_n27218_), .ZN(new_n27249_));
  NAND2_X1   g24026(.A1(new_n27239_), .A2(new_n14204_), .ZN(new_n27250_));
  NAND4_X1   g24027(.A1(new_n27249_), .A2(pi0790), .A3(new_n27250_), .A4(new_n27245_), .ZN(new_n27251_));
  NAND2_X1   g24028(.A1(new_n27251_), .A2(new_n7240_), .ZN(new_n27252_));
  OAI21_X1   g24029(.A1(new_n27252_), .A2(new_n27248_), .B(new_n26963_), .ZN(po0356));
  NOR2_X1    g24030(.A1(new_n14428_), .A2(new_n8555_), .ZN(new_n27254_));
  NOR2_X1    g24031(.A1(new_n19327_), .A2(new_n8555_), .ZN(new_n27255_));
  NOR2_X1    g24032(.A1(new_n3259_), .A2(new_n8555_), .ZN(new_n27256_));
  XOR2_X1    g24033(.A1(new_n27255_), .A2(new_n27256_), .Z(new_n27257_));
  NAND2_X1   g24034(.A1(new_n27257_), .A2(new_n26975_), .ZN(new_n27258_));
  AOI21_X1   g24035(.A1(new_n27258_), .A2(new_n8555_), .B(new_n19641_), .ZN(new_n27259_));
  AND3_X2    g24036(.A1(new_n27259_), .A2(pi0606), .A3(new_n3289_), .Z(new_n27260_));
  INV_X1     g24037(.I(pi0606), .ZN(new_n27261_));
  NOR3_X1    g24038(.A1(new_n27259_), .A2(new_n27261_), .A3(new_n3289_), .ZN(new_n27262_));
  OAI21_X1   g24039(.A1(new_n27260_), .A2(new_n27262_), .B(pi0200), .ZN(new_n27263_));
  INV_X1     g24040(.I(new_n27254_), .ZN(new_n27264_));
  NAND2_X1   g24041(.A1(new_n27264_), .A2(new_n27261_), .ZN(new_n27265_));
  NAND3_X1   g24042(.A1(new_n27263_), .A2(new_n13776_), .A3(new_n27265_), .ZN(new_n27266_));
  NOR2_X1    g24043(.A1(new_n27264_), .A2(new_n13776_), .ZN(new_n27267_));
  INV_X1     g24044(.I(new_n27267_), .ZN(new_n27268_));
  NAND2_X1   g24045(.A1(new_n27266_), .A2(new_n27268_), .ZN(new_n27269_));
  NAND3_X1   g24046(.A1(new_n27269_), .A2(pi0609), .A3(pi1155), .ZN(new_n27270_));
  NOR3_X1    g24047(.A1(new_n27269_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n27271_));
  INV_X1     g24048(.I(new_n27271_), .ZN(new_n27272_));
  AOI21_X1   g24049(.A1(new_n27272_), .A2(new_n27270_), .B(new_n27264_), .ZN(new_n27273_));
  NAND3_X1   g24050(.A1(new_n27269_), .A2(pi0609), .A3(pi1155), .ZN(new_n27274_));
  INV_X1     g24051(.I(new_n27269_), .ZN(new_n27275_));
  NAND3_X1   g24052(.A1(new_n27275_), .A2(pi1155), .A3(new_n14694_), .ZN(new_n27276_));
  AOI21_X1   g24053(.A1(new_n27276_), .A2(new_n27274_), .B(new_n27264_), .ZN(new_n27277_));
  NAND4_X1   g24054(.A1(new_n27273_), .A2(new_n27277_), .A3(pi0785), .A4(new_n27269_), .ZN(new_n27278_));
  NOR2_X1    g24055(.A1(new_n27273_), .A2(new_n13801_), .ZN(new_n27279_));
  NAND3_X1   g24056(.A1(new_n27277_), .A2(pi0785), .A3(new_n27269_), .ZN(new_n27280_));
  NAND2_X1   g24057(.A1(new_n27279_), .A2(new_n27280_), .ZN(new_n27281_));
  NAND2_X1   g24058(.A1(new_n27281_), .A2(new_n27278_), .ZN(new_n27282_));
  INV_X1     g24059(.I(new_n27282_), .ZN(new_n27283_));
  NOR2_X1    g24060(.A1(new_n27283_), .A2(pi0781), .ZN(new_n27284_));
  NAND3_X1   g24061(.A1(new_n27282_), .A2(new_n16689_), .A3(new_n27254_), .ZN(new_n27285_));
  NAND4_X1   g24062(.A1(new_n27281_), .A2(new_n16689_), .A3(new_n27264_), .A4(new_n27278_), .ZN(new_n27286_));
  AOI21_X1   g24063(.A1(new_n27285_), .A2(new_n27286_), .B(new_n13855_), .ZN(new_n27287_));
  NOR2_X1    g24064(.A1(new_n27287_), .A2(new_n27284_), .ZN(new_n27288_));
  AOI21_X1   g24065(.A1(new_n27288_), .A2(pi0619), .B(new_n13904_), .ZN(new_n27289_));
  NOR4_X1    g24066(.A1(new_n27287_), .A2(new_n13860_), .A3(pi1159), .A4(new_n27284_), .ZN(new_n27290_));
  OAI21_X1   g24067(.A1(new_n27289_), .A2(new_n27290_), .B(new_n27254_), .ZN(new_n27291_));
  INV_X1     g24068(.I(new_n27291_), .ZN(new_n27292_));
  NOR2_X1    g24069(.A1(new_n27254_), .A2(new_n13880_), .ZN(new_n27293_));
  NOR2_X1    g24070(.A1(new_n27264_), .A2(new_n13805_), .ZN(new_n27294_));
  INV_X1     g24071(.I(pi0643), .ZN(new_n27295_));
  NOR2_X1    g24072(.A1(new_n16149_), .A2(new_n8555_), .ZN(new_n27296_));
  INV_X1     g24073(.I(new_n27296_), .ZN(new_n27297_));
  NOR2_X1    g24074(.A1(new_n8555_), .A2(new_n3098_), .ZN(new_n27298_));
  INV_X1     g24075(.I(new_n27298_), .ZN(new_n27299_));
  AOI21_X1   g24076(.A1(new_n13699_), .A2(new_n3090_), .B(new_n13703_), .ZN(new_n27300_));
  NOR2_X1    g24077(.A1(new_n27300_), .A2(new_n8555_), .ZN(new_n27301_));
  XOR2_X1    g24078(.A1(new_n27301_), .A2(new_n27299_), .Z(new_n27302_));
  OAI21_X1   g24079(.A1(new_n14414_), .A2(new_n14415_), .B(new_n14418_), .ZN(new_n27303_));
  NAND4_X1   g24080(.A1(new_n13197_), .A2(pi0039), .A3(new_n13165_), .A4(pi0200), .ZN(new_n27304_));
  OAI21_X1   g24081(.A1(new_n27302_), .A2(new_n27303_), .B(new_n27304_), .ZN(new_n27305_));
  OAI21_X1   g24082(.A1(new_n13710_), .A2(pi0215), .B(new_n13713_), .ZN(new_n27306_));
  NAND2_X1   g24083(.A1(new_n27306_), .A2(pi0299), .ZN(new_n27307_));
  XOR2_X1    g24084(.A1(new_n27307_), .A2(new_n27299_), .Z(new_n27308_));
  NAND2_X1   g24085(.A1(new_n14406_), .A2(new_n14407_), .ZN(new_n27309_));
  NAND4_X1   g24086(.A1(new_n27305_), .A2(new_n13683_), .A3(new_n27308_), .A4(new_n27309_), .ZN(new_n27310_));
  NAND2_X1   g24087(.A1(new_n27310_), .A2(new_n3259_), .ZN(new_n27311_));
  AOI21_X1   g24088(.A1(new_n27311_), .A2(new_n27297_), .B(new_n27295_), .ZN(new_n27312_));
  NOR2_X1    g24089(.A1(new_n3290_), .A2(new_n27295_), .ZN(new_n27313_));
  XNOR2_X1   g24090(.A1(new_n27312_), .A2(new_n27313_), .ZN(new_n27314_));
  OAI22_X1   g24091(.A1(new_n27314_), .A2(new_n8555_), .B1(pi0643), .B2(new_n27254_), .ZN(new_n27315_));
  AOI21_X1   g24092(.A1(new_n27315_), .A2(pi0625), .B(new_n13620_), .ZN(new_n27316_));
  INV_X1     g24093(.I(new_n27315_), .ZN(new_n27317_));
  NOR3_X1    g24094(.A1(new_n27317_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n27318_));
  OAI21_X1   g24095(.A1(new_n27318_), .A2(new_n27316_), .B(new_n27254_), .ZN(new_n27319_));
  AOI21_X1   g24096(.A1(new_n27315_), .A2(pi1153), .B(new_n13620_), .ZN(new_n27320_));
  NAND3_X1   g24097(.A1(new_n27315_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n27321_));
  INV_X1     g24098(.I(new_n27321_), .ZN(new_n27322_));
  OAI21_X1   g24099(.A1(new_n27322_), .A2(new_n27320_), .B(new_n27254_), .ZN(new_n27323_));
  NOR4_X1    g24100(.A1(new_n27319_), .A2(new_n27323_), .A3(new_n13748_), .A4(new_n27315_), .ZN(new_n27324_));
  NAND2_X1   g24101(.A1(new_n27319_), .A2(pi0778), .ZN(new_n27325_));
  NOR3_X1    g24102(.A1(new_n27323_), .A2(new_n13748_), .A3(new_n27315_), .ZN(new_n27326_));
  NOR2_X1    g24103(.A1(new_n27326_), .A2(new_n27325_), .ZN(new_n27327_));
  NOR2_X1    g24104(.A1(new_n27327_), .A2(new_n27324_), .ZN(new_n27328_));
  AOI21_X1   g24105(.A1(new_n27328_), .A2(new_n13805_), .B(new_n27294_), .ZN(new_n27329_));
  AOI21_X1   g24106(.A1(new_n27329_), .A2(new_n13880_), .B(new_n27293_), .ZN(new_n27330_));
  NAND2_X1   g24107(.A1(new_n27263_), .A2(new_n27265_), .ZN(new_n27331_));
  INV_X1     g24108(.I(new_n27331_), .ZN(new_n27332_));
  INV_X1     g24109(.I(new_n19651_), .ZN(new_n27333_));
  NAND2_X1   g24110(.A1(new_n27010_), .A2(pi0200), .ZN(new_n27334_));
  XOR2_X1    g24111(.A1(new_n27334_), .A2(new_n27256_), .Z(new_n27335_));
  NOR3_X1    g24112(.A1(new_n27335_), .A2(new_n27333_), .A3(new_n27297_), .ZN(new_n27336_));
  NOR2_X1    g24113(.A1(new_n27336_), .A2(new_n13213_), .ZN(new_n27337_));
  AOI21_X1   g24114(.A1(pi0038), .A2(new_n15621_), .B(new_n15619_), .ZN(new_n27338_));
  INV_X1     g24115(.I(new_n27256_), .ZN(new_n27339_));
  NOR2_X1    g24116(.A1(new_n19657_), .A2(new_n8555_), .ZN(new_n27340_));
  XOR2_X1    g24117(.A1(new_n27340_), .A2(new_n27339_), .Z(new_n27341_));
  NOR4_X1    g24118(.A1(new_n19662_), .A2(new_n27261_), .A3(new_n3290_), .A4(new_n27339_), .ZN(new_n27342_));
  NAND3_X1   g24119(.A1(new_n13198_), .A2(new_n3183_), .A3(new_n27342_), .ZN(new_n27343_));
  NOR2_X1    g24120(.A1(new_n27341_), .A2(new_n27343_), .ZN(new_n27344_));
  OAI21_X1   g24121(.A1(new_n27344_), .A2(new_n27338_), .B(new_n3289_), .ZN(new_n27345_));
  NAND2_X1   g24122(.A1(new_n27338_), .A2(pi0200), .ZN(new_n27346_));
  AND3_X2    g24123(.A1(new_n27346_), .A2(new_n27261_), .A3(new_n3290_), .Z(new_n27347_));
  NAND2_X1   g24124(.A1(new_n27345_), .A2(new_n27347_), .ZN(new_n27348_));
  NOR2_X1    g24125(.A1(new_n13721_), .A2(new_n27295_), .ZN(new_n27349_));
  NAND2_X1   g24126(.A1(new_n27348_), .A2(new_n27349_), .ZN(new_n27350_));
  OAI22_X1   g24127(.A1(new_n27350_), .A2(new_n27337_), .B1(new_n27332_), .B2(pi0643), .ZN(new_n27351_));
  NOR2_X1    g24128(.A1(new_n27351_), .A2(new_n13613_), .ZN(new_n27352_));
  NOR2_X1    g24129(.A1(new_n27352_), .A2(new_n13620_), .ZN(new_n27353_));
  NAND2_X1   g24130(.A1(new_n27352_), .A2(new_n13620_), .ZN(new_n27354_));
  INV_X1     g24131(.I(new_n27354_), .ZN(new_n27355_));
  OAI21_X1   g24132(.A1(new_n27355_), .A2(new_n27353_), .B(new_n27332_), .ZN(new_n27356_));
  INV_X1     g24133(.I(new_n27320_), .ZN(new_n27357_));
  AOI21_X1   g24134(.A1(new_n27357_), .A2(new_n27321_), .B(new_n27264_), .ZN(new_n27358_));
  NOR2_X1    g24135(.A1(new_n27358_), .A2(pi0608), .ZN(new_n27359_));
  NAND2_X1   g24136(.A1(new_n27319_), .A2(new_n14081_), .ZN(new_n27360_));
  AOI21_X1   g24137(.A1(new_n27356_), .A2(new_n27359_), .B(new_n27360_), .ZN(new_n27361_));
  NAND3_X1   g24138(.A1(new_n27351_), .A2(pi0625), .A3(pi1153), .ZN(new_n27362_));
  NOR2_X1    g24139(.A1(new_n27351_), .A2(new_n13614_), .ZN(new_n27363_));
  NAND2_X1   g24140(.A1(new_n27363_), .A2(new_n13620_), .ZN(new_n27364_));
  NAND2_X1   g24141(.A1(new_n27364_), .A2(new_n27362_), .ZN(new_n27365_));
  NOR2_X1    g24142(.A1(new_n27331_), .A2(new_n13748_), .ZN(new_n27366_));
  NAND2_X1   g24143(.A1(new_n27365_), .A2(new_n27366_), .ZN(new_n27367_));
  OAI22_X1   g24144(.A1(new_n27361_), .A2(new_n27367_), .B1(pi0778), .B2(new_n27351_), .ZN(new_n27368_));
  NAND3_X1   g24145(.A1(new_n27368_), .A2(pi0609), .A3(pi1155), .ZN(new_n27369_));
  INV_X1     g24146(.I(new_n27351_), .ZN(new_n27370_));
  INV_X1     g24147(.I(new_n27353_), .ZN(new_n27371_));
  AOI21_X1   g24148(.A1(new_n27371_), .A2(new_n27354_), .B(new_n27331_), .ZN(new_n27372_));
  INV_X1     g24149(.I(new_n27359_), .ZN(new_n27373_));
  INV_X1     g24150(.I(new_n27360_), .ZN(new_n27374_));
  OAI21_X1   g24151(.A1(new_n27372_), .A2(new_n27373_), .B(new_n27374_), .ZN(new_n27375_));
  INV_X1     g24152(.I(new_n27367_), .ZN(new_n27376_));
  AOI22_X1   g24153(.A1(new_n27375_), .A2(new_n27376_), .B1(new_n13748_), .B2(new_n27370_), .ZN(new_n27377_));
  NAND3_X1   g24154(.A1(new_n27377_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n27378_));
  AOI21_X1   g24155(.A1(new_n27378_), .A2(new_n27369_), .B(new_n27328_), .ZN(new_n27379_));
  NOR2_X1    g24156(.A1(new_n27273_), .A2(new_n13783_), .ZN(new_n27380_));
  INV_X1     g24157(.I(new_n27380_), .ZN(new_n27381_));
  OAI21_X1   g24158(.A1(new_n27379_), .A2(new_n27381_), .B(pi0785), .ZN(new_n27382_));
  INV_X1     g24159(.I(new_n27328_), .ZN(new_n27383_));
  NAND3_X1   g24160(.A1(new_n27368_), .A2(pi0609), .A3(pi1155), .ZN(new_n27384_));
  NAND3_X1   g24161(.A1(new_n27377_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n27385_));
  NAND2_X1   g24162(.A1(new_n27385_), .A2(new_n27384_), .ZN(new_n27386_));
  INV_X1     g24163(.I(new_n27277_), .ZN(new_n27387_));
  NAND3_X1   g24164(.A1(new_n27368_), .A2(new_n16780_), .A3(new_n27387_), .ZN(new_n27388_));
  AOI21_X1   g24165(.A1(new_n27386_), .A2(new_n27383_), .B(new_n27388_), .ZN(new_n27389_));
  NAND2_X1   g24166(.A1(new_n27382_), .A2(new_n27389_), .ZN(new_n27390_));
  AOI21_X1   g24167(.A1(new_n27377_), .A2(pi1155), .B(new_n14694_), .ZN(new_n27391_));
  NOR3_X1    g24168(.A1(new_n27368_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n27392_));
  OAI21_X1   g24169(.A1(new_n27391_), .A2(new_n27392_), .B(new_n27383_), .ZN(new_n27393_));
  AOI21_X1   g24170(.A1(new_n27393_), .A2(new_n27380_), .B(new_n13801_), .ZN(new_n27394_));
  AOI21_X1   g24171(.A1(new_n27377_), .A2(pi0609), .B(new_n14694_), .ZN(new_n27395_));
  NOR3_X1    g24172(.A1(new_n27368_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n27396_));
  OAI21_X1   g24173(.A1(new_n27395_), .A2(new_n27396_), .B(new_n27383_), .ZN(new_n27397_));
  NAND4_X1   g24174(.A1(new_n27397_), .A2(new_n16780_), .A3(new_n27387_), .A4(new_n27368_), .ZN(new_n27398_));
  NAND2_X1   g24175(.A1(new_n27398_), .A2(new_n27394_), .ZN(new_n27399_));
  NAND2_X1   g24176(.A1(new_n27399_), .A2(new_n27390_), .ZN(new_n27400_));
  NAND2_X1   g24177(.A1(new_n27264_), .A2(pi0618), .ZN(new_n27401_));
  AOI21_X1   g24178(.A1(new_n13877_), .A2(new_n27401_), .B(new_n27282_), .ZN(new_n27402_));
  INV_X1     g24179(.I(new_n27402_), .ZN(new_n27403_));
  NOR2_X1    g24180(.A1(new_n13816_), .A2(new_n13817_), .ZN(new_n27404_));
  AOI21_X1   g24181(.A1(new_n27403_), .A2(new_n27404_), .B(pi0618), .ZN(new_n27405_));
  INV_X1     g24182(.I(new_n27405_), .ZN(new_n27406_));
  NAND2_X1   g24183(.A1(new_n27329_), .A2(pi0618), .ZN(new_n27407_));
  AOI21_X1   g24184(.A1(new_n27254_), .A2(new_n13824_), .B(pi0618), .ZN(new_n27408_));
  INV_X1     g24185(.I(new_n27408_), .ZN(new_n27409_));
  NAND4_X1   g24186(.A1(new_n27407_), .A2(new_n13817_), .A3(new_n27282_), .A4(new_n27409_), .ZN(new_n27410_));
  NAND2_X1   g24187(.A1(new_n27410_), .A2(new_n13816_), .ZN(new_n27411_));
  NAND4_X1   g24188(.A1(new_n27400_), .A2(pi0781), .A3(new_n27406_), .A4(new_n27411_), .ZN(new_n27412_));
  NOR2_X1    g24189(.A1(new_n27398_), .A2(new_n27394_), .ZN(new_n27413_));
  NOR2_X1    g24190(.A1(new_n27382_), .A2(new_n27389_), .ZN(new_n27414_));
  OAI21_X1   g24191(.A1(new_n27413_), .A2(new_n27414_), .B(new_n27406_), .ZN(new_n27415_));
  INV_X1     g24192(.I(new_n27411_), .ZN(new_n27416_));
  NOR2_X1    g24193(.A1(new_n27416_), .A2(new_n13855_), .ZN(new_n27417_));
  OAI21_X1   g24194(.A1(new_n27413_), .A2(new_n27414_), .B(new_n27417_), .ZN(new_n27418_));
  NAND3_X1   g24195(.A1(new_n27418_), .A2(new_n27415_), .A3(pi0781), .ZN(new_n27419_));
  NAND2_X1   g24196(.A1(new_n27419_), .A2(new_n27412_), .ZN(new_n27420_));
  NAND3_X1   g24197(.A1(new_n27420_), .A2(pi0619), .A3(pi1159), .ZN(new_n27421_));
  NAND4_X1   g24198(.A1(new_n27419_), .A2(new_n27412_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n27422_));
  AOI21_X1   g24199(.A1(new_n27421_), .A2(new_n27422_), .B(new_n27330_), .ZN(new_n27423_));
  OAI21_X1   g24200(.A1(new_n27423_), .A2(new_n20003_), .B(new_n27292_), .ZN(new_n27424_));
  AOI21_X1   g24201(.A1(new_n27288_), .A2(pi1159), .B(new_n13904_), .ZN(new_n27425_));
  NOR4_X1    g24202(.A1(new_n27287_), .A2(pi0619), .A3(new_n13868_), .A4(new_n27284_), .ZN(new_n27426_));
  OAI21_X1   g24203(.A1(new_n27425_), .A2(new_n27426_), .B(new_n27254_), .ZN(new_n27427_));
  NOR4_X1    g24204(.A1(new_n27291_), .A2(new_n27427_), .A3(new_n13896_), .A4(new_n27288_), .ZN(new_n27428_));
  NAND2_X1   g24205(.A1(new_n27291_), .A2(pi0789), .ZN(new_n27429_));
  OAI21_X1   g24206(.A1(new_n27287_), .A2(new_n27284_), .B(pi0789), .ZN(new_n27430_));
  NOR2_X1    g24207(.A1(new_n27427_), .A2(new_n27430_), .ZN(new_n27431_));
  NOR2_X1    g24208(.A1(new_n27431_), .A2(new_n27429_), .ZN(new_n27432_));
  NOR2_X1    g24209(.A1(new_n27432_), .A2(new_n27428_), .ZN(new_n27433_));
  AOI21_X1   g24210(.A1(new_n27433_), .A2(new_n13963_), .B(new_n19028_), .ZN(new_n27434_));
  NOR4_X1    g24211(.A1(new_n27432_), .A2(pi0626), .A3(new_n19208_), .A4(new_n27428_), .ZN(new_n27435_));
  OAI21_X1   g24212(.A1(new_n27434_), .A2(new_n27435_), .B(new_n27254_), .ZN(new_n27436_));
  AOI21_X1   g24213(.A1(new_n27433_), .A2(new_n13962_), .B(new_n18976_), .ZN(new_n27437_));
  NOR4_X1    g24214(.A1(new_n27432_), .A2(pi0626), .A3(new_n18974_), .A4(new_n27428_), .ZN(new_n27438_));
  OAI21_X1   g24215(.A1(new_n27437_), .A2(new_n27438_), .B(new_n27254_), .ZN(new_n27439_));
  NOR2_X1    g24216(.A1(new_n27264_), .A2(new_n13919_), .ZN(new_n27440_));
  AOI21_X1   g24217(.A1(new_n27330_), .A2(new_n13919_), .B(new_n27440_), .ZN(new_n27441_));
  OR2_X2     g24218(.A1(new_n27441_), .A2(new_n14162_), .Z(new_n27442_));
  AOI21_X1   g24219(.A1(new_n27436_), .A2(new_n27439_), .B(new_n27442_), .ZN(new_n27443_));
  NAND2_X1   g24220(.A1(new_n16424_), .A2(new_n14143_), .ZN(new_n27444_));
  AOI21_X1   g24221(.A1(new_n27420_), .A2(new_n13896_), .B(new_n27444_), .ZN(new_n27445_));
  OAI21_X1   g24222(.A1(new_n27443_), .A2(new_n13937_), .B(new_n27445_), .ZN(new_n27446_));
  NOR2_X1    g24223(.A1(new_n27413_), .A2(new_n27414_), .ZN(new_n27447_));
  NOR4_X1    g24224(.A1(new_n27447_), .A2(new_n13855_), .A3(new_n27405_), .A4(new_n27416_), .ZN(new_n27448_));
  AOI21_X1   g24225(.A1(new_n27399_), .A2(new_n27390_), .B(new_n27405_), .ZN(new_n27449_));
  INV_X1     g24226(.I(new_n27417_), .ZN(new_n27450_));
  AOI21_X1   g24227(.A1(new_n27399_), .A2(new_n27390_), .B(new_n27450_), .ZN(new_n27451_));
  NOR3_X1    g24228(.A1(new_n27449_), .A2(new_n27451_), .A3(new_n13855_), .ZN(new_n27452_));
  NOR3_X1    g24229(.A1(new_n27452_), .A2(new_n27448_), .A3(new_n13860_), .ZN(new_n27453_));
  NOR2_X1    g24230(.A1(new_n27453_), .A2(new_n13904_), .ZN(new_n27454_));
  NOR3_X1    g24231(.A1(new_n27420_), .A2(new_n13860_), .A3(pi1159), .ZN(new_n27455_));
  NOR2_X1    g24232(.A1(new_n27454_), .A2(new_n27455_), .ZN(new_n27456_));
  AND2_X2    g24233(.A1(new_n27427_), .A2(new_n13884_), .Z(new_n27457_));
  OAI21_X1   g24234(.A1(new_n27456_), .A2(new_n27330_), .B(new_n27457_), .ZN(new_n27458_));
  AOI21_X1   g24235(.A1(new_n27446_), .A2(new_n27424_), .B(new_n27458_), .ZN(new_n27459_));
  NOR2_X1    g24236(.A1(new_n27254_), .A2(new_n13966_), .ZN(new_n27460_));
  AOI21_X1   g24237(.A1(new_n27441_), .A2(new_n13966_), .B(new_n27460_), .ZN(new_n27461_));
  AOI21_X1   g24238(.A1(new_n27461_), .A2(pi0628), .B(new_n13971_), .ZN(new_n27462_));
  INV_X1     g24239(.I(new_n27460_), .ZN(new_n27463_));
  INV_X1     g24240(.I(new_n27440_), .ZN(new_n27464_));
  INV_X1     g24241(.I(new_n27293_), .ZN(new_n27465_));
  INV_X1     g24242(.I(new_n27294_), .ZN(new_n27466_));
  INV_X1     g24243(.I(new_n27324_), .ZN(new_n27467_));
  NAND3_X1   g24244(.A1(new_n27358_), .A2(pi0778), .A3(new_n27317_), .ZN(new_n27468_));
  NAND3_X1   g24245(.A1(new_n27468_), .A2(pi0778), .A3(new_n27319_), .ZN(new_n27469_));
  NAND3_X1   g24246(.A1(new_n27469_), .A2(new_n27467_), .A3(new_n13805_), .ZN(new_n27470_));
  NAND3_X1   g24247(.A1(new_n27470_), .A2(new_n13880_), .A3(new_n27466_), .ZN(new_n27471_));
  NAND3_X1   g24248(.A1(new_n27471_), .A2(new_n13919_), .A3(new_n27465_), .ZN(new_n27472_));
  NAND3_X1   g24249(.A1(new_n27472_), .A2(new_n13966_), .A3(new_n27464_), .ZN(new_n27473_));
  NAND2_X1   g24250(.A1(new_n27473_), .A2(new_n27463_), .ZN(new_n27474_));
  NOR3_X1    g24251(.A1(new_n27474_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n27475_));
  OAI21_X1   g24252(.A1(new_n27475_), .A2(new_n27462_), .B(new_n27254_), .ZN(new_n27476_));
  NAND2_X1   g24253(.A1(new_n27476_), .A2(pi0792), .ZN(new_n27477_));
  AOI21_X1   g24254(.A1(new_n27461_), .A2(pi1156), .B(new_n13971_), .ZN(new_n27478_));
  NOR3_X1    g24255(.A1(new_n27474_), .A2(pi0628), .A3(new_n13969_), .ZN(new_n27479_));
  OAI21_X1   g24256(.A1(new_n27479_), .A2(new_n27478_), .B(new_n27254_), .ZN(new_n27480_));
  NOR3_X1    g24257(.A1(new_n27480_), .A2(new_n12777_), .A3(new_n27461_), .ZN(new_n27481_));
  NAND2_X1   g24258(.A1(new_n27481_), .A2(new_n27477_), .ZN(new_n27482_));
  NAND3_X1   g24259(.A1(new_n27474_), .A2(pi0628), .A3(pi1156), .ZN(new_n27483_));
  NAND3_X1   g24260(.A1(new_n27461_), .A2(new_n13942_), .A3(pi1156), .ZN(new_n27484_));
  AOI21_X1   g24261(.A1(new_n27483_), .A2(new_n27484_), .B(new_n27264_), .ZN(new_n27485_));
  NAND3_X1   g24262(.A1(new_n27485_), .A2(pi0792), .A3(new_n27474_), .ZN(new_n27486_));
  NAND3_X1   g24263(.A1(new_n27486_), .A2(pi0792), .A3(new_n27476_), .ZN(new_n27487_));
  NAND2_X1   g24264(.A1(new_n27487_), .A2(new_n27482_), .ZN(new_n27488_));
  NOR2_X1    g24265(.A1(new_n27254_), .A2(pi0647), .ZN(new_n27489_));
  AOI21_X1   g24266(.A1(new_n27488_), .A2(pi0647), .B(new_n27489_), .ZN(new_n27490_));
  NOR4_X1    g24267(.A1(new_n27476_), .A2(new_n27480_), .A3(new_n12777_), .A4(new_n27461_), .ZN(new_n27491_));
  NOR2_X1    g24268(.A1(new_n27481_), .A2(new_n27477_), .ZN(new_n27492_));
  NOR2_X1    g24269(.A1(new_n27492_), .A2(new_n27491_), .ZN(new_n27493_));
  AOI21_X1   g24270(.A1(new_n27493_), .A2(pi0647), .B(new_n14008_), .ZN(new_n27494_));
  NOR3_X1    g24271(.A1(new_n27488_), .A2(new_n14005_), .A3(new_n14007_), .ZN(new_n27495_));
  OAI21_X1   g24272(.A1(new_n27495_), .A2(new_n27494_), .B(new_n27254_), .ZN(new_n27496_));
  NOR4_X1    g24273(.A1(new_n27496_), .A2(new_n14010_), .A3(new_n14006_), .A4(new_n27490_), .ZN(new_n27497_));
  NAND2_X1   g24274(.A1(new_n27490_), .A2(pi0630), .ZN(new_n27498_));
  NAND3_X1   g24275(.A1(new_n27488_), .A2(pi0647), .A3(pi1157), .ZN(new_n27499_));
  NAND3_X1   g24276(.A1(new_n27493_), .A2(pi0647), .A3(new_n14008_), .ZN(new_n27500_));
  AOI21_X1   g24277(.A1(new_n27499_), .A2(new_n27500_), .B(new_n27264_), .ZN(new_n27501_));
  AOI21_X1   g24278(.A1(new_n27501_), .A2(new_n14011_), .B(new_n27498_), .ZN(new_n27502_));
  OAI21_X1   g24279(.A1(new_n27497_), .A2(new_n27502_), .B(pi0787), .ZN(new_n27503_));
  NOR2_X1    g24280(.A1(new_n27433_), .A2(new_n14142_), .ZN(new_n27504_));
  AOI21_X1   g24281(.A1(new_n14142_), .A2(new_n27264_), .B(new_n27504_), .ZN(new_n27505_));
  NOR2_X1    g24282(.A1(new_n27505_), .A2(new_n13993_), .ZN(new_n27506_));
  NOR2_X1    g24283(.A1(new_n27254_), .A2(new_n13994_), .ZN(new_n27507_));
  OAI21_X1   g24284(.A1(new_n27506_), .A2(new_n27507_), .B(new_n16574_), .ZN(new_n27508_));
  AOI21_X1   g24285(.A1(new_n27503_), .A2(new_n16867_), .B(new_n27508_), .ZN(new_n27509_));
  AND2_X2    g24286(.A1(new_n27476_), .A2(pi0629), .Z(new_n27510_));
  NOR2_X1    g24287(.A1(new_n27485_), .A2(pi0629), .ZN(new_n27511_));
  OAI21_X1   g24288(.A1(new_n27510_), .A2(new_n27511_), .B(pi0792), .ZN(new_n27512_));
  AOI21_X1   g24289(.A1(new_n16875_), .A2(new_n27512_), .B(new_n27505_), .ZN(new_n27513_));
  OAI21_X1   g24290(.A1(new_n27509_), .A2(new_n27459_), .B(new_n27513_), .ZN(new_n27514_));
  AOI21_X1   g24291(.A1(new_n27490_), .A2(pi1157), .B(new_n12776_), .ZN(new_n27515_));
  AOI22_X1   g24292(.A1(new_n27496_), .A2(new_n27515_), .B1(new_n12776_), .B2(new_n27488_), .ZN(new_n27516_));
  OAI21_X1   g24293(.A1(new_n27506_), .A2(new_n27507_), .B(new_n14211_), .ZN(new_n27517_));
  NOR2_X1    g24294(.A1(new_n27254_), .A2(new_n14211_), .ZN(new_n27518_));
  INV_X1     g24295(.I(new_n27518_), .ZN(new_n27519_));
  NAND2_X1   g24296(.A1(pi0644), .A2(pi0715), .ZN(new_n27520_));
  AOI21_X1   g24297(.A1(new_n27517_), .A2(new_n27519_), .B(new_n27520_), .ZN(new_n27521_));
  AOI21_X1   g24298(.A1(new_n27521_), .A2(new_n27516_), .B(pi0644), .ZN(new_n27522_));
  NOR4_X1    g24299(.A1(new_n27514_), .A2(new_n14204_), .A3(new_n12775_), .A4(new_n27522_), .ZN(new_n27527_));
  OAI21_X1   g24300(.A1(new_n27514_), .A2(new_n27522_), .B(pi0790), .ZN(new_n27528_));
  INV_X1     g24301(.I(new_n19379_), .ZN(new_n27529_));
  NOR2_X1    g24302(.A1(new_n27514_), .A2(new_n27529_), .ZN(new_n27530_));
  NOR2_X1    g24303(.A1(new_n27528_), .A2(new_n27530_), .ZN(new_n27531_));
  OAI21_X1   g24304(.A1(new_n27531_), .A2(new_n27527_), .B(new_n7240_), .ZN(new_n27532_));
  NAND2_X1   g24305(.A1(po1038), .A2(pi0200), .ZN(new_n27533_));
  NAND2_X1   g24306(.A1(new_n27532_), .A2(new_n27533_), .ZN(po0357));
  NOR2_X1    g24307(.A1(pi0032), .A2(pi0070), .ZN(new_n27535_));
  AOI21_X1   g24308(.A1(new_n27535_), .A2(new_n2955_), .B(new_n2755_), .ZN(new_n27536_));
  NOR3_X1    g24309(.A1(new_n2794_), .A2(pi0070), .A3(pi0841), .ZN(new_n27537_));
  AOI21_X1   g24310(.A1(new_n2794_), .A2(pi0070), .B(new_n27537_), .ZN(new_n27538_));
  OAI21_X1   g24311(.A1(new_n27538_), .A2(pi0210), .B(new_n27536_), .ZN(new_n27539_));
  NAND3_X1   g24312(.A1(new_n27539_), .A2(new_n2777_), .A3(new_n2955_), .ZN(new_n27540_));
  NAND2_X1   g24313(.A1(new_n27540_), .A2(pi0096), .ZN(new_n27541_));
  NOR2_X1    g24314(.A1(new_n27541_), .A2(new_n5373_), .ZN(new_n27542_));
  NAND2_X1   g24315(.A1(new_n27541_), .A2(pi0947), .ZN(new_n27543_));
  NAND2_X1   g24316(.A1(new_n5383_), .A2(pi0947), .ZN(new_n27544_));
  XNOR2_X1   g24317(.A1(new_n27543_), .A2(new_n27544_), .ZN(new_n27545_));
  NOR2_X1    g24318(.A1(new_n5383_), .A2(pi0332), .ZN(new_n27546_));
  NOR2_X1    g24319(.A1(new_n27546_), .A2(pi0947), .ZN(new_n27547_));
  NOR2_X1    g24320(.A1(new_n27539_), .A2(pi0468), .ZN(new_n27548_));
  NOR2_X1    g24321(.A1(new_n9439_), .A2(pi0332), .ZN(new_n27549_));
  OAI21_X1   g24322(.A1(new_n27548_), .A2(new_n27549_), .B(new_n27547_), .ZN(new_n27550_));
  OAI21_X1   g24323(.A1(new_n27545_), .A2(new_n27550_), .B(new_n5796_), .ZN(new_n27551_));
  NAND2_X1   g24324(.A1(new_n27551_), .A2(new_n27542_), .ZN(new_n27552_));
  INV_X1     g24325(.I(new_n27552_), .ZN(new_n27553_));
  OAI21_X1   g24326(.A1(pi0070), .A2(pi0841), .B(pi0032), .ZN(new_n27554_));
  NAND3_X1   g24327(.A1(new_n2959_), .A2(new_n2436_), .A3(new_n27554_), .ZN(new_n27555_));
  NOR2_X1    g24328(.A1(new_n27538_), .A2(new_n2474_), .ZN(new_n27556_));
  AOI21_X1   g24329(.A1(new_n2697_), .A2(new_n27556_), .B(new_n27555_), .ZN(new_n27557_));
  OAI21_X1   g24330(.A1(new_n2855_), .A2(pi0095), .B(new_n2707_), .ZN(new_n27558_));
  NOR2_X1    g24331(.A1(pi0032), .A2(pi0096), .ZN(new_n27559_));
  NAND2_X1   g24332(.A1(new_n27558_), .A2(new_n27559_), .ZN(new_n27560_));
  AOI21_X1   g24333(.A1(new_n2777_), .A2(new_n2955_), .B(new_n2755_), .ZN(new_n27562_));
  INV_X1     g24334(.I(new_n27562_), .ZN(new_n27563_));
  NOR2_X1    g24335(.A1(new_n27563_), .A2(new_n5373_), .ZN(new_n27564_));
  NOR2_X1    g24336(.A1(new_n27562_), .A2(new_n5800_), .ZN(new_n27565_));
  XNOR2_X1   g24337(.A1(new_n27544_), .A2(new_n27565_), .ZN(new_n27566_));
  INV_X1     g24338(.I(new_n27549_), .ZN(new_n27567_));
  NAND2_X1   g24339(.A1(new_n27560_), .A2(pi0210), .ZN(new_n27568_));
  NAND2_X1   g24340(.A1(pi0210), .A2(pi0332), .ZN(new_n27569_));
  XOR2_X1    g24341(.A1(new_n27568_), .A2(new_n27569_), .Z(new_n27570_));
  NAND3_X1   g24342(.A1(new_n27570_), .A2(new_n9439_), .A3(new_n27557_), .ZN(new_n27571_));
  NAND2_X1   g24343(.A1(new_n27571_), .A2(new_n27567_), .ZN(new_n27572_));
  AND3_X2    g24344(.A1(new_n27572_), .A2(new_n27547_), .A3(new_n27566_), .Z(new_n27573_));
  OAI21_X1   g24345(.A1(new_n27573_), .A2(new_n5383_), .B(new_n27564_), .ZN(new_n27574_));
  NAND2_X1   g24346(.A1(new_n27574_), .A2(new_n3291_), .ZN(new_n27575_));
  OAI21_X1   g24347(.A1(new_n3291_), .A2(new_n27553_), .B(new_n27575_), .ZN(new_n27576_));
  NOR2_X1    g24348(.A1(new_n27576_), .A2(new_n3229_), .ZN(new_n27577_));
  NAND2_X1   g24349(.A1(new_n9163_), .A2(pi0059), .ZN(new_n27578_));
  XNOR2_X1   g24350(.A1(new_n27577_), .A2(new_n27578_), .ZN(new_n27579_));
  AOI21_X1   g24351(.A1(new_n27579_), .A2(new_n27553_), .B(new_n5371_), .ZN(new_n27580_));
  NAND2_X1   g24352(.A1(new_n27574_), .A2(new_n12116_), .ZN(new_n27581_));
  NAND2_X1   g24353(.A1(new_n12116_), .A2(pi0299), .ZN(new_n27582_));
  XOR2_X1    g24354(.A1(new_n27581_), .A2(new_n27582_), .Z(new_n27583_));
  NOR2_X1    g24355(.A1(new_n2755_), .A2(new_n3072_), .ZN(new_n27584_));
  INV_X1     g24356(.I(new_n27584_), .ZN(new_n27585_));
  NOR2_X1    g24357(.A1(new_n27585_), .A2(new_n2955_), .ZN(new_n27586_));
  INV_X1     g24358(.I(new_n27586_), .ZN(new_n27587_));
  NOR2_X1    g24359(.A1(new_n27538_), .A2(new_n2795_), .ZN(new_n27588_));
  AOI21_X1   g24360(.A1(new_n2905_), .A2(new_n27588_), .B(new_n27555_), .ZN(new_n27589_));
  NAND2_X1   g24361(.A1(pi0198), .A2(pi0332), .ZN(new_n27590_));
  NAND3_X1   g24362(.A1(new_n2734_), .A2(pi0070), .A3(pi0095), .ZN(new_n27591_));
  NOR4_X1    g24363(.A1(new_n2905_), .A2(new_n2796_), .A3(new_n27559_), .A4(new_n27591_), .ZN(new_n27592_));
  NOR2_X1    g24364(.A1(new_n27592_), .A2(new_n3072_), .ZN(new_n27593_));
  XNOR2_X1   g24365(.A1(new_n27593_), .A2(new_n27590_), .ZN(new_n27594_));
  NAND2_X1   g24366(.A1(new_n27594_), .A2(new_n27589_), .ZN(new_n27595_));
  AND3_X2    g24367(.A1(new_n27595_), .A2(new_n5383_), .A3(new_n27587_), .Z(new_n27599_));
  NOR2_X1    g24368(.A1(new_n27592_), .A2(new_n2777_), .ZN(new_n27600_));
  XNOR2_X1   g24369(.A1(new_n27600_), .A2(new_n27569_), .ZN(new_n27601_));
  NAND3_X1   g24370(.A1(new_n27601_), .A2(new_n9439_), .A3(new_n27589_), .ZN(new_n27602_));
  NAND2_X1   g24371(.A1(new_n27602_), .A2(new_n27567_), .ZN(new_n27603_));
  OAI21_X1   g24372(.A1(pi0210), .A2(pi0332), .B(pi0096), .ZN(new_n27604_));
  NAND2_X1   g24373(.A1(new_n27604_), .A2(pi0947), .ZN(new_n27605_));
  XOR2_X1    g24374(.A1(new_n27544_), .A2(new_n27605_), .Z(new_n27606_));
  NOR2_X1    g24375(.A1(new_n27604_), .A2(new_n5373_), .ZN(new_n27607_));
  OAI21_X1   g24376(.A1(new_n5796_), .A2(new_n27607_), .B(new_n27547_), .ZN(new_n27608_));
  NAND3_X1   g24377(.A1(new_n27608_), .A2(pi0299), .A3(new_n6325_), .ZN(new_n27609_));
  AOI21_X1   g24378(.A1(new_n27603_), .A2(new_n27606_), .B(new_n27609_), .ZN(new_n27610_));
  NAND2_X1   g24379(.A1(new_n27595_), .A2(new_n27587_), .ZN(new_n27611_));
  NOR3_X1    g24380(.A1(new_n27546_), .A2(pi0587), .A3(new_n5796_), .ZN(new_n27612_));
  INV_X1     g24381(.I(new_n27612_), .ZN(new_n27613_));
  AOI21_X1   g24382(.A1(new_n27611_), .A2(new_n27613_), .B(new_n5386_), .ZN(new_n27614_));
  OAI21_X1   g24383(.A1(new_n27610_), .A2(new_n27599_), .B(new_n27614_), .ZN(new_n27615_));
  OAI21_X1   g24384(.A1(new_n27538_), .A2(pi0198), .B(new_n27536_), .ZN(new_n27616_));
  OR3_X2     g24385(.A1(new_n5807_), .A2(new_n27546_), .A3(new_n27616_), .Z(new_n27617_));
  NOR2_X1    g24386(.A1(new_n3196_), .A2(pi0074), .ZN(new_n27618_));
  NAND3_X1   g24387(.A1(new_n27618_), .A2(pi0587), .A3(new_n5373_), .ZN(new_n27619_));
  AOI21_X1   g24388(.A1(new_n27617_), .A2(new_n3098_), .B(new_n27619_), .ZN(new_n27620_));
  NAND2_X1   g24389(.A1(new_n27616_), .A2(new_n27587_), .ZN(new_n27621_));
  NOR2_X1    g24390(.A1(new_n27621_), .A2(new_n3258_), .ZN(new_n27622_));
  OAI21_X1   g24391(.A1(new_n27620_), .A2(new_n5383_), .B(new_n27622_), .ZN(new_n27623_));
  AOI21_X1   g24392(.A1(new_n27623_), .A2(new_n3098_), .B(new_n3175_), .ZN(new_n27624_));
  NAND2_X1   g24393(.A1(new_n27553_), .A2(new_n27624_), .ZN(new_n27625_));
  NAND2_X1   g24394(.A1(new_n27560_), .A2(pi0198), .ZN(new_n27626_));
  XOR2_X1    g24395(.A1(new_n27626_), .A2(new_n27590_), .Z(new_n27627_));
  NAND2_X1   g24396(.A1(new_n27627_), .A2(new_n27557_), .ZN(new_n27628_));
  AOI21_X1   g24397(.A1(new_n27627_), .A2(new_n27557_), .B(new_n27586_), .ZN(new_n27629_));
  NAND3_X1   g24398(.A1(new_n27628_), .A2(new_n5383_), .A3(new_n27587_), .ZN(new_n27632_));
  AOI21_X1   g24399(.A1(new_n27615_), .A2(new_n27625_), .B(new_n27632_), .ZN(new_n27633_));
  NAND2_X1   g24400(.A1(new_n27583_), .A2(new_n27633_), .ZN(new_n27634_));
  NAND2_X1   g24401(.A1(new_n27576_), .A2(pi0055), .ZN(new_n27635_));
  AOI21_X1   g24402(.A1(new_n27634_), .A2(new_n3226_), .B(new_n27635_), .ZN(new_n27636_));
  NOR3_X1    g24403(.A1(new_n27552_), .A2(new_n5371_), .A3(new_n3226_), .ZN(new_n27637_));
  OAI21_X1   g24404(.A1(new_n27636_), .A2(pi0059), .B(new_n27637_), .ZN(new_n27638_));
  INV_X1     g24405(.I(pi0233), .ZN(new_n27639_));
  INV_X1     g24406(.I(pi0237), .ZN(new_n27640_));
  NOR2_X1    g24407(.A1(new_n27639_), .A2(new_n27640_), .ZN(new_n27641_));
  OAI21_X1   g24408(.A1(new_n27580_), .A2(new_n27638_), .B(new_n27641_), .ZN(new_n27642_));
  AOI21_X1   g24409(.A1(new_n27580_), .A2(new_n27638_), .B(new_n27642_), .ZN(new_n27643_));
  NAND3_X1   g24410(.A1(new_n3145_), .A2(new_n2955_), .A3(new_n5798_), .ZN(new_n27644_));
  AOI21_X1   g24411(.A1(new_n27644_), .A2(new_n3291_), .B(new_n3229_), .ZN(new_n27645_));
  XNOR2_X1   g24412(.A1(new_n27645_), .A2(new_n27578_), .ZN(new_n27646_));
  AOI21_X1   g24413(.A1(new_n27646_), .A2(pi0332), .B(new_n5371_), .ZN(new_n27647_));
  NOR3_X1    g24414(.A1(new_n3145_), .A2(new_n3098_), .A3(new_n5798_), .ZN(new_n27648_));
  NOR3_X1    g24415(.A1(new_n3145_), .A2(pi0299), .A3(new_n5802_), .ZN(new_n27649_));
  OAI21_X1   g24416(.A1(new_n27648_), .A2(new_n27649_), .B(new_n5809_), .ZN(new_n27650_));
  INV_X1     g24417(.I(new_n6325_), .ZN(new_n27651_));
  NOR4_X1    g24418(.A1(new_n27651_), .A2(new_n3196_), .A3(pi0054), .A4(pi0332), .ZN(new_n27652_));
  AOI21_X1   g24419(.A1(new_n27650_), .A2(new_n27652_), .B(pi0332), .ZN(new_n27653_));
  NOR2_X1    g24420(.A1(pi0299), .A2(pi0587), .ZN(new_n27654_));
  NOR2_X1    g24421(.A1(new_n2905_), .A2(new_n9173_), .ZN(new_n27655_));
  NAND3_X1   g24422(.A1(new_n27655_), .A2(pi0468), .A3(new_n5383_), .ZN(new_n27656_));
  NAND3_X1   g24423(.A1(new_n27655_), .A2(new_n9439_), .A3(new_n5796_), .ZN(new_n27657_));
  NAND2_X1   g24424(.A1(new_n27656_), .A2(new_n27657_), .ZN(new_n27658_));
  OAI21_X1   g24425(.A1(new_n17067_), .A2(new_n27654_), .B(new_n27658_), .ZN(new_n27659_));
  OAI21_X1   g24426(.A1(new_n27659_), .A2(new_n27653_), .B(pi0074), .ZN(new_n27660_));
  XOR2_X1    g24427(.A1(new_n27660_), .A2(new_n6327_), .Z(new_n27661_));
  OAI21_X1   g24428(.A1(new_n27661_), .A2(new_n2955_), .B(new_n3226_), .ZN(new_n27662_));
  NAND4_X1   g24429(.A1(new_n27662_), .A2(pi0055), .A3(new_n3291_), .A4(new_n27644_), .ZN(new_n27663_));
  NOR3_X1    g24430(.A1(new_n3226_), .A2(new_n5371_), .A3(new_n2955_), .ZN(new_n27664_));
  INV_X1     g24431(.I(new_n27664_), .ZN(new_n27665_));
  AOI21_X1   g24432(.A1(new_n27663_), .A2(new_n3229_), .B(new_n27665_), .ZN(new_n27666_));
  XOR2_X1    g24433(.A1(new_n27666_), .A2(new_n27647_), .Z(new_n27667_));
  NAND2_X1   g24434(.A1(new_n27667_), .A2(new_n27641_), .ZN(new_n27668_));
  XOR2_X1    g24435(.A1(new_n27643_), .A2(new_n27668_), .Z(new_n27669_));
  INV_X1     g24436(.I(new_n27641_), .ZN(new_n27670_));
  OAI21_X1   g24437(.A1(new_n12655_), .A2(new_n5798_), .B(new_n27585_), .ZN(new_n27672_));
  NAND2_X1   g24438(.A1(new_n27672_), .A2(new_n5809_), .ZN(new_n27673_));
  NOR2_X1    g24439(.A1(new_n27673_), .A2(new_n27670_), .ZN(new_n27674_));
  NAND2_X1   g24440(.A1(new_n27674_), .A2(pi0201), .ZN(new_n27675_));
  OAI21_X1   g24441(.A1(new_n27669_), .A2(pi0201), .B(new_n27675_), .ZN(po0358));
  INV_X1     g24442(.I(new_n27673_), .ZN(new_n27677_));
  NOR2_X1    g24443(.A1(new_n27640_), .A2(pi0233), .ZN(new_n27678_));
  NAND2_X1   g24444(.A1(new_n27677_), .A2(new_n27678_), .ZN(new_n27679_));
  INV_X1     g24445(.I(new_n27679_), .ZN(new_n27680_));
  NAND2_X1   g24446(.A1(new_n27680_), .A2(pi0202), .ZN(new_n27681_));
  OAI21_X1   g24447(.A1(new_n27669_), .A2(pi0202), .B(new_n27681_), .ZN(po0359));
  NOR3_X1    g24448(.A1(new_n27673_), .A2(pi0233), .A3(pi0237), .ZN(new_n27683_));
  NAND2_X1   g24449(.A1(new_n27683_), .A2(pi0203), .ZN(new_n27684_));
  OAI21_X1   g24450(.A1(new_n27669_), .A2(pi0203), .B(new_n27684_), .ZN(po0360));
  NAND2_X1   g24451(.A1(new_n27541_), .A2(pi0907), .ZN(new_n27686_));
  NOR2_X1    g24452(.A1(new_n5636_), .A2(new_n5741_), .ZN(new_n27687_));
  XOR2_X1    g24453(.A1(new_n27686_), .A2(new_n27687_), .Z(new_n27688_));
  AOI21_X1   g24454(.A1(new_n5636_), .A2(new_n2955_), .B(pi0907), .ZN(new_n27689_));
  OAI21_X1   g24455(.A1(new_n27548_), .A2(new_n27549_), .B(new_n27689_), .ZN(new_n27690_));
  OAI21_X1   g24456(.A1(new_n27688_), .A2(new_n27690_), .B(new_n5636_), .ZN(new_n27691_));
  NAND2_X1   g24457(.A1(new_n27691_), .A2(new_n27542_), .ZN(new_n27692_));
  INV_X1     g24458(.I(new_n27692_), .ZN(new_n27693_));
  NOR2_X1    g24459(.A1(new_n27562_), .A2(new_n5741_), .ZN(new_n27694_));
  XOR2_X1    g24460(.A1(new_n27687_), .A2(new_n27694_), .Z(new_n27695_));
  OAI21_X1   g24461(.A1(new_n27563_), .A2(new_n5373_), .B(new_n5375_), .ZN(new_n27696_));
  NOR2_X1    g24462(.A1(new_n12845_), .A2(new_n2955_), .ZN(new_n27697_));
  NAND2_X1   g24463(.A1(new_n27697_), .A2(new_n27696_), .ZN(new_n27698_));
  AOI22_X1   g24464(.A1(new_n27572_), .A2(new_n27695_), .B1(new_n27689_), .B2(new_n27698_), .ZN(new_n27699_));
  NAND2_X1   g24465(.A1(new_n27692_), .A2(new_n3292_), .ZN(new_n27700_));
  OAI21_X1   g24466(.A1(new_n27699_), .A2(new_n3292_), .B(new_n27700_), .ZN(new_n27701_));
  NOR2_X1    g24467(.A1(new_n27701_), .A2(new_n3229_), .ZN(new_n27702_));
  XNOR2_X1   g24468(.A1(new_n27702_), .A2(new_n27578_), .ZN(new_n27703_));
  AOI21_X1   g24469(.A1(new_n27703_), .A2(new_n27693_), .B(new_n5371_), .ZN(new_n27704_));
  NAND2_X1   g24470(.A1(new_n27604_), .A2(pi0907), .ZN(new_n27705_));
  XOR2_X1    g24471(.A1(new_n27687_), .A2(new_n27705_), .Z(new_n27706_));
  AOI21_X1   g24472(.A1(new_n27602_), .A2(new_n27567_), .B(new_n27706_), .ZN(new_n27707_));
  AOI21_X1   g24473(.A1(new_n5378_), .A2(new_n27584_), .B(new_n2955_), .ZN(new_n27708_));
  OAI21_X1   g24474(.A1(pi0299), .A2(new_n27708_), .B(new_n5555_), .ZN(new_n27709_));
  OAI21_X1   g24475(.A1(new_n27611_), .A2(new_n27709_), .B(new_n3098_), .ZN(new_n27710_));
  NOR2_X1    g24476(.A1(new_n5636_), .A2(new_n27607_), .ZN(new_n27711_));
  NAND2_X1   g24477(.A1(new_n12116_), .A2(new_n27689_), .ZN(new_n27712_));
  NOR2_X1    g24478(.A1(new_n27712_), .A2(new_n27711_), .ZN(new_n27713_));
  OAI21_X1   g24479(.A1(new_n27710_), .A2(new_n27707_), .B(new_n27713_), .ZN(new_n27714_));
  AOI21_X1   g24480(.A1(new_n27629_), .A2(new_n5555_), .B(new_n3098_), .ZN(new_n27715_));
  NAND3_X1   g24481(.A1(new_n27699_), .A2(pi0299), .A3(new_n27708_), .ZN(new_n27716_));
  XOR2_X1    g24482(.A1(new_n27716_), .A2(new_n27715_), .Z(new_n27717_));
  OAI21_X1   g24483(.A1(new_n27717_), .A2(new_n27651_), .B(new_n27714_), .ZN(new_n27718_));
  NAND2_X1   g24484(.A1(new_n27692_), .A2(pi0299), .ZN(new_n27719_));
  NAND2_X1   g24485(.A1(new_n27618_), .A2(pi0299), .ZN(new_n27720_));
  XNOR2_X1   g24486(.A1(new_n27719_), .A2(new_n27720_), .ZN(new_n27721_));
  NOR2_X1    g24487(.A1(pi0468), .A2(pi0602), .ZN(new_n27722_));
  AOI21_X1   g24488(.A1(new_n5636_), .A2(pi0468), .B(new_n27722_), .ZN(new_n27723_));
  INV_X1     g24489(.I(new_n27723_), .ZN(new_n27724_));
  NOR2_X1    g24490(.A1(new_n27724_), .A2(new_n27621_), .ZN(new_n27725_));
  OR3_X2     g24491(.A1(new_n27721_), .A2(new_n27708_), .A3(new_n27725_), .Z(new_n27726_));
  AOI21_X1   g24492(.A1(new_n27726_), .A2(new_n3258_), .B(new_n3175_), .ZN(new_n27727_));
  AOI21_X1   g24493(.A1(new_n27718_), .A2(new_n27727_), .B(new_n3225_), .ZN(new_n27728_));
  NAND2_X1   g24494(.A1(new_n27701_), .A2(pi0055), .ZN(new_n27729_));
  OAI21_X1   g24495(.A1(new_n27728_), .A2(new_n27729_), .B(new_n3229_), .ZN(new_n27730_));
  NAND4_X1   g24496(.A1(new_n27730_), .A2(pi0057), .A3(new_n3225_), .A4(new_n27693_), .ZN(new_n27731_));
  OAI21_X1   g24497(.A1(new_n27731_), .A2(new_n27704_), .B(new_n27641_), .ZN(new_n27732_));
  AOI21_X1   g24498(.A1(new_n27704_), .A2(new_n27731_), .B(new_n27732_), .ZN(new_n27733_));
  NAND3_X1   g24499(.A1(new_n5652_), .A2(new_n3145_), .A3(new_n2955_), .ZN(new_n27734_));
  NAND2_X1   g24500(.A1(new_n27734_), .A2(new_n3291_), .ZN(new_n27735_));
  NAND2_X1   g24501(.A1(new_n27735_), .A2(pi0059), .ZN(new_n27736_));
  XOR2_X1    g24502(.A1(new_n27736_), .A2(new_n27578_), .Z(new_n27737_));
  AOI21_X1   g24503(.A1(new_n27737_), .A2(pi0332), .B(new_n5371_), .ZN(new_n27738_));
  NOR3_X1    g24504(.A1(new_n5652_), .A2(new_n3145_), .A3(new_n3098_), .ZN(new_n27739_));
  NOR3_X1    g24505(.A1(new_n3145_), .A2(pi0299), .A3(new_n5656_), .ZN(new_n27740_));
  OAI21_X1   g24506(.A1(new_n27739_), .A2(new_n27740_), .B(new_n27724_), .ZN(new_n27741_));
  NAND2_X1   g24507(.A1(new_n12116_), .A2(new_n6325_), .ZN(new_n27742_));
  OAI21_X1   g24508(.A1(new_n27741_), .A2(new_n27742_), .B(new_n2955_), .ZN(new_n27743_));
  AOI21_X1   g24509(.A1(pi0055), .A2(pi0332), .B(new_n3195_), .ZN(new_n27744_));
  NOR3_X1    g24510(.A1(new_n27744_), .A2(new_n3175_), .A3(new_n3226_), .ZN(new_n27745_));
  OAI21_X1   g24511(.A1(new_n27735_), .A2(new_n3258_), .B(new_n27745_), .ZN(new_n27746_));
  NOR3_X1    g24512(.A1(new_n3098_), .A2(new_n9439_), .A3(new_n5741_), .ZN(new_n27747_));
  NOR3_X1    g24513(.A1(new_n3098_), .A2(pi0468), .A3(pi0907), .ZN(new_n27748_));
  NOR2_X1    g24514(.A1(new_n27747_), .A2(new_n27748_), .ZN(new_n27749_));
  NOR4_X1    g24515(.A1(new_n2905_), .A2(new_n5393_), .A3(new_n9173_), .A4(new_n27749_), .ZN(new_n27750_));
  OAI21_X1   g24516(.A1(new_n27750_), .A2(pi0468), .B(new_n5378_), .ZN(new_n27751_));
  AOI21_X1   g24517(.A1(new_n3175_), .A2(new_n27746_), .B(new_n27751_), .ZN(new_n27752_));
  NAND2_X1   g24518(.A1(new_n27752_), .A2(new_n27743_), .ZN(new_n27753_));
  AOI21_X1   g24519(.A1(new_n27753_), .A2(new_n3229_), .B(new_n27665_), .ZN(new_n27754_));
  XOR2_X1    g24520(.A1(new_n27754_), .A2(new_n27738_), .Z(new_n27755_));
  NAND2_X1   g24521(.A1(new_n27755_), .A2(new_n27641_), .ZN(new_n27756_));
  XOR2_X1    g24522(.A1(new_n27733_), .A2(new_n27756_), .Z(new_n27757_));
  OAI21_X1   g24523(.A1(new_n5652_), .A2(new_n12655_), .B(new_n27585_), .ZN(new_n27758_));
  NAND2_X1   g24524(.A1(new_n27758_), .A2(new_n5555_), .ZN(new_n27759_));
  NOR2_X1    g24525(.A1(new_n27759_), .A2(new_n27670_), .ZN(new_n27760_));
  NAND2_X1   g24526(.A1(new_n27760_), .A2(pi0204), .ZN(new_n27761_));
  OAI21_X1   g24527(.A1(new_n27757_), .A2(pi0204), .B(new_n27761_), .ZN(po0361));
  INV_X1     g24528(.I(new_n27759_), .ZN(new_n27763_));
  NAND3_X1   g24529(.A1(new_n27763_), .A2(pi0205), .A3(new_n27678_), .ZN(new_n27764_));
  OAI21_X1   g24530(.A1(new_n27757_), .A2(pi0205), .B(new_n27764_), .ZN(po0362));
  NOR2_X1    g24531(.A1(new_n27639_), .A2(pi0237), .ZN(new_n27766_));
  NAND3_X1   g24532(.A1(new_n27763_), .A2(pi0206), .A3(new_n27766_), .ZN(new_n27767_));
  OAI21_X1   g24533(.A1(new_n27757_), .A2(pi0206), .B(new_n27767_), .ZN(po0363));
  NAND2_X1   g24534(.A1(po1038), .A2(new_n8545_), .ZN(new_n27769_));
  NOR2_X1    g24535(.A1(new_n14428_), .A2(new_n13614_), .ZN(new_n27770_));
  XOR2_X1    g24536(.A1(new_n27770_), .A2(new_n13615_), .Z(new_n27771_));
  NOR2_X1    g24537(.A1(new_n15639_), .A2(new_n3290_), .ZN(new_n27772_));
  NAND2_X1   g24538(.A1(new_n27771_), .A2(new_n27772_), .ZN(new_n27773_));
  XOR2_X1    g24539(.A1(new_n19280_), .A2(new_n16146_), .Z(new_n27774_));
  NOR2_X1    g24540(.A1(new_n27774_), .A2(new_n3290_), .ZN(new_n27775_));
  NOR2_X1    g24541(.A1(new_n14428_), .A2(new_n13613_), .ZN(new_n27776_));
  XOR2_X1    g24542(.A1(new_n27776_), .A2(new_n13615_), .Z(new_n27777_));
  NAND2_X1   g24543(.A1(new_n27777_), .A2(new_n27775_), .ZN(new_n27778_));
  NAND3_X1   g24544(.A1(new_n27773_), .A2(new_n27778_), .A3(pi0608), .ZN(new_n27779_));
  NAND2_X1   g24545(.A1(new_n27779_), .A2(pi0778), .ZN(new_n27780_));
  INV_X1     g24546(.I(new_n27777_), .ZN(new_n27781_));
  NAND2_X1   g24547(.A1(new_n27771_), .A2(new_n27775_), .ZN(new_n27782_));
  NAND4_X1   g24548(.A1(new_n27782_), .A2(new_n27781_), .A3(new_n13749_), .A4(new_n27772_), .ZN(new_n27783_));
  INV_X1     g24549(.I(new_n27783_), .ZN(new_n27784_));
  XOR2_X1    g24550(.A1(new_n27780_), .A2(new_n27784_), .Z(new_n27785_));
  NAND4_X1   g24551(.A1(new_n27771_), .A2(new_n27777_), .A3(pi0778), .A4(new_n27775_), .ZN(new_n27786_));
  NAND3_X1   g24552(.A1(new_n27771_), .A2(pi0778), .A3(new_n27775_), .ZN(new_n27787_));
  NAND3_X1   g24553(.A1(new_n27787_), .A2(new_n27778_), .A3(pi0778), .ZN(new_n27788_));
  NAND2_X1   g24554(.A1(new_n27788_), .A2(new_n27786_), .ZN(new_n27789_));
  AOI21_X1   g24555(.A1(new_n27789_), .A2(new_n13766_), .B(new_n13783_), .ZN(new_n27790_));
  OAI21_X1   g24556(.A1(new_n27785_), .A2(new_n13766_), .B(new_n27790_), .ZN(new_n27791_));
  NAND2_X1   g24557(.A1(new_n27791_), .A2(new_n13784_), .ZN(new_n27792_));
  NAND2_X1   g24558(.A1(new_n27780_), .A2(new_n27784_), .ZN(new_n27793_));
  INV_X1     g24559(.I(new_n27793_), .ZN(new_n27794_));
  NOR2_X1    g24560(.A1(new_n27780_), .A2(new_n27784_), .ZN(new_n27795_));
  OAI21_X1   g24561(.A1(new_n27794_), .A2(new_n27795_), .B(pi0609), .ZN(new_n27796_));
  NAND3_X1   g24562(.A1(new_n27796_), .A2(new_n13785_), .A3(new_n27790_), .ZN(new_n27797_));
  AOI21_X1   g24563(.A1(new_n27792_), .A2(new_n27797_), .B(new_n13627_), .ZN(new_n27798_));
  INV_X1     g24564(.I(new_n27795_), .ZN(new_n27799_));
  AOI21_X1   g24565(.A1(new_n27799_), .A2(new_n27793_), .B(pi0609), .ZN(new_n27800_));
  AOI21_X1   g24566(.A1(new_n27789_), .A2(pi0609), .B(new_n13778_), .ZN(new_n27801_));
  INV_X1     g24567(.I(new_n27801_), .ZN(new_n27802_));
  OAI21_X1   g24568(.A1(new_n27800_), .A2(new_n27802_), .B(new_n13784_), .ZN(new_n27803_));
  OAI21_X1   g24569(.A1(new_n27794_), .A2(new_n27795_), .B(new_n13766_), .ZN(new_n27804_));
  NAND3_X1   g24570(.A1(new_n27804_), .A2(new_n13785_), .A3(new_n27801_), .ZN(new_n27805_));
  NOR2_X1    g24571(.A1(new_n13627_), .A2(new_n13801_), .ZN(new_n27806_));
  OAI21_X1   g24572(.A1(new_n27794_), .A2(new_n27795_), .B(new_n27806_), .ZN(new_n27807_));
  AOI21_X1   g24573(.A1(new_n27803_), .A2(new_n27805_), .B(new_n27807_), .ZN(new_n27808_));
  OAI21_X1   g24574(.A1(new_n27798_), .A2(new_n13801_), .B(new_n27808_), .ZN(new_n27809_));
  AOI21_X1   g24575(.A1(new_n27796_), .A2(new_n27790_), .B(new_n13785_), .ZN(new_n27810_));
  NOR2_X1    g24576(.A1(new_n27791_), .A2(new_n13784_), .ZN(new_n27811_));
  OAI21_X1   g24577(.A1(new_n27811_), .A2(new_n27810_), .B(new_n14428_), .ZN(new_n27812_));
  AOI21_X1   g24578(.A1(new_n27804_), .A2(new_n27801_), .B(new_n13785_), .ZN(new_n27813_));
  NOR3_X1    g24579(.A1(new_n27800_), .A2(new_n13784_), .A3(new_n27802_), .ZN(new_n27814_));
  INV_X1     g24580(.I(new_n27807_), .ZN(new_n27815_));
  OAI21_X1   g24581(.A1(new_n27814_), .A2(new_n27813_), .B(new_n27815_), .ZN(new_n27816_));
  NAND3_X1   g24582(.A1(new_n27812_), .A2(pi0785), .A3(new_n27816_), .ZN(new_n27817_));
  NAND3_X1   g24583(.A1(new_n27809_), .A2(new_n27817_), .A3(pi0618), .ZN(new_n27818_));
  NOR2_X1    g24584(.A1(new_n13627_), .A2(new_n13805_), .ZN(new_n27819_));
  AOI21_X1   g24585(.A1(new_n27789_), .A2(new_n13805_), .B(new_n27819_), .ZN(new_n27820_));
  INV_X1     g24586(.I(new_n27820_), .ZN(new_n27821_));
  AOI21_X1   g24587(.A1(new_n27821_), .A2(new_n13816_), .B(new_n13823_), .ZN(new_n27822_));
  AOI21_X1   g24588(.A1(new_n27818_), .A2(new_n27822_), .B(new_n14501_), .ZN(new_n27823_));
  AOI21_X1   g24589(.A1(new_n27812_), .A2(pi0785), .B(new_n27816_), .ZN(new_n27824_));
  NOR3_X1    g24590(.A1(new_n27798_), .A2(new_n27808_), .A3(new_n13801_), .ZN(new_n27825_));
  NOR3_X1    g24591(.A1(new_n27824_), .A2(new_n27825_), .A3(new_n13816_), .ZN(new_n27826_));
  INV_X1     g24592(.I(new_n27822_), .ZN(new_n27827_));
  NOR3_X1    g24593(.A1(new_n27826_), .A2(new_n13824_), .A3(new_n27827_), .ZN(new_n27828_));
  OAI21_X1   g24594(.A1(new_n27828_), .A2(new_n27823_), .B(new_n14428_), .ZN(new_n27829_));
  NAND3_X1   g24595(.A1(new_n27809_), .A2(new_n27817_), .A3(new_n13816_), .ZN(new_n27830_));
  AOI21_X1   g24596(.A1(new_n27821_), .A2(pi0618), .B(new_n13817_), .ZN(new_n27831_));
  AOI21_X1   g24597(.A1(new_n27830_), .A2(new_n27831_), .B(new_n14501_), .ZN(new_n27832_));
  NOR3_X1    g24598(.A1(new_n27824_), .A2(new_n27825_), .A3(pi0618), .ZN(new_n27833_));
  INV_X1     g24599(.I(new_n27831_), .ZN(new_n27834_));
  NOR3_X1    g24600(.A1(new_n27833_), .A2(new_n13824_), .A3(new_n27834_), .ZN(new_n27835_));
  NOR2_X1    g24601(.A1(new_n13627_), .A2(new_n13855_), .ZN(new_n27836_));
  OAI21_X1   g24602(.A1(new_n27824_), .A2(new_n27825_), .B(new_n27836_), .ZN(new_n27837_));
  INV_X1     g24603(.I(new_n27837_), .ZN(new_n27838_));
  OAI21_X1   g24604(.A1(new_n27835_), .A2(new_n27832_), .B(new_n27838_), .ZN(new_n27839_));
  AOI21_X1   g24605(.A1(pi0781), .A2(new_n27829_), .B(new_n27839_), .ZN(new_n27840_));
  OAI21_X1   g24606(.A1(new_n27826_), .A2(new_n27827_), .B(new_n13824_), .ZN(new_n27841_));
  NAND3_X1   g24607(.A1(new_n27818_), .A2(new_n14501_), .A3(new_n27822_), .ZN(new_n27842_));
  AOI21_X1   g24608(.A1(new_n27841_), .A2(new_n27842_), .B(new_n13627_), .ZN(new_n27843_));
  OAI21_X1   g24609(.A1(new_n27833_), .A2(new_n27834_), .B(new_n13824_), .ZN(new_n27844_));
  NAND3_X1   g24610(.A1(new_n27830_), .A2(new_n14501_), .A3(new_n27831_), .ZN(new_n27845_));
  AOI21_X1   g24611(.A1(new_n27844_), .A2(new_n27845_), .B(new_n27837_), .ZN(new_n27846_));
  NOR3_X1    g24612(.A1(new_n27843_), .A2(new_n27846_), .A3(new_n13855_), .ZN(new_n27847_));
  NOR3_X1    g24613(.A1(new_n27840_), .A2(new_n27847_), .A3(new_n13860_), .ZN(new_n27848_));
  NOR2_X1    g24614(.A1(new_n14428_), .A2(new_n13880_), .ZN(new_n27849_));
  AOI21_X1   g24615(.A1(new_n27820_), .A2(new_n13880_), .B(new_n27849_), .ZN(new_n27850_));
  AOI21_X1   g24616(.A1(new_n27850_), .A2(new_n13860_), .B(new_n13884_), .ZN(new_n27851_));
  INV_X1     g24617(.I(new_n27851_), .ZN(new_n27852_));
  OAI21_X1   g24618(.A1(new_n27848_), .A2(new_n27852_), .B(new_n13885_), .ZN(new_n27853_));
  OAI21_X1   g24619(.A1(new_n13855_), .A2(new_n27843_), .B(new_n27846_), .ZN(new_n27854_));
  NAND3_X1   g24620(.A1(new_n27829_), .A2(new_n27839_), .A3(pi0781), .ZN(new_n27855_));
  NAND3_X1   g24621(.A1(new_n27854_), .A2(new_n27855_), .A3(pi0619), .ZN(new_n27856_));
  NAND3_X1   g24622(.A1(new_n27856_), .A2(new_n14538_), .A3(new_n27851_), .ZN(new_n27857_));
  AOI21_X1   g24623(.A1(new_n27853_), .A2(new_n27857_), .B(new_n13627_), .ZN(new_n27858_));
  NOR3_X1    g24624(.A1(new_n27840_), .A2(new_n27847_), .A3(pi0619), .ZN(new_n27859_));
  AOI21_X1   g24625(.A1(new_n27850_), .A2(pi0619), .B(new_n13868_), .ZN(new_n27860_));
  INV_X1     g24626(.I(new_n27860_), .ZN(new_n27861_));
  OAI21_X1   g24627(.A1(new_n27859_), .A2(new_n27861_), .B(new_n13885_), .ZN(new_n27862_));
  NAND3_X1   g24628(.A1(new_n27854_), .A2(new_n27855_), .A3(new_n13860_), .ZN(new_n27863_));
  NAND3_X1   g24629(.A1(new_n27863_), .A2(new_n14538_), .A3(new_n27860_), .ZN(new_n27864_));
  NOR2_X1    g24630(.A1(new_n13627_), .A2(new_n13896_), .ZN(new_n27865_));
  OAI21_X1   g24631(.A1(new_n27840_), .A2(new_n27847_), .B(new_n27865_), .ZN(new_n27866_));
  AOI21_X1   g24632(.A1(new_n27862_), .A2(new_n27864_), .B(new_n27866_), .ZN(new_n27867_));
  OAI21_X1   g24633(.A1(new_n13896_), .A2(new_n27858_), .B(new_n27867_), .ZN(new_n27868_));
  AOI21_X1   g24634(.A1(new_n27856_), .A2(new_n27851_), .B(new_n14538_), .ZN(new_n27869_));
  NOR3_X1    g24635(.A1(new_n27848_), .A2(new_n13885_), .A3(new_n27852_), .ZN(new_n27870_));
  OAI21_X1   g24636(.A1(new_n27870_), .A2(new_n27869_), .B(new_n14428_), .ZN(new_n27871_));
  AOI21_X1   g24637(.A1(new_n27863_), .A2(new_n27860_), .B(new_n14538_), .ZN(new_n27872_));
  NOR3_X1    g24638(.A1(new_n27859_), .A2(new_n13885_), .A3(new_n27861_), .ZN(new_n27873_));
  INV_X1     g24639(.I(new_n27866_), .ZN(new_n27874_));
  OAI21_X1   g24640(.A1(new_n27873_), .A2(new_n27872_), .B(new_n27874_), .ZN(new_n27875_));
  NAND3_X1   g24641(.A1(new_n27871_), .A2(new_n27875_), .A3(pi0789), .ZN(new_n27876_));
  NOR2_X1    g24642(.A1(new_n13627_), .A2(new_n13919_), .ZN(new_n27877_));
  AOI21_X1   g24643(.A1(new_n27850_), .A2(new_n13919_), .B(new_n27877_), .ZN(new_n27878_));
  AOI21_X1   g24644(.A1(new_n13922_), .A2(new_n13929_), .B(pi0626), .ZN(new_n27879_));
  AOI21_X1   g24645(.A1(new_n27868_), .A2(new_n27876_), .B(new_n27879_), .ZN(new_n27880_));
  NOR2_X1    g24646(.A1(new_n16423_), .A2(new_n13937_), .ZN(new_n27883_));
  NOR2_X1    g24647(.A1(new_n13922_), .A2(new_n13929_), .ZN(new_n27884_));
  AOI21_X1   g24648(.A1(new_n27878_), .A2(new_n27884_), .B(pi0626), .ZN(new_n27885_));
  AOI21_X1   g24649(.A1(new_n27868_), .A2(new_n27876_), .B(new_n27885_), .ZN(new_n27886_));
  OAI21_X1   g24650(.A1(new_n27880_), .A2(new_n27883_), .B(new_n27886_), .ZN(new_n27887_));
  INV_X1     g24651(.I(new_n27887_), .ZN(new_n27888_));
  NOR2_X1    g24652(.A1(new_n19287_), .A2(new_n15392_), .ZN(new_n27889_));
  INV_X1     g24653(.I(new_n27889_), .ZN(new_n27890_));
  NOR3_X1    g24654(.A1(new_n27890_), .A2(new_n13766_), .A3(new_n13793_), .ZN(new_n27891_));
  NOR2_X1    g24655(.A1(new_n19390_), .A2(new_n3290_), .ZN(new_n27892_));
  AOI21_X1   g24656(.A1(new_n19287_), .A2(new_n14083_), .B(new_n13613_), .ZN(new_n27893_));
  AND2_X2    g24657(.A1(new_n27893_), .A2(pi1153), .Z(new_n27894_));
  OAI21_X1   g24658(.A1(new_n27894_), .A2(new_n27892_), .B(pi0625), .ZN(new_n27895_));
  OAI21_X1   g24659(.A1(new_n27895_), .A2(new_n27892_), .B(pi0778), .ZN(new_n27896_));
  AOI21_X1   g24660(.A1(new_n27896_), .A2(pi0609), .B(new_n27891_), .ZN(new_n27897_));
  INV_X1     g24661(.I(new_n27896_), .ZN(new_n27898_));
  NOR2_X1    g24662(.A1(new_n27898_), .A2(new_n13766_), .ZN(new_n27899_));
  OAI21_X1   g24663(.A1(new_n27899_), .A2(new_n27891_), .B(pi0785), .ZN(new_n27900_));
  NOR2_X1    g24664(.A1(new_n27900_), .A2(new_n27897_), .ZN(new_n27901_));
  NOR2_X1    g24665(.A1(new_n27898_), .A2(pi0785), .ZN(new_n27902_));
  OAI21_X1   g24666(.A1(new_n27901_), .A2(new_n27902_), .B(new_n13855_), .ZN(new_n27903_));
  INV_X1     g24667(.I(new_n15437_), .ZN(new_n27904_));
  NOR2_X1    g24668(.A1(new_n27890_), .A2(new_n27904_), .ZN(new_n27905_));
  INV_X1     g24669(.I(new_n27905_), .ZN(new_n27906_));
  NOR2_X1    g24670(.A1(new_n27906_), .A2(new_n18856_), .ZN(new_n27907_));
  NAND2_X1   g24671(.A1(new_n27903_), .A2(new_n27907_), .ZN(new_n27908_));
  NOR2_X1    g24672(.A1(new_n27890_), .A2(new_n13803_), .ZN(new_n27909_));
  INV_X1     g24673(.I(new_n27909_), .ZN(new_n27910_));
  NOR2_X1    g24674(.A1(new_n27901_), .A2(new_n27902_), .ZN(new_n27913_));
  INV_X1     g24675(.I(new_n13917_), .ZN(new_n27914_));
  XOR2_X1    g24676(.A1(pi0648), .A2(pi0789), .Z(new_n27915_));
  NAND4_X1   g24677(.A1(new_n27914_), .A2(pi0618), .A3(pi0619), .A4(new_n27915_), .ZN(new_n27916_));
  OAI21_X1   g24678(.A1(new_n27913_), .A2(new_n27916_), .B(new_n27908_), .ZN(new_n27917_));
  NOR2_X1    g24679(.A1(new_n27906_), .A2(new_n13918_), .ZN(new_n27918_));
  INV_X1     g24680(.I(new_n27918_), .ZN(new_n27919_));
  OAI21_X1   g24681(.A1(pi0641), .A2(pi1158), .B(new_n14577_), .ZN(new_n27920_));
  OAI21_X1   g24682(.A1(new_n27919_), .A2(new_n27920_), .B(new_n13901_), .ZN(new_n27921_));
  NAND2_X1   g24683(.A1(new_n27917_), .A2(new_n13937_), .ZN(new_n27922_));
  NOR2_X1    g24684(.A1(new_n27890_), .A2(new_n15396_), .ZN(new_n27923_));
  XOR2_X1    g24685(.A1(new_n27923_), .A2(new_n13994_), .Z(new_n27924_));
  NOR3_X1    g24686(.A1(new_n27924_), .A2(new_n13971_), .A3(new_n16423_), .ZN(new_n27925_));
  AOI22_X1   g24687(.A1(new_n27922_), .A2(new_n27925_), .B1(new_n27917_), .B2(new_n27921_), .ZN(new_n27926_));
  OAI21_X1   g24688(.A1(new_n27918_), .A2(new_n13901_), .B(new_n13922_), .ZN(new_n27927_));
  AOI21_X1   g24689(.A1(new_n27927_), .A2(new_n13929_), .B(new_n13901_), .ZN(new_n27928_));
  NAND2_X1   g24690(.A1(new_n27917_), .A2(new_n27928_), .ZN(new_n27929_));
  NOR2_X1    g24691(.A1(new_n27926_), .A2(new_n27929_), .ZN(new_n27930_));
  INV_X1     g24692(.I(new_n27930_), .ZN(new_n27931_));
  NOR3_X1    g24693(.A1(new_n27931_), .A2(new_n8545_), .A3(pi0623), .ZN(new_n27932_));
  INV_X1     g24694(.I(new_n27878_), .ZN(new_n27933_));
  NAND2_X1   g24695(.A1(new_n13627_), .A2(new_n13965_), .ZN(new_n27934_));
  OAI21_X1   g24696(.A1(new_n27933_), .A2(new_n13965_), .B(new_n27934_), .ZN(new_n27935_));
  NAND2_X1   g24697(.A1(new_n27935_), .A2(new_n14428_), .ZN(new_n27936_));
  NOR2_X1    g24698(.A1(new_n27936_), .A2(new_n13942_), .ZN(new_n27937_));
  XNOR2_X1   g24699(.A1(new_n27937_), .A2(new_n16420_), .ZN(new_n27938_));
  NOR2_X1    g24700(.A1(new_n27935_), .A2(new_n19484_), .ZN(new_n27939_));
  XOR2_X1    g24701(.A1(new_n27939_), .A2(new_n19486_), .Z(new_n27940_));
  NOR2_X1    g24702(.A1(new_n27940_), .A2(new_n13627_), .ZN(new_n27941_));
  INV_X1     g24703(.I(new_n27941_), .ZN(new_n27942_));
  NAND3_X1   g24704(.A1(new_n27942_), .A2(new_n13942_), .A3(new_n13969_), .ZN(new_n27943_));
  NOR2_X1    g24705(.A1(new_n13627_), .A2(new_n12777_), .ZN(new_n27944_));
  AOI21_X1   g24706(.A1(new_n27943_), .A2(new_n27944_), .B(pi1156), .ZN(new_n27945_));
  NOR2_X1    g24707(.A1(new_n27945_), .A2(new_n27938_), .ZN(new_n27946_));
  INV_X1     g24708(.I(new_n27946_), .ZN(new_n27947_));
  INV_X1     g24709(.I(new_n27789_), .ZN(new_n27948_));
  NOR2_X1    g24710(.A1(new_n22974_), .A2(new_n3290_), .ZN(new_n27949_));
  NOR2_X1    g24711(.A1(new_n19329_), .A2(new_n3290_), .ZN(new_n27950_));
  NOR2_X1    g24712(.A1(new_n27950_), .A2(new_n13613_), .ZN(new_n27951_));
  XOR2_X1    g24713(.A1(new_n27951_), .A2(new_n13615_), .Z(new_n27952_));
  AOI21_X1   g24714(.A1(new_n27952_), .A2(new_n27949_), .B(pi0608), .ZN(new_n27953_));
  AOI21_X1   g24715(.A1(new_n27782_), .A2(new_n27953_), .B(new_n13748_), .ZN(new_n27954_));
  NOR2_X1    g24716(.A1(new_n27950_), .A2(new_n13614_), .ZN(new_n27955_));
  XOR2_X1    g24717(.A1(new_n27955_), .A2(new_n13620_), .Z(new_n27956_));
  NOR2_X1    g24718(.A1(new_n14081_), .A2(new_n13748_), .ZN(new_n27957_));
  NAND3_X1   g24719(.A1(new_n27956_), .A2(new_n27949_), .A3(new_n27957_), .ZN(new_n27958_));
  AOI21_X1   g24720(.A1(new_n27777_), .A2(new_n27775_), .B(new_n27958_), .ZN(new_n27959_));
  INV_X1     g24721(.I(new_n27959_), .ZN(new_n27960_));
  NOR2_X1    g24722(.A1(new_n27954_), .A2(new_n27960_), .ZN(new_n27961_));
  XOR2_X1    g24723(.A1(new_n27770_), .A2(new_n13620_), .Z(new_n27962_));
  NAND2_X1   g24724(.A1(new_n19281_), .A2(new_n3289_), .ZN(new_n27963_));
  NOR2_X1    g24725(.A1(new_n27962_), .A2(new_n27963_), .ZN(new_n27964_));
  INV_X1     g24726(.I(new_n27953_), .ZN(new_n27965_));
  OAI21_X1   g24727(.A1(new_n27964_), .A2(new_n27965_), .B(pi0778), .ZN(new_n27966_));
  NOR2_X1    g24728(.A1(new_n27966_), .A2(new_n27959_), .ZN(new_n27967_));
  NOR2_X1    g24729(.A1(new_n27967_), .A2(new_n27961_), .ZN(new_n27968_));
  NAND2_X1   g24730(.A1(new_n27968_), .A2(pi1155), .ZN(new_n27969_));
  XOR2_X1    g24731(.A1(new_n27969_), .A2(new_n14090_), .Z(new_n27970_));
  NOR2_X1    g24732(.A1(new_n27950_), .A2(new_n13775_), .ZN(new_n27971_));
  AOI21_X1   g24733(.A1(new_n27971_), .A2(new_n16373_), .B(new_n13779_), .ZN(new_n27972_));
  NOR2_X1    g24734(.A1(new_n27972_), .A2(new_n13627_), .ZN(new_n27973_));
  NOR2_X1    g24735(.A1(new_n27973_), .A2(new_n13783_), .ZN(new_n27974_));
  OAI21_X1   g24736(.A1(new_n27970_), .A2(new_n27948_), .B(new_n27974_), .ZN(new_n27975_));
  NOR3_X1    g24737(.A1(new_n27950_), .A2(new_n13775_), .A3(new_n14694_), .ZN(new_n27976_));
  OAI21_X1   g24738(.A1(new_n14101_), .A2(new_n27976_), .B(new_n14428_), .ZN(new_n27977_));
  NAND3_X1   g24739(.A1(new_n27975_), .A2(new_n13783_), .A3(new_n27977_), .ZN(new_n27978_));
  NAND2_X1   g24740(.A1(new_n27968_), .A2(pi0609), .ZN(new_n27979_));
  XOR2_X1    g24741(.A1(new_n27979_), .A2(new_n14694_), .Z(new_n27980_));
  NAND4_X1   g24742(.A1(new_n27978_), .A2(pi0785), .A3(new_n27789_), .A4(new_n27980_), .ZN(new_n27981_));
  NAND2_X1   g24743(.A1(new_n27968_), .A2(new_n13801_), .ZN(new_n27982_));
  NAND2_X1   g24744(.A1(new_n27981_), .A2(new_n27982_), .ZN(new_n27983_));
  INV_X1     g24745(.I(new_n27983_), .ZN(new_n27984_));
  NAND3_X1   g24746(.A1(new_n27983_), .A2(pi0618), .A3(pi1154), .ZN(new_n27985_));
  INV_X1     g24747(.I(new_n27985_), .ZN(new_n27986_));
  NOR3_X1    g24748(.A1(new_n27983_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n27987_));
  OAI21_X1   g24749(.A1(new_n27986_), .A2(new_n27987_), .B(new_n27821_), .ZN(new_n27988_));
  NOR2_X1    g24750(.A1(new_n27973_), .A2(new_n13801_), .ZN(new_n27989_));
  NOR2_X1    g24751(.A1(new_n13627_), .A2(new_n13776_), .ZN(new_n27990_));
  AOI21_X1   g24752(.A1(new_n13776_), .A2(new_n27950_), .B(new_n27990_), .ZN(new_n27991_));
  NOR3_X1    g24753(.A1(new_n27991_), .A2(new_n27977_), .A3(new_n13801_), .ZN(new_n27992_));
  XNOR2_X1   g24754(.A1(new_n27992_), .A2(new_n27989_), .ZN(new_n27993_));
  NAND2_X1   g24755(.A1(new_n27993_), .A2(pi1154), .ZN(new_n27994_));
  XOR2_X1    g24756(.A1(new_n27994_), .A2(new_n13819_), .Z(new_n27995_));
  NAND2_X1   g24757(.A1(new_n27995_), .A2(new_n14428_), .ZN(new_n27996_));
  NAND2_X1   g24758(.A1(new_n27996_), .A2(new_n13823_), .ZN(new_n27997_));
  INV_X1     g24759(.I(new_n27997_), .ZN(new_n27998_));
  NAND2_X1   g24760(.A1(new_n27993_), .A2(pi0618), .ZN(new_n27999_));
  XOR2_X1    g24761(.A1(new_n27999_), .A2(new_n13819_), .Z(new_n28000_));
  NAND2_X1   g24762(.A1(new_n28000_), .A2(new_n14428_), .ZN(new_n28001_));
  NAND2_X1   g24763(.A1(new_n28001_), .A2(new_n13823_), .ZN(new_n28002_));
  AOI21_X1   g24764(.A1(new_n27988_), .A2(new_n27998_), .B(new_n28002_), .ZN(new_n28003_));
  NOR2_X1    g24765(.A1(new_n27983_), .A2(new_n13817_), .ZN(new_n28004_));
  NOR2_X1    g24766(.A1(new_n28004_), .A2(new_n13819_), .ZN(new_n28005_));
  NAND2_X1   g24767(.A1(new_n28004_), .A2(new_n13819_), .ZN(new_n28006_));
  INV_X1     g24768(.I(new_n28006_), .ZN(new_n28007_));
  OAI21_X1   g24769(.A1(new_n28007_), .A2(new_n28005_), .B(new_n27821_), .ZN(new_n28008_));
  NOR2_X1    g24770(.A1(new_n28003_), .A2(new_n28008_), .ZN(new_n28009_));
  NAND3_X1   g24771(.A1(new_n28009_), .A2(pi0619), .A3(pi0781), .ZN(new_n28010_));
  INV_X1     g24772(.I(new_n27987_), .ZN(new_n28011_));
  AOI21_X1   g24773(.A1(new_n28011_), .A2(new_n27985_), .B(new_n27820_), .ZN(new_n28012_));
  INV_X1     g24774(.I(new_n28002_), .ZN(new_n28013_));
  OAI21_X1   g24775(.A1(new_n28012_), .A2(new_n27997_), .B(new_n28013_), .ZN(new_n28014_));
  INV_X1     g24776(.I(new_n28005_), .ZN(new_n28015_));
  AOI21_X1   g24777(.A1(new_n28015_), .A2(new_n28006_), .B(new_n27820_), .ZN(new_n28016_));
  NAND2_X1   g24778(.A1(new_n28014_), .A2(new_n28016_), .ZN(new_n28017_));
  NAND3_X1   g24779(.A1(new_n28017_), .A2(pi0619), .A3(new_n13855_), .ZN(new_n28018_));
  AOI21_X1   g24780(.A1(new_n28018_), .A2(new_n28010_), .B(new_n27984_), .ZN(new_n28019_));
  NAND2_X1   g24781(.A1(new_n27996_), .A2(pi0781), .ZN(new_n28020_));
  NOR3_X1    g24782(.A1(new_n28001_), .A2(new_n13855_), .A3(new_n27993_), .ZN(new_n28021_));
  XOR2_X1    g24783(.A1(new_n28021_), .A2(new_n28020_), .Z(new_n28022_));
  NAND2_X1   g24784(.A1(new_n28022_), .A2(pi0619), .ZN(new_n28023_));
  NAND2_X1   g24785(.A1(new_n28023_), .A2(new_n13903_), .ZN(new_n28024_));
  XNOR2_X1   g24786(.A1(new_n28021_), .A2(new_n28020_), .ZN(new_n28025_));
  NOR2_X1    g24787(.A1(new_n28025_), .A2(new_n13860_), .ZN(new_n28026_));
  NAND2_X1   g24788(.A1(new_n28026_), .A2(new_n13904_), .ZN(new_n28027_));
  AOI21_X1   g24789(.A1(new_n28027_), .A2(new_n28024_), .B(new_n13627_), .ZN(new_n28028_));
  NOR2_X1    g24790(.A1(new_n28028_), .A2(new_n14538_), .ZN(new_n28029_));
  NOR2_X1    g24791(.A1(new_n27850_), .A2(pi0619), .ZN(new_n28030_));
  OAI21_X1   g24792(.A1(new_n28019_), .A2(new_n28029_), .B(new_n28030_), .ZN(new_n28031_));
  NAND2_X1   g24793(.A1(new_n28031_), .A2(new_n13896_), .ZN(new_n28032_));
  NOR2_X1    g24794(.A1(new_n27984_), .A2(pi0781), .ZN(new_n28033_));
  INV_X1     g24795(.I(new_n28033_), .ZN(new_n28034_));
  NAND3_X1   g24796(.A1(new_n28014_), .A2(pi0781), .A3(new_n28016_), .ZN(new_n28035_));
  AOI21_X1   g24797(.A1(new_n28035_), .A2(new_n28034_), .B(pi0789), .ZN(new_n28036_));
  NOR2_X1    g24798(.A1(new_n14428_), .A2(new_n16372_), .ZN(new_n28037_));
  INV_X1     g24799(.I(new_n28037_), .ZN(new_n28038_));
  NOR2_X1    g24800(.A1(new_n28025_), .A2(new_n13868_), .ZN(new_n28039_));
  NOR2_X1    g24801(.A1(new_n28039_), .A2(new_n13904_), .ZN(new_n28040_));
  NAND2_X1   g24802(.A1(new_n28022_), .A2(pi1159), .ZN(new_n28041_));
  NOR2_X1    g24803(.A1(new_n28041_), .A2(new_n13903_), .ZN(new_n28042_));
  OAI21_X1   g24804(.A1(new_n28040_), .A2(new_n28042_), .B(new_n14428_), .ZN(new_n28043_));
  NAND2_X1   g24805(.A1(new_n28043_), .A2(pi0789), .ZN(new_n28044_));
  NOR2_X1    g24806(.A1(new_n28026_), .A2(new_n13904_), .ZN(new_n28045_));
  NOR2_X1    g24807(.A1(new_n28023_), .A2(new_n13903_), .ZN(new_n28046_));
  NOR2_X1    g24808(.A1(new_n28045_), .A2(new_n28046_), .ZN(new_n28047_));
  NOR4_X1    g24809(.A1(new_n28047_), .A2(new_n13896_), .A3(new_n13627_), .A4(new_n28022_), .ZN(new_n28048_));
  NAND2_X1   g24810(.A1(new_n28048_), .A2(new_n28044_), .ZN(new_n28049_));
  NAND2_X1   g24811(.A1(new_n28041_), .A2(new_n13903_), .ZN(new_n28050_));
  NAND2_X1   g24812(.A1(new_n28039_), .A2(new_n13904_), .ZN(new_n28051_));
  AOI21_X1   g24813(.A1(new_n28051_), .A2(new_n28050_), .B(new_n13627_), .ZN(new_n28052_));
  NOR2_X1    g24814(.A1(new_n28052_), .A2(new_n13896_), .ZN(new_n28053_));
  NAND3_X1   g24815(.A1(new_n28028_), .A2(pi0789), .A3(new_n28025_), .ZN(new_n28054_));
  NAND2_X1   g24816(.A1(new_n28054_), .A2(new_n28053_), .ZN(new_n28055_));
  NAND2_X1   g24817(.A1(new_n28049_), .A2(new_n28055_), .ZN(new_n28056_));
  OAI21_X1   g24818(.A1(new_n28056_), .A2(new_n14142_), .B(new_n28038_), .ZN(new_n28057_));
  NAND2_X1   g24819(.A1(new_n27942_), .A2(new_n13985_), .ZN(new_n28058_));
  NOR2_X1    g24820(.A1(new_n13627_), .A2(pi0628), .ZN(new_n28059_));
  NOR2_X1    g24821(.A1(new_n27935_), .A2(new_n13942_), .ZN(new_n28060_));
  OAI21_X1   g24822(.A1(new_n28060_), .A2(new_n28059_), .B(pi0792), .ZN(new_n28061_));
  INV_X1     g24823(.I(new_n28061_), .ZN(new_n28062_));
  AOI21_X1   g24824(.A1(new_n28058_), .A2(new_n28062_), .B(new_n28057_), .ZN(new_n28063_));
  NOR2_X1    g24825(.A1(new_n28054_), .A2(new_n28053_), .ZN(new_n28064_));
  NOR2_X1    g24826(.A1(new_n28048_), .A2(new_n28044_), .ZN(new_n28065_));
  NOR2_X1    g24827(.A1(new_n28065_), .A2(new_n28064_), .ZN(new_n28066_));
  NOR2_X1    g24828(.A1(new_n28066_), .A2(pi1158), .ZN(new_n28067_));
  NOR2_X1    g24829(.A1(new_n28056_), .A2(new_n13929_), .ZN(new_n28068_));
  OAI21_X1   g24830(.A1(new_n14428_), .A2(pi0641), .B(new_n14139_), .ZN(new_n28069_));
  INV_X1     g24831(.I(new_n14140_), .ZN(new_n28070_));
  AOI21_X1   g24832(.A1(new_n13627_), .A2(pi0641), .B(new_n28070_), .ZN(new_n28071_));
  INV_X1     g24833(.I(new_n28071_), .ZN(new_n28072_));
  OAI22_X1   g24834(.A1(new_n27933_), .A2(new_n13922_), .B1(new_n28069_), .B2(new_n28072_), .ZN(new_n28073_));
  NOR2_X1    g24835(.A1(new_n28073_), .A2(new_n19203_), .ZN(new_n28074_));
  NOR4_X1    g24836(.A1(new_n28074_), .A2(new_n13901_), .A3(new_n13964_), .A4(new_n16875_), .ZN(new_n28075_));
  OAI21_X1   g24837(.A1(new_n28067_), .A2(new_n28068_), .B(new_n28075_), .ZN(new_n28076_));
  OAI22_X1   g24838(.A1(new_n28063_), .A2(new_n28076_), .B1(new_n28036_), .B2(new_n15479_), .ZN(new_n28077_));
  INV_X1     g24839(.I(new_n28077_), .ZN(new_n28078_));
  AOI21_X1   g24840(.A1(new_n28009_), .A2(pi0781), .B(new_n28033_), .ZN(new_n28079_));
  AOI21_X1   g24841(.A1(new_n28079_), .A2(pi0619), .B(new_n13904_), .ZN(new_n28080_));
  NAND3_X1   g24842(.A1(new_n28035_), .A2(pi0619), .A3(new_n28034_), .ZN(new_n28081_));
  NOR2_X1    g24843(.A1(new_n28081_), .A2(new_n13903_), .ZN(new_n28082_));
  NOR3_X1    g24844(.A1(new_n28052_), .A2(pi0648), .A3(new_n27850_), .ZN(new_n28083_));
  OAI21_X1   g24845(.A1(new_n28080_), .A2(new_n28082_), .B(new_n28083_), .ZN(new_n28084_));
  NOR2_X1    g24846(.A1(new_n28078_), .A2(new_n28084_), .ZN(new_n28085_));
  INV_X1     g24847(.I(new_n19323_), .ZN(new_n28086_));
  NAND3_X1   g24848(.A1(new_n15628_), .A2(pi0625), .A3(new_n3289_), .ZN(new_n28088_));
  NAND2_X1   g24849(.A1(new_n28088_), .A2(pi0778), .ZN(new_n28089_));
  AND3_X2    g24850(.A1(new_n15628_), .A2(new_n3289_), .A3(new_n20409_), .Z(new_n28091_));
  XOR2_X1    g24851(.A1(new_n28089_), .A2(new_n28091_), .Z(new_n28092_));
  NAND2_X1   g24852(.A1(new_n28092_), .A2(pi1155), .ZN(new_n28093_));
  XOR2_X1    g24853(.A1(new_n28093_), .A2(new_n14694_), .Z(new_n28094_));
  NAND2_X1   g24854(.A1(new_n28094_), .A2(new_n27889_), .ZN(new_n28095_));
  NOR3_X1    g24855(.A1(new_n28086_), .A2(new_n3290_), .A3(new_n13775_), .ZN(new_n28096_));
  INV_X1     g24856(.I(new_n28096_), .ZN(new_n28097_));
  AOI21_X1   g24857(.A1(new_n28097_), .A2(new_n13793_), .B(new_n13766_), .ZN(new_n28098_));
  AOI21_X1   g24858(.A1(new_n28095_), .A2(new_n28098_), .B(new_n13801_), .ZN(new_n28099_));
  INV_X1     g24859(.I(new_n28092_), .ZN(new_n28100_));
  NAND2_X1   g24860(.A1(new_n28092_), .A2(pi0609), .ZN(new_n28101_));
  XOR2_X1    g24861(.A1(new_n28101_), .A2(new_n14694_), .Z(new_n28102_));
  NAND2_X1   g24862(.A1(new_n28102_), .A2(new_n27889_), .ZN(new_n28103_));
  NAND4_X1   g24863(.A1(new_n28103_), .A2(pi0785), .A3(new_n28100_), .A4(new_n28098_), .ZN(new_n28104_));
  XNOR2_X1   g24864(.A1(new_n28104_), .A2(new_n28099_), .ZN(new_n28105_));
  NAND3_X1   g24865(.A1(new_n28105_), .A2(pi0618), .A3(pi1154), .ZN(new_n28106_));
  XOR2_X1    g24866(.A1(new_n28104_), .A2(new_n28099_), .Z(new_n28107_));
  NAND3_X1   g24867(.A1(new_n28107_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n28108_));
  OAI21_X1   g24868(.A1(new_n28097_), .A2(new_n16376_), .B(new_n13836_), .ZN(new_n28109_));
  NAND2_X1   g24869(.A1(new_n28109_), .A2(pi0618), .ZN(new_n28110_));
  OAI21_X1   g24870(.A1(new_n28110_), .A2(new_n13817_), .B(new_n13816_), .ZN(new_n28111_));
  NAND3_X1   g24871(.A1(new_n28111_), .A2(pi0781), .A3(new_n27909_), .ZN(new_n28112_));
  AOI21_X1   g24872(.A1(new_n28112_), .A2(new_n28110_), .B(new_n27910_), .ZN(new_n28113_));
  INV_X1     g24873(.I(new_n28113_), .ZN(new_n28114_));
  AOI21_X1   g24874(.A1(new_n28106_), .A2(new_n28108_), .B(new_n28114_), .ZN(new_n28115_));
  NOR3_X1    g24875(.A1(new_n28097_), .A2(new_n16376_), .A3(new_n16382_), .ZN(new_n28116_));
  NAND2_X1   g24876(.A1(new_n13860_), .A2(new_n13884_), .ZN(new_n28117_));
  NAND4_X1   g24877(.A1(new_n27905_), .A2(pi0789), .A3(pi1159), .A4(new_n28117_), .ZN(new_n28118_));
  NAND4_X1   g24878(.A1(new_n27905_), .A2(pi1159), .A3(new_n28116_), .A4(new_n28117_), .ZN(new_n28119_));
  OAI21_X1   g24879(.A1(new_n28118_), .A2(new_n28119_), .B(new_n13868_), .ZN(new_n28120_));
  NAND2_X1   g24880(.A1(new_n28120_), .A2(new_n28116_), .ZN(new_n28121_));
  NOR2_X1    g24881(.A1(new_n16697_), .A2(new_n18868_), .ZN(new_n28122_));
  NOR2_X1    g24882(.A1(new_n28121_), .A2(new_n28122_), .ZN(new_n28123_));
  OAI21_X1   g24883(.A1(new_n28107_), .A2(new_n13855_), .B(new_n13823_), .ZN(new_n28124_));
  AOI21_X1   g24884(.A1(new_n28124_), .A2(pi0618), .B(new_n28123_), .ZN(new_n28125_));
  INV_X1     g24885(.I(new_n28125_), .ZN(new_n28126_));
  NAND2_X1   g24886(.A1(new_n28121_), .A2(pi0789), .ZN(new_n28127_));
  OAI21_X1   g24887(.A1(new_n28126_), .A2(new_n28115_), .B(new_n28127_), .ZN(new_n28128_));
  NOR2_X1    g24888(.A1(new_n28128_), .A2(pi0788), .ZN(new_n28129_));
  INV_X1     g24889(.I(new_n28129_), .ZN(new_n28130_));
  AOI21_X1   g24890(.A1(new_n13942_), .A2(new_n13976_), .B(new_n13969_), .ZN(new_n28131_));
  NAND2_X1   g24891(.A1(new_n27923_), .A2(new_n28131_), .ZN(new_n28132_));
  INV_X1     g24892(.I(new_n28132_), .ZN(new_n28133_));
  AOI21_X1   g24893(.A1(new_n28116_), .A2(new_n13868_), .B(pi0619), .ZN(new_n28134_));
  OAI21_X1   g24894(.A1(new_n13868_), .A2(new_n28116_), .B(new_n28134_), .ZN(new_n28135_));
  NAND2_X1   g24895(.A1(new_n28135_), .A2(pi0789), .ZN(new_n28136_));
  NOR2_X1    g24896(.A1(new_n28136_), .A2(new_n14142_), .ZN(new_n28137_));
  INV_X1     g24897(.I(new_n28137_), .ZN(new_n28138_));
  AOI21_X1   g24898(.A1(new_n28138_), .A2(pi1156), .B(new_n28133_), .ZN(new_n28139_));
  AOI21_X1   g24899(.A1(new_n28138_), .A2(pi1156), .B(new_n28133_), .ZN(new_n28140_));
  NOR3_X1    g24900(.A1(new_n28139_), .A2(new_n28140_), .A3(new_n16423_), .ZN(new_n28141_));
  NOR2_X1    g24901(.A1(pi0626), .A2(pi1158), .ZN(new_n28142_));
  AOI21_X1   g24902(.A1(new_n28136_), .A2(new_n28142_), .B(new_n13922_), .ZN(new_n28143_));
  INV_X1     g24903(.I(new_n28143_), .ZN(new_n28144_));
  AOI21_X1   g24904(.A1(new_n28107_), .A2(pi1154), .B(new_n13819_), .ZN(new_n28145_));
  NOR3_X1    g24905(.A1(new_n28105_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n28146_));
  OAI21_X1   g24906(.A1(new_n28146_), .A2(new_n28145_), .B(new_n28113_), .ZN(new_n28147_));
  AOI22_X1   g24907(.A1(new_n28147_), .A2(new_n28125_), .B1(pi0789), .B2(new_n28121_), .ZN(new_n28148_));
  NAND3_X1   g24908(.A1(new_n27918_), .A2(pi0626), .A3(new_n13922_), .ZN(new_n28149_));
  AOI21_X1   g24909(.A1(new_n14160_), .A2(new_n28136_), .B(new_n28149_), .ZN(new_n28150_));
  OAI21_X1   g24910(.A1(new_n28148_), .A2(new_n28150_), .B(new_n14577_), .ZN(new_n28151_));
  NAND2_X1   g24911(.A1(new_n28151_), .A2(new_n28144_), .ZN(new_n28152_));
  NAND3_X1   g24912(.A1(new_n28148_), .A2(pi0626), .A3(pi0641), .ZN(new_n28153_));
  NAND3_X1   g24913(.A1(new_n28128_), .A2(new_n13901_), .A3(pi0641), .ZN(new_n28154_));
  NOR2_X1    g24914(.A1(new_n27919_), .A2(new_n12777_), .ZN(new_n28155_));
  INV_X1     g24915(.I(new_n28155_), .ZN(new_n28156_));
  AOI21_X1   g24916(.A1(new_n28154_), .A2(new_n28153_), .B(new_n28156_), .ZN(new_n28157_));
  AOI22_X1   g24917(.A1(new_n28157_), .A2(new_n28152_), .B1(new_n28130_), .B2(new_n28141_), .ZN(new_n28158_));
  AOI21_X1   g24918(.A1(pi0623), .A2(pi0710), .B(pi0207), .ZN(new_n28159_));
  INV_X1     g24919(.I(new_n28159_), .ZN(new_n28160_));
  NAND3_X1   g24920(.A1(new_n28085_), .A2(new_n28032_), .A3(new_n28160_), .ZN(new_n28161_));
  NOR2_X1    g24921(.A1(new_n28138_), .A2(new_n13993_), .ZN(new_n28162_));
  INV_X1     g24922(.I(new_n28162_), .ZN(new_n28163_));
  NOR3_X1    g24923(.A1(new_n28065_), .A2(new_n28064_), .A3(new_n14142_), .ZN(new_n28164_));
  OAI21_X1   g24924(.A1(new_n28164_), .A2(new_n28037_), .B(new_n13994_), .ZN(new_n28165_));
  NOR2_X1    g24925(.A1(new_n14428_), .A2(new_n13994_), .ZN(new_n28166_));
  INV_X1     g24926(.I(new_n28166_), .ZN(new_n28167_));
  NAND2_X1   g24927(.A1(new_n28165_), .A2(new_n28167_), .ZN(new_n28168_));
  NAND3_X1   g24928(.A1(new_n28168_), .A2(pi0207), .A3(pi0623), .ZN(new_n28169_));
  AOI21_X1   g24929(.A1(new_n28057_), .A2(new_n13994_), .B(new_n28166_), .ZN(new_n28170_));
  NAND3_X1   g24930(.A1(new_n28170_), .A2(new_n8545_), .A3(pi0623), .ZN(new_n28171_));
  AOI21_X1   g24931(.A1(new_n28171_), .A2(new_n28169_), .B(new_n28163_), .ZN(new_n28172_));
  NOR2_X1    g24932(.A1(new_n14428_), .A2(pi0207), .ZN(new_n28173_));
  INV_X1     g24933(.I(new_n28173_), .ZN(new_n28174_));
  NOR2_X1    g24934(.A1(new_n28174_), .A2(pi0623), .ZN(new_n28175_));
  INV_X1     g24935(.I(pi0710), .ZN(new_n28176_));
  NAND2_X1   g24936(.A1(new_n27936_), .A2(new_n14059_), .ZN(new_n28177_));
  NAND2_X1   g24937(.A1(new_n28177_), .A2(new_n8545_), .ZN(new_n28178_));
  NAND2_X1   g24938(.A1(new_n27923_), .A2(new_n14059_), .ZN(new_n28179_));
  INV_X1     g24939(.I(new_n28179_), .ZN(new_n28180_));
  NAND2_X1   g24940(.A1(new_n28180_), .A2(pi0207), .ZN(new_n28181_));
  AOI21_X1   g24941(.A1(new_n28178_), .A2(new_n28181_), .B(new_n28176_), .ZN(new_n28182_));
  AOI21_X1   g24942(.A1(new_n28176_), .A2(new_n28173_), .B(new_n28182_), .ZN(new_n28183_));
  AOI21_X1   g24943(.A1(new_n28183_), .A2(pi0647), .B(new_n14008_), .ZN(new_n28184_));
  NAND2_X1   g24944(.A1(new_n28183_), .A2(pi0647), .ZN(new_n28185_));
  NOR2_X1    g24945(.A1(new_n28185_), .A2(new_n14007_), .ZN(new_n28186_));
  OR2_X2     g24946(.A1(new_n28186_), .A2(new_n28184_), .Z(new_n28187_));
  AOI21_X1   g24947(.A1(new_n28187_), .A2(new_n28173_), .B(new_n14010_), .ZN(new_n28188_));
  NAND2_X1   g24948(.A1(new_n28183_), .A2(pi1157), .ZN(new_n28189_));
  XOR2_X1    g24949(.A1(new_n28189_), .A2(new_n14008_), .Z(new_n28190_));
  AOI21_X1   g24950(.A1(new_n28190_), .A2(new_n28173_), .B(pi0630), .ZN(new_n28191_));
  NOR2_X1    g24951(.A1(new_n28188_), .A2(new_n28191_), .ZN(new_n28192_));
  OAI22_X1   g24952(.A1(new_n28172_), .A2(new_n28175_), .B1(new_n12776_), .B2(new_n28192_), .ZN(new_n28193_));
  OAI21_X1   g24953(.A1(new_n28172_), .A2(new_n28175_), .B(new_n28176_), .ZN(new_n28194_));
  NOR2_X1    g24954(.A1(new_n16574_), .A2(new_n16867_), .ZN(new_n28195_));
  NAND3_X1   g24955(.A1(new_n28193_), .A2(new_n28194_), .A3(new_n28195_), .ZN(new_n28196_));
  AOI21_X1   g24956(.A1(new_n28196_), .A2(new_n28161_), .B(new_n27947_), .ZN(new_n28197_));
  OAI21_X1   g24957(.A1(new_n27888_), .A2(new_n27932_), .B(new_n28197_), .ZN(new_n28198_));
  INV_X1     g24958(.I(new_n28169_), .ZN(new_n28199_));
  INV_X1     g24959(.I(pi0623), .ZN(new_n28200_));
  NOR3_X1    g24960(.A1(new_n28168_), .A2(pi0207), .A3(new_n28200_), .ZN(new_n28201_));
  OAI21_X1   g24961(.A1(new_n28199_), .A2(new_n28201_), .B(new_n28162_), .ZN(new_n28202_));
  INV_X1     g24962(.I(new_n28175_), .ZN(new_n28203_));
  NAND2_X1   g24963(.A1(new_n28202_), .A2(new_n28203_), .ZN(new_n28204_));
  NOR2_X1    g24964(.A1(new_n28174_), .A2(new_n14211_), .ZN(new_n28205_));
  AOI21_X1   g24965(.A1(new_n28204_), .A2(new_n14211_), .B(new_n28205_), .ZN(new_n28206_));
  OAI21_X1   g24966(.A1(new_n28174_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n28207_));
  NAND2_X1   g24967(.A1(new_n28206_), .A2(new_n28207_), .ZN(new_n28208_));
  AOI21_X1   g24968(.A1(new_n28190_), .A2(new_n28173_), .B(new_n12776_), .ZN(new_n28209_));
  NAND2_X1   g24969(.A1(new_n28187_), .A2(new_n28173_), .ZN(new_n28210_));
  NOR3_X1    g24970(.A1(new_n28210_), .A2(new_n12776_), .A3(new_n28183_), .ZN(new_n28211_));
  XNOR2_X1   g24971(.A1(new_n28211_), .A2(new_n28209_), .ZN(new_n28212_));
  NAND4_X1   g24972(.A1(new_n28208_), .A2(pi0644), .A3(new_n14200_), .A4(new_n28212_), .ZN(new_n28213_));
  AOI21_X1   g24973(.A1(new_n28198_), .A2(new_n28213_), .B(new_n14204_), .ZN(new_n28214_));
  NAND2_X1   g24974(.A1(pi0644), .A2(pi0715), .ZN(new_n28215_));
  NOR2_X1    g24975(.A1(new_n28206_), .A2(new_n28215_), .ZN(new_n28216_));
  OAI21_X1   g24976(.A1(new_n28216_), .A2(pi0644), .B(pi0790), .ZN(new_n28217_));
  NOR2_X1    g24977(.A1(new_n28198_), .A2(new_n28217_), .ZN(new_n28218_));
  NOR3_X1    g24978(.A1(new_n28214_), .A2(new_n28218_), .A3(new_n12775_), .ZN(new_n28219_));
  NOR2_X1    g24979(.A1(new_n27888_), .A2(new_n27932_), .ZN(new_n28220_));
  INV_X1     g24980(.I(new_n28161_), .ZN(new_n28221_));
  INV_X1     g24981(.I(new_n28192_), .ZN(new_n28222_));
  AOI22_X1   g24982(.A1(new_n28202_), .A2(new_n28203_), .B1(pi0787), .B2(new_n28222_), .ZN(new_n28223_));
  NAND2_X1   g24983(.A1(new_n28194_), .A2(new_n28195_), .ZN(new_n28224_));
  NOR2_X1    g24984(.A1(new_n28224_), .A2(new_n28223_), .ZN(new_n28225_));
  OAI21_X1   g24985(.A1(new_n28225_), .A2(new_n28221_), .B(new_n27946_), .ZN(new_n28226_));
  NOR2_X1    g24986(.A1(new_n28226_), .A2(new_n28220_), .ZN(new_n28227_));
  NAND3_X1   g24987(.A1(new_n28227_), .A2(pi0644), .A3(pi0790), .ZN(new_n28229_));
  NAND2_X1   g24988(.A1(new_n28229_), .A2(new_n7240_), .ZN(new_n28230_));
  OAI21_X1   g24989(.A1(new_n28219_), .A2(new_n28230_), .B(new_n27769_), .ZN(po0364));
  NAND2_X1   g24990(.A1(po1038), .A2(new_n8546_), .ZN(new_n28232_));
  NOR3_X1    g24991(.A1(new_n27931_), .A2(new_n8546_), .A3(pi0607), .ZN(new_n28233_));
  AOI21_X1   g24992(.A1(pi0607), .A2(pi0638), .B(pi0208), .ZN(new_n28234_));
  INV_X1     g24993(.I(new_n28234_), .ZN(new_n28235_));
  NAND3_X1   g24994(.A1(new_n28085_), .A2(new_n28032_), .A3(new_n28235_), .ZN(new_n28236_));
  NAND3_X1   g24995(.A1(new_n28168_), .A2(pi0208), .A3(pi0607), .ZN(new_n28237_));
  NAND3_X1   g24996(.A1(new_n28170_), .A2(new_n8546_), .A3(pi0607), .ZN(new_n28238_));
  AOI21_X1   g24997(.A1(new_n28238_), .A2(new_n28237_), .B(new_n28163_), .ZN(new_n28239_));
  NOR2_X1    g24998(.A1(new_n14428_), .A2(pi0208), .ZN(new_n28240_));
  INV_X1     g24999(.I(new_n28240_), .ZN(new_n28241_));
  NOR2_X1    g25000(.A1(new_n28241_), .A2(pi0607), .ZN(new_n28242_));
  INV_X1     g25001(.I(pi0638), .ZN(new_n28243_));
  NAND2_X1   g25002(.A1(new_n28177_), .A2(new_n8546_), .ZN(new_n28244_));
  NAND2_X1   g25003(.A1(new_n28180_), .A2(pi0208), .ZN(new_n28245_));
  AOI21_X1   g25004(.A1(new_n28244_), .A2(new_n28245_), .B(new_n28243_), .ZN(new_n28246_));
  AOI21_X1   g25005(.A1(new_n28243_), .A2(new_n28240_), .B(new_n28246_), .ZN(new_n28247_));
  AOI21_X1   g25006(.A1(new_n28247_), .A2(pi0647), .B(new_n14008_), .ZN(new_n28248_));
  NAND2_X1   g25007(.A1(new_n28247_), .A2(pi0647), .ZN(new_n28249_));
  NOR2_X1    g25008(.A1(new_n28249_), .A2(new_n14007_), .ZN(new_n28250_));
  OR2_X2     g25009(.A1(new_n28250_), .A2(new_n28248_), .Z(new_n28251_));
  AOI21_X1   g25010(.A1(new_n28251_), .A2(new_n28240_), .B(new_n14010_), .ZN(new_n28252_));
  NAND2_X1   g25011(.A1(new_n28247_), .A2(pi1157), .ZN(new_n28253_));
  XOR2_X1    g25012(.A1(new_n28253_), .A2(new_n14008_), .Z(new_n28254_));
  AOI21_X1   g25013(.A1(new_n28254_), .A2(new_n28240_), .B(pi0630), .ZN(new_n28255_));
  NOR2_X1    g25014(.A1(new_n28252_), .A2(new_n28255_), .ZN(new_n28256_));
  OAI22_X1   g25015(.A1(new_n28239_), .A2(new_n28242_), .B1(new_n12776_), .B2(new_n28256_), .ZN(new_n28257_));
  OAI21_X1   g25016(.A1(new_n28239_), .A2(new_n28242_), .B(new_n28243_), .ZN(new_n28258_));
  NAND3_X1   g25017(.A1(new_n28257_), .A2(new_n28258_), .A3(new_n28195_), .ZN(new_n28259_));
  AOI21_X1   g25018(.A1(new_n28259_), .A2(new_n28236_), .B(new_n27947_), .ZN(new_n28260_));
  OAI21_X1   g25019(.A1(new_n27888_), .A2(new_n28233_), .B(new_n28260_), .ZN(new_n28261_));
  INV_X1     g25020(.I(new_n28237_), .ZN(new_n28262_));
  INV_X1     g25021(.I(pi0607), .ZN(new_n28263_));
  NOR3_X1    g25022(.A1(new_n28168_), .A2(pi0208), .A3(new_n28263_), .ZN(new_n28264_));
  OAI21_X1   g25023(.A1(new_n28262_), .A2(new_n28264_), .B(new_n28162_), .ZN(new_n28265_));
  INV_X1     g25024(.I(new_n28242_), .ZN(new_n28266_));
  NAND2_X1   g25025(.A1(new_n28265_), .A2(new_n28266_), .ZN(new_n28267_));
  NOR2_X1    g25026(.A1(new_n28241_), .A2(new_n14211_), .ZN(new_n28268_));
  AOI21_X1   g25027(.A1(new_n28267_), .A2(new_n14211_), .B(new_n28268_), .ZN(new_n28269_));
  OAI21_X1   g25028(.A1(new_n28241_), .A2(new_n14204_), .B(new_n14243_), .ZN(new_n28270_));
  NAND2_X1   g25029(.A1(new_n28269_), .A2(new_n28270_), .ZN(new_n28271_));
  AOI21_X1   g25030(.A1(new_n28254_), .A2(new_n28240_), .B(new_n12776_), .ZN(new_n28272_));
  NAND2_X1   g25031(.A1(new_n28251_), .A2(new_n28240_), .ZN(new_n28273_));
  NOR3_X1    g25032(.A1(new_n28273_), .A2(new_n12776_), .A3(new_n28247_), .ZN(new_n28274_));
  XNOR2_X1   g25033(.A1(new_n28274_), .A2(new_n28272_), .ZN(new_n28275_));
  NAND4_X1   g25034(.A1(new_n28271_), .A2(pi0644), .A3(new_n14200_), .A4(new_n28275_), .ZN(new_n28276_));
  AOI21_X1   g25035(.A1(new_n28261_), .A2(new_n28276_), .B(new_n14204_), .ZN(new_n28277_));
  NAND2_X1   g25036(.A1(pi0644), .A2(pi0715), .ZN(new_n28278_));
  NOR2_X1    g25037(.A1(new_n28269_), .A2(new_n28278_), .ZN(new_n28279_));
  OAI21_X1   g25038(.A1(new_n28279_), .A2(pi0644), .B(pi0790), .ZN(new_n28280_));
  NOR2_X1    g25039(.A1(new_n28261_), .A2(new_n28280_), .ZN(new_n28281_));
  NOR3_X1    g25040(.A1(new_n28277_), .A2(new_n28281_), .A3(new_n12775_), .ZN(new_n28282_));
  NOR2_X1    g25041(.A1(new_n27888_), .A2(new_n28233_), .ZN(new_n28283_));
  INV_X1     g25042(.I(new_n28236_), .ZN(new_n28284_));
  INV_X1     g25043(.I(new_n28256_), .ZN(new_n28285_));
  AOI22_X1   g25044(.A1(new_n28265_), .A2(new_n28266_), .B1(pi0787), .B2(new_n28285_), .ZN(new_n28286_));
  NAND2_X1   g25045(.A1(new_n28258_), .A2(new_n28195_), .ZN(new_n28287_));
  NOR2_X1    g25046(.A1(new_n28287_), .A2(new_n28286_), .ZN(new_n28288_));
  OAI21_X1   g25047(.A1(new_n28288_), .A2(new_n28284_), .B(new_n27946_), .ZN(new_n28289_));
  NOR2_X1    g25048(.A1(new_n28289_), .A2(new_n28283_), .ZN(new_n28290_));
  NAND3_X1   g25049(.A1(new_n28290_), .A2(pi0644), .A3(pi0790), .ZN(new_n28292_));
  NAND2_X1   g25050(.A1(new_n28292_), .A2(new_n7240_), .ZN(new_n28293_));
  OAI21_X1   g25051(.A1(new_n28282_), .A2(new_n28293_), .B(new_n28232_), .ZN(po0365));
  NOR2_X1    g25052(.A1(new_n14396_), .A2(new_n8345_), .ZN(new_n28295_));
  INV_X1     g25053(.I(pi0622), .ZN(new_n28296_));
  INV_X1     g25054(.I(pi0639), .ZN(new_n28297_));
  AOI21_X1   g25055(.A1(new_n14428_), .A2(pi0647), .B(new_n14209_), .ZN(new_n28298_));
  OAI21_X1   g25056(.A1(new_n28177_), .A2(pi0647), .B(new_n28298_), .ZN(new_n28299_));
  NOR2_X1    g25057(.A1(pi0647), .A2(pi1157), .ZN(new_n28300_));
  NAND2_X1   g25058(.A1(new_n28299_), .A2(new_n28300_), .ZN(new_n28301_));
  NOR2_X1    g25059(.A1(new_n13627_), .A2(new_n12776_), .ZN(new_n28302_));
  AOI21_X1   g25060(.A1(new_n28301_), .A2(new_n28302_), .B(pi1157), .ZN(new_n28303_));
  INV_X1     g25061(.I(new_n28177_), .ZN(new_n28304_));
  NOR3_X1    g25062(.A1(new_n28304_), .A2(new_n14010_), .A3(new_n14005_), .ZN(new_n28305_));
  NOR3_X1    g25063(.A1(new_n28177_), .A2(pi0630), .A3(new_n14005_), .ZN(new_n28306_));
  OAI21_X1   g25064(.A1(new_n28305_), .A2(new_n28306_), .B(new_n14428_), .ZN(new_n28307_));
  INV_X1     g25065(.I(new_n28307_), .ZN(new_n28308_));
  NOR2_X1    g25066(.A1(new_n14428_), .A2(pi0647), .ZN(new_n28309_));
  NOR4_X1    g25067(.A1(new_n28308_), .A2(new_n16419_), .A3(new_n28303_), .A4(new_n28309_), .ZN(new_n28310_));
  INV_X1     g25068(.I(new_n28310_), .ZN(new_n28311_));
  AOI21_X1   g25069(.A1(new_n27887_), .A2(new_n28311_), .B(new_n27947_), .ZN(new_n28312_));
  NOR2_X1    g25070(.A1(new_n13627_), .A2(new_n15402_), .ZN(new_n28313_));
  AOI21_X1   g25071(.A1(new_n28304_), .A2(new_n15402_), .B(new_n28313_), .ZN(new_n28314_));
  OAI21_X1   g25072(.A1(pi0715), .A2(pi1160), .B(new_n14204_), .ZN(new_n28315_));
  AOI22_X1   g25073(.A1(new_n28312_), .A2(new_n28315_), .B1(pi0790), .B2(new_n7240_), .ZN(new_n28316_));
  AOI21_X1   g25074(.A1(new_n28314_), .A2(new_n14204_), .B(new_n14200_), .ZN(new_n28317_));
  AOI21_X1   g25075(.A1(new_n14428_), .A2(new_n14200_), .B(new_n14203_), .ZN(new_n28318_));
  AOI21_X1   g25076(.A1(new_n28317_), .A2(new_n28318_), .B(pi0644), .ZN(new_n28319_));
  INV_X1     g25077(.I(new_n28319_), .ZN(new_n28320_));
  NAND2_X1   g25078(.A1(new_n28312_), .A2(new_n28320_), .ZN(new_n28321_));
  NOR4_X1    g25079(.A1(new_n28316_), .A2(new_n28296_), .A3(new_n28297_), .A4(new_n28321_), .ZN(new_n28322_));
  NOR2_X1    g25080(.A1(new_n28316_), .A2(new_n28321_), .ZN(new_n28323_));
  NOR3_X1    g25081(.A1(new_n28323_), .A2(pi0622), .A3(new_n28297_), .ZN(new_n28324_));
  OAI21_X1   g25082(.A1(new_n28324_), .A2(new_n28322_), .B(new_n28295_), .ZN(new_n28325_));
  AOI21_X1   g25083(.A1(new_n28158_), .A2(pi1157), .B(new_n14008_), .ZN(new_n28326_));
  INV_X1     g25084(.I(new_n28141_), .ZN(new_n28327_));
  INV_X1     g25085(.I(new_n28152_), .ZN(new_n28328_));
  NOR3_X1    g25086(.A1(new_n28128_), .A2(new_n13901_), .A3(new_n13922_), .ZN(new_n28329_));
  NOR3_X1    g25087(.A1(new_n28148_), .A2(pi0626), .A3(new_n13922_), .ZN(new_n28330_));
  OAI21_X1   g25088(.A1(new_n28329_), .A2(new_n28330_), .B(new_n28155_), .ZN(new_n28331_));
  OAI22_X1   g25089(.A1(new_n28328_), .A2(new_n28331_), .B1(new_n28129_), .B2(new_n28327_), .ZN(new_n28332_));
  NOR3_X1    g25090(.A1(new_n28332_), .A2(pi0647), .A3(new_n14006_), .ZN(new_n28333_));
  OAI21_X1   g25091(.A1(new_n28333_), .A2(new_n28326_), .B(new_n28162_), .ZN(new_n28334_));
  AOI21_X1   g25092(.A1(new_n28179_), .A2(new_n14012_), .B(new_n14005_), .ZN(new_n28335_));
  AOI21_X1   g25093(.A1(new_n28334_), .A2(new_n28335_), .B(new_n12776_), .ZN(new_n28336_));
  NAND3_X1   g25094(.A1(new_n28332_), .A2(pi0647), .A3(pi1157), .ZN(new_n28337_));
  NAND3_X1   g25095(.A1(new_n28158_), .A2(pi0647), .A3(new_n14006_), .ZN(new_n28338_));
  AOI21_X1   g25096(.A1(new_n28337_), .A2(new_n28338_), .B(new_n28163_), .ZN(new_n28339_));
  INV_X1     g25097(.I(new_n28335_), .ZN(new_n28340_));
  NOR3_X1    g25098(.A1(new_n28158_), .A2(new_n12776_), .A3(new_n28340_), .ZN(new_n28341_));
  INV_X1     g25099(.I(new_n28341_), .ZN(new_n28342_));
  NOR3_X1    g25100(.A1(new_n28336_), .A2(new_n28339_), .A3(new_n28342_), .ZN(new_n28343_));
  NAND3_X1   g25101(.A1(new_n28332_), .A2(pi0647), .A3(pi1157), .ZN(new_n28344_));
  NAND3_X1   g25102(.A1(new_n28158_), .A2(new_n14005_), .A3(pi1157), .ZN(new_n28345_));
  AOI21_X1   g25103(.A1(new_n28344_), .A2(new_n28345_), .B(new_n28163_), .ZN(new_n28346_));
  OAI21_X1   g25104(.A1(new_n28346_), .A2(new_n28340_), .B(pi0787), .ZN(new_n28347_));
  NAND2_X1   g25105(.A1(new_n28337_), .A2(new_n28338_), .ZN(new_n28348_));
  AOI21_X1   g25106(.A1(new_n28348_), .A2(new_n28162_), .B(new_n28342_), .ZN(new_n28349_));
  NOR2_X1    g25107(.A1(new_n28347_), .A2(new_n28349_), .ZN(new_n28350_));
  NAND2_X1   g25108(.A1(new_n28137_), .A2(new_n18804_), .ZN(new_n28351_));
  AOI21_X1   g25109(.A1(new_n28179_), .A2(new_n14217_), .B(new_n15402_), .ZN(new_n28352_));
  NAND2_X1   g25110(.A1(new_n28352_), .A2(pi0644), .ZN(new_n28353_));
  AOI21_X1   g25111(.A1(new_n28351_), .A2(new_n15385_), .B(new_n28353_), .ZN(new_n28354_));
  NOR3_X1    g25112(.A1(new_n28343_), .A2(new_n28350_), .A3(new_n28354_), .ZN(new_n28355_));
  NOR2_X1    g25113(.A1(new_n28343_), .A2(new_n28350_), .ZN(new_n28356_));
  NAND2_X1   g25114(.A1(new_n7240_), .A2(pi0790), .ZN(new_n28357_));
  OAI21_X1   g25115(.A1(new_n28355_), .A2(new_n14204_), .B(new_n28357_), .ZN(new_n28358_));
  NAND3_X1   g25116(.A1(new_n28351_), .A2(new_n14204_), .A3(new_n14203_), .ZN(new_n28359_));
  INV_X1     g25117(.I(new_n28352_), .ZN(new_n28360_));
  NOR2_X1    g25118(.A1(new_n28360_), .A2(new_n14200_), .ZN(new_n28361_));
  AOI21_X1   g25119(.A1(new_n28359_), .A2(new_n28361_), .B(pi0644), .ZN(new_n28362_));
  NOR2_X1    g25120(.A1(new_n28356_), .A2(new_n28362_), .ZN(new_n28363_));
  INV_X1     g25121(.I(pi0209), .ZN(new_n28364_));
  OAI21_X1   g25122(.A1(new_n14007_), .A2(new_n28300_), .B(new_n14210_), .ZN(new_n28365_));
  OAI22_X1   g25123(.A1(new_n27931_), .A2(new_n28179_), .B1(new_n16419_), .B2(new_n28365_), .ZN(new_n28366_));
  AOI21_X1   g25124(.A1(new_n28360_), .A2(new_n14203_), .B(new_n14204_), .ZN(new_n28367_));
  NAND2_X1   g25125(.A1(new_n28366_), .A2(new_n28367_), .ZN(new_n28368_));
  NAND2_X1   g25126(.A1(new_n28366_), .A2(new_n12775_), .ZN(new_n28369_));
  NAND2_X1   g25127(.A1(new_n28369_), .A2(new_n7240_), .ZN(new_n28370_));
  AOI21_X1   g25128(.A1(new_n28366_), .A2(new_n28367_), .B(pi0790), .ZN(new_n28371_));
  AOI21_X1   g25129(.A1(new_n28370_), .A2(new_n28371_), .B(new_n28368_), .ZN(new_n28372_));
  NAND2_X1   g25130(.A1(new_n14204_), .A2(pi1160), .ZN(new_n28373_));
  NAND2_X1   g25131(.A1(new_n14203_), .A2(pi0644), .ZN(new_n28374_));
  AOI21_X1   g25132(.A1(new_n28373_), .A2(new_n28374_), .B(new_n12775_), .ZN(new_n28375_));
  NOR3_X1    g25133(.A1(new_n28351_), .A2(po1038), .A3(new_n28375_), .ZN(new_n28376_));
  AOI21_X1   g25134(.A1(new_n28296_), .A2(new_n28297_), .B(new_n28364_), .ZN(new_n28377_));
  NAND3_X1   g25135(.A1(new_n28358_), .A2(new_n28363_), .A3(new_n28377_), .ZN(new_n28378_));
  NOR2_X1    g25136(.A1(new_n13627_), .A2(pi0644), .ZN(new_n28379_));
  NAND2_X1   g25137(.A1(new_n14428_), .A2(new_n14210_), .ZN(new_n28380_));
  OAI21_X1   g25138(.A1(new_n28168_), .A2(new_n14210_), .B(new_n28380_), .ZN(new_n28381_));
  AOI21_X1   g25139(.A1(new_n28381_), .A2(pi0644), .B(new_n28379_), .ZN(new_n28382_));
  INV_X1     g25140(.I(new_n28382_), .ZN(new_n28383_));
  NOR2_X1    g25141(.A1(new_n13627_), .A2(new_n14204_), .ZN(new_n28384_));
  AOI21_X1   g25142(.A1(new_n28381_), .A2(new_n14204_), .B(new_n28384_), .ZN(new_n28385_));
  NOR3_X1    g25143(.A1(new_n28385_), .A2(new_n12775_), .A3(new_n14203_), .ZN(new_n28386_));
  AND3_X2    g25144(.A1(new_n28385_), .A2(pi0790), .A3(new_n14203_), .Z(new_n28387_));
  OAI21_X1   g25145(.A1(new_n28387_), .A2(new_n28386_), .B(new_n28383_), .ZN(new_n28388_));
  NAND2_X1   g25146(.A1(new_n28381_), .A2(pi0790), .ZN(new_n28389_));
  AOI21_X1   g25147(.A1(new_n28388_), .A2(new_n7240_), .B(new_n28389_), .ZN(new_n28390_));
  NAND2_X1   g25148(.A1(new_n28299_), .A2(new_n16574_), .ZN(new_n28391_));
  AOI21_X1   g25149(.A1(new_n28308_), .A2(pi1157), .B(new_n28391_), .ZN(new_n28392_));
  OAI21_X1   g25150(.A1(new_n28170_), .A2(new_n16576_), .B(new_n28392_), .ZN(new_n28393_));
  NAND3_X1   g25151(.A1(new_n28085_), .A2(new_n28032_), .A3(pi0787), .ZN(new_n28394_));
  NAND2_X1   g25152(.A1(new_n28394_), .A2(new_n28393_), .ZN(new_n28395_));
  OAI21_X1   g25153(.A1(pi0715), .A2(pi1160), .B(new_n14204_), .ZN(new_n28396_));
  NOR2_X1    g25154(.A1(po1038), .A2(new_n12775_), .ZN(new_n28398_));
  AOI21_X1   g25155(.A1(new_n28395_), .A2(new_n28396_), .B(new_n28398_), .ZN(new_n28399_));
  INV_X1     g25156(.I(new_n28393_), .ZN(new_n28400_));
  NOR3_X1    g25157(.A1(new_n28017_), .A2(new_n13860_), .A3(new_n13855_), .ZN(new_n28401_));
  NOR3_X1    g25158(.A1(new_n28009_), .A2(new_n13860_), .A3(pi0781), .ZN(new_n28402_));
  NOR2_X1    g25159(.A1(new_n28401_), .A2(new_n28402_), .ZN(new_n28403_));
  OAI22_X1   g25160(.A1(new_n28403_), .A2(new_n27984_), .B1(new_n14538_), .B2(new_n28028_), .ZN(new_n28404_));
  AOI21_X1   g25161(.A1(new_n28404_), .A2(new_n28030_), .B(pi0789), .ZN(new_n28405_));
  NAND2_X1   g25162(.A1(new_n28081_), .A2(new_n13903_), .ZN(new_n28406_));
  NAND3_X1   g25163(.A1(new_n28079_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n28407_));
  NAND2_X1   g25164(.A1(new_n28407_), .A2(new_n28406_), .ZN(new_n28408_));
  NAND3_X1   g25165(.A1(new_n28408_), .A2(new_n28077_), .A3(new_n28083_), .ZN(new_n28409_));
  NOR3_X1    g25166(.A1(new_n28405_), .A2(new_n28409_), .A3(new_n12776_), .ZN(new_n28410_));
  NAND2_X1   g25167(.A1(new_n28314_), .A2(new_n14204_), .ZN(new_n28411_));
  NAND3_X1   g25168(.A1(new_n28411_), .A2(pi0715), .A3(pi1160), .ZN(new_n28412_));
  NAND2_X1   g25169(.A1(new_n28412_), .A2(new_n14204_), .ZN(new_n28413_));
  OAI21_X1   g25170(.A1(new_n28410_), .A2(new_n28400_), .B(new_n28413_), .ZN(new_n28414_));
  NOR4_X1    g25171(.A1(new_n28399_), .A2(new_n28296_), .A3(new_n28297_), .A4(new_n28414_), .ZN(new_n28415_));
  OAI21_X1   g25172(.A1(new_n28410_), .A2(new_n28400_), .B(new_n28396_), .ZN(new_n28416_));
  INV_X1     g25173(.I(new_n28398_), .ZN(new_n28417_));
  AOI21_X1   g25174(.A1(new_n28416_), .A2(new_n28417_), .B(new_n28414_), .ZN(new_n28418_));
  NOR3_X1    g25175(.A1(new_n28418_), .A2(new_n28296_), .A3(pi0639), .ZN(new_n28419_));
  OAI21_X1   g25176(.A1(new_n28419_), .A2(new_n28415_), .B(new_n28390_), .ZN(new_n28420_));
  AOI21_X1   g25177(.A1(new_n28325_), .A2(new_n28378_), .B(new_n28420_), .ZN(po0366));
  NOR2_X1    g25178(.A1(new_n5800_), .A2(pi0634), .ZN(new_n28422_));
  NAND3_X1   g25179(.A1(pi0633), .A2(pi0907), .A3(pi0947), .ZN(new_n28423_));
  XOR2_X1    g25180(.A1(new_n28422_), .A2(new_n28423_), .Z(new_n28424_));
  INV_X1     g25181(.I(new_n28424_), .ZN(new_n28425_));
  NOR2_X1    g25182(.A1(new_n28425_), .A2(new_n3259_), .ZN(new_n28426_));
  XOR2_X1    g25183(.A1(new_n13723_), .A2(new_n28426_), .Z(new_n28427_));
  AOI21_X1   g25184(.A1(new_n28427_), .A2(pi0210), .B(new_n8345_), .ZN(new_n28428_));
  NOR2_X1    g25185(.A1(new_n12784_), .A2(pi0210), .ZN(new_n28429_));
  AOI21_X1   g25186(.A1(new_n12784_), .A2(new_n28425_), .B(new_n28429_), .ZN(new_n28430_));
  NOR2_X1    g25187(.A1(new_n14316_), .A2(new_n2777_), .ZN(new_n28431_));
  NAND2_X1   g25188(.A1(new_n28431_), .A2(new_n5741_), .ZN(new_n28432_));
  INV_X1     g25189(.I(new_n28429_), .ZN(new_n28433_));
  OAI21_X1   g25190(.A1(pi0633), .A2(new_n12809_), .B(new_n28433_), .ZN(new_n28434_));
  NOR2_X1    g25191(.A1(new_n12818_), .A2(pi0210), .ZN(new_n28435_));
  AOI21_X1   g25192(.A1(new_n26463_), .A2(new_n12818_), .B(new_n28435_), .ZN(new_n28436_));
  NAND2_X1   g25193(.A1(new_n28436_), .A2(pi0947), .ZN(new_n28437_));
  NOR2_X1    g25194(.A1(new_n7611_), .A2(new_n5800_), .ZN(new_n28438_));
  XNOR2_X1   g25195(.A1(new_n28437_), .A2(new_n28438_), .ZN(new_n28439_));
  NAND2_X1   g25196(.A1(new_n28439_), .A2(new_n28434_), .ZN(new_n28440_));
  AOI21_X1   g25197(.A1(new_n26624_), .A2(new_n12784_), .B(new_n28429_), .ZN(new_n28441_));
  INV_X1     g25198(.I(new_n28441_), .ZN(new_n28442_));
  NOR2_X1    g25199(.A1(new_n28435_), .A2(new_n5741_), .ZN(new_n28443_));
  OAI21_X1   g25200(.A1(pi0634), .A2(new_n12806_), .B(new_n28443_), .ZN(new_n28444_));
  NOR2_X1    g25201(.A1(new_n7611_), .A2(new_n5741_), .ZN(new_n28445_));
  INV_X1     g25202(.I(new_n28445_), .ZN(new_n28446_));
  XOR2_X1    g25203(.A1(new_n28444_), .A2(new_n28446_), .Z(new_n28447_));
  NAND2_X1   g25204(.A1(new_n28447_), .A2(new_n28442_), .ZN(new_n28448_));
  NAND2_X1   g25205(.A1(new_n28448_), .A2(pi0947), .ZN(new_n28449_));
  AOI21_X1   g25206(.A1(new_n28440_), .A2(new_n5397_), .B(new_n28449_), .ZN(new_n28450_));
  OAI21_X1   g25207(.A1(new_n28434_), .A2(new_n5386_), .B(po1101), .ZN(new_n28451_));
  AOI21_X1   g25208(.A1(new_n28434_), .A2(new_n5384_), .B(new_n5800_), .ZN(new_n28452_));
  AOI21_X1   g25209(.A1(new_n28452_), .A2(new_n28451_), .B(new_n5373_), .ZN(new_n28453_));
  OAI21_X1   g25210(.A1(new_n28453_), .A2(new_n28436_), .B(new_n5397_), .ZN(new_n28454_));
  AOI21_X1   g25211(.A1(new_n28450_), .A2(new_n28432_), .B(new_n28454_), .ZN(new_n28455_));
  NOR2_X1    g25212(.A1(new_n6448_), .A2(new_n5741_), .ZN(new_n28456_));
  XOR2_X1    g25213(.A1(new_n28444_), .A2(new_n28456_), .Z(new_n28457_));
  OAI21_X1   g25214(.A1(new_n28457_), .A2(new_n28441_), .B(new_n5800_), .ZN(new_n28458_));
  NAND3_X1   g25215(.A1(new_n12949_), .A2(pi0210), .A3(po1101), .ZN(new_n28459_));
  NAND3_X1   g25216(.A1(new_n12945_), .A2(pi0210), .A3(new_n5384_), .ZN(new_n28460_));
  AOI21_X1   g25217(.A1(new_n28459_), .A2(new_n28460_), .B(new_n12809_), .ZN(new_n28461_));
  NAND3_X1   g25218(.A1(new_n28458_), .A2(pi0907), .A3(new_n28461_), .ZN(new_n28462_));
  OAI21_X1   g25219(.A1(new_n28455_), .A2(new_n28462_), .B(new_n3091_), .ZN(new_n28463_));
  XOR2_X1    g25220(.A1(new_n28463_), .A2(new_n13412_), .Z(new_n28464_));
  NOR2_X1    g25221(.A1(new_n28464_), .A2(new_n28430_), .ZN(new_n28465_));
  NOR2_X1    g25222(.A1(new_n5398_), .A2(pi0223), .ZN(new_n28466_));
  NOR2_X1    g25223(.A1(new_n12878_), .A2(pi0634), .ZN(new_n28467_));
  NOR2_X1    g25224(.A1(new_n12862_), .A2(pi0210), .ZN(new_n28468_));
  NOR3_X1    g25225(.A1(new_n28467_), .A2(new_n28468_), .A3(new_n5741_), .ZN(new_n28469_));
  XOR2_X1    g25226(.A1(new_n28469_), .A2(new_n28456_), .Z(new_n28470_));
  AOI21_X1   g25227(.A1(new_n28470_), .A2(new_n28442_), .B(pi0947), .ZN(new_n28471_));
  NAND3_X1   g25228(.A1(new_n13334_), .A2(pi0210), .A3(po1101), .ZN(new_n28472_));
  NAND3_X1   g25229(.A1(new_n12890_), .A2(pi0210), .A3(new_n5384_), .ZN(new_n28473_));
  NAND2_X1   g25230(.A1(new_n28472_), .A2(new_n28473_), .ZN(new_n28474_));
  NAND3_X1   g25231(.A1(new_n28474_), .A2(pi0907), .A3(new_n12784_), .ZN(new_n28475_));
  OAI21_X1   g25232(.A1(new_n28471_), .A2(new_n28475_), .B(new_n28466_), .ZN(new_n28476_));
  AOI21_X1   g25233(.A1(new_n26463_), .A2(new_n12862_), .B(new_n28468_), .ZN(new_n28477_));
  NOR2_X1    g25234(.A1(new_n28453_), .A2(new_n28477_), .ZN(new_n28478_));
  NAND2_X1   g25235(.A1(new_n28477_), .A2(pi0947), .ZN(new_n28479_));
  XNOR2_X1   g25236(.A1(new_n28479_), .A2(new_n28438_), .ZN(new_n28480_));
  NAND2_X1   g25237(.A1(new_n28480_), .A2(new_n28434_), .ZN(new_n28481_));
  NAND2_X1   g25238(.A1(new_n28481_), .A2(new_n5397_), .ZN(new_n28482_));
  AOI21_X1   g25239(.A1(new_n28476_), .A2(new_n28478_), .B(new_n28482_), .ZN(new_n28483_));
  OR2_X2     g25240(.A1(new_n28469_), .A2(new_n28446_), .Z(new_n28484_));
  NAND2_X1   g25241(.A1(new_n28469_), .A2(new_n28446_), .ZN(new_n28485_));
  AOI21_X1   g25242(.A1(new_n28484_), .A2(new_n28485_), .B(new_n28441_), .ZN(new_n28486_));
  INV_X1     g25243(.I(new_n28486_), .ZN(new_n28487_));
  NOR2_X1    g25244(.A1(new_n7611_), .A2(new_n2723_), .ZN(new_n28488_));
  AOI21_X1   g25245(.A1(new_n28488_), .A2(new_n13677_), .B(new_n2777_), .ZN(new_n28489_));
  NAND2_X1   g25246(.A1(new_n12878_), .A2(new_n28489_), .ZN(new_n28490_));
  NAND2_X1   g25247(.A1(new_n28487_), .A2(new_n28490_), .ZN(new_n28491_));
  NAND2_X1   g25248(.A1(new_n28491_), .A2(new_n5800_), .ZN(new_n28492_));
  OAI21_X1   g25249(.A1(new_n28483_), .A2(new_n28492_), .B(new_n3098_), .ZN(new_n28493_));
  NAND2_X1   g25250(.A1(new_n13162_), .A2(new_n28424_), .ZN(new_n28494_));
  XNOR2_X1   g25251(.A1(new_n13163_), .A2(new_n28494_), .ZN(new_n28495_));
  OAI21_X1   g25252(.A1(new_n28495_), .A2(new_n2777_), .B(new_n3211_), .ZN(new_n28496_));
  AOI21_X1   g25253(.A1(pi0299), .A2(new_n28425_), .B(new_n13063_), .ZN(new_n28497_));
  NOR3_X1    g25254(.A1(new_n28497_), .A2(new_n2777_), .A3(new_n13176_), .ZN(new_n28498_));
  AOI21_X1   g25255(.A1(new_n28496_), .A2(new_n28498_), .B(pi0039), .ZN(new_n28499_));
  OAI21_X1   g25256(.A1(new_n28465_), .A2(new_n28493_), .B(new_n28499_), .ZN(new_n28500_));
  OAI21_X1   g25257(.A1(new_n28448_), .A2(pi0907), .B(new_n5451_), .ZN(new_n28501_));
  NAND2_X1   g25258(.A1(new_n28440_), .A2(new_n3313_), .ZN(new_n28502_));
  NAND4_X1   g25259(.A1(new_n28501_), .A2(new_n28502_), .A3(pi0947), .A4(new_n28431_), .ZN(new_n28503_));
  NAND2_X1   g25260(.A1(new_n28503_), .A2(new_n3111_), .ZN(new_n28504_));
  NOR2_X1    g25261(.A1(new_n28430_), .A2(new_n3313_), .ZN(new_n28505_));
  NAND2_X1   g25262(.A1(new_n28504_), .A2(new_n28505_), .ZN(new_n28506_));
  NAND2_X1   g25263(.A1(new_n28506_), .A2(new_n3098_), .ZN(new_n28507_));
  AOI21_X1   g25264(.A1(new_n28474_), .A2(new_n12784_), .B(new_n5451_), .ZN(new_n28508_));
  NAND2_X1   g25265(.A1(new_n13077_), .A2(pi0907), .ZN(new_n28509_));
  XOR2_X1    g25266(.A1(new_n28508_), .A2(new_n28509_), .Z(new_n28510_));
  OAI22_X1   g25267(.A1(new_n28510_), .A2(new_n28490_), .B1(new_n5800_), .B2(new_n28481_), .ZN(new_n28511_));
  NOR4_X1    g25268(.A1(new_n28487_), .A2(new_n2777_), .A3(new_n3111_), .A4(new_n8345_), .ZN(new_n28512_));
  NAND4_X1   g25269(.A1(new_n28500_), .A2(new_n28507_), .A3(new_n28511_), .A4(new_n28512_), .ZN(new_n28513_));
  XNOR2_X1   g25270(.A1(new_n28513_), .A2(new_n28428_), .ZN(po0367));
  NOR2_X1    g25271(.A1(new_n17466_), .A2(new_n3290_), .ZN(new_n28515_));
  NOR2_X1    g25272(.A1(new_n17464_), .A2(new_n3290_), .ZN(new_n28516_));
  INV_X1     g25273(.I(new_n28516_), .ZN(new_n28517_));
  NOR3_X1    g25274(.A1(new_n28517_), .A2(new_n27261_), .A3(new_n27295_), .ZN(new_n28518_));
  NOR3_X1    g25275(.A1(new_n28516_), .A2(pi0606), .A3(new_n27295_), .ZN(new_n28519_));
  OAI21_X1   g25276(.A1(new_n28518_), .A2(new_n28519_), .B(new_n28515_), .ZN(new_n28520_));
  NAND2_X1   g25277(.A1(new_n17098_), .A2(new_n3289_), .ZN(new_n28521_));
  NAND3_X1   g25278(.A1(new_n28520_), .A2(new_n27261_), .A3(new_n28521_), .ZN(new_n28522_));
  AOI21_X1   g25279(.A1(new_n28522_), .A2(pi0643), .B(new_n8684_), .ZN(po0368));
  NOR3_X1    g25280(.A1(new_n28517_), .A2(new_n28263_), .A3(new_n28243_), .ZN(new_n28524_));
  NOR3_X1    g25281(.A1(new_n28516_), .A2(pi0607), .A3(new_n28243_), .ZN(new_n28525_));
  OAI21_X1   g25282(.A1(new_n28524_), .A2(new_n28525_), .B(new_n28515_), .ZN(new_n28526_));
  NAND3_X1   g25283(.A1(new_n28526_), .A2(new_n28263_), .A3(new_n28521_), .ZN(new_n28527_));
  AOI21_X1   g25284(.A1(new_n28527_), .A2(pi0638), .B(new_n8739_), .ZN(po0369));
  INV_X1     g25285(.I(pi0213), .ZN(new_n28529_));
  NOR3_X1    g25286(.A1(new_n28517_), .A2(new_n28296_), .A3(new_n28297_), .ZN(new_n28530_));
  NOR3_X1    g25287(.A1(new_n28516_), .A2(pi0622), .A3(new_n28297_), .ZN(new_n28531_));
  OAI21_X1   g25288(.A1(new_n28530_), .A2(new_n28531_), .B(new_n28515_), .ZN(new_n28532_));
  NAND3_X1   g25289(.A1(new_n28532_), .A2(new_n28296_), .A3(new_n28521_), .ZN(new_n28533_));
  AOI21_X1   g25290(.A1(new_n28533_), .A2(pi0639), .B(new_n28529_), .ZN(po0370));
  NOR3_X1    g25291(.A1(new_n28517_), .A2(new_n28200_), .A3(new_n28176_), .ZN(new_n28535_));
  NOR3_X1    g25292(.A1(new_n28516_), .A2(pi0623), .A3(new_n28176_), .ZN(new_n28536_));
  OAI21_X1   g25293(.A1(new_n28535_), .A2(new_n28536_), .B(new_n28515_), .ZN(new_n28537_));
  NAND3_X1   g25294(.A1(new_n28537_), .A2(new_n28200_), .A3(new_n28521_), .ZN(new_n28538_));
  AOI21_X1   g25295(.A1(new_n28538_), .A2(pi0710), .B(new_n8685_), .ZN(po0371));
  NOR2_X1    g25296(.A1(new_n5632_), .A2(new_n5741_), .ZN(new_n28540_));
  NOR2_X1    g25297(.A1(new_n28540_), .A2(pi0947), .ZN(new_n28541_));
  AOI21_X1   g25298(.A1(new_n5379_), .A2(pi0947), .B(new_n28541_), .ZN(new_n28542_));
  NAND2_X1   g25299(.A1(new_n28542_), .A2(pi0038), .ZN(new_n28543_));
  XNOR2_X1   g25300(.A1(new_n13723_), .A2(new_n28543_), .ZN(new_n28544_));
  AOI21_X1   g25301(.A1(new_n28544_), .A2(pi0215), .B(new_n8345_), .ZN(new_n28545_));
  NAND2_X1   g25302(.A1(new_n12809_), .A2(new_n13464_), .ZN(new_n28546_));
  INV_X1     g25303(.I(new_n28546_), .ZN(new_n28547_));
  OAI21_X1   g25304(.A1(new_n12931_), .A2(pi0947), .B(new_n12930_), .ZN(new_n28548_));
  NAND2_X1   g25305(.A1(new_n28548_), .A2(new_n5397_), .ZN(new_n28549_));
  INV_X1     g25306(.I(new_n12864_), .ZN(new_n28550_));
  AOI21_X1   g25307(.A1(new_n5379_), .A2(new_n12845_), .B(new_n12848_), .ZN(new_n28551_));
  OAI21_X1   g25308(.A1(new_n12846_), .A2(new_n5379_), .B(new_n5800_), .ZN(new_n28552_));
  NAND3_X1   g25309(.A1(new_n28550_), .A2(new_n28551_), .A3(new_n28552_), .ZN(new_n28553_));
  AND3_X2    g25310(.A1(new_n28549_), .A2(new_n3090_), .A3(new_n28553_), .Z(new_n28554_));
  INV_X1     g25311(.I(new_n28540_), .ZN(new_n28555_));
  NOR2_X1    g25312(.A1(new_n12927_), .A2(new_n5397_), .ZN(new_n28556_));
  OAI21_X1   g25313(.A1(new_n28556_), .A2(new_n28555_), .B(new_n17067_), .ZN(new_n28557_));
  OAI22_X1   g25314(.A1(new_n28554_), .A2(new_n28557_), .B1(new_n28542_), .B2(new_n28547_), .ZN(new_n28558_));
  NOR2_X1    g25315(.A1(new_n12949_), .A2(new_n5375_), .ZN(new_n28559_));
  NOR3_X1    g25316(.A1(new_n12846_), .A2(new_n5379_), .A3(new_n5800_), .ZN(new_n28560_));
  OAI21_X1   g25317(.A1(new_n28551_), .A2(new_n28560_), .B(new_n28559_), .ZN(new_n28561_));
  NAND2_X1   g25318(.A1(new_n28540_), .A2(new_n5800_), .ZN(new_n28562_));
  AOI21_X1   g25319(.A1(new_n28561_), .A2(new_n5397_), .B(new_n28562_), .ZN(new_n28563_));
  AOI21_X1   g25320(.A1(new_n28563_), .A2(new_n12960_), .B(new_n3091_), .ZN(new_n28564_));
  AOI21_X1   g25321(.A1(new_n13262_), .A2(new_n5636_), .B(new_n13416_), .ZN(new_n28565_));
  NOR3_X1    g25322(.A1(new_n28565_), .A2(new_n5379_), .A3(new_n12845_), .ZN(new_n28566_));
  NOR2_X1    g25323(.A1(new_n28566_), .A2(new_n5800_), .ZN(new_n28567_));
  NOR4_X1    g25324(.A1(new_n12844_), .A2(new_n28555_), .A3(new_n5379_), .A4(new_n5800_), .ZN(new_n28568_));
  NAND3_X1   g25325(.A1(new_n12826_), .A2(new_n13262_), .A3(new_n28568_), .ZN(new_n28569_));
  XNOR2_X1   g25326(.A1(new_n28567_), .A2(new_n28569_), .ZN(new_n28570_));
  NAND2_X1   g25327(.A1(new_n28570_), .A2(new_n5398_), .ZN(new_n28571_));
  NOR2_X1    g25328(.A1(new_n28571_), .A2(new_n28564_), .ZN(new_n28572_));
  AOI21_X1   g25329(.A1(new_n28572_), .A2(new_n28558_), .B(new_n3111_), .ZN(new_n28573_));
  OAI21_X1   g25330(.A1(new_n13413_), .A2(new_n28542_), .B(new_n3092_), .ZN(new_n28574_));
  AOI21_X1   g25331(.A1(new_n17298_), .A2(new_n28541_), .B(new_n28574_), .ZN(new_n28575_));
  NAND4_X1   g25332(.A1(new_n12949_), .A2(pi0642), .A3(pi0947), .A4(new_n5397_), .ZN(new_n28576_));
  OAI21_X1   g25333(.A1(new_n28575_), .A2(new_n28576_), .B(pi0299), .ZN(new_n28577_));
  NOR2_X1    g25334(.A1(new_n12843_), .A2(new_n5634_), .ZN(new_n28578_));
  NAND2_X1   g25335(.A1(new_n12878_), .A2(new_n28578_), .ZN(new_n28579_));
  NAND2_X1   g25336(.A1(new_n28579_), .A2(new_n5379_), .ZN(new_n28580_));
  NAND2_X1   g25337(.A1(new_n28580_), .A2(new_n5378_), .ZN(new_n28581_));
  OAI21_X1   g25338(.A1(new_n12932_), .A2(new_n28581_), .B(pi0947), .ZN(new_n28582_));
  NOR3_X1    g25339(.A1(new_n13080_), .A2(pi0947), .A3(new_n16977_), .ZN(new_n28583_));
  NAND2_X1   g25340(.A1(new_n28583_), .A2(pi0947), .ZN(new_n28584_));
  XOR2_X1    g25341(.A1(new_n28584_), .A2(new_n28582_), .Z(new_n28585_));
  NAND2_X1   g25342(.A1(new_n5398_), .A2(pi0947), .ZN(new_n28586_));
  XOR2_X1    g25343(.A1(new_n28582_), .A2(new_n28586_), .Z(new_n28587_));
  NAND3_X1   g25344(.A1(new_n12927_), .A2(pi0642), .A3(new_n5378_), .ZN(new_n28588_));
  NAND3_X1   g25345(.A1(new_n12898_), .A2(new_n5379_), .A3(new_n5378_), .ZN(new_n28589_));
  NAND2_X1   g25346(.A1(new_n28540_), .A2(pi0299), .ZN(new_n28590_));
  AOI21_X1   g25347(.A1(new_n3090_), .A2(new_n28562_), .B(new_n28590_), .ZN(new_n28591_));
  NAND2_X1   g25348(.A1(new_n13334_), .A2(new_n28591_), .ZN(new_n28592_));
  AOI21_X1   g25349(.A1(new_n28589_), .A2(new_n28588_), .B(new_n28592_), .ZN(new_n28593_));
  NAND4_X1   g25350(.A1(new_n28585_), .A2(new_n17046_), .A3(new_n28587_), .A4(new_n28593_), .ZN(new_n28594_));
  XOR2_X1    g25351(.A1(new_n28594_), .A2(new_n28577_), .Z(new_n28595_));
  NAND2_X1   g25352(.A1(new_n28570_), .A2(new_n3313_), .ZN(new_n28596_));
  NAND2_X1   g25353(.A1(new_n13343_), .A2(new_n28542_), .ZN(new_n28597_));
  NAND4_X1   g25354(.A1(new_n28595_), .A2(new_n3695_), .A3(new_n28596_), .A4(new_n28597_), .ZN(new_n28598_));
  AND2_X2    g25355(.A1(new_n28598_), .A2(new_n28573_), .Z(new_n28599_));
  OAI21_X1   g25356(.A1(new_n28598_), .A2(new_n28573_), .B(pi0039), .ZN(new_n28600_));
  NAND2_X1   g25357(.A1(new_n28542_), .A2(pi0299), .ZN(new_n28601_));
  XOR2_X1    g25358(.A1(new_n13069_), .A2(new_n28601_), .Z(new_n28602_));
  AOI21_X1   g25359(.A1(new_n28602_), .A2(pi0215), .B(new_n3212_), .ZN(new_n28603_));
  NAND2_X1   g25360(.A1(new_n13162_), .A2(new_n28542_), .ZN(new_n28604_));
  XNOR2_X1   g25361(.A1(new_n13163_), .A2(new_n28604_), .ZN(new_n28605_));
  NOR4_X1    g25362(.A1(new_n28603_), .A2(new_n3111_), .A3(new_n8345_), .A4(new_n28605_), .ZN(new_n28606_));
  OAI21_X1   g25363(.A1(new_n28599_), .A2(new_n28600_), .B(new_n28606_), .ZN(new_n28607_));
  XNOR2_X1   g25364(.A1(new_n28607_), .A2(new_n28545_), .ZN(po0372));
  NOR2_X1    g25365(.A1(new_n16969_), .A2(new_n5633_), .ZN(new_n28609_));
  NOR2_X1    g25366(.A1(new_n12868_), .A2(new_n5800_), .ZN(new_n28610_));
  NOR2_X1    g25367(.A1(new_n28609_), .A2(new_n28610_), .ZN(new_n28611_));
  NOR2_X1    g25368(.A1(new_n28611_), .A2(new_n3259_), .ZN(new_n28612_));
  XOR2_X1    g25369(.A1(new_n13723_), .A2(new_n28612_), .Z(new_n28613_));
  AOI21_X1   g25370(.A1(new_n28613_), .A2(pi0216), .B(new_n8345_), .ZN(new_n28614_));
  INV_X1     g25371(.I(new_n28583_), .ZN(new_n28615_));
  NAND4_X1   g25372(.A1(new_n12930_), .A2(new_n12868_), .A3(new_n12841_), .A4(new_n5795_), .ZN(new_n28616_));
  NOR2_X1    g25373(.A1(new_n28616_), .A2(new_n12862_), .ZN(new_n28617_));
  INV_X1     g25374(.I(new_n28617_), .ZN(new_n28618_));
  NOR3_X1    g25375(.A1(new_n28618_), .A2(new_n12868_), .A3(new_n5636_), .ZN(new_n28619_));
  NOR3_X1    g25376(.A1(new_n28617_), .A2(pi0614), .A3(new_n5636_), .ZN(new_n28620_));
  OAI21_X1   g25377(.A1(new_n28619_), .A2(new_n28620_), .B(new_n12878_), .ZN(new_n28621_));
  OAI21_X1   g25378(.A1(new_n28609_), .A2(pi0216), .B(pi0947), .ZN(new_n28622_));
  NOR2_X1    g25379(.A1(new_n28621_), .A2(new_n28622_), .ZN(new_n28623_));
  NAND2_X1   g25380(.A1(pi0662), .A2(pi0907), .ZN(new_n28624_));
  OAI21_X1   g25381(.A1(new_n12932_), .A2(new_n28624_), .B(pi0947), .ZN(new_n28625_));
  NOR2_X1    g25382(.A1(new_n12809_), .A2(new_n5375_), .ZN(new_n28626_));
  NAND2_X1   g25383(.A1(new_n12961_), .A2(new_n5800_), .ZN(new_n28627_));
  NAND4_X1   g25384(.A1(new_n28550_), .A2(new_n28626_), .A3(new_n12962_), .A4(new_n28627_), .ZN(new_n28628_));
  NOR2_X1    g25385(.A1(new_n28628_), .A2(new_n5800_), .ZN(new_n28629_));
  XOR2_X1    g25386(.A1(new_n28625_), .A2(new_n28629_), .Z(new_n28630_));
  OAI21_X1   g25387(.A1(new_n28630_), .A2(new_n12930_), .B(new_n3011_), .ZN(new_n28631_));
  AOI21_X1   g25388(.A1(new_n28631_), .A2(new_n3695_), .B(new_n28623_), .ZN(new_n28632_));
  OAI21_X1   g25389(.A1(new_n13417_), .A2(pi0614), .B(pi0947), .ZN(new_n28633_));
  NOR3_X1    g25390(.A1(new_n5398_), .A2(new_n28609_), .A3(new_n3092_), .ZN(new_n28634_));
  AOI21_X1   g25391(.A1(new_n28633_), .A2(new_n28634_), .B(pi0947), .ZN(new_n28635_));
  NOR3_X1    g25392(.A1(new_n28609_), .A2(new_n3011_), .A3(new_n3090_), .ZN(new_n28636_));
  NOR2_X1    g25393(.A1(new_n17046_), .A2(new_n28636_), .ZN(new_n28637_));
  NAND2_X1   g25394(.A1(new_n28621_), .A2(pi0947), .ZN(new_n28638_));
  XOR2_X1    g25395(.A1(new_n28638_), .A2(new_n28586_), .Z(new_n28639_));
  NOR2_X1    g25396(.A1(new_n12884_), .A2(new_n12841_), .ZN(new_n28640_));
  NAND2_X1   g25397(.A1(new_n5378_), .A2(pi0616), .ZN(new_n28641_));
  XOR2_X1    g25398(.A1(new_n28640_), .A2(new_n28641_), .Z(new_n28642_));
  OAI21_X1   g25399(.A1(new_n28642_), .A2(new_n12809_), .B(new_n12868_), .ZN(new_n28643_));
  INV_X1     g25400(.I(new_n28611_), .ZN(new_n28644_));
  NOR4_X1    g25401(.A1(new_n12890_), .A2(new_n5636_), .A3(new_n13413_), .A4(new_n28644_), .ZN(new_n28645_));
  NAND3_X1   g25402(.A1(new_n28639_), .A2(new_n28643_), .A3(new_n28645_), .ZN(new_n28646_));
  OAI22_X1   g25403(.A1(new_n28637_), .A2(new_n28646_), .B1(new_n13086_), .B2(new_n28635_), .ZN(new_n28647_));
  NOR2_X1    g25404(.A1(new_n12951_), .A2(new_n12953_), .ZN(new_n28648_));
  INV_X1     g25405(.I(new_n28648_), .ZN(new_n28649_));
  NOR2_X1    g25406(.A1(new_n5397_), .A2(new_n28624_), .ZN(new_n28650_));
  AOI21_X1   g25407(.A1(new_n12973_), .A2(new_n28650_), .B(pi0947), .ZN(new_n28651_));
  NOR2_X1    g25408(.A1(new_n28651_), .A2(new_n28649_), .ZN(new_n28652_));
  AOI21_X1   g25409(.A1(new_n28647_), .A2(new_n28652_), .B(new_n15098_), .ZN(new_n28653_));
  NOR2_X1    g25410(.A1(new_n28611_), .A2(new_n3098_), .ZN(new_n28654_));
  XOR2_X1    g25411(.A1(new_n13069_), .A2(new_n28654_), .Z(new_n28655_));
  OAI21_X1   g25412(.A1(new_n28655_), .A2(new_n3011_), .B(new_n3211_), .ZN(new_n28656_));
  NAND3_X1   g25413(.A1(new_n28549_), .A2(new_n3090_), .A3(new_n28628_), .ZN(new_n28657_));
  NAND3_X1   g25414(.A1(new_n5633_), .A2(new_n5741_), .A3(new_n5800_), .ZN(new_n28658_));
  NAND3_X1   g25415(.A1(new_n28657_), .A2(new_n28556_), .A3(new_n28658_), .ZN(new_n28659_));
  INV_X1     g25416(.I(new_n28565_), .ZN(new_n28660_));
  AOI22_X1   g25417(.A1(new_n28660_), .A2(new_n28610_), .B1(new_n12826_), .B2(new_n28609_), .ZN(new_n28661_));
  NOR4_X1    g25418(.A1(new_n28547_), .A2(new_n3011_), .A3(new_n5397_), .A4(new_n28644_), .ZN(new_n28662_));
  NAND2_X1   g25419(.A1(new_n28661_), .A2(new_n28662_), .ZN(new_n28663_));
  AOI21_X1   g25420(.A1(new_n28659_), .A2(new_n3011_), .B(new_n28663_), .ZN(new_n28664_));
  INV_X1     g25421(.I(new_n28609_), .ZN(new_n28665_));
  NAND2_X1   g25422(.A1(new_n12963_), .A2(new_n12961_), .ZN(new_n28666_));
  AOI21_X1   g25423(.A1(new_n28666_), .A2(pi0947), .B(new_n5397_), .ZN(new_n28667_));
  OAI21_X1   g25424(.A1(new_n12971_), .A2(new_n28665_), .B(new_n28667_), .ZN(new_n28668_));
  NAND2_X1   g25425(.A1(new_n28668_), .A2(new_n3092_), .ZN(new_n28669_));
  NAND2_X1   g25426(.A1(new_n13162_), .A2(new_n28644_), .ZN(new_n28670_));
  XOR2_X1    g25427(.A1(new_n13163_), .A2(new_n28670_), .Z(new_n28671_));
  NAND4_X1   g25428(.A1(new_n28656_), .A2(new_n28664_), .A3(new_n28669_), .A4(new_n28671_), .ZN(new_n28672_));
  OAI22_X1   g25429(.A1(new_n28653_), .A2(new_n28672_), .B1(new_n28615_), .B2(new_n28632_), .ZN(new_n28673_));
  NOR3_X1    g25430(.A1(new_n28661_), .A2(pi0216), .A3(new_n3121_), .ZN(new_n28674_));
  OAI21_X1   g25431(.A1(new_n16996_), .A2(new_n28611_), .B(pi0215), .ZN(new_n28675_));
  OAI21_X1   g25432(.A1(new_n28674_), .A2(new_n28675_), .B(new_n3011_), .ZN(new_n28676_));
  NAND2_X1   g25433(.A1(new_n28633_), .A2(new_n28665_), .ZN(new_n28677_));
  NAND4_X1   g25434(.A1(new_n28676_), .A2(pi0216), .A3(new_n8297_), .A4(new_n28677_), .ZN(new_n28678_));
  NOR3_X1    g25435(.A1(new_n17068_), .A2(new_n5800_), .A3(new_n28678_), .ZN(new_n28679_));
  NAND2_X1   g25436(.A1(new_n28673_), .A2(new_n28679_), .ZN(new_n28680_));
  XNOR2_X1   g25437(.A1(new_n28680_), .A2(new_n28614_), .ZN(po0373));
  INV_X1     g25438(.I(pi0695), .ZN(new_n28682_));
  INV_X1     g25439(.I(pi0612), .ZN(new_n28683_));
  NOR2_X1    g25440(.A1(new_n10168_), .A2(new_n28683_), .ZN(new_n28684_));
  NOR2_X1    g25441(.A1(new_n28372_), .A2(new_n28684_), .ZN(new_n28685_));
  NAND3_X1   g25442(.A1(new_n28295_), .A2(new_n10168_), .A3(pi0695), .ZN(new_n28686_));
  OAI21_X1   g25443(.A1(new_n28685_), .A2(new_n28686_), .B(new_n28682_), .ZN(new_n28687_));
  NAND2_X1   g25444(.A1(new_n28323_), .A2(new_n28687_), .ZN(new_n28688_));
  NAND4_X1   g25445(.A1(new_n28358_), .A2(pi0217), .A3(new_n28363_), .A4(pi0695), .ZN(new_n28689_));
  NAND2_X1   g25446(.A1(new_n28358_), .A2(new_n28363_), .ZN(new_n28690_));
  NAND3_X1   g25447(.A1(new_n28690_), .A2(pi0217), .A3(new_n28682_), .ZN(new_n28691_));
  NAND2_X1   g25448(.A1(new_n28691_), .A2(new_n28689_), .ZN(new_n28692_));
  AOI21_X1   g25449(.A1(new_n28692_), .A2(new_n28376_), .B(pi0612), .ZN(new_n28693_));
  NOR4_X1    g25450(.A1(new_n28399_), .A2(new_n10168_), .A3(new_n28682_), .A4(new_n28414_), .ZN(new_n28694_));
  NOR3_X1    g25451(.A1(new_n28418_), .A2(pi0217), .A3(new_n28682_), .ZN(new_n28695_));
  OAI21_X1   g25452(.A1(new_n28695_), .A2(new_n28694_), .B(new_n28390_), .ZN(new_n28696_));
  AOI21_X1   g25453(.A1(new_n28693_), .A2(new_n28688_), .B(new_n28696_), .ZN(po0374));
  NOR3_X1    g25454(.A1(new_n27759_), .A2(pi0233), .A3(pi0237), .ZN(new_n28698_));
  NAND2_X1   g25455(.A1(new_n28698_), .A2(pi0218), .ZN(new_n28699_));
  OAI21_X1   g25456(.A1(new_n27757_), .A2(pi0218), .B(new_n28699_), .ZN(po0375));
  NOR3_X1    g25457(.A1(new_n28517_), .A2(new_n26964_), .A3(new_n26983_), .ZN(new_n28701_));
  NOR3_X1    g25458(.A1(new_n28516_), .A2(pi0617), .A3(new_n26983_), .ZN(new_n28702_));
  OAI21_X1   g25459(.A1(new_n28701_), .A2(new_n28702_), .B(new_n28515_), .ZN(new_n28703_));
  NAND3_X1   g25460(.A1(new_n28703_), .A2(new_n26964_), .A3(new_n28521_), .ZN(new_n28704_));
  AOI21_X1   g25461(.A1(new_n28704_), .A2(pi0637), .B(new_n8683_), .ZN(po0376));
  NAND3_X1   g25462(.A1(new_n27677_), .A2(pi0220), .A3(new_n27766_), .ZN(new_n28706_));
  OAI21_X1   g25463(.A1(new_n27669_), .A2(pi0220), .B(new_n28706_), .ZN(po0377));
  NOR2_X1    g25464(.A1(new_n16969_), .A2(new_n5374_), .ZN(new_n28708_));
  NOR2_X1    g25465(.A1(new_n12841_), .A2(new_n5800_), .ZN(new_n28709_));
  NOR2_X1    g25466(.A1(new_n28708_), .A2(new_n28709_), .ZN(new_n28710_));
  NOR2_X1    g25467(.A1(new_n28710_), .A2(new_n3259_), .ZN(new_n28711_));
  XOR2_X1    g25468(.A1(new_n13723_), .A2(new_n28711_), .Z(new_n28712_));
  AOI21_X1   g25469(.A1(new_n28712_), .A2(pi0221), .B(new_n8345_), .ZN(new_n28713_));
  NOR2_X1    g25470(.A1(new_n12809_), .A2(new_n12868_), .ZN(new_n28714_));
  AOI21_X1   g25471(.A1(new_n12967_), .A2(new_n12868_), .B(new_n28714_), .ZN(new_n28715_));
  INV_X1     g25472(.I(new_n28715_), .ZN(new_n28716_));
  AOI21_X1   g25473(.A1(new_n28648_), .A2(new_n12963_), .B(new_n12845_), .ZN(new_n28717_));
  NOR2_X1    g25474(.A1(new_n12845_), .A2(new_n12841_), .ZN(new_n28718_));
  XOR2_X1    g25475(.A1(new_n28717_), .A2(new_n28718_), .Z(new_n28719_));
  AOI21_X1   g25476(.A1(new_n28719_), .A2(new_n28716_), .B(new_n5397_), .ZN(new_n28720_));
  XOR2_X1    g25477(.A1(new_n28720_), .A2(new_n28586_), .Z(new_n28721_));
  NOR2_X1    g25478(.A1(new_n28721_), .A2(new_n12980_), .ZN(new_n28722_));
  INV_X1     g25479(.I(new_n28708_), .ZN(new_n28723_));
  NOR2_X1    g25480(.A1(new_n12818_), .A2(new_n5386_), .ZN(new_n28724_));
  AOI21_X1   g25481(.A1(new_n28715_), .A2(new_n5386_), .B(new_n28724_), .ZN(new_n28725_));
  NOR2_X1    g25482(.A1(new_n13417_), .A2(pi0642), .ZN(new_n28726_));
  NOR3_X1    g25483(.A1(new_n12845_), .A2(pi0616), .A3(new_n5800_), .ZN(new_n28727_));
  OAI21_X1   g25484(.A1(new_n28726_), .A2(new_n28727_), .B(new_n28566_), .ZN(new_n28728_));
  AOI21_X1   g25485(.A1(new_n28725_), .A2(new_n12849_), .B(new_n28728_), .ZN(new_n28729_));
  AOI21_X1   g25486(.A1(new_n28729_), .A2(new_n5398_), .B(pi0947), .ZN(new_n28730_));
  OAI21_X1   g25487(.A1(new_n28730_), .A2(new_n13086_), .B(new_n28723_), .ZN(new_n28731_));
  INV_X1     g25488(.I(new_n28710_), .ZN(new_n28732_));
  NOR2_X1    g25489(.A1(new_n28547_), .A2(new_n28732_), .ZN(new_n28733_));
  OAI21_X1   g25490(.A1(new_n28722_), .A2(new_n28731_), .B(new_n28733_), .ZN(new_n28734_));
  NAND2_X1   g25491(.A1(new_n28733_), .A2(new_n3091_), .ZN(new_n28735_));
  XOR2_X1    g25492(.A1(new_n28734_), .A2(new_n28735_), .Z(new_n28736_));
  NOR2_X1    g25493(.A1(new_n12911_), .A2(new_n5397_), .ZN(new_n28737_));
  XOR2_X1    g25494(.A1(new_n28737_), .A2(new_n28586_), .Z(new_n28738_));
  OAI21_X1   g25495(.A1(new_n12923_), .A2(new_n12922_), .B(new_n5636_), .ZN(new_n28739_));
  NOR2_X1    g25496(.A1(pi0616), .A2(pi0947), .ZN(new_n28740_));
  AOI21_X1   g25497(.A1(new_n28739_), .A2(new_n28740_), .B(new_n28579_), .ZN(new_n28741_));
  AOI21_X1   g25498(.A1(new_n28741_), .A2(new_n5398_), .B(pi0947), .ZN(new_n28742_));
  NAND3_X1   g25499(.A1(new_n12895_), .A2(pi0223), .A3(new_n28708_), .ZN(new_n28743_));
  NOR4_X1    g25500(.A1(new_n28738_), .A2(new_n12935_), .A3(new_n28742_), .A4(new_n28743_), .ZN(new_n28744_));
  INV_X1     g25501(.I(new_n28556_), .ZN(new_n28745_));
  INV_X1     g25502(.I(new_n28549_), .ZN(new_n28746_));
  NOR2_X1    g25503(.A1(new_n12865_), .A2(new_n5800_), .ZN(new_n28747_));
  AOI21_X1   g25504(.A1(new_n28746_), .A2(new_n28747_), .B(new_n28708_), .ZN(new_n28748_));
  OAI21_X1   g25505(.A1(new_n28748_), .A2(new_n28745_), .B(pi0223), .ZN(new_n28749_));
  NOR2_X1    g25506(.A1(new_n3098_), .A2(pi0221), .ZN(new_n28750_));
  AOI21_X1   g25507(.A1(new_n28749_), .A2(new_n28750_), .B(new_n28733_), .ZN(new_n28751_));
  AOI21_X1   g25508(.A1(pi0947), .A2(new_n12847_), .B(new_n12850_), .ZN(new_n28752_));
  NOR3_X1    g25509(.A1(new_n28752_), .A2(new_n12949_), .A3(new_n5375_), .ZN(new_n28753_));
  OAI21_X1   g25510(.A1(new_n28753_), .A2(new_n5398_), .B(new_n28708_), .ZN(new_n28754_));
  OAI21_X1   g25511(.A1(new_n12971_), .A2(new_n28754_), .B(new_n3092_), .ZN(new_n28755_));
  AOI22_X1   g25512(.A1(new_n28660_), .A2(new_n28709_), .B1(new_n12826_), .B2(new_n28708_), .ZN(new_n28756_));
  NAND3_X1   g25513(.A1(new_n28755_), .A2(new_n5398_), .A3(new_n28756_), .ZN(new_n28757_));
  OAI21_X1   g25514(.A1(new_n28751_), .A2(new_n28757_), .B(new_n3121_), .ZN(new_n28758_));
  NOR2_X1    g25515(.A1(new_n28744_), .A2(new_n28758_), .ZN(new_n28759_));
  NOR2_X1    g25516(.A1(new_n28759_), .A2(new_n12809_), .ZN(new_n28760_));
  NAND2_X1   g25517(.A1(new_n28732_), .A2(pi0299), .ZN(new_n28761_));
  XOR2_X1    g25518(.A1(new_n13069_), .A2(new_n28761_), .Z(new_n28762_));
  AOI21_X1   g25519(.A1(new_n28762_), .A2(pi0221), .B(new_n3212_), .ZN(new_n28763_));
  NAND2_X1   g25520(.A1(new_n13162_), .A2(new_n28732_), .ZN(new_n28764_));
  XOR2_X1    g25521(.A1(new_n13163_), .A2(new_n28764_), .Z(new_n28765_));
  NAND2_X1   g25522(.A1(new_n28765_), .A2(pi0221), .ZN(new_n28766_));
  OAI21_X1   g25523(.A1(new_n28766_), .A2(new_n28763_), .B(new_n3183_), .ZN(new_n28767_));
  AOI21_X1   g25524(.A1(new_n28736_), .A2(new_n28760_), .B(new_n28767_), .ZN(new_n28768_));
  NAND2_X1   g25525(.A1(new_n5741_), .A2(new_n5800_), .ZN(new_n28769_));
  NAND2_X1   g25526(.A1(new_n28769_), .A2(pi0661), .ZN(new_n28770_));
  NAND2_X1   g25527(.A1(new_n28710_), .A2(pi0215), .ZN(new_n28771_));
  AOI21_X1   g25528(.A1(new_n12809_), .A2(new_n3312_), .B(new_n28771_), .ZN(new_n28772_));
  OAI21_X1   g25529(.A1(pi0216), .A2(new_n28772_), .B(new_n28756_), .ZN(new_n28773_));
  NAND3_X1   g25530(.A1(new_n28773_), .A2(new_n3121_), .A3(new_n28770_), .ZN(new_n28774_));
  AOI21_X1   g25531(.A1(new_n28774_), .A2(new_n28729_), .B(pi0299), .ZN(new_n28775_));
  NOR2_X1    g25532(.A1(new_n28747_), .A2(new_n28708_), .ZN(new_n28776_));
  OAI21_X1   g25533(.A1(new_n28776_), .A2(new_n28548_), .B(new_n3121_), .ZN(new_n28777_));
  NOR2_X1    g25534(.A1(new_n28723_), .A2(new_n3178_), .ZN(new_n28778_));
  NAND4_X1   g25535(.A1(new_n28777_), .A2(new_n8297_), .A3(new_n28741_), .A4(new_n28778_), .ZN(new_n28779_));
  NOR4_X1    g25536(.A1(new_n28768_), .A2(new_n28615_), .A3(new_n28775_), .A4(new_n28779_), .ZN(new_n28780_));
  XOR2_X1    g25537(.A1(new_n28780_), .A2(new_n28713_), .Z(po0378));
  NOR2_X1    g25538(.A1(new_n17298_), .A2(new_n3090_), .ZN(new_n28782_));
  XOR2_X1    g25539(.A1(new_n28782_), .A2(new_n3512_), .Z(new_n28783_));
  AOI21_X1   g25540(.A1(new_n28783_), .A2(new_n17052_), .B(new_n3183_), .ZN(new_n28784_));
  NOR2_X1    g25541(.A1(new_n3289_), .A2(pi0038), .ZN(new_n28785_));
  INV_X1     g25542(.I(new_n28785_), .ZN(new_n28786_));
  AOI21_X1   g25543(.A1(new_n28784_), .A2(new_n13085_), .B(new_n28786_), .ZN(new_n28787_));
  OAI21_X1   g25544(.A1(new_n28787_), .A2(new_n14300_), .B(pi0222), .ZN(new_n28788_));
  INV_X1     g25545(.I(new_n28788_), .ZN(new_n28789_));
  NOR2_X1    g25546(.A1(new_n28715_), .A2(pi0616), .ZN(new_n28790_));
  AOI21_X1   g25547(.A1(pi0616), .A2(new_n13275_), .B(new_n28790_), .ZN(new_n28791_));
  NOR2_X1    g25548(.A1(new_n13103_), .A2(new_n12841_), .ZN(new_n28792_));
  INV_X1     g25549(.I(new_n28792_), .ZN(new_n28793_));
  AOI21_X1   g25550(.A1(new_n12945_), .A2(new_n5634_), .B(new_n28793_), .ZN(new_n28794_));
  OAI21_X1   g25551(.A1(new_n28794_), .A2(new_n12842_), .B(new_n5376_), .ZN(new_n28795_));
  NOR2_X1    g25552(.A1(new_n28791_), .A2(new_n28795_), .ZN(new_n28796_));
  AOI21_X1   g25553(.A1(new_n12843_), .A2(new_n28791_), .B(new_n28796_), .ZN(new_n28797_));
  INV_X1     g25554(.I(new_n28797_), .ZN(new_n28798_));
  NOR2_X1    g25555(.A1(new_n14317_), .A2(new_n12841_), .ZN(new_n28799_));
  INV_X1     g25556(.I(new_n28799_), .ZN(new_n28800_));
  NAND2_X1   g25557(.A1(new_n28725_), .A2(new_n12841_), .ZN(new_n28801_));
  NAND2_X1   g25558(.A1(new_n28801_), .A2(new_n28800_), .ZN(new_n28802_));
  NAND3_X1   g25559(.A1(new_n28802_), .A2(new_n5376_), .A3(new_n12842_), .ZN(new_n28803_));
  AOI21_X1   g25560(.A1(new_n28725_), .A2(new_n12841_), .B(new_n28799_), .ZN(new_n28804_));
  NAND3_X1   g25561(.A1(new_n28804_), .A2(new_n5634_), .A3(new_n12842_), .ZN(new_n28805_));
  NAND2_X1   g25562(.A1(new_n28803_), .A2(new_n28805_), .ZN(new_n28806_));
  NOR4_X1    g25563(.A1(new_n13253_), .A2(new_n13142_), .A3(new_n2726_), .A4(new_n12813_), .ZN(new_n28807_));
  OAI21_X1   g25564(.A1(new_n28807_), .A2(pi0616), .B(new_n13203_), .ZN(new_n28808_));
  INV_X1     g25565(.I(new_n28808_), .ZN(new_n28809_));
  NOR2_X1    g25566(.A1(new_n28802_), .A2(new_n12842_), .ZN(new_n28810_));
  AOI21_X1   g25567(.A1(new_n28806_), .A2(new_n28809_), .B(new_n28810_), .ZN(new_n28811_));
  NAND3_X1   g25568(.A1(new_n28811_), .A2(pi0222), .A3(new_n5454_), .ZN(new_n28812_));
  NAND2_X1   g25569(.A1(new_n5454_), .A2(pi0222), .ZN(new_n28813_));
  NOR2_X1    g25570(.A1(new_n28811_), .A2(new_n3099_), .ZN(new_n28814_));
  NAND2_X1   g25571(.A1(new_n28814_), .A2(new_n28813_), .ZN(new_n28815_));
  AOI21_X1   g25572(.A1(new_n28815_), .A2(new_n28812_), .B(new_n28798_), .ZN(new_n28816_));
  NOR2_X1    g25573(.A1(new_n13364_), .A2(new_n12841_), .ZN(new_n28818_));
  NOR2_X1    g25574(.A1(new_n3312_), .A2(new_n3111_), .ZN(new_n28819_));
  INV_X1     g25575(.I(new_n28819_), .ZN(new_n28820_));
  AOI21_X1   g25576(.A1(new_n13368_), .A2(pi0616), .B(new_n28641_), .ZN(new_n28821_));
  NOR3_X1    g25577(.A1(new_n13372_), .A2(new_n12841_), .A3(new_n5378_), .ZN(new_n28822_));
  OAI21_X1   g25578(.A1(new_n28821_), .A2(new_n28822_), .B(new_n13363_), .ZN(new_n28823_));
  NOR2_X1    g25579(.A1(new_n13263_), .A2(new_n13103_), .ZN(new_n28824_));
  NAND2_X1   g25580(.A1(new_n28824_), .A2(pi0616), .ZN(new_n28825_));
  INV_X1     g25581(.I(new_n28825_), .ZN(new_n28826_));
  NOR2_X1    g25582(.A1(new_n12842_), .A2(pi0616), .ZN(new_n28827_));
  AOI21_X1   g25583(.A1(new_n13542_), .A2(new_n28827_), .B(new_n5634_), .ZN(new_n28828_));
  OAI21_X1   g25584(.A1(new_n28825_), .A2(new_n5376_), .B(new_n28828_), .ZN(new_n28829_));
  OAI21_X1   g25585(.A1(new_n12842_), .A2(new_n28826_), .B(new_n28829_), .ZN(new_n28830_));
  NAND2_X1   g25586(.A1(new_n28830_), .A2(new_n5454_), .ZN(new_n28831_));
  XNOR2_X1   g25587(.A1(new_n28831_), .A2(new_n28813_), .ZN(new_n28832_));
  NOR2_X1    g25588(.A1(new_n28832_), .A2(new_n28823_), .ZN(new_n28833_));
  OAI21_X1   g25589(.A1(new_n28816_), .A2(new_n28820_), .B(new_n28833_), .ZN(new_n28834_));
  AOI22_X1   g25590(.A1(new_n12878_), .A2(pi0616), .B1(new_n5376_), .B2(new_n13310_), .ZN(new_n28835_));
  OAI21_X1   g25591(.A1(new_n28835_), .A2(new_n12843_), .B(new_n5634_), .ZN(new_n28836_));
  NAND2_X1   g25592(.A1(new_n12924_), .A2(new_n28836_), .ZN(new_n28837_));
  AOI21_X1   g25593(.A1(pi0616), .A2(new_n14304_), .B(new_n12932_), .ZN(new_n28838_));
  OR2_X2     g25594(.A1(new_n28838_), .A2(new_n12842_), .Z(new_n28839_));
  AOI21_X1   g25595(.A1(new_n28839_), .A2(new_n28837_), .B(new_n3099_), .ZN(new_n28840_));
  XNOR2_X1   g25596(.A1(new_n28840_), .A2(new_n28813_), .ZN(new_n28841_));
  NOR2_X1    g25597(.A1(new_n13386_), .A2(new_n5636_), .ZN(new_n28842_));
  INV_X1     g25598(.I(new_n28842_), .ZN(new_n28843_));
  AOI21_X1   g25599(.A1(new_n12841_), .A2(new_n13364_), .B(new_n28843_), .ZN(new_n28844_));
  AND2_X2    g25600(.A1(new_n28844_), .A2(new_n3099_), .Z(new_n28845_));
  AOI21_X1   g25601(.A1(pi0616), .A2(new_n13276_), .B(new_n12903_), .ZN(new_n28846_));
  OAI21_X1   g25602(.A1(new_n13334_), .A2(new_n5376_), .B(new_n28792_), .ZN(new_n28847_));
  AOI21_X1   g25603(.A1(new_n28847_), .A2(new_n12843_), .B(new_n5634_), .ZN(new_n28848_));
  NAND2_X1   g25604(.A1(new_n28846_), .A2(new_n28848_), .ZN(new_n28849_));
  OAI21_X1   g25605(.A1(new_n12842_), .A2(new_n28846_), .B(new_n28849_), .ZN(new_n28850_));
  INV_X1     g25606(.I(new_n28850_), .ZN(new_n28851_));
  NAND3_X1   g25607(.A1(new_n28841_), .A2(new_n28845_), .A3(new_n28851_), .ZN(new_n28852_));
  AOI21_X1   g25608(.A1(new_n28852_), .A2(new_n12930_), .B(new_n13309_), .ZN(new_n28853_));
  INV_X1     g25609(.I(new_n28853_), .ZN(new_n28854_));
  AOI21_X1   g25610(.A1(new_n28834_), .A2(new_n3098_), .B(new_n28854_), .ZN(new_n28855_));
  NAND3_X1   g25611(.A1(new_n28811_), .A2(pi0222), .A3(new_n5398_), .ZN(new_n28856_));
  NOR2_X1    g25612(.A1(new_n5397_), .A2(new_n3099_), .ZN(new_n28857_));
  INV_X1     g25613(.I(new_n28857_), .ZN(new_n28858_));
  NAND2_X1   g25614(.A1(new_n28814_), .A2(new_n28858_), .ZN(new_n28859_));
  NAND2_X1   g25615(.A1(new_n28859_), .A2(new_n28856_), .ZN(new_n28860_));
  NAND2_X1   g25616(.A1(new_n28860_), .A2(new_n28797_), .ZN(new_n28861_));
  NAND4_X1   g25617(.A1(new_n28839_), .A2(pi0222), .A3(new_n5398_), .A4(new_n28837_), .ZN(new_n28862_));
  NAND2_X1   g25618(.A1(new_n28840_), .A2(new_n28858_), .ZN(new_n28863_));
  AOI21_X1   g25619(.A1(new_n28863_), .A2(new_n28862_), .B(new_n28850_), .ZN(new_n28864_));
  NAND2_X1   g25620(.A1(new_n28845_), .A2(new_n13700_), .ZN(new_n28865_));
  INV_X1     g25621(.I(new_n28865_), .ZN(new_n28866_));
  AOI21_X1   g25622(.A1(new_n28864_), .A2(new_n28866_), .B(pi0223), .ZN(new_n28867_));
  NOR3_X1    g25623(.A1(new_n13180_), .A2(new_n3183_), .A3(new_n12841_), .ZN(new_n28868_));
  NOR3_X1    g25624(.A1(new_n13180_), .A2(pi0039), .A3(pi0616), .ZN(new_n28869_));
  NOR2_X1    g25625(.A1(new_n3259_), .A2(new_n3099_), .ZN(new_n28870_));
  OAI21_X1   g25626(.A1(new_n28868_), .A2(new_n28869_), .B(new_n28870_), .ZN(new_n28871_));
  AOI21_X1   g25627(.A1(new_n28871_), .A2(new_n3099_), .B(new_n14338_), .ZN(new_n28872_));
  AOI21_X1   g25628(.A1(new_n13109_), .A2(pi0222), .B(new_n16715_), .ZN(new_n28873_));
  NOR2_X1    g25629(.A1(new_n3289_), .A2(new_n3099_), .ZN(new_n28874_));
  INV_X1     g25630(.I(new_n28874_), .ZN(new_n28875_));
  NOR2_X1    g25631(.A1(new_n13107_), .A2(new_n28875_), .ZN(new_n28876_));
  OAI21_X1   g25632(.A1(new_n28873_), .A2(pi0616), .B(new_n28876_), .ZN(new_n28877_));
  INV_X1     g25633(.I(new_n28877_), .ZN(new_n28878_));
  INV_X1     g25634(.I(new_n28818_), .ZN(new_n28879_));
  INV_X1     g25635(.I(new_n28823_), .ZN(new_n28880_));
  NAND2_X1   g25636(.A1(new_n28830_), .A2(pi0224), .ZN(new_n28881_));
  NOR2_X1    g25637(.A1(new_n5397_), .A2(new_n3100_), .ZN(new_n28882_));
  INV_X1     g25638(.I(new_n28882_), .ZN(new_n28883_));
  XOR2_X1    g25639(.A1(new_n28881_), .A2(new_n28883_), .Z(new_n28884_));
  AOI21_X1   g25640(.A1(new_n28884_), .A2(new_n28880_), .B(pi0222), .ZN(new_n28885_));
  NOR4_X1    g25641(.A1(new_n28885_), .A2(new_n3100_), .A3(new_n3098_), .A4(new_n28879_), .ZN(new_n28886_));
  OAI21_X1   g25642(.A1(new_n28872_), .A2(new_n28878_), .B(new_n28886_), .ZN(new_n28887_));
  AOI21_X1   g25643(.A1(new_n28861_), .A2(new_n28867_), .B(new_n28887_), .ZN(new_n28888_));
  OAI21_X1   g25644(.A1(new_n28855_), .A2(pi0039), .B(new_n28888_), .ZN(new_n28889_));
  NAND2_X1   g25645(.A1(new_n28788_), .A2(new_n13775_), .ZN(new_n28890_));
  OAI21_X1   g25646(.A1(new_n28889_), .A2(new_n13775_), .B(new_n28890_), .ZN(new_n28891_));
  NOR2_X1    g25647(.A1(new_n28891_), .A2(new_n13766_), .ZN(new_n28892_));
  NOR2_X1    g25648(.A1(new_n28892_), .A2(new_n14694_), .ZN(new_n28893_));
  NOR3_X1    g25649(.A1(new_n28891_), .A2(new_n13766_), .A3(new_n14090_), .ZN(new_n28894_));
  OAI21_X1   g25650(.A1(new_n28893_), .A2(new_n28894_), .B(new_n28789_), .ZN(new_n28895_));
  NAND2_X1   g25651(.A1(new_n28895_), .A2(pi0785), .ZN(new_n28896_));
  INV_X1     g25652(.I(new_n28891_), .ZN(new_n28897_));
  NAND3_X1   g25653(.A1(new_n28891_), .A2(pi0609), .A3(pi1155), .ZN(new_n28898_));
  INV_X1     g25654(.I(new_n28898_), .ZN(new_n28899_));
  NOR3_X1    g25655(.A1(new_n28891_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n28900_));
  OAI21_X1   g25656(.A1(new_n28899_), .A2(new_n28900_), .B(new_n28789_), .ZN(new_n28901_));
  NOR3_X1    g25657(.A1(new_n28901_), .A2(new_n13801_), .A3(new_n28897_), .ZN(new_n28902_));
  NAND2_X1   g25658(.A1(new_n28902_), .A2(new_n28896_), .ZN(new_n28903_));
  INV_X1     g25659(.I(new_n28900_), .ZN(new_n28904_));
  AOI21_X1   g25660(.A1(new_n28904_), .A2(new_n28898_), .B(new_n28788_), .ZN(new_n28905_));
  NAND3_X1   g25661(.A1(new_n28905_), .A2(pi0785), .A3(new_n28891_), .ZN(new_n28906_));
  NAND3_X1   g25662(.A1(new_n28906_), .A2(pi0785), .A3(new_n28895_), .ZN(new_n28907_));
  NAND2_X1   g25663(.A1(new_n28907_), .A2(new_n28903_), .ZN(new_n28908_));
  NAND3_X1   g25664(.A1(new_n28908_), .A2(pi0618), .A3(pi1154), .ZN(new_n28909_));
  NOR3_X1    g25665(.A1(new_n28908_), .A2(new_n13816_), .A3(new_n13818_), .ZN(new_n28910_));
  INV_X1     g25666(.I(new_n28910_), .ZN(new_n28911_));
  AOI21_X1   g25667(.A1(new_n28911_), .A2(new_n28909_), .B(new_n28788_), .ZN(new_n28912_));
  NAND3_X1   g25668(.A1(new_n28908_), .A2(pi0618), .A3(pi1154), .ZN(new_n28913_));
  AOI21_X1   g25669(.A1(pi0785), .A2(new_n28895_), .B(new_n28906_), .ZN(new_n28914_));
  NOR2_X1    g25670(.A1(new_n28902_), .A2(new_n28896_), .ZN(new_n28915_));
  NOR2_X1    g25671(.A1(new_n28914_), .A2(new_n28915_), .ZN(new_n28916_));
  NAND3_X1   g25672(.A1(new_n28916_), .A2(pi1154), .A3(new_n13819_), .ZN(new_n28917_));
  AOI21_X1   g25673(.A1(new_n28917_), .A2(new_n28913_), .B(new_n28788_), .ZN(new_n28918_));
  NAND4_X1   g25674(.A1(new_n28912_), .A2(new_n28918_), .A3(pi0781), .A4(new_n28908_), .ZN(new_n28919_));
  AOI21_X1   g25675(.A1(new_n28916_), .A2(pi0618), .B(new_n13819_), .ZN(new_n28920_));
  OAI21_X1   g25676(.A1(new_n28920_), .A2(new_n28910_), .B(new_n28789_), .ZN(new_n28921_));
  NOR2_X1    g25677(.A1(new_n28916_), .A2(new_n13855_), .ZN(new_n28922_));
  NAND2_X1   g25678(.A1(new_n28918_), .A2(new_n28922_), .ZN(new_n28923_));
  NAND3_X1   g25679(.A1(new_n28923_), .A2(pi0781), .A3(new_n28921_), .ZN(new_n28924_));
  NAND2_X1   g25680(.A1(new_n28924_), .A2(new_n28919_), .ZN(new_n28925_));
  NAND3_X1   g25681(.A1(new_n28925_), .A2(pi0619), .A3(pi1159), .ZN(new_n28926_));
  AOI21_X1   g25682(.A1(new_n28916_), .A2(pi1154), .B(new_n13819_), .ZN(new_n28927_));
  NOR3_X1    g25683(.A1(new_n28908_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n28928_));
  OAI21_X1   g25684(.A1(new_n28927_), .A2(new_n28928_), .B(new_n28789_), .ZN(new_n28929_));
  NOR4_X1    g25685(.A1(new_n28929_), .A2(new_n28921_), .A3(new_n13855_), .A4(new_n28916_), .ZN(new_n28930_));
  NAND2_X1   g25686(.A1(new_n28921_), .A2(pi0781), .ZN(new_n28931_));
  NOR3_X1    g25687(.A1(new_n28929_), .A2(new_n13855_), .A3(new_n28916_), .ZN(new_n28932_));
  NOR2_X1    g25688(.A1(new_n28932_), .A2(new_n28931_), .ZN(new_n28933_));
  NOR2_X1    g25689(.A1(new_n28933_), .A2(new_n28930_), .ZN(new_n28934_));
  NAND3_X1   g25690(.A1(new_n28934_), .A2(pi0619), .A3(new_n13868_), .ZN(new_n28935_));
  AOI21_X1   g25691(.A1(new_n28935_), .A2(new_n28926_), .B(new_n28788_), .ZN(new_n28936_));
  NOR2_X1    g25692(.A1(new_n5374_), .A2(new_n5375_), .ZN(new_n28937_));
  OAI21_X1   g25693(.A1(new_n13159_), .A2(new_n3099_), .B(new_n3098_), .ZN(new_n28938_));
  NOR2_X1    g25694(.A1(new_n28938_), .A2(new_n28937_), .ZN(new_n28939_));
  NOR2_X1    g25695(.A1(new_n15066_), .A2(new_n28938_), .ZN(new_n28940_));
  XOR2_X1    g25696(.A1(new_n28940_), .A2(new_n28939_), .Z(new_n28941_));
  AOI21_X1   g25697(.A1(new_n28941_), .A2(pi0222), .B(new_n3183_), .ZN(new_n28942_));
  INV_X1     g25698(.I(new_n28942_), .ZN(new_n28943_));
  OAI21_X1   g25699(.A1(pi0680), .A2(new_n12821_), .B(new_n13646_), .ZN(new_n28944_));
  INV_X1     g25700(.I(new_n28944_), .ZN(new_n28945_));
  NOR2_X1    g25701(.A1(new_n28945_), .A2(new_n5374_), .ZN(new_n28946_));
  AOI21_X1   g25702(.A1(new_n12974_), .A2(new_n5374_), .B(new_n28946_), .ZN(new_n28947_));
  NOR2_X1    g25703(.A1(new_n12960_), .A2(new_n5374_), .ZN(new_n28948_));
  NOR2_X1    g25704(.A1(new_n13538_), .A2(new_n13643_), .ZN(new_n28949_));
  NAND2_X1   g25705(.A1(new_n28949_), .A2(new_n12920_), .ZN(new_n28950_));
  XOR2_X1    g25706(.A1(new_n28950_), .A2(new_n28948_), .Z(new_n28951_));
  NOR2_X1    g25707(.A1(new_n5633_), .A2(new_n5375_), .ZN(new_n28952_));
  INV_X1     g25708(.I(new_n28952_), .ZN(new_n28953_));
  NOR3_X1    g25709(.A1(new_n12960_), .A2(new_n12949_), .A3(new_n28953_), .ZN(new_n28954_));
  NOR3_X1    g25710(.A1(new_n12971_), .A2(new_n12945_), .A3(new_n28953_), .ZN(new_n28955_));
  NOR3_X1    g25711(.A1(new_n28955_), .A2(new_n28954_), .A3(new_n12843_), .ZN(new_n28956_));
  OAI21_X1   g25712(.A1(new_n28951_), .A2(new_n28956_), .B(pi0222), .ZN(new_n28957_));
  XNOR2_X1   g25713(.A1(new_n28957_), .A2(new_n28813_), .ZN(new_n28958_));
  OAI21_X1   g25714(.A1(new_n12784_), .A2(new_n3099_), .B(new_n3312_), .ZN(new_n28959_));
  OAI21_X1   g25715(.A1(new_n28959_), .A2(new_n3111_), .B(new_n5374_), .ZN(new_n28960_));
  AOI21_X1   g25716(.A1(new_n28960_), .A2(new_n13707_), .B(new_n3312_), .ZN(new_n28961_));
  OAI21_X1   g25717(.A1(new_n28958_), .A2(new_n28947_), .B(new_n28961_), .ZN(new_n28962_));
  NAND2_X1   g25718(.A1(new_n12826_), .A2(new_n13206_), .ZN(new_n28963_));
  NAND2_X1   g25719(.A1(new_n13691_), .A2(new_n28937_), .ZN(new_n28964_));
  NAND2_X1   g25720(.A1(new_n28964_), .A2(new_n5454_), .ZN(new_n28965_));
  XNOR2_X1   g25721(.A1(new_n28965_), .A2(new_n28813_), .ZN(new_n28966_));
  NOR3_X1    g25722(.A1(new_n28966_), .A2(new_n5374_), .A3(new_n28963_), .ZN(new_n28967_));
  AOI21_X1   g25723(.A1(new_n28962_), .A2(new_n28967_), .B(new_n3098_), .ZN(new_n28968_));
  XOR2_X1    g25724(.A1(new_n28957_), .A2(new_n28857_), .Z(new_n28969_));
  OAI21_X1   g25725(.A1(new_n28969_), .A2(new_n28947_), .B(new_n3090_), .ZN(new_n28970_));
  NAND2_X1   g25726(.A1(new_n28964_), .A2(pi0224), .ZN(new_n28971_));
  XOR2_X1    g25727(.A1(new_n28971_), .A2(new_n28882_), .Z(new_n28972_));
  OAI21_X1   g25728(.A1(pi0661), .A2(new_n3101_), .B(new_n13707_), .ZN(new_n28973_));
  NOR4_X1    g25729(.A1(new_n28972_), .A2(new_n5374_), .A3(new_n28963_), .A4(new_n28973_), .ZN(new_n28974_));
  NAND2_X1   g25730(.A1(new_n28970_), .A2(new_n28974_), .ZN(new_n28975_));
  AOI22_X1   g25731(.A1(new_n12927_), .A2(new_n13641_), .B1(pi0680), .B2(new_n13470_), .ZN(new_n28976_));
  NOR2_X1    g25732(.A1(new_n28976_), .A2(new_n5374_), .ZN(new_n28977_));
  AOI21_X1   g25733(.A1(new_n12911_), .A2(new_n5374_), .B(new_n28977_), .ZN(new_n28978_));
  INV_X1     g25734(.I(new_n28978_), .ZN(new_n28979_));
  NOR2_X1    g25735(.A1(new_n12924_), .A2(new_n5374_), .ZN(new_n28980_));
  NAND2_X1   g25736(.A1(new_n13658_), .A2(new_n13661_), .ZN(new_n28981_));
  NAND2_X1   g25737(.A1(new_n28981_), .A2(new_n12920_), .ZN(new_n28982_));
  XOR2_X1    g25738(.A1(new_n28982_), .A2(new_n28980_), .Z(new_n28983_));
  NOR2_X1    g25739(.A1(new_n12919_), .A2(new_n12843_), .ZN(new_n28984_));
  OAI21_X1   g25740(.A1(new_n28983_), .A2(new_n28984_), .B(pi0222), .ZN(new_n28985_));
  XOR2_X1    g25741(.A1(new_n28985_), .A2(new_n28813_), .Z(new_n28986_));
  NAND2_X1   g25742(.A1(new_n28986_), .A2(new_n28979_), .ZN(new_n28987_));
  NOR2_X1    g25743(.A1(new_n13712_), .A2(pi0661), .ZN(new_n28988_));
  AOI21_X1   g25744(.A1(new_n28987_), .A2(new_n28988_), .B(new_n3099_), .ZN(new_n28989_));
  XOR2_X1    g25745(.A1(new_n28985_), .A2(new_n28857_), .Z(new_n28990_));
  NOR2_X1    g25746(.A1(new_n28990_), .A2(new_n28978_), .ZN(new_n28991_));
  NAND3_X1   g25747(.A1(new_n13702_), .A2(new_n3090_), .A3(new_n5374_), .ZN(new_n28992_));
  NAND2_X1   g25748(.A1(new_n28992_), .A2(pi0222), .ZN(new_n28993_));
  OAI21_X1   g25749(.A1(new_n28991_), .A2(new_n28993_), .B(new_n3695_), .ZN(new_n28994_));
  NOR2_X1    g25750(.A1(new_n28994_), .A2(new_n28989_), .ZN(new_n28995_));
  NAND2_X1   g25751(.A1(new_n28995_), .A2(new_n28975_), .ZN(new_n28996_));
  XNOR2_X1   g25752(.A1(new_n28996_), .A2(new_n28968_), .ZN(new_n28997_));
  INV_X1     g25753(.I(new_n28937_), .ZN(new_n28998_));
  OAI21_X1   g25754(.A1(new_n13155_), .A2(new_n3099_), .B(pi0299), .ZN(new_n28999_));
  NOR3_X1    g25755(.A1(new_n28999_), .A2(new_n13141_), .A3(new_n28998_), .ZN(new_n29000_));
  INV_X1     g25756(.I(new_n13141_), .ZN(new_n29001_));
  NOR3_X1    g25757(.A1(new_n28999_), .A2(new_n29001_), .A3(new_n28937_), .ZN(new_n29002_));
  NOR2_X1    g25758(.A1(new_n29000_), .A2(new_n29002_), .ZN(new_n29003_));
  NOR3_X1    g25759(.A1(new_n29003_), .A2(new_n3183_), .A3(new_n3099_), .ZN(new_n29004_));
  NAND3_X1   g25760(.A1(new_n28997_), .A2(new_n28943_), .A3(new_n29004_), .ZN(new_n29005_));
  NAND2_X1   g25761(.A1(new_n28997_), .A2(new_n29004_), .ZN(new_n29006_));
  NAND2_X1   g25762(.A1(new_n29006_), .A2(new_n28942_), .ZN(new_n29007_));
  NOR2_X1    g25763(.A1(new_n28873_), .A2(pi0661), .ZN(new_n29008_));
  INV_X1     g25764(.I(new_n29008_), .ZN(new_n29009_));
  INV_X1     g25765(.I(new_n13719_), .ZN(new_n29010_));
  NOR2_X1    g25766(.A1(new_n29010_), .A2(new_n28875_), .ZN(new_n29011_));
  AOI21_X1   g25767(.A1(new_n29009_), .A2(new_n29011_), .B(pi0038), .ZN(new_n29012_));
  AOI21_X1   g25768(.A1(new_n29007_), .A2(new_n29005_), .B(new_n29012_), .ZN(new_n29013_));
  NAND3_X1   g25769(.A1(new_n29013_), .A2(pi0625), .A3(pi1153), .ZN(new_n29014_));
  INV_X1     g25770(.I(new_n29013_), .ZN(new_n29015_));
  NAND3_X1   g25771(.A1(new_n29015_), .A2(pi0625), .A3(new_n13614_), .ZN(new_n29016_));
  NAND2_X1   g25772(.A1(new_n29016_), .A2(new_n29014_), .ZN(new_n29017_));
  NAND2_X1   g25773(.A1(new_n29017_), .A2(new_n28789_), .ZN(new_n29018_));
  NAND2_X1   g25774(.A1(new_n29018_), .A2(pi0778), .ZN(new_n29019_));
  NAND3_X1   g25775(.A1(new_n29013_), .A2(pi0625), .A3(pi1153), .ZN(new_n29020_));
  NAND3_X1   g25776(.A1(new_n29015_), .A2(new_n13613_), .A3(pi1153), .ZN(new_n29021_));
  AOI21_X1   g25777(.A1(new_n29021_), .A2(new_n29020_), .B(new_n28788_), .ZN(new_n29022_));
  NAND3_X1   g25778(.A1(new_n29022_), .A2(pi0778), .A3(new_n29013_), .ZN(new_n29023_));
  XOR2_X1    g25779(.A1(new_n29019_), .A2(new_n29023_), .Z(new_n29024_));
  NOR2_X1    g25780(.A1(new_n28789_), .A2(new_n13805_), .ZN(new_n29025_));
  AOI21_X1   g25781(.A1(new_n29024_), .A2(new_n13805_), .B(new_n29025_), .ZN(new_n29026_));
  NAND2_X1   g25782(.A1(new_n28788_), .A2(new_n13879_), .ZN(new_n29027_));
  OAI21_X1   g25783(.A1(new_n29026_), .A2(new_n13879_), .B(new_n29027_), .ZN(new_n29028_));
  INV_X1     g25784(.I(new_n29028_), .ZN(new_n29029_));
  AOI21_X1   g25785(.A1(pi0778), .A2(new_n29018_), .B(new_n29023_), .ZN(new_n29030_));
  INV_X1     g25786(.I(new_n29023_), .ZN(new_n29031_));
  NOR2_X1    g25787(.A1(new_n29031_), .A2(new_n29019_), .ZN(new_n29032_));
  NOR2_X1    g25788(.A1(new_n29032_), .A2(new_n29030_), .ZN(new_n29033_));
  NOR2_X1    g25789(.A1(new_n12841_), .A2(pi0039), .ZN(new_n29034_));
  NOR2_X1    g25790(.A1(new_n28998_), .A2(new_n3099_), .ZN(new_n29035_));
  NAND2_X1   g25791(.A1(new_n29035_), .A2(pi0616), .ZN(new_n29036_));
  XOR2_X1    g25792(.A1(new_n29036_), .A2(new_n29034_), .Z(new_n29037_));
  NOR2_X1    g25793(.A1(new_n14291_), .A2(new_n13378_), .ZN(new_n29038_));
  OAI21_X1   g25794(.A1(new_n13203_), .A2(new_n28937_), .B(new_n13213_), .ZN(new_n29039_));
  NAND3_X1   g25795(.A1(new_n13108_), .A2(new_n28793_), .A3(new_n29039_), .ZN(new_n29040_));
  OAI21_X1   g25796(.A1(pi0222), .A2(new_n13108_), .B(new_n29040_), .ZN(new_n29041_));
  AOI21_X1   g25797(.A1(new_n29041_), .A2(pi0038), .B(new_n29038_), .ZN(new_n29042_));
  OAI21_X1   g25798(.A1(new_n29042_), .A2(new_n29037_), .B(new_n3289_), .ZN(new_n29043_));
  INV_X1     g25799(.I(new_n13570_), .ZN(new_n29044_));
  NOR2_X1    g25800(.A1(new_n29044_), .A2(pi0680), .ZN(new_n29045_));
  NAND3_X1   g25801(.A1(new_n13480_), .A2(pi0616), .A3(new_n13379_), .ZN(new_n29046_));
  OAI21_X1   g25802(.A1(new_n29045_), .A2(new_n29046_), .B(new_n5374_), .ZN(new_n29047_));
  NAND3_X1   g25803(.A1(new_n29047_), .A2(pi0680), .A3(new_n28838_), .ZN(new_n29048_));
  NOR2_X1    g25804(.A1(new_n5632_), .A2(pi0661), .ZN(new_n29049_));
  NAND2_X1   g25805(.A1(new_n28838_), .A2(new_n29049_), .ZN(new_n29050_));
  AOI21_X1   g25806(.A1(new_n29048_), .A2(new_n28837_), .B(new_n29050_), .ZN(new_n29051_));
  AOI21_X1   g25807(.A1(new_n13494_), .A2(pi0616), .B(new_n5375_), .ZN(new_n29052_));
  INV_X1     g25808(.I(new_n29052_), .ZN(new_n29053_));
  AOI21_X1   g25809(.A1(new_n28846_), .A2(new_n5375_), .B(new_n5374_), .ZN(new_n29054_));
  OAI21_X1   g25810(.A1(new_n13560_), .A2(new_n29053_), .B(new_n29054_), .ZN(new_n29055_));
  NAND2_X1   g25811(.A1(new_n29055_), .A2(new_n28849_), .ZN(new_n29056_));
  NAND3_X1   g25812(.A1(new_n29056_), .A2(new_n28846_), .A3(new_n29049_), .ZN(new_n29057_));
  NAND2_X1   g25813(.A1(new_n29057_), .A2(pi0222), .ZN(new_n29058_));
  XOR2_X1    g25814(.A1(new_n29058_), .A2(new_n28813_), .Z(new_n29059_));
  NAND2_X1   g25815(.A1(new_n29059_), .A2(new_n29051_), .ZN(new_n29060_));
  NOR2_X1    g25816(.A1(pi0215), .A2(pi0299), .ZN(new_n29061_));
  NAND2_X1   g25817(.A1(new_n29060_), .A2(new_n29061_), .ZN(new_n29062_));
  NOR3_X1    g25818(.A1(new_n28844_), .A2(new_n13210_), .A3(new_n28937_), .ZN(new_n29063_));
  NAND2_X1   g25819(.A1(new_n13323_), .A2(new_n5375_), .ZN(new_n29064_));
  NOR2_X1    g25820(.A1(new_n26505_), .A2(new_n13398_), .ZN(new_n29065_));
  NAND3_X1   g25821(.A1(new_n29064_), .A2(pi0616), .A3(new_n29065_), .ZN(new_n29066_));
  NOR2_X1    g25822(.A1(pi0616), .A2(pi0661), .ZN(new_n29067_));
  AOI21_X1   g25823(.A1(new_n13390_), .A2(new_n29067_), .B(new_n5375_), .ZN(new_n29068_));
  NAND2_X1   g25824(.A1(new_n29066_), .A2(new_n29068_), .ZN(new_n29069_));
  NOR2_X1    g25825(.A1(new_n5636_), .A2(new_n5374_), .ZN(new_n29070_));
  OAI21_X1   g25826(.A1(new_n28879_), .A2(new_n12878_), .B(new_n29070_), .ZN(new_n29071_));
  AOI21_X1   g25827(.A1(new_n29071_), .A2(new_n13390_), .B(new_n12841_), .ZN(new_n29072_));
  NAND2_X1   g25828(.A1(new_n29069_), .A2(new_n29072_), .ZN(new_n29073_));
  NAND2_X1   g25829(.A1(new_n29073_), .A2(new_n5454_), .ZN(new_n29074_));
  XNOR2_X1   g25830(.A1(new_n29074_), .A2(new_n28813_), .ZN(new_n29075_));
  NOR3_X1    g25831(.A1(new_n29075_), .A2(new_n13478_), .A3(new_n29063_), .ZN(new_n29076_));
  NOR2_X1    g25832(.A1(new_n13381_), .A2(new_n12841_), .ZN(new_n29077_));
  INV_X1     g25833(.I(new_n29077_), .ZN(new_n29078_));
  OAI21_X1   g25834(.A1(pi0616), .A2(new_n13297_), .B(new_n29078_), .ZN(new_n29079_));
  NAND2_X1   g25835(.A1(new_n29079_), .A2(new_n28937_), .ZN(new_n29080_));
  AOI21_X1   g25836(.A1(new_n29080_), .A2(new_n12841_), .B(new_n13103_), .ZN(new_n29081_));
  OAI21_X1   g25837(.A1(new_n29081_), .A2(new_n28959_), .B(new_n3111_), .ZN(new_n29082_));
  AOI21_X1   g25838(.A1(new_n29062_), .A2(new_n29076_), .B(new_n29082_), .ZN(new_n29083_));
  XOR2_X1    g25839(.A1(new_n29058_), .A2(new_n28858_), .Z(new_n29084_));
  NAND2_X1   g25840(.A1(new_n29084_), .A2(new_n29051_), .ZN(new_n29085_));
  INV_X1     g25841(.I(new_n29063_), .ZN(new_n29086_));
  NAND2_X1   g25842(.A1(new_n29073_), .A2(new_n5398_), .ZN(new_n29087_));
  XOR2_X1    g25843(.A1(new_n29087_), .A2(new_n28858_), .Z(new_n29088_));
  NAND4_X1   g25844(.A1(new_n29088_), .A2(pi0039), .A3(new_n13340_), .A4(new_n29086_), .ZN(new_n29089_));
  AOI21_X1   g25845(.A1(new_n29085_), .A2(new_n3381_), .B(new_n29089_), .ZN(new_n29090_));
  NOR2_X1    g25846(.A1(new_n29090_), .A2(pi0223), .ZN(new_n29091_));
  NOR2_X1    g25847(.A1(new_n29079_), .A2(new_n28998_), .ZN(new_n29092_));
  XNOR2_X1   g25848(.A1(new_n29092_), .A2(new_n29035_), .ZN(new_n29093_));
  NAND4_X1   g25849(.A1(new_n28818_), .A2(pi0222), .A3(new_n3289_), .A4(new_n3313_), .ZN(new_n29094_));
  NOR4_X1    g25850(.A1(new_n29091_), .A2(new_n29083_), .A3(new_n29093_), .A4(new_n29094_), .ZN(new_n29095_));
  INV_X1     g25851(.I(new_n13281_), .ZN(new_n29096_));
  NAND3_X1   g25852(.A1(new_n29096_), .A2(pi0661), .A3(pi0680), .ZN(new_n29097_));
  AOI21_X1   g25853(.A1(new_n29097_), .A2(new_n12841_), .B(new_n13381_), .ZN(new_n29098_));
  NOR3_X1    g25854(.A1(new_n5376_), .A2(pi0616), .A3(new_n12842_), .ZN(new_n29099_));
  NOR2_X1    g25855(.A1(new_n13368_), .A2(new_n29099_), .ZN(new_n29100_));
  NOR3_X1    g25856(.A1(new_n28879_), .A2(pi0661), .A3(new_n5632_), .ZN(new_n29101_));
  OAI21_X1   g25857(.A1(new_n29098_), .A2(new_n29100_), .B(new_n29101_), .ZN(new_n29102_));
  NAND2_X1   g25858(.A1(new_n13264_), .A2(new_n13250_), .ZN(new_n29103_));
  XNOR2_X1   g25859(.A1(new_n29103_), .A2(new_n13252_), .ZN(new_n29104_));
  AOI21_X1   g25860(.A1(new_n29104_), .A2(new_n13249_), .B(pi0680), .ZN(new_n29105_));
  NOR3_X1    g25861(.A1(new_n29105_), .A2(new_n12841_), .A3(new_n13420_), .ZN(new_n29106_));
  NOR2_X1    g25862(.A1(new_n29106_), .A2(pi0661), .ZN(new_n29107_));
  NAND2_X1   g25863(.A1(new_n28826_), .A2(pi0680), .ZN(new_n29108_));
  OAI21_X1   g25864(.A1(new_n29107_), .A2(new_n29108_), .B(new_n28829_), .ZN(new_n29109_));
  NAND3_X1   g25865(.A1(new_n29109_), .A2(new_n28826_), .A3(new_n29049_), .ZN(new_n29110_));
  NAND2_X1   g25866(.A1(new_n29110_), .A2(new_n5454_), .ZN(new_n29111_));
  XNOR2_X1   g25867(.A1(new_n29111_), .A2(new_n28813_), .ZN(new_n29112_));
  OAI21_X1   g25868(.A1(new_n13535_), .A2(new_n13524_), .B(new_n29052_), .ZN(new_n29113_));
  INV_X1     g25869(.I(new_n28791_), .ZN(new_n29114_));
  AOI21_X1   g25870(.A1(new_n29114_), .A2(new_n5375_), .B(new_n5374_), .ZN(new_n29115_));
  AOI21_X1   g25871(.A1(new_n29113_), .A2(new_n29115_), .B(new_n28796_), .ZN(new_n29116_));
  NOR4_X1    g25872(.A1(new_n29116_), .A2(pi0661), .A3(new_n5632_), .A4(new_n28791_), .ZN(new_n29117_));
  NAND2_X1   g25873(.A1(new_n28806_), .A2(new_n28809_), .ZN(new_n29118_));
  OAI21_X1   g25874(.A1(new_n13290_), .A2(new_n5386_), .B(new_n13479_), .ZN(new_n29119_));
  INV_X1     g25875(.I(new_n29119_), .ZN(new_n29120_));
  OAI21_X1   g25876(.A1(new_n13103_), .A2(new_n13263_), .B(new_n29120_), .ZN(new_n29121_));
  INV_X1     g25877(.I(new_n29121_), .ZN(new_n29122_));
  NAND2_X1   g25878(.A1(new_n29119_), .A2(pi0603), .ZN(new_n29123_));
  NAND2_X1   g25879(.A1(new_n13287_), .A2(pi0603), .ZN(new_n29124_));
  XOR2_X1    g25880(.A1(new_n29123_), .A2(new_n29124_), .Z(new_n29125_));
  AOI21_X1   g25881(.A1(new_n29125_), .A2(new_n12806_), .B(new_n5382_), .ZN(new_n29126_));
  XOR2_X1    g25882(.A1(new_n29126_), .A2(new_n26490_), .Z(new_n29127_));
  NAND2_X1   g25883(.A1(new_n29127_), .A2(new_n29122_), .ZN(new_n29128_));
  NOR2_X1    g25884(.A1(new_n29120_), .A2(new_n13378_), .ZN(new_n29129_));
  OAI21_X1   g25885(.A1(new_n29129_), .A2(new_n12841_), .B(pi0680), .ZN(new_n29130_));
  NAND3_X1   g25886(.A1(new_n29122_), .A2(pi0614), .A3(new_n12841_), .ZN(new_n29131_));
  AOI21_X1   g25887(.A1(new_n29128_), .A2(new_n29130_), .B(new_n29131_), .ZN(new_n29132_));
  NOR2_X1    g25888(.A1(new_n28804_), .A2(new_n5375_), .ZN(new_n29133_));
  OAI21_X1   g25889(.A1(new_n29132_), .A2(pi0661), .B(new_n29133_), .ZN(new_n29134_));
  NAND2_X1   g25890(.A1(new_n29134_), .A2(new_n29118_), .ZN(new_n29135_));
  NAND3_X1   g25891(.A1(new_n29135_), .A2(new_n28802_), .A3(new_n29049_), .ZN(new_n29136_));
  NAND2_X1   g25892(.A1(new_n29136_), .A2(pi0222), .ZN(new_n29137_));
  XOR2_X1    g25893(.A1(new_n29137_), .A2(new_n28813_), .Z(new_n29138_));
  NAND2_X1   g25894(.A1(new_n29138_), .A2(new_n29117_), .ZN(new_n29139_));
  OAI21_X1   g25895(.A1(new_n29102_), .A2(new_n29112_), .B(new_n29139_), .ZN(new_n29140_));
  INV_X1     g25896(.I(new_n13149_), .ZN(new_n29141_));
  NAND2_X1   g25897(.A1(new_n29141_), .A2(new_n13147_), .ZN(new_n29142_));
  NAND2_X1   g25898(.A1(new_n13145_), .A2(pi0603), .ZN(new_n29143_));
  NOR3_X1    g25899(.A1(new_n13155_), .A2(new_n5794_), .A3(new_n13124_), .ZN(new_n29144_));
  XOR2_X1    g25900(.A1(new_n29144_), .A2(new_n29143_), .Z(new_n29145_));
  AOI21_X1   g25901(.A1(new_n13192_), .A2(new_n12841_), .B(new_n3099_), .ZN(new_n29146_));
  AOI21_X1   g25902(.A1(new_n29145_), .A2(new_n29146_), .B(new_n29142_), .ZN(new_n29147_));
  NAND2_X1   g25903(.A1(new_n28937_), .A2(new_n3099_), .ZN(new_n29148_));
  NOR2_X1    g25904(.A1(new_n13178_), .A2(new_n12841_), .ZN(new_n29149_));
  OR3_X2     g25905(.A1(new_n29147_), .A2(new_n29148_), .A3(new_n29149_), .Z(new_n29150_));
  NAND2_X1   g25906(.A1(new_n29150_), .A2(new_n5374_), .ZN(new_n29151_));
  AOI21_X1   g25907(.A1(new_n29151_), .A2(new_n15052_), .B(new_n3098_), .ZN(new_n29152_));
  XOR2_X1    g25908(.A1(new_n29152_), .A2(new_n11324_), .Z(new_n29153_));
  NOR2_X1    g25909(.A1(new_n13123_), .A2(new_n5794_), .ZN(new_n29154_));
  NOR3_X1    g25910(.A1(new_n13159_), .A2(new_n5794_), .A3(new_n13124_), .ZN(new_n29155_));
  XOR2_X1    g25911(.A1(new_n29155_), .A2(new_n29154_), .Z(new_n29156_));
  OAI21_X1   g25912(.A1(new_n13173_), .A2(pi0616), .B(pi0222), .ZN(new_n29157_));
  NOR2_X1    g25913(.A1(new_n29156_), .A2(new_n29157_), .ZN(new_n29158_));
  AOI21_X1   g25914(.A1(new_n13174_), .A2(pi0616), .B(new_n29148_), .ZN(new_n29159_));
  OAI21_X1   g25915(.A1(new_n29158_), .A2(new_n13136_), .B(new_n29159_), .ZN(new_n29160_));
  NAND2_X1   g25916(.A1(new_n29160_), .A2(new_n5374_), .ZN(new_n29161_));
  NAND2_X1   g25917(.A1(new_n29161_), .A2(new_n13138_), .ZN(new_n29162_));
  OAI21_X1   g25918(.A1(new_n29153_), .A2(new_n29162_), .B(new_n3259_), .ZN(new_n29163_));
  XOR2_X1    g25919(.A1(new_n29137_), .A2(new_n28857_), .Z(new_n29164_));
  INV_X1     g25920(.I(new_n29102_), .ZN(new_n29165_));
  NAND2_X1   g25921(.A1(new_n29110_), .A2(pi0224), .ZN(new_n29166_));
  XOR2_X1    g25922(.A1(new_n29166_), .A2(new_n28883_), .Z(new_n29167_));
  NAND3_X1   g25923(.A1(new_n29167_), .A2(new_n29165_), .A3(new_n29117_), .ZN(new_n29168_));
  OAI22_X1   g25924(.A1(new_n29164_), .A2(new_n29168_), .B1(pi0222), .B2(new_n3100_), .ZN(new_n29169_));
  NAND4_X1   g25925(.A1(new_n29163_), .A2(new_n29095_), .A3(new_n29140_), .A4(new_n29169_), .ZN(new_n29170_));
  XNOR2_X1   g25926(.A1(new_n29170_), .A2(new_n29043_), .ZN(new_n29171_));
  NAND2_X1   g25927(.A1(new_n28889_), .A2(pi0625), .ZN(new_n29172_));
  XOR2_X1    g25928(.A1(new_n29172_), .A2(new_n13615_), .Z(new_n29173_));
  OAI21_X1   g25929(.A1(new_n29171_), .A2(new_n29173_), .B(new_n14081_), .ZN(new_n29174_));
  NAND2_X1   g25930(.A1(new_n28889_), .A2(pi1153), .ZN(new_n29175_));
  XOR2_X1    g25931(.A1(new_n29175_), .A2(new_n13615_), .Z(new_n29176_));
  OAI21_X1   g25932(.A1(new_n29171_), .A2(new_n29176_), .B(new_n14081_), .ZN(new_n29177_));
  INV_X1     g25933(.I(new_n29177_), .ZN(new_n29178_));
  OAI21_X1   g25934(.A1(new_n29022_), .A2(new_n29174_), .B(new_n29178_), .ZN(new_n29179_));
  INV_X1     g25935(.I(new_n29179_), .ZN(new_n29180_));
  NAND3_X1   g25936(.A1(new_n29017_), .A2(pi0778), .A3(new_n28789_), .ZN(new_n29181_));
  NAND2_X1   g25937(.A1(new_n29171_), .A2(new_n13748_), .ZN(new_n29182_));
  OAI21_X1   g25938(.A1(new_n29180_), .A2(new_n29181_), .B(new_n29182_), .ZN(new_n29183_));
  NAND3_X1   g25939(.A1(new_n29183_), .A2(pi0609), .A3(pi1155), .ZN(new_n29184_));
  INV_X1     g25940(.I(new_n29181_), .ZN(new_n29185_));
  AOI22_X1   g25941(.A1(new_n29185_), .A2(new_n29179_), .B1(new_n13748_), .B2(new_n29171_), .ZN(new_n29186_));
  NAND3_X1   g25942(.A1(new_n29186_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n29187_));
  AOI21_X1   g25943(.A1(new_n29184_), .A2(new_n29187_), .B(new_n29033_), .ZN(new_n29188_));
  INV_X1     g25944(.I(new_n28895_), .ZN(new_n29189_));
  NOR2_X1    g25945(.A1(new_n29189_), .A2(new_n13783_), .ZN(new_n29190_));
  INV_X1     g25946(.I(new_n29190_), .ZN(new_n29191_));
  OAI21_X1   g25947(.A1(new_n29188_), .A2(new_n29191_), .B(pi0785), .ZN(new_n29192_));
  INV_X1     g25948(.I(new_n16780_), .ZN(new_n29193_));
  NAND3_X1   g25949(.A1(new_n29183_), .A2(pi0609), .A3(pi1155), .ZN(new_n29194_));
  NAND3_X1   g25950(.A1(new_n29186_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n29195_));
  AOI21_X1   g25951(.A1(new_n29194_), .A2(new_n29195_), .B(new_n29033_), .ZN(new_n29196_));
  NOR4_X1    g25952(.A1(new_n29196_), .A2(new_n29193_), .A3(new_n28905_), .A4(new_n29186_), .ZN(new_n29197_));
  NAND2_X1   g25953(.A1(new_n29197_), .A2(new_n29192_), .ZN(new_n29198_));
  AOI21_X1   g25954(.A1(new_n29186_), .A2(pi1155), .B(new_n14694_), .ZN(new_n29199_));
  NOR3_X1    g25955(.A1(new_n29183_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n29200_));
  OAI21_X1   g25956(.A1(new_n29200_), .A2(new_n29199_), .B(new_n29024_), .ZN(new_n29201_));
  AOI21_X1   g25957(.A1(new_n29201_), .A2(new_n29190_), .B(new_n13801_), .ZN(new_n29202_));
  AOI21_X1   g25958(.A1(new_n29186_), .A2(pi0609), .B(new_n14694_), .ZN(new_n29203_));
  NOR3_X1    g25959(.A1(new_n29183_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n29204_));
  OAI21_X1   g25960(.A1(new_n29204_), .A2(new_n29203_), .B(new_n29024_), .ZN(new_n29205_));
  NAND4_X1   g25961(.A1(new_n29205_), .A2(new_n16780_), .A3(new_n28901_), .A4(new_n29183_), .ZN(new_n29206_));
  NAND2_X1   g25962(.A1(new_n29206_), .A2(new_n29202_), .ZN(new_n29207_));
  NAND2_X1   g25963(.A1(new_n29207_), .A2(new_n29198_), .ZN(new_n29208_));
  OAI21_X1   g25964(.A1(new_n29026_), .A2(pi0618), .B(new_n13824_), .ZN(new_n29209_));
  OAI21_X1   g25965(.A1(new_n29209_), .A2(new_n28912_), .B(new_n13816_), .ZN(new_n29210_));
  AOI21_X1   g25966(.A1(new_n28929_), .A2(new_n13836_), .B(pi0618), .ZN(new_n29211_));
  INV_X1     g25967(.I(new_n29211_), .ZN(new_n29212_));
  NAND4_X1   g25968(.A1(new_n29208_), .A2(pi0781), .A3(new_n29210_), .A4(new_n29212_), .ZN(new_n29213_));
  NOR2_X1    g25969(.A1(new_n29206_), .A2(new_n29202_), .ZN(new_n29214_));
  NOR2_X1    g25970(.A1(new_n29197_), .A2(new_n29192_), .ZN(new_n29215_));
  OAI21_X1   g25971(.A1(new_n29214_), .A2(new_n29215_), .B(new_n29210_), .ZN(new_n29216_));
  NOR2_X1    g25972(.A1(new_n29211_), .A2(new_n13855_), .ZN(new_n29217_));
  OAI21_X1   g25973(.A1(new_n29214_), .A2(new_n29215_), .B(new_n29217_), .ZN(new_n29218_));
  NAND3_X1   g25974(.A1(new_n29216_), .A2(new_n29218_), .A3(pi0781), .ZN(new_n29219_));
  NAND2_X1   g25975(.A1(new_n29219_), .A2(new_n29213_), .ZN(new_n29220_));
  NAND3_X1   g25976(.A1(new_n29220_), .A2(pi0619), .A3(pi1159), .ZN(new_n29221_));
  NAND4_X1   g25977(.A1(new_n29219_), .A2(new_n29213_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n29222_));
  AOI21_X1   g25978(.A1(new_n29221_), .A2(new_n29222_), .B(new_n29029_), .ZN(new_n29223_));
  OAI21_X1   g25979(.A1(new_n29223_), .A2(new_n20003_), .B(new_n28936_), .ZN(new_n29224_));
  NAND3_X1   g25980(.A1(new_n28925_), .A2(pi0619), .A3(pi1159), .ZN(new_n29225_));
  NAND4_X1   g25981(.A1(new_n28924_), .A2(new_n13860_), .A3(new_n28919_), .A4(pi1159), .ZN(new_n29226_));
  AOI21_X1   g25982(.A1(new_n29225_), .A2(new_n29226_), .B(new_n28788_), .ZN(new_n29227_));
  NAND4_X1   g25983(.A1(new_n28936_), .A2(new_n29227_), .A3(pi0789), .A4(new_n28925_), .ZN(new_n29228_));
  INV_X1     g25984(.I(new_n29228_), .ZN(new_n29229_));
  AOI21_X1   g25985(.A1(new_n28934_), .A2(pi0619), .B(new_n13904_), .ZN(new_n29230_));
  NOR3_X1    g25986(.A1(new_n28925_), .A2(new_n13860_), .A3(new_n13903_), .ZN(new_n29231_));
  OAI21_X1   g25987(.A1(new_n29230_), .A2(new_n29231_), .B(new_n28789_), .ZN(new_n29232_));
  NAND2_X1   g25988(.A1(new_n29232_), .A2(pi0789), .ZN(new_n29233_));
  AOI21_X1   g25989(.A1(new_n28934_), .A2(pi1159), .B(new_n13904_), .ZN(new_n29234_));
  INV_X1     g25990(.I(new_n29226_), .ZN(new_n29235_));
  OAI21_X1   g25991(.A1(new_n29234_), .A2(new_n29235_), .B(new_n28789_), .ZN(new_n29236_));
  NOR3_X1    g25992(.A1(new_n29236_), .A2(new_n13896_), .A3(new_n28934_), .ZN(new_n29237_));
  NOR2_X1    g25993(.A1(new_n29237_), .A2(new_n29233_), .ZN(new_n29238_));
  NOR2_X1    g25994(.A1(new_n29238_), .A2(new_n29229_), .ZN(new_n29239_));
  AOI21_X1   g25995(.A1(new_n29239_), .A2(new_n13962_), .B(new_n18976_), .ZN(new_n29240_));
  NOR2_X1    g25996(.A1(new_n28934_), .A2(new_n13896_), .ZN(new_n29241_));
  NAND2_X1   g25997(.A1(new_n29227_), .A2(new_n29241_), .ZN(new_n29242_));
  NAND3_X1   g25998(.A1(new_n29242_), .A2(pi0789), .A3(new_n29232_), .ZN(new_n29243_));
  NAND4_X1   g25999(.A1(new_n29243_), .A2(new_n13901_), .A3(new_n13962_), .A4(new_n29228_), .ZN(new_n29244_));
  INV_X1     g26000(.I(new_n29244_), .ZN(new_n29245_));
  OAI21_X1   g26001(.A1(new_n29240_), .A2(new_n29245_), .B(new_n28789_), .ZN(new_n29246_));
  NOR2_X1    g26002(.A1(new_n29028_), .A2(new_n14162_), .ZN(new_n29247_));
  XOR2_X1    g26003(.A1(new_n29247_), .A2(new_n16829_), .Z(new_n29248_));
  NOR2_X1    g26004(.A1(new_n29248_), .A2(new_n28788_), .ZN(new_n29249_));
  INV_X1     g26005(.I(new_n29249_), .ZN(new_n29250_));
  AOI21_X1   g26006(.A1(new_n29239_), .A2(new_n13963_), .B(new_n19028_), .ZN(new_n29251_));
  NAND4_X1   g26007(.A1(new_n29243_), .A2(new_n13901_), .A3(new_n13963_), .A4(new_n29228_), .ZN(new_n29252_));
  INV_X1     g26008(.I(new_n29252_), .ZN(new_n29253_));
  OAI21_X1   g26009(.A1(new_n29251_), .A2(new_n29253_), .B(new_n28789_), .ZN(new_n29254_));
  NAND4_X1   g26010(.A1(new_n29246_), .A2(new_n29254_), .A3(new_n29220_), .A4(new_n29250_), .ZN(new_n29255_));
  NAND2_X1   g26011(.A1(pi0788), .A2(pi0789), .ZN(new_n29256_));
  NAND2_X1   g26012(.A1(new_n29255_), .A2(new_n29256_), .ZN(new_n29257_));
  NAND2_X1   g26013(.A1(new_n29243_), .A2(new_n29228_), .ZN(new_n29258_));
  NAND3_X1   g26014(.A1(new_n29258_), .A2(pi0626), .A3(new_n13962_), .ZN(new_n29259_));
  AOI21_X1   g26015(.A1(new_n29259_), .A2(new_n29244_), .B(new_n28788_), .ZN(new_n29260_));
  NAND3_X1   g26016(.A1(new_n29258_), .A2(pi0626), .A3(new_n13963_), .ZN(new_n29261_));
  AOI21_X1   g26017(.A1(new_n29261_), .A2(new_n29252_), .B(new_n28788_), .ZN(new_n29262_));
  NOR3_X1    g26018(.A1(new_n29260_), .A2(new_n29262_), .A3(new_n29249_), .ZN(new_n29263_));
  AOI21_X1   g26019(.A1(new_n29263_), .A2(new_n15479_), .B(new_n16423_), .ZN(new_n29264_));
  NAND2_X1   g26020(.A1(new_n29257_), .A2(new_n29264_), .ZN(new_n29265_));
  AND3_X2    g26021(.A1(new_n29220_), .A2(pi0619), .A3(pi1159), .Z(new_n29266_));
  NOR3_X1    g26022(.A1(new_n29220_), .A2(new_n13860_), .A3(pi1159), .ZN(new_n29267_));
  OAI21_X1   g26023(.A1(new_n29266_), .A2(new_n29267_), .B(new_n29028_), .ZN(new_n29268_));
  NOR2_X1    g26024(.A1(new_n29227_), .A2(pi0648), .ZN(new_n29269_));
  NAND2_X1   g26025(.A1(new_n29268_), .A2(new_n29269_), .ZN(new_n29270_));
  AOI21_X1   g26026(.A1(new_n29265_), .A2(new_n29224_), .B(new_n29270_), .ZN(new_n29271_));
  NOR2_X1    g26027(.A1(new_n28789_), .A2(new_n13994_), .ZN(new_n29272_));
  NOR2_X1    g26028(.A1(new_n28788_), .A2(new_n16372_), .ZN(new_n29273_));
  AOI21_X1   g26029(.A1(new_n29239_), .A2(new_n16372_), .B(new_n29273_), .ZN(new_n29274_));
  AOI21_X1   g26030(.A1(new_n29274_), .A2(new_n13994_), .B(new_n29272_), .ZN(new_n29275_));
  NOR2_X1    g26031(.A1(new_n28788_), .A2(new_n14059_), .ZN(new_n29276_));
  INV_X1     g26032(.I(new_n29025_), .ZN(new_n29277_));
  OAI21_X1   g26033(.A1(new_n29033_), .A2(new_n13803_), .B(new_n29277_), .ZN(new_n29278_));
  NAND4_X1   g26034(.A1(new_n29278_), .A2(new_n13880_), .A3(new_n15395_), .A4(new_n28789_), .ZN(new_n29279_));
  NAND4_X1   g26035(.A1(new_n29026_), .A2(new_n13880_), .A3(new_n15395_), .A4(new_n28788_), .ZN(new_n29280_));
  AOI21_X1   g26036(.A1(new_n29280_), .A2(new_n29279_), .B(new_n14059_), .ZN(new_n29281_));
  NOR2_X1    g26037(.A1(new_n29281_), .A2(new_n29276_), .ZN(new_n29282_));
  AOI21_X1   g26038(.A1(new_n29282_), .A2(pi0647), .B(new_n14008_), .ZN(new_n29283_));
  NOR4_X1    g26039(.A1(new_n29281_), .A2(new_n14005_), .A3(pi1157), .A4(new_n29276_), .ZN(new_n29284_));
  OAI21_X1   g26040(.A1(new_n29283_), .A2(new_n29284_), .B(new_n28789_), .ZN(new_n29285_));
  NAND2_X1   g26041(.A1(new_n29285_), .A2(pi0630), .ZN(new_n29286_));
  AOI21_X1   g26042(.A1(new_n29282_), .A2(pi1157), .B(new_n14008_), .ZN(new_n29287_));
  NOR4_X1    g26043(.A1(new_n29281_), .A2(pi0647), .A3(new_n14006_), .A4(new_n29276_), .ZN(new_n29288_));
  OAI21_X1   g26044(.A1(new_n29287_), .A2(new_n29288_), .B(new_n28789_), .ZN(new_n29289_));
  NAND2_X1   g26045(.A1(new_n29289_), .A2(new_n14010_), .ZN(new_n29290_));
  AOI21_X1   g26046(.A1(new_n29286_), .A2(new_n29290_), .B(new_n12776_), .ZN(new_n29291_));
  OAI21_X1   g26047(.A1(new_n29291_), .A2(new_n16576_), .B(new_n16574_), .ZN(new_n29292_));
  NOR2_X1    g26048(.A1(new_n29292_), .A2(new_n29275_), .ZN(new_n29293_));
  NAND2_X1   g26049(.A1(new_n29280_), .A2(new_n29279_), .ZN(new_n29294_));
  INV_X1     g26050(.I(new_n29294_), .ZN(new_n29295_));
  NAND2_X1   g26051(.A1(new_n28788_), .A2(pi0628), .ZN(new_n29296_));
  AOI22_X1   g26052(.A1(new_n29295_), .A2(pi0628), .B1(new_n13991_), .B2(new_n29296_), .ZN(new_n29297_));
  NOR2_X1    g26053(.A1(new_n13985_), .A2(new_n13942_), .ZN(new_n29298_));
  AOI22_X1   g26054(.A1(new_n29295_), .A2(pi0628), .B1(new_n28789_), .B2(new_n29298_), .ZN(new_n29299_));
  OR3_X2     g26055(.A1(new_n29297_), .A2(new_n29299_), .A3(new_n12777_), .Z(new_n29300_));
  AOI21_X1   g26056(.A1(new_n29300_), .A2(new_n29274_), .B(new_n16875_), .ZN(new_n29301_));
  OAI21_X1   g26057(.A1(new_n29271_), .A2(new_n29293_), .B(new_n29301_), .ZN(new_n29302_));
  NOR2_X1    g26058(.A1(new_n28788_), .A2(new_n14211_), .ZN(new_n29303_));
  INV_X1     g26059(.I(new_n29303_), .ZN(new_n29304_));
  INV_X1     g26060(.I(new_n29272_), .ZN(new_n29305_));
  INV_X1     g26061(.I(new_n29273_), .ZN(new_n29306_));
  NAND3_X1   g26062(.A1(new_n29243_), .A2(new_n16372_), .A3(new_n29228_), .ZN(new_n29307_));
  NAND3_X1   g26063(.A1(new_n29307_), .A2(new_n13994_), .A3(new_n29306_), .ZN(new_n29308_));
  NAND3_X1   g26064(.A1(new_n29308_), .A2(new_n14211_), .A3(new_n29305_), .ZN(new_n29309_));
  NAND3_X1   g26065(.A1(new_n29309_), .A2(pi0715), .A3(new_n29304_), .ZN(new_n29310_));
  XOR2_X1    g26066(.A1(new_n29310_), .A2(new_n14205_), .Z(new_n29311_));
  OR4_X2     g26067(.A1(new_n12776_), .A2(new_n29285_), .A3(new_n29289_), .A4(new_n29282_), .Z(new_n29312_));
  INV_X1     g26068(.I(new_n29282_), .ZN(new_n29313_));
  INV_X1     g26069(.I(new_n29289_), .ZN(new_n29314_));
  NAND3_X1   g26070(.A1(new_n29314_), .A2(pi0787), .A3(new_n29313_), .ZN(new_n29315_));
  NAND3_X1   g26071(.A1(new_n29315_), .A2(pi0787), .A3(new_n29285_), .ZN(new_n29316_));
  NAND2_X1   g26072(.A1(new_n29316_), .A2(new_n29312_), .ZN(new_n29317_));
  AOI21_X1   g26073(.A1(new_n29317_), .A2(pi0644), .B(new_n15386_), .ZN(new_n29318_));
  OAI21_X1   g26074(.A1(new_n28788_), .A2(new_n29311_), .B(new_n29318_), .ZN(new_n29319_));
  AOI21_X1   g26075(.A1(new_n29275_), .A2(new_n14211_), .B(new_n29303_), .ZN(new_n29321_));
  AOI21_X1   g26076(.A1(new_n29321_), .A2(pi0644), .B(new_n14217_), .ZN(new_n29322_));
  AND4_X2    g26077(.A1(pi0644), .A2(new_n29309_), .A3(new_n14200_), .A4(new_n29304_), .Z(new_n29323_));
  OAI21_X1   g26078(.A1(new_n29322_), .A2(new_n29323_), .B(new_n28789_), .ZN(new_n29324_));
  AOI21_X1   g26079(.A1(new_n29317_), .A2(new_n14204_), .B(new_n19370_), .ZN(new_n29325_));
  NOR3_X1    g26080(.A1(new_n29302_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n29327_));
  AOI21_X1   g26081(.A1(new_n29302_), .A2(new_n29319_), .B(new_n14204_), .ZN(new_n29328_));
  AOI22_X1   g26082(.A1(new_n29263_), .A2(new_n29220_), .B1(pi0788), .B2(pi0789), .ZN(new_n29329_));
  NAND4_X1   g26083(.A1(new_n29246_), .A2(new_n29254_), .A3(new_n15479_), .A4(new_n29250_), .ZN(new_n29330_));
  NAND2_X1   g26084(.A1(new_n29330_), .A2(new_n16424_), .ZN(new_n29331_));
  OAI21_X1   g26085(.A1(new_n29329_), .A2(new_n29331_), .B(new_n29224_), .ZN(new_n29332_));
  INV_X1     g26086(.I(new_n29270_), .ZN(new_n29333_));
  AOI21_X1   g26087(.A1(new_n29332_), .A2(new_n29333_), .B(new_n29293_), .ZN(new_n29334_));
  INV_X1     g26088(.I(new_n29301_), .ZN(new_n29335_));
  AOI21_X1   g26089(.A1(new_n29325_), .A2(new_n29324_), .B(pi0644), .ZN(new_n29336_));
  NOR4_X1    g26090(.A1(new_n29334_), .A2(new_n29336_), .A3(new_n12775_), .A4(new_n29335_), .ZN(new_n29337_));
  NOR3_X1    g26091(.A1(new_n29328_), .A2(new_n12775_), .A3(new_n29337_), .ZN(new_n29338_));
  OAI21_X1   g26092(.A1(new_n29338_), .A2(new_n29327_), .B(new_n7240_), .ZN(new_n29339_));
  NAND2_X1   g26093(.A1(po1038), .A2(pi0222), .ZN(new_n29340_));
  NAND2_X1   g26094(.A1(new_n29339_), .A2(new_n29340_), .ZN(po0379));
  NOR2_X1    g26095(.A1(new_n12977_), .A2(pi0039), .ZN(new_n29342_));
  AOI22_X1   g26096(.A1(new_n14300_), .A2(new_n11543_), .B1(pi0223), .B2(new_n14906_), .ZN(new_n29343_));
  OR3_X2     g26097(.A1(new_n29343_), .A2(new_n3098_), .A3(new_n17045_), .Z(new_n29344_));
  NOR2_X1    g26098(.A1(new_n29344_), .A2(new_n29342_), .ZN(new_n29345_));
  INV_X1     g26099(.I(new_n29345_), .ZN(new_n29346_));
  NOR2_X1    g26100(.A1(new_n29346_), .A2(new_n13776_), .ZN(new_n29347_));
  INV_X1     g26101(.I(new_n29347_), .ZN(new_n29348_));
  AOI21_X1   g26102(.A1(pi0039), .A2(pi0223), .B(new_n3259_), .ZN(new_n29349_));
  AOI21_X1   g26103(.A1(new_n14291_), .A2(new_n3090_), .B(pi0039), .ZN(new_n29350_));
  NOR2_X1    g26104(.A1(new_n13103_), .A2(new_n5379_), .ZN(new_n29351_));
  NOR2_X1    g26105(.A1(new_n14291_), .A2(new_n29351_), .ZN(new_n29352_));
  INV_X1     g26106(.I(new_n29352_), .ZN(new_n29353_));
  NAND2_X1   g26107(.A1(new_n29353_), .A2(new_n29350_), .ZN(new_n29354_));
  AOI21_X1   g26108(.A1(new_n29354_), .A2(new_n29349_), .B(new_n3290_), .ZN(new_n29355_));
  INV_X1     g26109(.I(new_n29355_), .ZN(new_n29356_));
  NOR3_X1    g26110(.A1(new_n12809_), .A2(new_n5381_), .A3(new_n29351_), .ZN(new_n29357_));
  INV_X1     g26111(.I(new_n29357_), .ZN(new_n29358_));
  NOR2_X1    g26112(.A1(new_n13530_), .A2(new_n5382_), .ZN(new_n29359_));
  XNOR2_X1   g26113(.A1(new_n29359_), .A2(new_n26490_), .ZN(new_n29360_));
  OAI21_X1   g26114(.A1(new_n29360_), .A2(new_n13276_), .B(new_n29358_), .ZN(new_n29361_));
  NOR2_X1    g26115(.A1(new_n29361_), .A2(new_n5632_), .ZN(new_n29362_));
  AOI21_X1   g26116(.A1(new_n13273_), .A2(pi0642), .B(new_n12945_), .ZN(new_n29363_));
  NAND2_X1   g26117(.A1(new_n29361_), .A2(new_n5635_), .ZN(new_n29364_));
  XNOR2_X1   g26118(.A1(new_n29364_), .A2(new_n12822_), .ZN(new_n29365_));
  NOR2_X1    g26119(.A1(new_n29365_), .A2(new_n29363_), .ZN(new_n29366_));
  NOR3_X1    g26120(.A1(new_n29366_), .A2(new_n5455_), .A3(new_n29362_), .ZN(new_n29367_));
  NOR2_X1    g26121(.A1(new_n14317_), .A2(new_n5379_), .ZN(new_n29368_));
  AOI21_X1   g26122(.A1(new_n5379_), .A2(new_n12826_), .B(new_n29368_), .ZN(new_n29369_));
  NOR2_X1    g26123(.A1(new_n5635_), .A2(pi0681), .ZN(new_n29370_));
  NAND2_X1   g26124(.A1(new_n12818_), .A2(new_n29370_), .ZN(new_n29371_));
  NAND3_X1   g26125(.A1(new_n29371_), .A2(new_n5454_), .A3(new_n29351_), .ZN(new_n29372_));
  AOI21_X1   g26126(.A1(new_n29369_), .A2(new_n29372_), .B(new_n5377_), .ZN(new_n29373_));
  NAND2_X1   g26127(.A1(new_n29369_), .A2(pi0681), .ZN(new_n29374_));
  AOI21_X1   g26128(.A1(new_n29373_), .A2(new_n29374_), .B(new_n3090_), .ZN(new_n29375_));
  INV_X1     g26129(.I(new_n29375_), .ZN(new_n29376_));
  AOI21_X1   g26130(.A1(new_n12809_), .A2(pi0223), .B(new_n3313_), .ZN(new_n29377_));
  AOI21_X1   g26131(.A1(new_n29377_), .A2(pi0215), .B(pi0642), .ZN(new_n29378_));
  OAI21_X1   g26132(.A1(new_n29378_), .A2(new_n13364_), .B(new_n3313_), .ZN(new_n29379_));
  INV_X1     g26133(.I(new_n29379_), .ZN(new_n29380_));
  OAI21_X1   g26134(.A1(new_n29367_), .A2(new_n29376_), .B(new_n29380_), .ZN(new_n29381_));
  NOR2_X1    g26135(.A1(pi0642), .A2(pi0681), .ZN(new_n29382_));
  AOI21_X1   g26136(.A1(new_n13203_), .A2(pi0642), .B(new_n5635_), .ZN(new_n29383_));
  NOR2_X1    g26137(.A1(new_n13262_), .A2(new_n29383_), .ZN(new_n29384_));
  AOI21_X1   g26138(.A1(new_n13262_), .A2(new_n29351_), .B(new_n5632_), .ZN(new_n29385_));
  NOR2_X1    g26139(.A1(new_n29385_), .A2(new_n29384_), .ZN(new_n29386_));
  NOR2_X1    g26140(.A1(new_n5635_), .A2(pi0642), .ZN(new_n29387_));
  OR3_X2     g26141(.A1(new_n13368_), .A2(new_n5632_), .A3(new_n29387_), .Z(new_n29388_));
  AOI21_X1   g26142(.A1(new_n29388_), .A2(new_n5379_), .B(new_n13364_), .ZN(new_n29389_));
  INV_X1     g26143(.I(new_n29389_), .ZN(new_n29390_));
  NOR2_X1    g26144(.A1(new_n29386_), .A2(new_n16921_), .ZN(new_n29391_));
  NAND2_X1   g26145(.A1(new_n16920_), .A2(pi0947), .ZN(new_n29392_));
  XOR2_X1    g26146(.A1(new_n29391_), .A2(new_n29392_), .Z(new_n29393_));
  OAI21_X1   g26147(.A1(new_n29393_), .A2(new_n29390_), .B(new_n3090_), .ZN(new_n29394_));
  AND3_X2    g26148(.A1(new_n29394_), .A2(pi0947), .A3(new_n29386_), .Z(new_n29395_));
  AOI21_X1   g26149(.A1(new_n29381_), .A2(new_n29395_), .B(pi0299), .ZN(new_n29396_));
  NAND2_X1   g26150(.A1(new_n14304_), .A2(pi0642), .ZN(new_n29397_));
  AOI21_X1   g26151(.A1(new_n12862_), .A2(new_n29370_), .B(new_n29397_), .ZN(new_n29398_));
  NOR2_X1    g26152(.A1(new_n14302_), .A2(new_n5379_), .ZN(new_n29399_));
  AOI21_X1   g26153(.A1(new_n12924_), .A2(new_n5379_), .B(new_n29399_), .ZN(new_n29400_));
  NAND2_X1   g26154(.A1(new_n29400_), .A2(new_n5632_), .ZN(new_n29401_));
  AOI22_X1   g26155(.A1(new_n29401_), .A2(new_n5635_), .B1(pi0681), .B2(new_n29398_), .ZN(new_n29402_));
  NOR2_X1    g26156(.A1(new_n5455_), .A2(new_n3090_), .ZN(new_n29403_));
  NAND2_X1   g26157(.A1(new_n13276_), .A2(pi0642), .ZN(new_n29404_));
  AND2_X2    g26158(.A1(new_n28846_), .A2(new_n29404_), .Z(new_n29405_));
  NOR2_X1    g26159(.A1(new_n29405_), .A2(new_n29357_), .ZN(new_n29406_));
  NOR3_X1    g26160(.A1(new_n12890_), .A2(new_n5377_), .A3(new_n29353_), .ZN(new_n29407_));
  NOR4_X1    g26161(.A1(new_n29406_), .A2(new_n5632_), .A3(new_n5635_), .A4(new_n29407_), .ZN(new_n29408_));
  OR2_X2     g26162(.A1(new_n29408_), .A2(new_n3090_), .Z(new_n29409_));
  XOR2_X1    g26163(.A1(new_n29409_), .A2(new_n29403_), .Z(new_n29410_));
  NOR2_X1    g26164(.A1(new_n13403_), .A2(new_n29387_), .ZN(new_n29411_));
  AOI21_X1   g26165(.A1(new_n12922_), .A2(new_n29398_), .B(new_n29411_), .ZN(new_n29412_));
  NAND2_X1   g26166(.A1(new_n29412_), .A2(pi0681), .ZN(new_n29413_));
  AOI21_X1   g26167(.A1(new_n29413_), .A2(new_n5379_), .B(new_n13390_), .ZN(new_n29414_));
  NOR2_X1    g26168(.A1(new_n29414_), .A2(new_n5800_), .ZN(new_n29415_));
  NOR2_X1    g26169(.A1(new_n29415_), .A2(pi0223), .ZN(new_n29416_));
  OAI21_X1   g26170(.A1(new_n29410_), .A2(new_n29402_), .B(new_n29416_), .ZN(new_n29417_));
  INV_X1     g26171(.I(new_n29411_), .ZN(new_n29418_));
  NAND2_X1   g26172(.A1(new_n29418_), .A2(new_n5454_), .ZN(new_n29419_));
  NAND2_X1   g26173(.A1(new_n13363_), .A2(pi0642), .ZN(new_n29420_));
  OAI21_X1   g26174(.A1(new_n29419_), .A2(new_n29420_), .B(new_n5800_), .ZN(new_n29421_));
  NAND4_X1   g26175(.A1(new_n29414_), .A2(pi0215), .A3(new_n16920_), .A4(new_n29421_), .ZN(new_n29422_));
  INV_X1     g26176(.I(new_n29422_), .ZN(new_n29423_));
  NAND2_X1   g26177(.A1(new_n29417_), .A2(new_n29423_), .ZN(new_n29424_));
  NAND2_X1   g26178(.A1(new_n26522_), .A2(new_n5795_), .ZN(new_n29425_));
  INV_X1     g26179(.I(new_n29425_), .ZN(new_n29426_));
  NOR2_X1    g26180(.A1(pi0299), .A2(pi0642), .ZN(new_n29427_));
  NAND2_X1   g26181(.A1(new_n13178_), .A2(new_n29427_), .ZN(new_n29428_));
  NAND2_X1   g26182(.A1(new_n14980_), .A2(new_n3090_), .ZN(new_n29430_));
  AOI21_X1   g26183(.A1(new_n29430_), .A2(new_n29426_), .B(new_n3212_), .ZN(new_n29431_));
  INV_X1     g26184(.I(new_n29431_), .ZN(new_n29432_));
  INV_X1     g26185(.I(new_n14973_), .ZN(new_n29433_));
  AOI21_X1   g26186(.A1(new_n13173_), .A2(new_n29427_), .B(new_n3090_), .ZN(new_n29434_));
  INV_X1     g26187(.I(new_n29434_), .ZN(new_n29435_));
  AOI21_X1   g26188(.A1(new_n13174_), .A2(new_n5379_), .B(new_n3090_), .ZN(new_n29436_));
  AOI21_X1   g26189(.A1(new_n29433_), .A2(new_n29436_), .B(new_n29435_), .ZN(new_n29437_));
  AOI21_X1   g26190(.A1(new_n29432_), .A2(new_n29437_), .B(pi0039), .ZN(new_n29438_));
  OAI21_X1   g26191(.A1(new_n29424_), .A2(new_n29396_), .B(new_n29438_), .ZN(new_n29439_));
  INV_X1     g26192(.I(new_n29402_), .ZN(new_n29440_));
  XOR2_X1    g26193(.A1(new_n29409_), .A2(new_n13466_), .Z(new_n29441_));
  NAND2_X1   g26194(.A1(new_n29441_), .A2(new_n29440_), .ZN(new_n29442_));
  NAND2_X1   g26195(.A1(new_n29442_), .A2(new_n3098_), .ZN(new_n29443_));
  NOR2_X1    g26196(.A1(new_n29386_), .A2(new_n5397_), .ZN(new_n29444_));
  XOR2_X1    g26197(.A1(new_n29444_), .A2(new_n12982_), .Z(new_n29445_));
  NOR2_X1    g26198(.A1(new_n3290_), .A2(new_n3090_), .ZN(new_n29446_));
  OAI21_X1   g26199(.A1(pi0642), .A2(new_n13412_), .B(new_n29446_), .ZN(new_n29447_));
  NOR4_X1    g26200(.A1(new_n29445_), .A2(new_n13364_), .A3(new_n29390_), .A4(new_n29447_), .ZN(new_n29448_));
  NAND2_X1   g26201(.A1(new_n29443_), .A2(new_n29448_), .ZN(new_n29449_));
  INV_X1     g26202(.I(new_n29449_), .ZN(new_n29450_));
  NAND3_X1   g26203(.A1(new_n29450_), .A2(new_n29356_), .A3(new_n29439_), .ZN(new_n29451_));
  AOI21_X1   g26204(.A1(new_n29450_), .A2(new_n29439_), .B(new_n29356_), .ZN(new_n29452_));
  INV_X1     g26205(.I(new_n29452_), .ZN(new_n29453_));
  NAND3_X1   g26206(.A1(new_n29453_), .A2(new_n13776_), .A3(new_n29451_), .ZN(new_n29454_));
  NAND2_X1   g26207(.A1(new_n29454_), .A2(new_n29348_), .ZN(new_n29455_));
  INV_X1     g26208(.I(new_n29451_), .ZN(new_n29456_));
  NOR2_X1    g26209(.A1(new_n29456_), .A2(new_n29452_), .ZN(new_n29457_));
  AOI21_X1   g26210(.A1(new_n29457_), .A2(new_n13776_), .B(new_n29347_), .ZN(new_n29458_));
  AOI21_X1   g26211(.A1(new_n29458_), .A2(pi0609), .B(new_n14694_), .ZN(new_n29459_));
  INV_X1     g26212(.I(new_n29459_), .ZN(new_n29460_));
  NAND3_X1   g26213(.A1(new_n29458_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n29461_));
  AOI21_X1   g26214(.A1(new_n29460_), .A2(new_n29461_), .B(new_n29346_), .ZN(new_n29462_));
  NAND3_X1   g26215(.A1(new_n29455_), .A2(pi0609), .A3(pi1155), .ZN(new_n29463_));
  NAND3_X1   g26216(.A1(new_n29458_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n29464_));
  AOI21_X1   g26217(.A1(new_n29464_), .A2(new_n29463_), .B(new_n29346_), .ZN(new_n29465_));
  NAND4_X1   g26218(.A1(new_n29462_), .A2(pi0785), .A3(new_n29455_), .A4(new_n29465_), .ZN(new_n29466_));
  INV_X1     g26219(.I(new_n29461_), .ZN(new_n29467_));
  OAI21_X1   g26220(.A1(new_n29467_), .A2(new_n29459_), .B(new_n29345_), .ZN(new_n29468_));
  NAND3_X1   g26221(.A1(new_n29465_), .A2(pi0785), .A3(new_n29455_), .ZN(new_n29469_));
  NAND3_X1   g26222(.A1(new_n29469_), .A2(pi0785), .A3(new_n29468_), .ZN(new_n29470_));
  NAND2_X1   g26223(.A1(new_n29470_), .A2(new_n29466_), .ZN(new_n29471_));
  NAND3_X1   g26224(.A1(new_n29471_), .A2(pi0618), .A3(pi1154), .ZN(new_n29472_));
  AOI21_X1   g26225(.A1(new_n29458_), .A2(pi1155), .B(new_n14694_), .ZN(new_n29473_));
  NOR3_X1    g26226(.A1(new_n29455_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n29474_));
  OAI21_X1   g26227(.A1(new_n29473_), .A2(new_n29474_), .B(new_n29345_), .ZN(new_n29475_));
  NOR4_X1    g26228(.A1(new_n29468_), .A2(new_n29475_), .A3(new_n13801_), .A4(new_n29458_), .ZN(new_n29476_));
  NOR3_X1    g26229(.A1(new_n29475_), .A2(new_n13801_), .A3(new_n29458_), .ZN(new_n29477_));
  NOR3_X1    g26230(.A1(new_n29477_), .A2(new_n13801_), .A3(new_n29462_), .ZN(new_n29478_));
  NOR2_X1    g26231(.A1(new_n29478_), .A2(new_n29476_), .ZN(new_n29479_));
  NAND3_X1   g26232(.A1(new_n29479_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n29480_));
  AOI21_X1   g26233(.A1(new_n29480_), .A2(new_n29472_), .B(new_n29346_), .ZN(new_n29481_));
  NAND3_X1   g26234(.A1(new_n29471_), .A2(pi0618), .A3(pi1154), .ZN(new_n29482_));
  NAND4_X1   g26235(.A1(new_n29470_), .A2(new_n29466_), .A3(new_n13816_), .A4(pi1154), .ZN(new_n29483_));
  AOI21_X1   g26236(.A1(new_n29482_), .A2(new_n29483_), .B(new_n29346_), .ZN(new_n29484_));
  NAND4_X1   g26237(.A1(new_n29481_), .A2(new_n29484_), .A3(pi0781), .A4(new_n29471_), .ZN(new_n29485_));
  INV_X1     g26238(.I(new_n29485_), .ZN(new_n29486_));
  AOI21_X1   g26239(.A1(new_n29479_), .A2(pi0618), .B(new_n13819_), .ZN(new_n29487_));
  NOR3_X1    g26240(.A1(new_n29471_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n29488_));
  OAI21_X1   g26241(.A1(new_n29487_), .A2(new_n29488_), .B(new_n29345_), .ZN(new_n29489_));
  NAND2_X1   g26242(.A1(new_n29489_), .A2(pi0781), .ZN(new_n29490_));
  AOI21_X1   g26243(.A1(new_n29479_), .A2(pi1154), .B(new_n13819_), .ZN(new_n29491_));
  INV_X1     g26244(.I(new_n29483_), .ZN(new_n29492_));
  OAI21_X1   g26245(.A1(new_n29491_), .A2(new_n29492_), .B(new_n29345_), .ZN(new_n29493_));
  NOR3_X1    g26246(.A1(new_n29493_), .A2(new_n13855_), .A3(new_n29479_), .ZN(new_n29494_));
  NOR2_X1    g26247(.A1(new_n29494_), .A2(new_n29490_), .ZN(new_n29495_));
  NOR2_X1    g26248(.A1(new_n29495_), .A2(new_n29486_), .ZN(new_n29496_));
  AOI21_X1   g26249(.A1(new_n29496_), .A2(pi0619), .B(new_n13904_), .ZN(new_n29497_));
  NOR2_X1    g26250(.A1(new_n29479_), .A2(new_n13855_), .ZN(new_n29498_));
  NAND2_X1   g26251(.A1(new_n29484_), .A2(new_n29498_), .ZN(new_n29499_));
  NAND3_X1   g26252(.A1(new_n29499_), .A2(pi0781), .A3(new_n29489_), .ZN(new_n29500_));
  NAND2_X1   g26253(.A1(new_n29500_), .A2(new_n29485_), .ZN(new_n29501_));
  NOR3_X1    g26254(.A1(new_n29501_), .A2(new_n13860_), .A3(pi1159), .ZN(new_n29502_));
  OAI21_X1   g26255(.A1(new_n29497_), .A2(new_n29502_), .B(new_n29345_), .ZN(new_n29503_));
  NOR2_X1    g26256(.A1(new_n29345_), .A2(new_n13880_), .ZN(new_n29504_));
  NOR2_X1    g26257(.A1(new_n29346_), .A2(new_n13805_), .ZN(new_n29505_));
  NOR2_X1    g26258(.A1(new_n29010_), .A2(new_n5632_), .ZN(new_n29506_));
  INV_X1     g26259(.I(new_n29506_), .ZN(new_n29507_));
  AOI21_X1   g26260(.A1(new_n13109_), .A2(pi0223), .B(new_n3259_), .ZN(new_n29508_));
  AOI21_X1   g26261(.A1(new_n29507_), .A2(new_n29508_), .B(new_n3290_), .ZN(new_n29509_));
  INV_X1     g26262(.I(new_n12920_), .ZN(new_n29510_));
  XOR2_X1    g26263(.A1(new_n28980_), .A2(new_n29510_), .Z(new_n29511_));
  OAI22_X1   g26264(.A1(new_n29511_), .A2(new_n12919_), .B1(new_n28981_), .B2(new_n5632_), .ZN(new_n29512_));
  NAND2_X1   g26265(.A1(new_n29512_), .A2(pi0223), .ZN(new_n29513_));
  XOR2_X1    g26266(.A1(new_n29513_), .A2(new_n13466_), .Z(new_n29514_));
  NOR3_X1    g26267(.A1(new_n12908_), .A2(new_n5632_), .A3(new_n28976_), .ZN(new_n29515_));
  XOR2_X1    g26268(.A1(new_n29515_), .A2(new_n12867_), .Z(new_n29516_));
  NAND2_X1   g26269(.A1(new_n13707_), .A2(pi0681), .ZN(new_n29517_));
  INV_X1     g26270(.I(new_n29517_), .ZN(new_n29518_));
  NOR2_X1    g26271(.A1(new_n5375_), .A2(new_n5632_), .ZN(new_n29519_));
  NAND2_X1   g26272(.A1(new_n13691_), .A2(new_n29519_), .ZN(new_n29520_));
  NAND2_X1   g26273(.A1(new_n29520_), .A2(new_n5398_), .ZN(new_n29521_));
  XOR2_X1    g26274(.A1(new_n29521_), .A2(new_n12981_), .Z(new_n29522_));
  NOR4_X1    g26275(.A1(new_n29522_), .A2(new_n3090_), .A3(new_n5632_), .A4(new_n28963_), .ZN(new_n29523_));
  OAI21_X1   g26276(.A1(new_n29523_), .A2(new_n3091_), .B(new_n29518_), .ZN(new_n29524_));
  AOI21_X1   g26277(.A1(new_n29524_), .A2(new_n3097_), .B(new_n29516_), .ZN(new_n29525_));
  INV_X1     g26278(.I(new_n29519_), .ZN(new_n29526_));
  OAI21_X1   g26279(.A1(new_n13155_), .A2(new_n3090_), .B(pi0299), .ZN(new_n29527_));
  NOR3_X1    g26280(.A1(new_n29527_), .A2(new_n13141_), .A3(new_n29526_), .ZN(new_n29528_));
  NOR3_X1    g26281(.A1(new_n29527_), .A2(new_n29001_), .A3(new_n29519_), .ZN(new_n29529_));
  OAI21_X1   g26282(.A1(new_n29529_), .A2(new_n29528_), .B(pi0223), .ZN(new_n29530_));
  OAI21_X1   g26283(.A1(new_n13159_), .A2(new_n3090_), .B(new_n3098_), .ZN(new_n29531_));
  NOR3_X1    g26284(.A1(new_n15066_), .A2(new_n29526_), .A3(new_n29531_), .ZN(new_n29532_));
  NOR3_X1    g26285(.A1(new_n29531_), .A2(new_n13134_), .A3(new_n29519_), .ZN(new_n29533_));
  NOR2_X1    g26286(.A1(new_n29532_), .A2(new_n29533_), .ZN(new_n29534_));
  NOR2_X1    g26287(.A1(new_n29534_), .A2(new_n3090_), .ZN(new_n29535_));
  NOR2_X1    g26288(.A1(new_n29535_), .A2(new_n15600_), .ZN(new_n29536_));
  AOI22_X1   g26289(.A1(new_n29536_), .A2(new_n29530_), .B1(new_n29514_), .B2(new_n29525_), .ZN(new_n29537_));
  NOR2_X1    g26290(.A1(new_n28949_), .A2(new_n5632_), .ZN(new_n29538_));
  NOR2_X1    g26291(.A1(new_n5454_), .A2(new_n3090_), .ZN(new_n29539_));
  AOI21_X1   g26292(.A1(new_n12828_), .A2(new_n29539_), .B(pi0681), .ZN(new_n29540_));
  OAI21_X1   g26293(.A1(new_n29540_), .A2(new_n28945_), .B(new_n5455_), .ZN(new_n29541_));
  NOR3_X1    g26294(.A1(new_n28649_), .A2(pi0681), .A3(new_n28666_), .ZN(new_n29542_));
  OAI21_X1   g26295(.A1(new_n29538_), .A2(new_n29541_), .B(new_n29542_), .ZN(new_n29543_));
  NOR2_X1    g26296(.A1(new_n28963_), .A2(new_n5632_), .ZN(new_n29544_));
  NAND2_X1   g26297(.A1(new_n29520_), .A2(new_n5454_), .ZN(new_n29545_));
  XNOR2_X1   g26298(.A1(new_n29545_), .A2(new_n29403_), .ZN(new_n29546_));
  NAND2_X1   g26299(.A1(new_n3313_), .A2(pi0215), .ZN(new_n29547_));
  AOI21_X1   g26300(.A1(new_n29546_), .A2(new_n29544_), .B(new_n29547_), .ZN(new_n29548_));
  AOI21_X1   g26301(.A1(new_n29548_), .A2(new_n29543_), .B(new_n29377_), .ZN(new_n29549_));
  OAI21_X1   g26302(.A1(new_n29549_), .A2(new_n29517_), .B(new_n3098_), .ZN(new_n29550_));
  XNOR2_X1   g26303(.A1(new_n29513_), .A2(new_n29403_), .ZN(new_n29551_));
  NOR2_X1    g26304(.A1(new_n5632_), .A2(pi0223), .ZN(new_n29552_));
  NAND2_X1   g26305(.A1(new_n13712_), .A2(new_n29552_), .ZN(new_n29553_));
  NAND4_X1   g26306(.A1(new_n29553_), .A2(pi0215), .A3(pi0223), .A4(new_n3289_), .ZN(new_n29554_));
  NOR2_X1    g26307(.A1(new_n29516_), .A2(new_n29554_), .ZN(new_n29555_));
  NAND3_X1   g26308(.A1(new_n29551_), .A2(new_n29550_), .A3(new_n29555_), .ZN(new_n29556_));
  OR3_X2     g26309(.A1(new_n29537_), .A2(new_n29509_), .A3(new_n29556_), .Z(new_n29557_));
  OAI21_X1   g26310(.A1(new_n29537_), .A2(new_n29556_), .B(new_n29509_), .ZN(new_n29558_));
  NAND2_X1   g26311(.A1(new_n29557_), .A2(new_n29558_), .ZN(new_n29559_));
  NOR2_X1    g26312(.A1(new_n29559_), .A2(new_n13613_), .ZN(new_n29560_));
  XOR2_X1    g26313(.A1(new_n29560_), .A2(new_n13615_), .Z(new_n29561_));
  NAND2_X1   g26314(.A1(new_n29561_), .A2(new_n29345_), .ZN(new_n29562_));
  NAND2_X1   g26315(.A1(new_n29562_), .A2(pi0778), .ZN(new_n29563_));
  NOR2_X1    g26316(.A1(new_n29559_), .A2(new_n13614_), .ZN(new_n29564_));
  XOR2_X1    g26317(.A1(new_n29564_), .A2(new_n13615_), .Z(new_n29565_));
  NAND4_X1   g26318(.A1(new_n29565_), .A2(pi0778), .A3(new_n29345_), .A4(new_n29559_), .ZN(new_n29566_));
  XNOR2_X1   g26319(.A1(new_n29563_), .A2(new_n29566_), .ZN(new_n29567_));
  AOI21_X1   g26320(.A1(new_n29567_), .A2(new_n13805_), .B(new_n29505_), .ZN(new_n29568_));
  AOI21_X1   g26321(.A1(new_n29568_), .A2(new_n13880_), .B(new_n29504_), .ZN(new_n29569_));
  INV_X1     g26322(.I(new_n29569_), .ZN(new_n29570_));
  NOR3_X1    g26323(.A1(new_n14291_), .A2(new_n5379_), .A3(new_n13212_), .ZN(new_n29571_));
  NOR3_X1    g26324(.A1(new_n14291_), .A2(pi0642), .A3(new_n13211_), .ZN(new_n29572_));
  OAI21_X1   g26325(.A1(new_n29571_), .A2(new_n29572_), .B(new_n13379_), .ZN(new_n29573_));
  INV_X1     g26326(.I(new_n29573_), .ZN(new_n29574_));
  NOR3_X1    g26327(.A1(new_n29353_), .A2(new_n3090_), .A3(new_n29526_), .ZN(new_n29575_));
  NOR3_X1    g26328(.A1(new_n29352_), .A2(new_n3090_), .A3(new_n29519_), .ZN(new_n29576_));
  OAI21_X1   g26329(.A1(new_n29575_), .A2(new_n29576_), .B(new_n29574_), .ZN(new_n29577_));
  AOI21_X1   g26330(.A1(new_n13212_), .A2(new_n5379_), .B(new_n29526_), .ZN(new_n29578_));
  NAND3_X1   g26331(.A1(new_n29038_), .A2(new_n29351_), .A3(new_n29519_), .ZN(new_n29579_));
  XOR2_X1    g26332(.A1(new_n29579_), .A2(new_n29578_), .Z(new_n29580_));
  INV_X1     g26333(.I(new_n29580_), .ZN(new_n29581_));
  AOI21_X1   g26334(.A1(new_n29349_), .A2(new_n29350_), .B(new_n29581_), .ZN(new_n29582_));
  OAI21_X1   g26335(.A1(new_n29582_), .A2(new_n29577_), .B(new_n3289_), .ZN(new_n29583_));
  INV_X1     g26336(.I(new_n13321_), .ZN(new_n29584_));
  INV_X1     g26337(.I(new_n29061_), .ZN(new_n29585_));
  NAND2_X1   g26338(.A1(new_n13480_), .A2(new_n13379_), .ZN(new_n29589_));
  NOR2_X1    g26339(.A1(new_n29400_), .A2(new_n5377_), .ZN(new_n29593_));
  NAND2_X1   g26340(.A1(new_n5381_), .A2(pi0680), .ZN(new_n29594_));
  AOI21_X1   g26341(.A1(new_n29573_), .A2(new_n29594_), .B(new_n15019_), .ZN(new_n29595_));
  OAI21_X1   g26342(.A1(new_n29406_), .A2(pi0680), .B(pi0681), .ZN(new_n29596_));
  NOR2_X1    g26343(.A1(new_n29407_), .A2(pi0681), .ZN(new_n29597_));
  NOR4_X1    g26344(.A1(new_n29405_), .A2(new_n5377_), .A3(new_n29357_), .A4(new_n29597_), .ZN(new_n29598_));
  AOI21_X1   g26345(.A1(new_n29596_), .A2(new_n29598_), .B(new_n29595_), .ZN(new_n29599_));
  NOR3_X1    g26346(.A1(new_n13554_), .A2(new_n13551_), .A3(new_n13470_), .ZN(new_n29600_));
  NAND2_X1   g26347(.A1(new_n13494_), .A2(pi0642), .ZN(new_n29601_));
  NOR2_X1    g26348(.A1(new_n29601_), .A2(new_n12841_), .ZN(new_n29602_));
  OAI21_X1   g26349(.A1(new_n29600_), .A2(new_n29602_), .B(pi0614), .ZN(new_n29603_));
  NOR2_X1    g26350(.A1(new_n29599_), .A2(new_n29603_), .ZN(new_n29604_));
  NOR2_X1    g26351(.A1(new_n29604_), .A2(new_n3090_), .ZN(new_n29605_));
  XOR2_X1    g26352(.A1(new_n29605_), .A2(new_n29403_), .Z(new_n29606_));
  AOI21_X1   g26353(.A1(new_n29606_), .A2(new_n29593_), .B(new_n29585_), .ZN(new_n29607_));
  NOR2_X1    g26354(.A1(new_n5381_), .A2(pi0642), .ZN(new_n29608_));
  AOI21_X1   g26355(.A1(new_n13311_), .A2(new_n29608_), .B(pi0680), .ZN(new_n29609_));
  NAND2_X1   g26356(.A1(new_n13390_), .A2(new_n29382_), .ZN(new_n29610_));
  NAND4_X1   g26357(.A1(new_n29065_), .A2(new_n29610_), .A3(pi0642), .A4(pi0680), .ZN(new_n29611_));
  OAI21_X1   g26358(.A1(new_n29611_), .A2(new_n29609_), .B(new_n13365_), .ZN(new_n29612_));
  NAND4_X1   g26359(.A1(new_n29612_), .A2(new_n13279_), .A3(new_n13320_), .A4(new_n13398_), .ZN(new_n29613_));
  NOR2_X1    g26360(.A1(new_n29412_), .A2(pi0223), .ZN(new_n29614_));
  NAND2_X1   g26361(.A1(new_n29613_), .A2(new_n29614_), .ZN(new_n29615_));
  NOR2_X1    g26362(.A1(new_n29411_), .A2(new_n5455_), .ZN(new_n29616_));
  AOI21_X1   g26363(.A1(new_n29615_), .A2(new_n29616_), .B(pi0681), .ZN(new_n29617_));
  AOI21_X1   g26364(.A1(new_n13381_), .A2(pi0642), .B(new_n5382_), .ZN(new_n29618_));
  AOI21_X1   g26365(.A1(new_n13363_), .A2(pi0642), .B(pi0680), .ZN(new_n29619_));
  NAND3_X1   g26366(.A1(new_n12784_), .A2(pi0680), .A3(new_n5382_), .ZN(new_n29620_));
  AOI21_X1   g26367(.A1(new_n13212_), .A2(new_n29620_), .B(new_n29601_), .ZN(new_n29621_));
  AOI21_X1   g26368(.A1(new_n29621_), .A2(new_n29619_), .B(new_n29618_), .ZN(new_n29622_));
  NOR4_X1    g26369(.A1(new_n29607_), .A2(new_n29584_), .A3(new_n29617_), .A4(new_n29622_), .ZN(new_n29623_));
  NAND2_X1   g26370(.A1(new_n15052_), .A2(new_n29552_), .ZN(new_n29624_));
  NAND4_X1   g26371(.A1(new_n29145_), .A2(pi0223), .A3(new_n29425_), .A4(new_n29428_), .ZN(new_n29625_));
  AOI21_X1   g26372(.A1(new_n29625_), .A2(new_n13150_), .B(new_n29526_), .ZN(new_n29626_));
  AOI21_X1   g26373(.A1(new_n29626_), .A2(new_n29624_), .B(new_n3212_), .ZN(new_n29627_));
  XOR2_X1    g26374(.A1(new_n29605_), .A2(new_n13466_), .Z(new_n29628_));
  AOI21_X1   g26375(.A1(new_n29621_), .A2(new_n29618_), .B(pi0642), .ZN(new_n29629_));
  NAND2_X1   g26376(.A1(new_n13274_), .A2(new_n13279_), .ZN(new_n29630_));
  OAI21_X1   g26377(.A1(new_n29630_), .A2(new_n29629_), .B(new_n29388_), .ZN(new_n29631_));
  NAND2_X1   g26378(.A1(new_n29631_), .A2(new_n29619_), .ZN(new_n29632_));
  INV_X1     g26379(.I(new_n29385_), .ZN(new_n29633_));
  INV_X1     g26380(.I(new_n29608_), .ZN(new_n29634_));
  NOR2_X1    g26381(.A1(new_n13420_), .A2(new_n5379_), .ZN(new_n29635_));
  OAI22_X1   g26382(.A1(new_n29635_), .A2(new_n5375_), .B1(new_n13265_), .B2(new_n29634_), .ZN(new_n29636_));
  NAND4_X1   g26383(.A1(new_n29636_), .A2(new_n13249_), .A3(new_n13336_), .A4(new_n29384_), .ZN(new_n29637_));
  AOI21_X1   g26384(.A1(new_n29637_), .A2(new_n29526_), .B(new_n29633_), .ZN(new_n29638_));
  NOR2_X1    g26385(.A1(new_n29638_), .A2(new_n5397_), .ZN(new_n29639_));
  XOR2_X1    g26386(.A1(new_n29639_), .A2(new_n12982_), .Z(new_n29640_));
  OAI21_X1   g26387(.A1(new_n29640_), .A2(new_n29632_), .B(new_n3090_), .ZN(new_n29641_));
  NOR3_X1    g26388(.A1(new_n29581_), .A2(new_n3092_), .A3(new_n12809_), .ZN(new_n29642_));
  AOI21_X1   g26389(.A1(new_n29641_), .A2(new_n29642_), .B(new_n15098_), .ZN(new_n29643_));
  NOR2_X1    g26390(.A1(new_n29156_), .A2(new_n29436_), .ZN(new_n29644_));
  NAND2_X1   g26391(.A1(new_n13136_), .A2(new_n29519_), .ZN(new_n29645_));
  OAI21_X1   g26392(.A1(new_n29645_), .A2(new_n29644_), .B(new_n29435_), .ZN(new_n29646_));
  NAND4_X1   g26393(.A1(new_n29646_), .A2(new_n13138_), .A3(new_n29552_), .A4(new_n29593_), .ZN(new_n29647_));
  NOR4_X1    g26394(.A1(new_n29647_), .A2(new_n29627_), .A3(new_n29628_), .A4(new_n29643_), .ZN(new_n29648_));
  NAND4_X1   g26395(.A1(new_n29595_), .A2(new_n13494_), .A3(pi0642), .A4(new_n5381_), .ZN(new_n29650_));
  NOR3_X1    g26396(.A1(new_n29366_), .A2(new_n5455_), .A3(new_n29650_), .ZN(new_n29651_));
  OAI21_X1   g26397(.A1(new_n29651_), .A2(new_n29519_), .B(new_n29362_), .ZN(new_n29652_));
  NOR2_X1    g26398(.A1(new_n3312_), .A2(pi0223), .ZN(new_n29653_));
  NOR2_X1    g26399(.A1(new_n29638_), .A2(new_n5455_), .ZN(new_n29654_));
  XOR2_X1    g26400(.A1(new_n29654_), .A2(new_n29403_), .Z(new_n29655_));
  NAND2_X1   g26401(.A1(new_n29125_), .A2(new_n12806_), .ZN(new_n29656_));
  NAND2_X1   g26402(.A1(new_n29656_), .A2(new_n13336_), .ZN(new_n29657_));
  AOI21_X1   g26403(.A1(new_n29122_), .A2(new_n29608_), .B(pi0680), .ZN(new_n29658_));
  NOR4_X1    g26404(.A1(new_n29658_), .A2(new_n5379_), .A3(new_n13378_), .A4(new_n29120_), .ZN(new_n29659_));
  NAND3_X1   g26405(.A1(new_n29659_), .A2(new_n29657_), .A3(new_n29373_), .ZN(new_n29660_));
  NAND2_X1   g26406(.A1(new_n29660_), .A2(new_n29526_), .ZN(new_n29661_));
  INV_X1     g26407(.I(new_n29377_), .ZN(new_n29662_));
  NAND3_X1   g26408(.A1(new_n29580_), .A2(pi0223), .A3(new_n12784_), .ZN(new_n29663_));
  AOI21_X1   g26409(.A1(new_n29662_), .A2(new_n29577_), .B(new_n29663_), .ZN(new_n29664_));
  OAI21_X1   g26410(.A1(new_n29664_), .A2(pi0215), .B(new_n29446_), .ZN(new_n29665_));
  NOR3_X1    g26411(.A1(new_n29632_), .A2(new_n29374_), .A3(new_n29665_), .ZN(new_n29666_));
  NAND3_X1   g26412(.A1(new_n29655_), .A2(new_n29661_), .A3(new_n29666_), .ZN(new_n29667_));
  AOI21_X1   g26413(.A1(new_n29652_), .A2(new_n29653_), .B(new_n29667_), .ZN(new_n29668_));
  OAI21_X1   g26414(.A1(new_n29623_), .A2(new_n29648_), .B(new_n29668_), .ZN(new_n29669_));
  XNOR2_X1   g26415(.A1(new_n29669_), .A2(new_n29583_), .ZN(new_n29670_));
  NAND2_X1   g26416(.A1(new_n29457_), .A2(pi0625), .ZN(new_n29671_));
  XOR2_X1    g26417(.A1(new_n29671_), .A2(new_n13615_), .Z(new_n29672_));
  NOR2_X1    g26418(.A1(new_n29672_), .A2(new_n29670_), .ZN(new_n29673_));
  NAND2_X1   g26419(.A1(new_n29565_), .A2(new_n29345_), .ZN(new_n29674_));
  NAND2_X1   g26420(.A1(new_n29674_), .A2(new_n14081_), .ZN(new_n29675_));
  NOR2_X1    g26421(.A1(new_n29673_), .A2(new_n29675_), .ZN(new_n29676_));
  NAND2_X1   g26422(.A1(new_n29457_), .A2(pi1153), .ZN(new_n29677_));
  XOR2_X1    g26423(.A1(new_n29677_), .A2(new_n13615_), .Z(new_n29678_));
  OAI21_X1   g26424(.A1(new_n29678_), .A2(new_n29670_), .B(new_n14081_), .ZN(new_n29679_));
  NOR2_X1    g26425(.A1(new_n29562_), .A2(new_n13748_), .ZN(new_n29680_));
  OAI21_X1   g26426(.A1(new_n29676_), .A2(new_n29679_), .B(new_n29680_), .ZN(new_n29681_));
  NAND2_X1   g26427(.A1(new_n29670_), .A2(new_n13748_), .ZN(new_n29682_));
  NAND2_X1   g26428(.A1(new_n29681_), .A2(new_n29682_), .ZN(new_n29683_));
  NAND3_X1   g26429(.A1(new_n29683_), .A2(pi0609), .A3(pi1155), .ZN(new_n29684_));
  NAND4_X1   g26430(.A1(new_n29681_), .A2(pi0609), .A3(new_n13778_), .A4(new_n29682_), .ZN(new_n29685_));
  AOI21_X1   g26431(.A1(new_n29684_), .A2(new_n29685_), .B(new_n29567_), .ZN(new_n29686_));
  NOR2_X1    g26432(.A1(new_n29465_), .A2(pi0660), .ZN(new_n29687_));
  INV_X1     g26433(.I(new_n29687_), .ZN(new_n29688_));
  NOR2_X1    g26434(.A1(new_n29462_), .A2(pi0660), .ZN(new_n29689_));
  OAI21_X1   g26435(.A1(new_n29686_), .A2(new_n29688_), .B(new_n29689_), .ZN(new_n29690_));
  INV_X1     g26436(.I(new_n29567_), .ZN(new_n29691_));
  NOR2_X1    g26437(.A1(new_n29683_), .A2(new_n13778_), .ZN(new_n29692_));
  XOR2_X1    g26438(.A1(new_n29692_), .A2(new_n14090_), .Z(new_n29693_));
  AND3_X2    g26439(.A1(new_n29693_), .A2(pi0785), .A3(new_n29691_), .Z(new_n29694_));
  AOI22_X1   g26440(.A1(new_n29694_), .A2(new_n29690_), .B1(new_n13801_), .B2(new_n29683_), .ZN(new_n29695_));
  AOI21_X1   g26441(.A1(new_n29568_), .A2(new_n13816_), .B(new_n14501_), .ZN(new_n29696_));
  AOI21_X1   g26442(.A1(new_n29489_), .A2(new_n29696_), .B(pi0618), .ZN(new_n29697_));
  AOI21_X1   g26443(.A1(new_n29493_), .A2(new_n13836_), .B(pi0618), .ZN(new_n29698_));
  NOR4_X1    g26444(.A1(new_n29695_), .A2(new_n13855_), .A3(new_n29697_), .A4(new_n29698_), .ZN(new_n29699_));
  OAI21_X1   g26445(.A1(new_n29695_), .A2(new_n29697_), .B(pi0781), .ZN(new_n29700_));
  NOR3_X1    g26446(.A1(new_n29695_), .A2(new_n13855_), .A3(new_n29698_), .ZN(new_n29701_));
  NOR2_X1    g26447(.A1(new_n29701_), .A2(new_n29700_), .ZN(new_n29702_));
  NOR2_X1    g26448(.A1(new_n29702_), .A2(new_n29699_), .ZN(new_n29703_));
  AOI21_X1   g26449(.A1(new_n29703_), .A2(pi1159), .B(new_n13904_), .ZN(new_n29704_));
  NOR4_X1    g26450(.A1(new_n29702_), .A2(pi0619), .A3(new_n13868_), .A4(new_n29699_), .ZN(new_n29705_));
  OAI21_X1   g26451(.A1(new_n29704_), .A2(new_n29705_), .B(new_n29570_), .ZN(new_n29706_));
  AOI21_X1   g26452(.A1(new_n29706_), .A2(new_n16474_), .B(new_n29503_), .ZN(new_n29707_));
  INV_X1     g26453(.I(new_n29707_), .ZN(new_n29708_));
  NAND3_X1   g26454(.A1(new_n29501_), .A2(pi0619), .A3(pi1159), .ZN(new_n29709_));
  NAND3_X1   g26455(.A1(new_n29496_), .A2(pi0619), .A3(new_n13904_), .ZN(new_n29710_));
  AOI21_X1   g26456(.A1(new_n29710_), .A2(new_n29709_), .B(new_n29346_), .ZN(new_n29711_));
  NAND3_X1   g26457(.A1(new_n29501_), .A2(pi0619), .A3(pi1159), .ZN(new_n29712_));
  NAND4_X1   g26458(.A1(new_n29500_), .A2(new_n13860_), .A3(pi1159), .A4(new_n29485_), .ZN(new_n29713_));
  AOI21_X1   g26459(.A1(new_n29712_), .A2(new_n29713_), .B(new_n29346_), .ZN(new_n29714_));
  NAND4_X1   g26460(.A1(new_n29711_), .A2(new_n29714_), .A3(pi0789), .A4(new_n29501_), .ZN(new_n29715_));
  NOR2_X1    g26461(.A1(new_n29496_), .A2(new_n13896_), .ZN(new_n29716_));
  NAND2_X1   g26462(.A1(new_n29714_), .A2(new_n29716_), .ZN(new_n29717_));
  NAND3_X1   g26463(.A1(new_n29717_), .A2(pi0789), .A3(new_n29503_), .ZN(new_n29718_));
  NAND3_X1   g26464(.A1(new_n29718_), .A2(new_n13962_), .A3(new_n29715_), .ZN(new_n29719_));
  NAND2_X1   g26465(.A1(new_n29719_), .A2(new_n18975_), .ZN(new_n29720_));
  AOI21_X1   g26466(.A1(pi0789), .A2(new_n29503_), .B(new_n29717_), .ZN(new_n29721_));
  NAND2_X1   g26467(.A1(new_n29503_), .A2(pi0789), .ZN(new_n29722_));
  AOI21_X1   g26468(.A1(new_n29496_), .A2(pi1159), .B(new_n13904_), .ZN(new_n29723_));
  INV_X1     g26469(.I(new_n29713_), .ZN(new_n29724_));
  OAI21_X1   g26470(.A1(new_n29723_), .A2(new_n29724_), .B(new_n29345_), .ZN(new_n29725_));
  NOR3_X1    g26471(.A1(new_n29725_), .A2(new_n13896_), .A3(new_n29496_), .ZN(new_n29726_));
  NOR2_X1    g26472(.A1(new_n29726_), .A2(new_n29722_), .ZN(new_n29727_));
  NOR2_X1    g26473(.A1(new_n29727_), .A2(new_n29721_), .ZN(new_n29728_));
  NAND3_X1   g26474(.A1(new_n29728_), .A2(new_n13901_), .A3(new_n13962_), .ZN(new_n29729_));
  AOI21_X1   g26475(.A1(new_n29729_), .A2(new_n29720_), .B(new_n29346_), .ZN(new_n29730_));
  NAND2_X1   g26476(.A1(new_n29569_), .A2(new_n16639_), .ZN(new_n29731_));
  XOR2_X1    g26477(.A1(new_n29731_), .A2(new_n16829_), .Z(new_n29732_));
  AOI21_X1   g26478(.A1(new_n29732_), .A2(new_n29345_), .B(pi0788), .ZN(new_n29733_));
  INV_X1     g26479(.I(new_n29733_), .ZN(new_n29734_));
  NAND2_X1   g26480(.A1(new_n29718_), .A2(new_n29715_), .ZN(new_n29735_));
  NAND3_X1   g26481(.A1(new_n29735_), .A2(pi0626), .A3(new_n13963_), .ZN(new_n29736_));
  NAND3_X1   g26482(.A1(new_n29728_), .A2(new_n13901_), .A3(new_n13963_), .ZN(new_n29737_));
  NOR2_X1    g26483(.A1(new_n29346_), .A2(new_n15479_), .ZN(new_n29738_));
  OAI21_X1   g26484(.A1(new_n29703_), .A2(pi0789), .B(new_n29738_), .ZN(new_n29739_));
  AOI21_X1   g26485(.A1(new_n29737_), .A2(new_n29736_), .B(new_n29739_), .ZN(new_n29740_));
  OAI21_X1   g26486(.A1(new_n29730_), .A2(new_n29734_), .B(new_n29740_), .ZN(new_n29741_));
  AOI21_X1   g26487(.A1(new_n29703_), .A2(pi0619), .B(new_n13904_), .ZN(new_n29742_));
  NOR4_X1    g26488(.A1(new_n29702_), .A2(new_n13860_), .A3(pi1159), .A4(new_n29699_), .ZN(new_n29743_));
  OAI21_X1   g26489(.A1(new_n29742_), .A2(new_n29743_), .B(new_n29570_), .ZN(new_n29744_));
  NAND3_X1   g26490(.A1(new_n29744_), .A2(new_n13884_), .A3(new_n29725_), .ZN(new_n29745_));
  AOI21_X1   g26491(.A1(new_n29708_), .A2(new_n29741_), .B(new_n29745_), .ZN(new_n29746_));
  NOR2_X1    g26492(.A1(new_n29346_), .A2(new_n16372_), .ZN(new_n29747_));
  AOI21_X1   g26493(.A1(new_n29728_), .A2(new_n16372_), .B(new_n29747_), .ZN(new_n29748_));
  AOI21_X1   g26494(.A1(new_n29346_), .A2(pi0628), .B(new_n19484_), .ZN(new_n29749_));
  INV_X1     g26495(.I(new_n29749_), .ZN(new_n29750_));
  NAND3_X1   g26496(.A1(new_n29570_), .A2(new_n15395_), .A3(new_n29345_), .ZN(new_n29751_));
  NAND3_X1   g26497(.A1(new_n29569_), .A2(new_n15395_), .A3(new_n29346_), .ZN(new_n29752_));
  NAND2_X1   g26498(.A1(new_n29751_), .A2(new_n29752_), .ZN(new_n29753_));
  NAND2_X1   g26499(.A1(new_n29345_), .A2(new_n29298_), .ZN(new_n29754_));
  OAI22_X1   g26500(.A1(new_n29753_), .A2(new_n13942_), .B1(new_n29750_), .B2(new_n29754_), .ZN(new_n29755_));
  OAI21_X1   g26501(.A1(new_n29748_), .A2(new_n16874_), .B(new_n29755_), .ZN(new_n29756_));
  NOR2_X1    g26502(.A1(new_n29345_), .A2(new_n13994_), .ZN(new_n29757_));
  INV_X1     g26503(.I(new_n29757_), .ZN(new_n29758_));
  INV_X1     g26504(.I(new_n29747_), .ZN(new_n29759_));
  NAND3_X1   g26505(.A1(new_n29718_), .A2(new_n16372_), .A3(new_n29715_), .ZN(new_n29760_));
  NAND3_X1   g26506(.A1(new_n29760_), .A2(new_n13994_), .A3(new_n29759_), .ZN(new_n29761_));
  OAI21_X1   g26507(.A1(new_n29753_), .A2(new_n29345_), .B(new_n14058_), .ZN(new_n29762_));
  AOI21_X1   g26508(.A1(new_n29762_), .A2(pi0647), .B(new_n14008_), .ZN(new_n29763_));
  INV_X1     g26509(.I(new_n29762_), .ZN(new_n29764_));
  NOR3_X1    g26510(.A1(new_n29764_), .A2(new_n14005_), .A3(new_n14007_), .ZN(new_n29765_));
  OAI21_X1   g26511(.A1(new_n29765_), .A2(new_n29763_), .B(new_n29345_), .ZN(new_n29766_));
  NAND2_X1   g26512(.A1(new_n29766_), .A2(pi0630), .ZN(new_n29767_));
  AOI21_X1   g26513(.A1(new_n29762_), .A2(pi1157), .B(new_n14008_), .ZN(new_n29768_));
  NOR3_X1    g26514(.A1(new_n29764_), .A2(new_n14006_), .A3(new_n14007_), .ZN(new_n29769_));
  OAI21_X1   g26515(.A1(new_n29769_), .A2(new_n29768_), .B(new_n29345_), .ZN(new_n29770_));
  NAND2_X1   g26516(.A1(new_n29770_), .A2(new_n14010_), .ZN(new_n29771_));
  AOI21_X1   g26517(.A1(new_n29767_), .A2(new_n29771_), .B(new_n12776_), .ZN(new_n29772_));
  OAI21_X1   g26518(.A1(new_n29772_), .A2(new_n16576_), .B(new_n16419_), .ZN(new_n29773_));
  AOI21_X1   g26519(.A1(new_n29761_), .A2(new_n29758_), .B(new_n29773_), .ZN(new_n29774_));
  OAI21_X1   g26520(.A1(new_n29756_), .A2(new_n16424_), .B(new_n29774_), .ZN(new_n29775_));
  INV_X1     g26521(.I(new_n29775_), .ZN(new_n29776_));
  AND2_X2    g26522(.A1(new_n29756_), .A2(pi0792), .Z(new_n29777_));
  OAI21_X1   g26523(.A1(new_n29746_), .A2(new_n29776_), .B(new_n29777_), .ZN(new_n29778_));
  NOR2_X1    g26524(.A1(new_n29346_), .A2(new_n14211_), .ZN(new_n29779_));
  INV_X1     g26525(.I(new_n29779_), .ZN(new_n29780_));
  NAND3_X1   g26526(.A1(new_n29761_), .A2(new_n14211_), .A3(new_n29758_), .ZN(new_n29781_));
  NAND3_X1   g26527(.A1(new_n29781_), .A2(pi0715), .A3(new_n29780_), .ZN(new_n29782_));
  XOR2_X1    g26528(.A1(new_n29782_), .A2(new_n14205_), .Z(new_n29783_));
  AND2_X2    g26529(.A1(new_n29766_), .A2(pi0787), .Z(new_n29784_));
  NOR3_X1    g26530(.A1(new_n29770_), .A2(new_n12776_), .A3(new_n29762_), .ZN(new_n29785_));
  XOR2_X1    g26531(.A1(new_n29784_), .A2(new_n29785_), .Z(new_n29786_));
  AOI21_X1   g26532(.A1(new_n29786_), .A2(pi0644), .B(new_n15386_), .ZN(new_n29787_));
  OAI21_X1   g26533(.A1(new_n29783_), .A2(new_n29346_), .B(new_n29787_), .ZN(new_n29788_));
  AOI21_X1   g26534(.A1(new_n29748_), .A2(new_n13994_), .B(new_n29757_), .ZN(new_n29790_));
  AOI21_X1   g26535(.A1(new_n29790_), .A2(new_n14211_), .B(new_n29779_), .ZN(new_n29791_));
  AOI21_X1   g26536(.A1(new_n29791_), .A2(pi0644), .B(new_n14217_), .ZN(new_n29792_));
  AND4_X2    g26537(.A1(pi0644), .A2(new_n29781_), .A3(new_n14200_), .A4(new_n29780_), .Z(new_n29793_));
  OAI21_X1   g26538(.A1(new_n29792_), .A2(new_n29793_), .B(new_n29345_), .ZN(new_n29794_));
  AOI21_X1   g26539(.A1(new_n29786_), .A2(new_n14204_), .B(new_n19370_), .ZN(new_n29795_));
  NOR3_X1    g26540(.A1(new_n29778_), .A2(new_n14204_), .A3(new_n12775_), .ZN(new_n29797_));
  AOI21_X1   g26541(.A1(new_n29788_), .A2(new_n29778_), .B(new_n14204_), .ZN(new_n29798_));
  AOI21_X1   g26542(.A1(new_n29794_), .A2(new_n29795_), .B(pi0644), .ZN(new_n29799_));
  XOR2_X1    g26543(.A1(new_n29719_), .A2(new_n18975_), .Z(new_n29800_));
  OAI21_X1   g26544(.A1(new_n29800_), .A2(new_n29346_), .B(new_n29733_), .ZN(new_n29801_));
  AOI21_X1   g26545(.A1(new_n29801_), .A2(new_n29740_), .B(new_n29707_), .ZN(new_n29802_));
  OAI21_X1   g26546(.A1(new_n29802_), .A2(new_n29745_), .B(new_n29775_), .ZN(new_n29803_));
  NAND3_X1   g26547(.A1(new_n29803_), .A2(pi0790), .A3(new_n29777_), .ZN(new_n29804_));
  NOR2_X1    g26548(.A1(new_n29799_), .A2(new_n29804_), .ZN(new_n29805_));
  NOR3_X1    g26549(.A1(new_n29805_), .A2(new_n29798_), .A3(new_n12775_), .ZN(new_n29806_));
  OAI21_X1   g26550(.A1(new_n29806_), .A2(new_n29797_), .B(new_n7240_), .ZN(new_n29807_));
  NAND2_X1   g26551(.A1(po1038), .A2(pi0223), .ZN(new_n29808_));
  NAND2_X1   g26552(.A1(new_n29807_), .A2(new_n29808_), .ZN(po0380));
  OR2_X2     g26553(.A1(new_n28787_), .A2(new_n14300_), .Z(new_n29810_));
  NAND2_X1   g26554(.A1(new_n29810_), .A2(pi0224), .ZN(new_n29811_));
  AOI21_X1   g26555(.A1(new_n13109_), .A2(pi0224), .B(new_n3259_), .ZN(new_n29812_));
  INV_X1     g26556(.I(new_n29812_), .ZN(new_n29813_));
  AOI21_X1   g26557(.A1(pi0614), .A2(new_n13106_), .B(new_n29813_), .ZN(new_n29814_));
  NOR2_X1    g26558(.A1(new_n29814_), .A2(new_n3290_), .ZN(new_n29815_));
  INV_X1     g26559(.I(new_n29815_), .ZN(new_n29816_));
  NOR2_X1    g26560(.A1(new_n13263_), .A2(new_n12868_), .ZN(new_n29817_));
  NAND2_X1   g26561(.A1(new_n28799_), .A2(pi0614), .ZN(new_n29818_));
  XOR2_X1    g26562(.A1(new_n29818_), .A2(new_n29817_), .Z(new_n29819_));
  NAND2_X1   g26563(.A1(new_n13261_), .A2(new_n5381_), .ZN(new_n29820_));
  OAI21_X1   g26564(.A1(new_n29819_), .A2(new_n29820_), .B(new_n12951_), .ZN(new_n29821_));
  NAND2_X1   g26565(.A1(new_n29821_), .A2(new_n5373_), .ZN(new_n29822_));
  NOR2_X1    g26566(.A1(new_n13103_), .A2(new_n12868_), .ZN(new_n29823_));
  INV_X1     g26567(.I(new_n29823_), .ZN(new_n29824_));
  NOR2_X1    g26568(.A1(new_n12818_), .A2(new_n29824_), .ZN(new_n29825_));
  AOI21_X1   g26569(.A1(new_n13541_), .A2(pi0614), .B(new_n5375_), .ZN(new_n29826_));
  AOI21_X1   g26570(.A1(new_n29825_), .A2(new_n12844_), .B(pi0680), .ZN(new_n29827_));
  NOR2_X1    g26571(.A1(new_n29822_), .A2(new_n29827_), .ZN(new_n29828_));
  AOI21_X1   g26572(.A1(new_n12845_), .A2(new_n29822_), .B(new_n29828_), .ZN(new_n29829_));
  NAND2_X1   g26573(.A1(new_n29824_), .A2(pi0680), .ZN(new_n29830_));
  AOI21_X1   g26574(.A1(new_n12784_), .A2(new_n29824_), .B(new_n5383_), .ZN(new_n29831_));
  AOI21_X1   g26575(.A1(new_n28715_), .A2(new_n12841_), .B(new_n29831_), .ZN(new_n29832_));
  NAND3_X1   g26576(.A1(new_n29832_), .A2(pi0680), .A3(new_n12949_), .ZN(new_n29833_));
  XOR2_X1    g26577(.A1(new_n29833_), .A2(new_n29830_), .Z(new_n29834_));
  NAND2_X1   g26578(.A1(new_n29834_), .A2(new_n12844_), .ZN(new_n29835_));
  AOI21_X1   g26579(.A1(new_n29832_), .A2(new_n12845_), .B(new_n3100_), .ZN(new_n29836_));
  NAND2_X1   g26580(.A1(new_n29835_), .A2(new_n29836_), .ZN(new_n29837_));
  NOR2_X1    g26581(.A1(new_n5455_), .A2(new_n3100_), .ZN(new_n29838_));
  NAND2_X1   g26582(.A1(new_n29837_), .A2(new_n29838_), .ZN(new_n29839_));
  INV_X1     g26583(.I(new_n29838_), .ZN(new_n29840_));
  NAND3_X1   g26584(.A1(new_n29835_), .A2(new_n29836_), .A3(new_n29840_), .ZN(new_n29841_));
  NAND2_X1   g26585(.A1(new_n29839_), .A2(new_n29841_), .ZN(new_n29842_));
  AND2_X2    g26586(.A1(new_n29842_), .A2(new_n29829_), .Z(new_n29843_));
  NOR2_X1    g26587(.A1(new_n13364_), .A2(new_n12868_), .ZN(new_n29844_));
  NOR2_X1    g26588(.A1(new_n12784_), .A2(new_n3100_), .ZN(new_n29845_));
  NOR2_X1    g26589(.A1(new_n3312_), .A2(new_n3111_), .ZN(new_n29846_));
  INV_X1     g26590(.I(new_n29846_), .ZN(new_n29847_));
  NOR3_X1    g26591(.A1(new_n13368_), .A2(new_n12868_), .A3(new_n5636_), .ZN(new_n29848_));
  NOR3_X1    g26592(.A1(new_n13372_), .A2(new_n12868_), .A3(new_n5378_), .ZN(new_n29849_));
  OAI21_X1   g26593(.A1(new_n29848_), .A2(new_n29849_), .B(new_n13363_), .ZN(new_n29850_));
  NOR2_X1    g26594(.A1(new_n13263_), .A2(new_n29824_), .ZN(new_n29851_));
  NOR2_X1    g26595(.A1(new_n29851_), .A2(pi0680), .ZN(new_n29852_));
  OAI21_X1   g26596(.A1(new_n29852_), .A2(new_n29826_), .B(new_n12844_), .ZN(new_n29853_));
  OAI21_X1   g26597(.A1(new_n12844_), .A2(new_n29851_), .B(new_n29853_), .ZN(new_n29854_));
  NAND2_X1   g26598(.A1(new_n29854_), .A2(new_n5454_), .ZN(new_n29855_));
  XOR2_X1    g26599(.A1(new_n29855_), .A2(new_n29838_), .Z(new_n29856_));
  NOR2_X1    g26600(.A1(new_n29856_), .A2(new_n29850_), .ZN(new_n29857_));
  OAI21_X1   g26601(.A1(new_n29843_), .A2(new_n29847_), .B(new_n29857_), .ZN(new_n29858_));
  NAND2_X1   g26602(.A1(new_n29858_), .A2(new_n3098_), .ZN(new_n29859_));
  NOR2_X1    g26603(.A1(new_n12903_), .A2(new_n29831_), .ZN(new_n29860_));
  NAND3_X1   g26604(.A1(new_n29860_), .A2(pi0680), .A3(new_n13334_), .ZN(new_n29861_));
  XOR2_X1    g26605(.A1(new_n29861_), .A2(new_n29830_), .Z(new_n29862_));
  NAND2_X1   g26606(.A1(new_n29862_), .A2(new_n12844_), .ZN(new_n29863_));
  AOI21_X1   g26607(.A1(new_n29860_), .A2(new_n12845_), .B(new_n3100_), .ZN(new_n29864_));
  NAND2_X1   g26608(.A1(new_n29863_), .A2(new_n29864_), .ZN(new_n29865_));
  XOR2_X1    g26609(.A1(new_n29865_), .A2(new_n29840_), .Z(new_n29866_));
  AOI21_X1   g26610(.A1(pi0614), .A2(new_n14302_), .B(new_n28617_), .ZN(new_n29867_));
  INV_X1     g26611(.I(new_n29867_), .ZN(new_n29868_));
  AOI21_X1   g26612(.A1(new_n12878_), .A2(pi0680), .B(pi0614), .ZN(new_n29869_));
  INV_X1     g26613(.I(new_n29869_), .ZN(new_n29870_));
  NOR2_X1    g26614(.A1(new_n14304_), .A2(new_n12845_), .ZN(new_n29871_));
  AOI21_X1   g26615(.A1(new_n29870_), .A2(new_n29871_), .B(pi0680), .ZN(new_n29872_));
  NOR2_X1    g26616(.A1(new_n29868_), .A2(new_n29872_), .ZN(new_n29873_));
  INV_X1     g26617(.I(new_n29873_), .ZN(new_n29874_));
  OAI21_X1   g26618(.A1(new_n12844_), .A2(new_n29867_), .B(new_n29874_), .ZN(new_n29875_));
  AOI21_X1   g26619(.A1(new_n12868_), .A2(new_n13364_), .B(new_n28843_), .ZN(new_n29876_));
  NAND2_X1   g26620(.A1(new_n29876_), .A2(new_n3100_), .ZN(new_n29877_));
  NOR2_X1    g26621(.A1(new_n29875_), .A2(new_n29877_), .ZN(new_n29878_));
  AOI21_X1   g26622(.A1(new_n29866_), .A2(new_n29878_), .B(new_n12922_), .ZN(new_n29879_));
  XOR2_X1    g26623(.A1(new_n29865_), .A2(new_n28882_), .Z(new_n29880_));
  OAI21_X1   g26624(.A1(new_n29880_), .A2(new_n29875_), .B(new_n3090_), .ZN(new_n29881_));
  NAND4_X1   g26625(.A1(new_n3289_), .A2(pi0215), .A3(new_n5454_), .A4(pi0224), .ZN(new_n29882_));
  NOR3_X1    g26626(.A1(new_n29877_), .A2(new_n13701_), .A3(new_n29882_), .ZN(new_n29883_));
  NAND2_X1   g26627(.A1(new_n29881_), .A2(new_n29883_), .ZN(new_n29884_));
  OAI21_X1   g26628(.A1(new_n13173_), .A2(pi0614), .B(pi0224), .ZN(new_n29885_));
  NOR2_X1    g26629(.A1(new_n14973_), .A2(new_n29885_), .ZN(new_n29886_));
  NAND2_X1   g26630(.A1(new_n13174_), .A2(pi0614), .ZN(new_n29887_));
  OAI21_X1   g26631(.A1(new_n29887_), .A2(pi0224), .B(new_n3098_), .ZN(new_n29888_));
  OAI21_X1   g26632(.A1(new_n29888_), .A2(new_n29886_), .B(new_n3183_), .ZN(new_n29889_));
  AOI21_X1   g26633(.A1(new_n13192_), .A2(pi0614), .B(new_n3100_), .ZN(new_n29890_));
  AOI21_X1   g26634(.A1(pi0224), .A2(new_n14336_), .B(new_n14979_), .ZN(new_n29891_));
  NAND2_X1   g26635(.A1(new_n29890_), .A2(new_n29891_), .ZN(new_n29892_));
  NOR2_X1    g26636(.A1(new_n29892_), .A2(new_n3098_), .ZN(new_n29893_));
  AOI21_X1   g26637(.A1(new_n29889_), .A2(new_n29893_), .B(pi0038), .ZN(new_n29894_));
  XOR2_X1    g26638(.A1(new_n29837_), .A2(new_n28883_), .Z(new_n29895_));
  NAND2_X1   g26639(.A1(new_n29854_), .A2(new_n5138_), .ZN(new_n29896_));
  NOR2_X1    g26640(.A1(new_n5397_), .A2(new_n5139_), .ZN(new_n29897_));
  INV_X1     g26641(.I(new_n29897_), .ZN(new_n29898_));
  XOR2_X1    g26642(.A1(new_n29896_), .A2(new_n29898_), .Z(new_n29899_));
  NAND4_X1   g26643(.A1(new_n12987_), .A2(pi0223), .A3(pi0614), .A4(new_n13203_), .ZN(new_n29900_));
  NOR2_X1    g26644(.A1(new_n29850_), .A2(new_n29900_), .ZN(new_n29901_));
  AND3_X2    g26645(.A1(new_n29829_), .A2(new_n29899_), .A3(new_n29901_), .Z(new_n29902_));
  AOI21_X1   g26646(.A1(new_n29902_), .A2(new_n29895_), .B(new_n5827_), .ZN(new_n29903_));
  NOR4_X1    g26647(.A1(new_n29903_), .A2(new_n29879_), .A3(new_n29884_), .A4(new_n29894_), .ZN(new_n29904_));
  NAND3_X1   g26648(.A1(new_n29859_), .A2(new_n29816_), .A3(new_n29904_), .ZN(new_n29905_));
  INV_X1     g26649(.I(new_n29905_), .ZN(new_n29906_));
  AOI21_X1   g26650(.A1(new_n29859_), .A2(new_n29904_), .B(new_n29816_), .ZN(new_n29907_));
  OAI21_X1   g26651(.A1(new_n29906_), .A2(new_n29907_), .B(new_n13776_), .ZN(new_n29908_));
  NAND2_X1   g26652(.A1(new_n29811_), .A2(new_n13775_), .ZN(new_n29909_));
  NAND2_X1   g26653(.A1(new_n29908_), .A2(new_n29909_), .ZN(new_n29910_));
  NAND3_X1   g26654(.A1(new_n29910_), .A2(pi0609), .A3(pi1155), .ZN(new_n29911_));
  INV_X1     g26655(.I(new_n29907_), .ZN(new_n29912_));
  AOI21_X1   g26656(.A1(new_n29912_), .A2(new_n29905_), .B(new_n13775_), .ZN(new_n29913_));
  INV_X1     g26657(.I(new_n29909_), .ZN(new_n29914_));
  NOR3_X1    g26658(.A1(new_n29913_), .A2(new_n13766_), .A3(new_n29914_), .ZN(new_n29915_));
  NAND2_X1   g26659(.A1(new_n29915_), .A2(new_n14694_), .ZN(new_n29916_));
  AOI21_X1   g26660(.A1(new_n29916_), .A2(new_n29911_), .B(new_n29811_), .ZN(new_n29917_));
  NAND3_X1   g26661(.A1(new_n29910_), .A2(pi0609), .A3(pi1155), .ZN(new_n29918_));
  NAND4_X1   g26662(.A1(new_n29908_), .A2(new_n13766_), .A3(pi1155), .A4(new_n29909_), .ZN(new_n29919_));
  AOI21_X1   g26663(.A1(new_n29918_), .A2(new_n29919_), .B(new_n29811_), .ZN(new_n29920_));
  NAND4_X1   g26664(.A1(new_n29917_), .A2(new_n29920_), .A3(pi0785), .A4(new_n29910_), .ZN(new_n29921_));
  INV_X1     g26665(.I(new_n29811_), .ZN(new_n29922_));
  NOR2_X1    g26666(.A1(new_n29915_), .A2(new_n14694_), .ZN(new_n29923_));
  NOR3_X1    g26667(.A1(new_n29910_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n29924_));
  OAI21_X1   g26668(.A1(new_n29923_), .A2(new_n29924_), .B(new_n29922_), .ZN(new_n29925_));
  INV_X1     g26669(.I(new_n29910_), .ZN(new_n29926_));
  NOR2_X1    g26670(.A1(new_n29926_), .A2(new_n13801_), .ZN(new_n29927_));
  NAND2_X1   g26671(.A1(new_n29920_), .A2(new_n29927_), .ZN(new_n29928_));
  NAND3_X1   g26672(.A1(new_n29928_), .A2(pi0785), .A3(new_n29925_), .ZN(new_n29929_));
  NAND2_X1   g26673(.A1(new_n29929_), .A2(new_n29921_), .ZN(new_n29930_));
  NAND3_X1   g26674(.A1(new_n29930_), .A2(pi0618), .A3(pi1154), .ZN(new_n29931_));
  NOR2_X1    g26675(.A1(new_n29917_), .A2(new_n13801_), .ZN(new_n29932_));
  XOR2_X1    g26676(.A1(new_n29932_), .A2(new_n29928_), .Z(new_n29933_));
  NAND3_X1   g26677(.A1(new_n29933_), .A2(pi0618), .A3(new_n13817_), .ZN(new_n29934_));
  AOI21_X1   g26678(.A1(new_n29934_), .A2(new_n29931_), .B(new_n29811_), .ZN(new_n29935_));
  NAND3_X1   g26679(.A1(new_n29930_), .A2(pi0618), .A3(pi1154), .ZN(new_n29936_));
  NAND4_X1   g26680(.A1(new_n29929_), .A2(new_n13816_), .A3(pi1154), .A4(new_n29921_), .ZN(new_n29937_));
  AOI21_X1   g26681(.A1(new_n29936_), .A2(new_n29937_), .B(new_n29811_), .ZN(new_n29938_));
  NAND4_X1   g26682(.A1(new_n29935_), .A2(pi0781), .A3(new_n29938_), .A4(new_n29930_), .ZN(new_n29939_));
  AOI21_X1   g26683(.A1(new_n29933_), .A2(pi0618), .B(new_n13819_), .ZN(new_n29940_));
  NOR3_X1    g26684(.A1(new_n29930_), .A2(new_n13816_), .A3(pi1154), .ZN(new_n29941_));
  OAI21_X1   g26685(.A1(new_n29940_), .A2(new_n29941_), .B(new_n29922_), .ZN(new_n29942_));
  NAND3_X1   g26686(.A1(new_n29938_), .A2(pi0781), .A3(new_n29930_), .ZN(new_n29943_));
  NAND3_X1   g26687(.A1(new_n29943_), .A2(pi0781), .A3(new_n29942_), .ZN(new_n29944_));
  NAND2_X1   g26688(.A1(new_n29944_), .A2(new_n29939_), .ZN(new_n29945_));
  NAND3_X1   g26689(.A1(new_n29945_), .A2(pi0619), .A3(pi1159), .ZN(new_n29946_));
  NAND4_X1   g26690(.A1(new_n29944_), .A2(pi0619), .A3(new_n29939_), .A4(new_n13868_), .ZN(new_n29947_));
  AOI21_X1   g26691(.A1(new_n29946_), .A2(new_n29947_), .B(new_n29811_), .ZN(new_n29948_));
  NOR2_X1    g26692(.A1(new_n29010_), .A2(new_n5633_), .ZN(new_n29949_));
  OAI21_X1   g26693(.A1(new_n29813_), .A2(new_n29949_), .B(new_n3289_), .ZN(new_n29950_));
  NOR2_X1    g26694(.A1(new_n3100_), .A2(new_n3098_), .ZN(new_n29951_));
  NAND2_X1   g26695(.A1(new_n13141_), .A2(pi0299), .ZN(new_n29952_));
  XNOR2_X1   g26696(.A1(new_n29952_), .A2(new_n29951_), .ZN(new_n29953_));
  NOR2_X1    g26697(.A1(new_n13155_), .A2(new_n3183_), .ZN(new_n29954_));
  AOI21_X1   g26698(.A1(new_n29953_), .A2(new_n29954_), .B(new_n29001_), .ZN(new_n29955_));
  NOR2_X1    g26699(.A1(new_n28963_), .A2(new_n5633_), .ZN(new_n29956_));
  NAND2_X1   g26700(.A1(new_n13691_), .A2(new_n28952_), .ZN(new_n29957_));
  NAND2_X1   g26701(.A1(new_n13695_), .A2(pi0662), .ZN(new_n29958_));
  NAND2_X1   g26702(.A1(new_n29958_), .A2(new_n6459_), .ZN(new_n29959_));
  AOI21_X1   g26703(.A1(new_n29957_), .A2(new_n5398_), .B(new_n29959_), .ZN(new_n29960_));
  OAI21_X1   g26704(.A1(new_n29960_), .A2(new_n5398_), .B(new_n29956_), .ZN(new_n29961_));
  NAND2_X1   g26705(.A1(new_n12911_), .A2(new_n5633_), .ZN(new_n29962_));
  OAI21_X1   g26706(.A1(new_n5633_), .A2(new_n28976_), .B(new_n29962_), .ZN(new_n29963_));
  AOI21_X1   g26707(.A1(new_n28981_), .A2(pi0662), .B(new_n3100_), .ZN(new_n29964_));
  OAI21_X1   g26708(.A1(pi0662), .A2(new_n12935_), .B(new_n29964_), .ZN(new_n29965_));
  XOR2_X1    g26709(.A1(new_n29965_), .A2(new_n28883_), .Z(new_n29966_));
  NAND3_X1   g26710(.A1(new_n13702_), .A2(new_n3090_), .A3(new_n5633_), .ZN(new_n29967_));
  NAND2_X1   g26711(.A1(new_n29967_), .A2(pi0224), .ZN(new_n29968_));
  AOI21_X1   g26712(.A1(new_n29966_), .A2(new_n29963_), .B(new_n29968_), .ZN(new_n29969_));
  NAND2_X1   g26713(.A1(new_n3098_), .A2(pi0039), .ZN(new_n29970_));
  OAI21_X1   g26714(.A1(new_n29969_), .A2(new_n29970_), .B(new_n29961_), .ZN(new_n29971_));
  XOR2_X1    g26715(.A1(new_n29965_), .A2(new_n29840_), .Z(new_n29972_));
  AOI21_X1   g26716(.A1(new_n29972_), .A2(new_n29963_), .B(new_n29585_), .ZN(new_n29973_));
  AOI21_X1   g26717(.A1(new_n28949_), .A2(pi0662), .B(new_n3100_), .ZN(new_n29974_));
  OAI21_X1   g26718(.A1(pi0662), .A2(new_n12980_), .B(new_n29974_), .ZN(new_n29975_));
  XOR2_X1    g26719(.A1(new_n29975_), .A2(new_n28883_), .Z(new_n29976_));
  AOI21_X1   g26720(.A1(new_n5634_), .A2(new_n28945_), .B(new_n13086_), .ZN(new_n29977_));
  NOR2_X1    g26721(.A1(new_n5633_), .A2(pi0224), .ZN(new_n29978_));
  NAND4_X1   g26722(.A1(new_n29976_), .A2(new_n13712_), .A3(new_n29977_), .A4(new_n29978_), .ZN(new_n29979_));
  NOR2_X1    g26723(.A1(new_n29979_), .A2(new_n29973_), .ZN(new_n29980_));
  AOI21_X1   g26724(.A1(new_n29980_), .A2(new_n29971_), .B(pi0215), .ZN(new_n29981_));
  INV_X1     g26725(.I(new_n29977_), .ZN(new_n29982_));
  XOR2_X1    g26726(.A1(new_n29975_), .A2(new_n29838_), .Z(new_n29983_));
  NOR2_X1    g26727(.A1(new_n29983_), .A2(new_n29982_), .ZN(new_n29984_));
  NOR2_X1    g26728(.A1(pi0216), .A2(pi0221), .ZN(new_n29985_));
  NAND2_X1   g26729(.A1(new_n29957_), .A2(new_n5454_), .ZN(new_n29986_));
  XOR2_X1    g26730(.A1(new_n29986_), .A2(new_n29838_), .Z(new_n29987_));
  NOR4_X1    g26731(.A1(new_n29987_), .A2(new_n3259_), .A3(new_n5633_), .A4(new_n28963_), .ZN(new_n29988_));
  OAI21_X1   g26732(.A1(new_n29984_), .A2(new_n29985_), .B(new_n29988_), .ZN(new_n29989_));
  OAI22_X1   g26733(.A1(new_n29981_), .A2(new_n29989_), .B1(new_n28953_), .B2(new_n29955_), .ZN(new_n29990_));
  OAI21_X1   g26734(.A1(new_n13159_), .A2(new_n3100_), .B(new_n3098_), .ZN(new_n29991_));
  NOR3_X1    g26735(.A1(new_n15066_), .A2(new_n28953_), .A3(new_n29991_), .ZN(new_n29992_));
  NOR3_X1    g26736(.A1(new_n29991_), .A2(new_n13134_), .A3(new_n28952_), .ZN(new_n29993_));
  NOR2_X1    g26737(.A1(new_n29992_), .A2(new_n29993_), .ZN(new_n29994_));
  NOR3_X1    g26738(.A1(new_n29994_), .A2(new_n3100_), .A3(new_n3290_), .ZN(new_n29995_));
  NAND2_X1   g26739(.A1(new_n29990_), .A2(new_n29995_), .ZN(new_n29996_));
  XOR2_X1    g26740(.A1(new_n29996_), .A2(new_n29950_), .Z(new_n29997_));
  NOR2_X1    g26741(.A1(new_n29997_), .A2(new_n13613_), .ZN(new_n29998_));
  XOR2_X1    g26742(.A1(new_n29998_), .A2(new_n13615_), .Z(new_n29999_));
  NAND2_X1   g26743(.A1(new_n29999_), .A2(new_n29922_), .ZN(new_n30000_));
  NAND2_X1   g26744(.A1(new_n30000_), .A2(pi0778), .ZN(new_n30001_));
  NOR2_X1    g26745(.A1(new_n29997_), .A2(new_n13614_), .ZN(new_n30002_));
  XOR2_X1    g26746(.A1(new_n30002_), .A2(new_n13615_), .Z(new_n30003_));
  NAND2_X1   g26747(.A1(new_n30003_), .A2(new_n29922_), .ZN(new_n30004_));
  NAND2_X1   g26748(.A1(new_n29997_), .A2(pi0778), .ZN(new_n30005_));
  NOR2_X1    g26749(.A1(new_n30004_), .A2(new_n30005_), .ZN(new_n30006_));
  XOR2_X1    g26750(.A1(new_n30006_), .A2(new_n30001_), .Z(new_n30007_));
  NOR2_X1    g26751(.A1(new_n29922_), .A2(new_n13805_), .ZN(new_n30008_));
  INV_X1     g26752(.I(new_n30008_), .ZN(new_n30009_));
  OAI21_X1   g26753(.A1(new_n30007_), .A2(new_n13803_), .B(new_n30009_), .ZN(new_n30010_));
  NOR2_X1    g26754(.A1(new_n29922_), .A2(new_n13880_), .ZN(new_n30011_));
  AOI21_X1   g26755(.A1(new_n30010_), .A2(new_n13880_), .B(new_n30011_), .ZN(new_n30012_));
  NOR3_X1    g26756(.A1(new_n29814_), .A2(pi0662), .A3(new_n13213_), .ZN(new_n30013_));
  OAI21_X1   g26757(.A1(new_n30013_), .A2(new_n13109_), .B(new_n3289_), .ZN(new_n30014_));
  AOI21_X1   g26758(.A1(new_n29096_), .A2(pi0680), .B(new_n29844_), .ZN(new_n30015_));
  NOR2_X1    g26759(.A1(new_n30015_), .A2(new_n5633_), .ZN(new_n30016_));
  AOI21_X1   g26760(.A1(new_n29078_), .A2(new_n12868_), .B(new_n13297_), .ZN(new_n30017_));
  NOR3_X1    g26761(.A1(new_n29850_), .A2(new_n28953_), .A3(new_n30017_), .ZN(new_n30018_));
  XNOR2_X1   g26762(.A1(new_n30016_), .A2(new_n30018_), .ZN(new_n30019_));
  NOR2_X1    g26763(.A1(new_n13351_), .A2(new_n5375_), .ZN(new_n30020_));
  NOR2_X1    g26764(.A1(new_n12868_), .A2(new_n5375_), .ZN(new_n30021_));
  XOR2_X1    g26765(.A1(new_n30020_), .A2(new_n30021_), .Z(new_n30022_));
  INV_X1     g26766(.I(new_n29852_), .ZN(new_n30023_));
  NAND2_X1   g26767(.A1(new_n12843_), .A2(new_n5633_), .ZN(new_n30024_));
  NAND3_X1   g26768(.A1(new_n29851_), .A2(pi0662), .A3(new_n30024_), .ZN(new_n30025_));
  AOI21_X1   g26769(.A1(new_n30023_), .A2(new_n30025_), .B(new_n13420_), .ZN(new_n30026_));
  NAND2_X1   g26770(.A1(new_n30022_), .A2(new_n30026_), .ZN(new_n30027_));
  NAND2_X1   g26771(.A1(new_n30027_), .A2(new_n5138_), .ZN(new_n30028_));
  XOR2_X1    g26772(.A1(new_n30028_), .A2(new_n29897_), .Z(new_n30029_));
  OAI21_X1   g26773(.A1(new_n30029_), .A2(new_n30019_), .B(new_n3090_), .ZN(new_n30030_));
  AOI21_X1   g26774(.A1(new_n29844_), .A2(pi0224), .B(new_n28952_), .ZN(new_n30031_));
  NOR2_X1    g26775(.A1(new_n30031_), .A2(new_n13297_), .ZN(new_n30032_));
  INV_X1     g26776(.I(new_n30032_), .ZN(new_n30033_));
  NOR2_X1    g26777(.A1(new_n30033_), .A2(new_n3099_), .ZN(new_n30034_));
  NOR4_X1    g26778(.A1(new_n30017_), .A2(new_n5633_), .A3(new_n5375_), .A4(new_n29844_), .ZN(new_n30035_));
  AOI22_X1   g26779(.A1(new_n13341_), .A2(new_n30035_), .B1(new_n5633_), .B2(new_n29876_), .ZN(new_n30036_));
  INV_X1     g26780(.I(new_n30036_), .ZN(new_n30037_));
  AND2_X2    g26781(.A1(new_n13559_), .A2(new_n13557_), .Z(new_n30038_));
  OAI21_X1   g26782(.A1(new_n30038_), .A2(new_n13494_), .B(pi0680), .ZN(new_n30039_));
  NOR3_X1    g26783(.A1(new_n14291_), .A2(pi0614), .A3(new_n13211_), .ZN(new_n30040_));
  AOI21_X1   g26784(.A1(pi0614), .A2(new_n29038_), .B(new_n30040_), .ZN(new_n30041_));
  NOR2_X1    g26785(.A1(new_n30041_), .A2(new_n13463_), .ZN(new_n30042_));
  OR3_X2     g26786(.A1(new_n30042_), .A2(new_n12841_), .A3(new_n5375_), .Z(new_n30043_));
  NOR3_X1    g26787(.A1(new_n12903_), .A2(new_n29831_), .A3(new_n30043_), .ZN(new_n30044_));
  XNOR2_X1   g26788(.A1(new_n30039_), .A2(new_n30044_), .ZN(new_n30045_));
  NOR2_X1    g26789(.A1(new_n12842_), .A2(pi0662), .ZN(new_n30046_));
  INV_X1     g26790(.I(new_n30046_), .ZN(new_n30047_));
  OAI22_X1   g26791(.A1(new_n29862_), .A2(new_n12845_), .B1(new_n29860_), .B2(new_n30047_), .ZN(new_n30048_));
  NAND3_X1   g26792(.A1(new_n30045_), .A2(pi0662), .A3(new_n30048_), .ZN(new_n30049_));
  NAND2_X1   g26793(.A1(new_n30049_), .A2(new_n5398_), .ZN(new_n30050_));
  XOR2_X1    g26794(.A1(new_n30050_), .A2(new_n28883_), .Z(new_n30051_));
  NAND2_X1   g26795(.A1(new_n30051_), .A2(new_n30037_), .ZN(new_n30052_));
  NOR4_X1    g26796(.A1(new_n13312_), .A2(new_n12868_), .A3(new_n12841_), .A4(new_n5375_), .ZN(new_n30053_));
  NOR3_X1    g26797(.A1(new_n13313_), .A2(pi0614), .A3(new_n5375_), .ZN(new_n30054_));
  OAI21_X1   g26798(.A1(new_n30054_), .A2(new_n30053_), .B(new_n29065_), .ZN(new_n30055_));
  NAND2_X1   g26799(.A1(new_n29876_), .A2(new_n12930_), .ZN(new_n30056_));
  NAND3_X1   g26800(.A1(new_n13390_), .A2(new_n12868_), .A3(new_n5633_), .ZN(new_n30057_));
  NAND3_X1   g26801(.A1(new_n30056_), .A2(new_n30057_), .A3(new_n5376_), .ZN(new_n30058_));
  OAI21_X1   g26802(.A1(new_n13321_), .A2(new_n13311_), .B(new_n5381_), .ZN(new_n30059_));
  AOI21_X1   g26803(.A1(new_n30055_), .A2(new_n30058_), .B(new_n30059_), .ZN(new_n30060_));
  NAND2_X1   g26804(.A1(new_n29589_), .A2(pi0614), .ZN(new_n30061_));
  AOI21_X1   g26805(.A1(new_n29044_), .A2(new_n30061_), .B(new_n5633_), .ZN(new_n30062_));
  XOR2_X1    g26806(.A1(new_n30062_), .A2(new_n28953_), .Z(new_n30063_));
  AOI21_X1   g26807(.A1(new_n29868_), .A2(new_n30046_), .B(new_n29873_), .ZN(new_n30064_));
  OAI21_X1   g26808(.A1(new_n30063_), .A2(new_n29868_), .B(new_n30064_), .ZN(new_n30065_));
  NAND2_X1   g26809(.A1(new_n30065_), .A2(pi0224), .ZN(new_n30066_));
  XOR2_X1    g26810(.A1(new_n30066_), .A2(new_n28883_), .Z(new_n30067_));
  AOI21_X1   g26811(.A1(new_n30067_), .A2(new_n30060_), .B(new_n3565_), .ZN(new_n30068_));
  AOI22_X1   g26812(.A1(new_n30052_), .A2(new_n30068_), .B1(new_n30030_), .B2(new_n30034_), .ZN(new_n30069_));
  NAND2_X1   g26813(.A1(new_n29128_), .A2(pi0680), .ZN(new_n30070_));
  NAND2_X1   g26814(.A1(new_n29121_), .A2(pi0614), .ZN(new_n30071_));
  NAND2_X1   g26815(.A1(new_n29129_), .A2(new_n12869_), .ZN(new_n30072_));
  XNOR2_X1   g26816(.A1(new_n30071_), .A2(new_n30072_), .ZN(new_n30073_));
  NOR3_X1    g26817(.A1(new_n29822_), .A2(new_n5375_), .A3(new_n30073_), .ZN(new_n30074_));
  XOR2_X1    g26818(.A1(new_n30074_), .A2(new_n30070_), .Z(new_n30075_));
  AOI21_X1   g26819(.A1(new_n29821_), .A2(new_n5373_), .B(new_n30047_), .ZN(new_n30076_));
  OAI21_X1   g26820(.A1(new_n29828_), .A2(new_n30076_), .B(pi0662), .ZN(new_n30077_));
  NOR2_X1    g26821(.A1(new_n30075_), .A2(new_n30077_), .ZN(new_n30078_));
  OAI21_X1   g26822(.A1(new_n13535_), .A2(new_n13494_), .B(pi0680), .ZN(new_n30079_));
  INV_X1     g26823(.I(new_n29832_), .ZN(new_n30080_));
  NOR2_X1    g26824(.A1(new_n30080_), .A2(new_n30043_), .ZN(new_n30081_));
  XNOR2_X1   g26825(.A1(new_n30079_), .A2(new_n30081_), .ZN(new_n30082_));
  OAI22_X1   g26826(.A1(new_n29834_), .A2(new_n12845_), .B1(new_n29832_), .B2(new_n30047_), .ZN(new_n30083_));
  AND2_X2    g26827(.A1(new_n30083_), .A2(pi0662), .Z(new_n30084_));
  NAND2_X1   g26828(.A1(new_n30084_), .A2(new_n30082_), .ZN(new_n30085_));
  NAND2_X1   g26829(.A1(new_n30085_), .A2(pi0224), .ZN(new_n30086_));
  XOR2_X1    g26830(.A1(new_n30086_), .A2(new_n28883_), .Z(new_n30087_));
  NAND2_X1   g26831(.A1(new_n30087_), .A2(new_n30078_), .ZN(new_n30088_));
  OAI21_X1   g26832(.A1(new_n30088_), .A2(new_n30069_), .B(new_n3183_), .ZN(new_n30089_));
  INV_X1     g26833(.I(new_n30089_), .ZN(new_n30090_));
  NAND4_X1   g26834(.A1(new_n30084_), .A2(pi0224), .A3(new_n5454_), .A4(new_n30082_), .ZN(new_n30091_));
  NAND3_X1   g26835(.A1(new_n30085_), .A2(new_n3100_), .A3(new_n5454_), .ZN(new_n30092_));
  AND2_X2    g26836(.A1(new_n30092_), .A2(new_n30091_), .Z(new_n30093_));
  NOR2_X1    g26837(.A1(new_n29845_), .A2(new_n3313_), .ZN(new_n30094_));
  OR3_X2     g26838(.A1(new_n30032_), .A2(pi0215), .A3(new_n30094_), .Z(new_n30095_));
  NAND3_X1   g26839(.A1(pi0224), .A2(pi0662), .A3(pi0680), .ZN(new_n30096_));
  NOR2_X1    g26840(.A1(new_n30041_), .A2(new_n30096_), .ZN(new_n30097_));
  AOI21_X1   g26841(.A1(new_n30095_), .A2(new_n30097_), .B(new_n3312_), .ZN(new_n30098_));
  OAI21_X1   g26842(.A1(new_n30093_), .A2(new_n30019_), .B(new_n30098_), .ZN(new_n30099_));
  NAND2_X1   g26843(.A1(new_n30049_), .A2(pi0224), .ZN(new_n30100_));
  XOR2_X1    g26844(.A1(new_n30100_), .A2(new_n29838_), .Z(new_n30101_));
  NOR2_X1    g26845(.A1(new_n30101_), .A2(new_n30065_), .ZN(new_n30102_));
  NOR2_X1    g26846(.A1(new_n30102_), .A2(new_n29585_), .ZN(new_n30103_));
  NAND2_X1   g26847(.A1(new_n30027_), .A2(pi0224), .ZN(new_n30104_));
  XOR2_X1    g26848(.A1(new_n30104_), .A2(new_n29840_), .Z(new_n30105_));
  NAND2_X1   g26849(.A1(new_n30036_), .A2(new_n5454_), .ZN(new_n30106_));
  XOR2_X1    g26850(.A1(new_n30106_), .A2(new_n29840_), .Z(new_n30107_));
  NAND4_X1   g26851(.A1(new_n30105_), .A2(new_n30060_), .A3(new_n30078_), .A4(new_n30107_), .ZN(new_n30108_));
  NOR2_X1    g26852(.A1(new_n30103_), .A2(new_n30108_), .ZN(new_n30109_));
  NAND2_X1   g26853(.A1(new_n30109_), .A2(new_n30099_), .ZN(new_n30110_));
  OAI21_X1   g26854(.A1(new_n30090_), .A2(new_n30110_), .B(new_n3259_), .ZN(new_n30111_));
  INV_X1     g26855(.I(new_n29156_), .ZN(new_n30112_));
  NAND2_X1   g26856(.A1(new_n30112_), .A2(new_n29885_), .ZN(new_n30113_));
  NAND3_X1   g26857(.A1(new_n30113_), .A2(new_n13136_), .A3(new_n28952_), .ZN(new_n30114_));
  NAND2_X1   g26858(.A1(new_n29892_), .A2(pi0299), .ZN(new_n30115_));
  NAND2_X1   g26859(.A1(new_n28952_), .A2(pi0299), .ZN(new_n30116_));
  XOR2_X1    g26860(.A1(new_n30115_), .A2(new_n30116_), .Z(new_n30117_));
  NAND2_X1   g26861(.A1(new_n13192_), .A2(new_n12868_), .ZN(new_n30118_));
  NAND4_X1   g26862(.A1(new_n29142_), .A2(pi0224), .A3(new_n29145_), .A4(new_n30118_), .ZN(new_n30119_));
  XNOR2_X1   g26863(.A1(new_n30119_), .A2(new_n29890_), .ZN(new_n30120_));
  NAND3_X1   g26864(.A1(new_n30120_), .A2(pi0299), .A3(new_n30117_), .ZN(new_n30121_));
  NAND2_X1   g26865(.A1(new_n30121_), .A2(new_n30114_), .ZN(new_n30122_));
  OAI21_X1   g26866(.A1(new_n29887_), .A2(new_n3100_), .B(new_n28953_), .ZN(new_n30123_));
  NOR3_X1    g26867(.A1(new_n3290_), .A2(new_n3183_), .A3(new_n3100_), .ZN(new_n30124_));
  NAND4_X1   g26868(.A1(new_n30122_), .A2(new_n13136_), .A3(new_n30123_), .A4(new_n30124_), .ZN(new_n30125_));
  INV_X1     g26869(.I(new_n30125_), .ZN(new_n30126_));
  NAND3_X1   g26870(.A1(new_n30111_), .A2(new_n30014_), .A3(new_n30126_), .ZN(new_n30127_));
  INV_X1     g26871(.I(new_n30014_), .ZN(new_n30128_));
  INV_X1     g26872(.I(new_n30110_), .ZN(new_n30129_));
  AOI21_X1   g26873(.A1(new_n30129_), .A2(new_n30089_), .B(pi0038), .ZN(new_n30130_));
  OAI21_X1   g26874(.A1(new_n30130_), .A2(new_n30125_), .B(new_n30128_), .ZN(new_n30131_));
  NAND2_X1   g26875(.A1(new_n30131_), .A2(new_n30127_), .ZN(new_n30132_));
  NAND2_X1   g26876(.A1(new_n29912_), .A2(new_n29905_), .ZN(new_n30133_));
  NOR3_X1    g26877(.A1(new_n30130_), .A2(new_n30128_), .A3(new_n30125_), .ZN(new_n30134_));
  AOI21_X1   g26878(.A1(new_n30111_), .A2(new_n30126_), .B(new_n30014_), .ZN(new_n30135_));
  NOR2_X1    g26879(.A1(new_n30134_), .A2(new_n30135_), .ZN(new_n30136_));
  AOI21_X1   g26880(.A1(new_n30136_), .A2(pi0625), .B(new_n13620_), .ZN(new_n30137_));
  NOR3_X1    g26881(.A1(new_n30132_), .A2(new_n13613_), .A3(new_n13615_), .ZN(new_n30138_));
  OAI21_X1   g26882(.A1(new_n30137_), .A2(new_n30138_), .B(new_n30133_), .ZN(new_n30139_));
  AOI21_X1   g26883(.A1(new_n30003_), .A2(new_n29922_), .B(pi0608), .ZN(new_n30140_));
  AOI21_X1   g26884(.A1(new_n29999_), .A2(new_n29922_), .B(pi0608), .ZN(new_n30141_));
  INV_X1     g26885(.I(new_n30141_), .ZN(new_n30142_));
  AOI21_X1   g26886(.A1(new_n30139_), .A2(new_n30140_), .B(new_n30142_), .ZN(new_n30143_));
  NOR2_X1    g26887(.A1(new_n30132_), .A2(new_n13614_), .ZN(new_n30144_));
  NOR2_X1    g26888(.A1(new_n30144_), .A2(new_n13620_), .ZN(new_n30145_));
  NAND2_X1   g26889(.A1(new_n30144_), .A2(new_n13620_), .ZN(new_n30146_));
  INV_X1     g26890(.I(new_n30146_), .ZN(new_n30147_));
  INV_X1     g26891(.I(new_n30133_), .ZN(new_n30148_));
  NOR2_X1    g26892(.A1(new_n30148_), .A2(new_n13748_), .ZN(new_n30149_));
  OAI21_X1   g26893(.A1(new_n30147_), .A2(new_n30145_), .B(new_n30149_), .ZN(new_n30150_));
  OAI22_X1   g26894(.A1(new_n30150_), .A2(new_n30143_), .B1(pi0778), .B2(new_n30132_), .ZN(new_n30151_));
  NAND3_X1   g26895(.A1(new_n30151_), .A2(pi0609), .A3(pi1155), .ZN(new_n30152_));
  NAND3_X1   g26896(.A1(new_n30132_), .A2(pi0625), .A3(pi1153), .ZN(new_n30153_));
  NAND3_X1   g26897(.A1(new_n30136_), .A2(pi0625), .A3(new_n13620_), .ZN(new_n30154_));
  AOI21_X1   g26898(.A1(new_n30154_), .A2(new_n30153_), .B(new_n30148_), .ZN(new_n30155_));
  INV_X1     g26899(.I(new_n30140_), .ZN(new_n30156_));
  OAI21_X1   g26900(.A1(new_n30155_), .A2(new_n30156_), .B(new_n30141_), .ZN(new_n30157_));
  INV_X1     g26901(.I(new_n30145_), .ZN(new_n30158_));
  INV_X1     g26902(.I(new_n30149_), .ZN(new_n30159_));
  AOI21_X1   g26903(.A1(new_n30158_), .A2(new_n30146_), .B(new_n30159_), .ZN(new_n30160_));
  AOI22_X1   g26904(.A1(new_n30160_), .A2(new_n30157_), .B1(new_n13748_), .B2(new_n30136_), .ZN(new_n30161_));
  NAND3_X1   g26905(.A1(new_n30161_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n30162_));
  AOI21_X1   g26906(.A1(new_n30162_), .A2(new_n30152_), .B(new_n30007_), .ZN(new_n30163_));
  NOR2_X1    g26907(.A1(new_n29917_), .A2(new_n13783_), .ZN(new_n30164_));
  INV_X1     g26908(.I(new_n30164_), .ZN(new_n30165_));
  OAI21_X1   g26909(.A1(new_n30163_), .A2(new_n30165_), .B(pi0785), .ZN(new_n30166_));
  INV_X1     g26910(.I(new_n30007_), .ZN(new_n30167_));
  NAND3_X1   g26911(.A1(new_n30151_), .A2(pi0609), .A3(pi1155), .ZN(new_n30168_));
  NAND3_X1   g26912(.A1(new_n30161_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n30169_));
  NAND2_X1   g26913(.A1(new_n30169_), .A2(new_n30168_), .ZN(new_n30170_));
  NOR3_X1    g26914(.A1(new_n30161_), .A2(new_n29193_), .A3(new_n29920_), .ZN(new_n30171_));
  INV_X1     g26915(.I(new_n30171_), .ZN(new_n30172_));
  AOI21_X1   g26916(.A1(new_n30170_), .A2(new_n30167_), .B(new_n30172_), .ZN(new_n30173_));
  NAND2_X1   g26917(.A1(new_n30166_), .A2(new_n30173_), .ZN(new_n30174_));
  AOI21_X1   g26918(.A1(new_n30161_), .A2(pi1155), .B(new_n14694_), .ZN(new_n30175_));
  NOR3_X1    g26919(.A1(new_n30151_), .A2(pi0609), .A3(new_n13778_), .ZN(new_n30176_));
  OAI21_X1   g26920(.A1(new_n30175_), .A2(new_n30176_), .B(new_n30167_), .ZN(new_n30177_));
  AOI21_X1   g26921(.A1(new_n30177_), .A2(new_n30164_), .B(new_n13801_), .ZN(new_n30178_));
  AOI21_X1   g26922(.A1(new_n30161_), .A2(pi0609), .B(new_n14694_), .ZN(new_n30179_));
  NOR3_X1    g26923(.A1(new_n30151_), .A2(new_n13766_), .A3(pi1155), .ZN(new_n30180_));
  OAI21_X1   g26924(.A1(new_n30179_), .A2(new_n30180_), .B(new_n30167_), .ZN(new_n30181_));
  NAND2_X1   g26925(.A1(new_n30181_), .A2(new_n30171_), .ZN(new_n30182_));
  NAND2_X1   g26926(.A1(new_n30178_), .A2(new_n30182_), .ZN(new_n30183_));
  NAND2_X1   g26927(.A1(new_n30183_), .A2(new_n30174_), .ZN(new_n30184_));
  INV_X1     g26928(.I(new_n30010_), .ZN(new_n30185_));
  NOR2_X1    g26929(.A1(new_n29935_), .A2(new_n14501_), .ZN(new_n30186_));
  AOI21_X1   g26930(.A1(new_n30186_), .A2(new_n30185_), .B(pi0618), .ZN(new_n30187_));
  INV_X1     g26931(.I(new_n30187_), .ZN(new_n30188_));
  AOI21_X1   g26932(.A1(new_n29933_), .A2(pi1154), .B(new_n13819_), .ZN(new_n30189_));
  INV_X1     g26933(.I(new_n29937_), .ZN(new_n30190_));
  OAI21_X1   g26934(.A1(new_n30189_), .A2(new_n30190_), .B(new_n29922_), .ZN(new_n30191_));
  AOI21_X1   g26935(.A1(new_n30191_), .A2(new_n13836_), .B(pi0618), .ZN(new_n30192_));
  INV_X1     g26936(.I(new_n30192_), .ZN(new_n30193_));
  NAND4_X1   g26937(.A1(new_n30184_), .A2(pi0781), .A3(new_n30188_), .A4(new_n30193_), .ZN(new_n30194_));
  NOR2_X1    g26938(.A1(new_n30178_), .A2(new_n30182_), .ZN(new_n30195_));
  NOR2_X1    g26939(.A1(new_n30166_), .A2(new_n30173_), .ZN(new_n30196_));
  OAI21_X1   g26940(.A1(new_n30195_), .A2(new_n30196_), .B(new_n30188_), .ZN(new_n30197_));
  NOR2_X1    g26941(.A1(new_n30192_), .A2(new_n13855_), .ZN(new_n30198_));
  OAI21_X1   g26942(.A1(new_n30195_), .A2(new_n30196_), .B(new_n30198_), .ZN(new_n30199_));
  NAND3_X1   g26943(.A1(new_n30197_), .A2(new_n30199_), .A3(pi0781), .ZN(new_n30200_));
  NAND2_X1   g26944(.A1(new_n30200_), .A2(new_n30194_), .ZN(new_n30201_));
  NAND3_X1   g26945(.A1(new_n30201_), .A2(pi0619), .A3(pi1159), .ZN(new_n30202_));
  NAND4_X1   g26946(.A1(new_n30200_), .A2(new_n30194_), .A3(new_n13860_), .A4(pi1159), .ZN(new_n30203_));
  AOI21_X1   g26947(.A1(new_n30202_), .A2(new_n30203_), .B(new_n30012_), .ZN(new_n30204_));
  OAI21_X1   g26948(.A1(new_n30204_), .A2(new_n20003_), .B(new_n29948_), .ZN(new_n30205_));
  NAND3_X1   g26949(.A1(new_n29945_), .A2(pi0619), .A3(pi1159), .ZN(new_n30206_));
  NAND4_X1   g26950(.A1(new_n29944_), .A2(new_n13860_), .A3(new_n29939_), .A4(pi1159), .ZN(new_n30207_));
  AOI21_X1   g26951(.A1(new_n30206_), .A2(new_n30207_), .B(new_n29811_), .ZN(new_n30208_));
  NAND4_X1   g26952(.A1(new_n29948_), .A2(new_n30208_), .A3(pi0789), .A4(new_n29945_), .ZN(new_n30209_));
  AOI21_X1   g26953(.A1(pi0781), .A2(new_n29942_), .B(new_n29943_), .ZN(new_n30210_));
  NAND2_X1   g26954(.A1(new_n29942_), .A2(pi0781), .ZN(new_n30211_));
  NOR3_X1    g26955(.A1(new_n30191_), .A2(new_n13855_), .A3(new_n29933_), .ZN(new_n30212_));
  NOR2_X1    g26956(.A1(new_n30212_), .A2(new_n30211_), .ZN(new_n30213_));
  NOR2_X1    g26957(.A1(new_n30213_), .A2(new_n30210_), .ZN(new_n30214_));
  AOI21_X1   g26958(.A1(new_n30214_), .A2(pi0619), .B(new_n13904_), .ZN(new_n30215_));
  INV_X1     g26959(.I(new_n29947_), .ZN(new_n30216_));
  OAI21_X1   g26960(.A1(new_n30215_), .A2(new_n30216_), .B(new_n29922_), .ZN(new_n30217_));
  NOR2_X1    g26961(.A1(new_n30214_), .A2(new_n13896_), .ZN(new_n30218_));
  NAND2_X1   g26962(.A1(new_n30208_), .A2(new_n30218_), .ZN(new_n30219_));
  NAND3_X1   g26963(.A1(new_n30219_), .A2(pi0789), .A3(new_n30217_), .ZN(new_n30220_));
  NAND3_X1   g26964(.A1(new_n30220_), .A2(new_n13962_), .A3(new_n30209_), .ZN(new_n30221_));
  NAND2_X1   g26965(.A1(new_n30221_), .A2(new_n18975_), .ZN(new_n30222_));
  NAND4_X1   g26966(.A1(new_n30220_), .A2(new_n13901_), .A3(new_n13962_), .A4(new_n30209_), .ZN(new_n30223_));
  NAND2_X1   g26967(.A1(new_n30222_), .A2(new_n30223_), .ZN(new_n30224_));
  NAND2_X1   g26968(.A1(new_n30201_), .A2(new_n13896_), .ZN(new_n30225_));
  INV_X1     g26969(.I(new_n30209_), .ZN(new_n30226_));
  NAND2_X1   g26970(.A1(new_n30217_), .A2(pi0789), .ZN(new_n30227_));
  INV_X1     g26971(.I(new_n30219_), .ZN(new_n30228_));
  NOR2_X1    g26972(.A1(new_n30228_), .A2(new_n30227_), .ZN(new_n30229_));
  AOI21_X1   g26973(.A1(new_n30012_), .A2(new_n16639_), .B(new_n16829_), .ZN(new_n30230_));
  INV_X1     g26974(.I(new_n30012_), .ZN(new_n30231_));
  NOR3_X1    g26975(.A1(new_n30231_), .A2(new_n14162_), .A3(new_n16828_), .ZN(new_n30232_));
  NOR3_X1    g26976(.A1(new_n29811_), .A2(pi0626), .A3(new_n19208_), .ZN(new_n30233_));
  OAI21_X1   g26977(.A1(new_n30232_), .A2(new_n30230_), .B(new_n30233_), .ZN(new_n30234_));
  NAND2_X1   g26978(.A1(new_n30234_), .A2(new_n13901_), .ZN(new_n30235_));
  OAI21_X1   g26979(.A1(new_n30229_), .A2(new_n30226_), .B(new_n30235_), .ZN(new_n30236_));
  NAND2_X1   g26980(.A1(new_n29922_), .A2(new_n14143_), .ZN(new_n30237_));
  AOI21_X1   g26981(.A1(new_n30236_), .A2(new_n19204_), .B(new_n30237_), .ZN(new_n30238_));
  NAND3_X1   g26982(.A1(new_n30224_), .A2(new_n30238_), .A3(new_n30225_), .ZN(new_n30239_));
  NOR2_X1    g26983(.A1(new_n30195_), .A2(new_n30196_), .ZN(new_n30240_));
  NOR4_X1    g26984(.A1(new_n30240_), .A2(new_n13855_), .A3(new_n30187_), .A4(new_n30192_), .ZN(new_n30241_));
  AOI21_X1   g26985(.A1(new_n30183_), .A2(new_n30174_), .B(new_n30187_), .ZN(new_n30242_));
  INV_X1     g26986(.I(new_n30198_), .ZN(new_n30243_));
  AOI21_X1   g26987(.A1(new_n30183_), .A2(new_n30174_), .B(new_n30243_), .ZN(new_n30244_));
  NOR3_X1    g26988(.A1(new_n30242_), .A2(new_n30244_), .A3(new_n13855_), .ZN(new_n30245_));
  NOR3_X1    g26989(.A1(new_n30245_), .A2(new_n30241_), .A3(new_n13860_), .ZN(new_n30246_));
  NOR2_X1    g26990(.A1(new_n30246_), .A2(new_n13904_), .ZN(new_n30247_));
  NOR3_X1    g26991(.A1(new_n30201_), .A2(new_n13860_), .A3(new_n13903_), .ZN(new_n30248_));
  OAI21_X1   g26992(.A1(new_n30247_), .A2(new_n30248_), .B(new_n30231_), .ZN(new_n30249_));
  NOR2_X1    g26993(.A1(new_n30208_), .A2(pi0648), .ZN(new_n30250_));
  NAND2_X1   g26994(.A1(new_n30249_), .A2(new_n30250_), .ZN(new_n30251_));
  AOI21_X1   g26995(.A1(new_n30239_), .A2(new_n30205_), .B(new_n30251_), .ZN(new_n30252_));
  NOR2_X1    g26996(.A1(new_n29811_), .A2(new_n14059_), .ZN(new_n30253_));
  NAND3_X1   g26997(.A1(new_n30231_), .A2(new_n15395_), .A3(new_n29922_), .ZN(new_n30254_));
  NAND3_X1   g26998(.A1(new_n30012_), .A2(new_n15395_), .A3(new_n29811_), .ZN(new_n30255_));
  AOI21_X1   g26999(.A1(new_n30254_), .A2(new_n30255_), .B(new_n14059_), .ZN(new_n30256_));
  NOR2_X1    g27000(.A1(new_n30256_), .A2(new_n30253_), .ZN(new_n30257_));
  AOI21_X1   g27001(.A1(new_n30257_), .A2(pi0647), .B(new_n14008_), .ZN(new_n30258_));
  NOR4_X1    g27002(.A1(new_n30256_), .A2(new_n14005_), .A3(pi1157), .A4(new_n30253_), .ZN(new_n30259_));
  OAI21_X1   g27003(.A1(new_n30258_), .A2(new_n30259_), .B(new_n29922_), .ZN(new_n30260_));
  NAND2_X1   g27004(.A1(new_n30260_), .A2(pi0630), .ZN(new_n30261_));
  AOI21_X1   g27005(.A1(new_n30257_), .A2(pi1157), .B(new_n14008_), .ZN(new_n30262_));
  NOR4_X1    g27006(.A1(new_n30256_), .A2(pi0647), .A3(new_n14006_), .A4(new_n30253_), .ZN(new_n30263_));
  OAI21_X1   g27007(.A1(new_n30262_), .A2(new_n30263_), .B(new_n29922_), .ZN(new_n30264_));
  NAND2_X1   g27008(.A1(new_n30264_), .A2(new_n14010_), .ZN(new_n30265_));
  NAND2_X1   g27009(.A1(new_n30261_), .A2(new_n30265_), .ZN(new_n30266_));
  AOI21_X1   g27010(.A1(new_n30266_), .A2(pi0787), .B(new_n16576_), .ZN(new_n30267_));
  NOR2_X1    g27011(.A1(new_n29922_), .A2(new_n13994_), .ZN(new_n30268_));
  NOR2_X1    g27012(.A1(new_n29811_), .A2(new_n16372_), .ZN(new_n30269_));
  INV_X1     g27013(.I(new_n30269_), .ZN(new_n30270_));
  NAND3_X1   g27014(.A1(new_n30220_), .A2(new_n16372_), .A3(new_n30209_), .ZN(new_n30271_));
  AND2_X2    g27015(.A1(new_n30271_), .A2(new_n30270_), .Z(new_n30272_));
  AOI21_X1   g27016(.A1(new_n30272_), .A2(new_n13994_), .B(new_n30268_), .ZN(new_n30273_));
  NOR3_X1    g27017(.A1(new_n30273_), .A2(new_n16419_), .A3(new_n30267_), .ZN(new_n30274_));
  NAND2_X1   g27018(.A1(new_n30254_), .A2(new_n30255_), .ZN(new_n30275_));
  NOR2_X1    g27019(.A1(new_n29922_), .A2(new_n13942_), .ZN(new_n30276_));
  OAI22_X1   g27020(.A1(new_n30275_), .A2(new_n13942_), .B1(new_n19484_), .B2(new_n30276_), .ZN(new_n30277_));
  NAND3_X1   g27021(.A1(new_n30254_), .A2(pi0628), .A3(new_n30255_), .ZN(new_n30278_));
  NAND2_X1   g27022(.A1(new_n29922_), .A2(new_n29298_), .ZN(new_n30279_));
  AOI21_X1   g27023(.A1(new_n30278_), .A2(new_n30279_), .B(new_n12777_), .ZN(new_n30280_));
  NAND2_X1   g27024(.A1(new_n30277_), .A2(new_n30280_), .ZN(new_n30281_));
  AOI21_X1   g27025(.A1(new_n30272_), .A2(new_n30281_), .B(new_n16875_), .ZN(new_n30282_));
  OAI21_X1   g27026(.A1(new_n30252_), .A2(new_n30274_), .B(new_n30282_), .ZN(new_n30283_));
  NAND2_X1   g27027(.A1(new_n29922_), .A2(new_n14210_), .ZN(new_n30284_));
  INV_X1     g27028(.I(new_n30268_), .ZN(new_n30285_));
  NAND3_X1   g27029(.A1(new_n30271_), .A2(new_n13994_), .A3(new_n30270_), .ZN(new_n30286_));
  NAND3_X1   g27030(.A1(new_n30286_), .A2(new_n14211_), .A3(new_n30285_), .ZN(new_n30287_));
  NAND3_X1   g27031(.A1(new_n30287_), .A2(pi0715), .A3(new_n30284_), .ZN(new_n30288_));
  NAND2_X1   g27032(.A1(new_n30288_), .A2(new_n14205_), .ZN(new_n30289_));
  NAND4_X1   g27033(.A1(new_n30287_), .A2(new_n14204_), .A3(pi0715), .A4(new_n30284_), .ZN(new_n30290_));
  AOI21_X1   g27034(.A1(new_n30289_), .A2(new_n30290_), .B(new_n29811_), .ZN(new_n30291_));
  NAND2_X1   g27035(.A1(new_n30260_), .A2(pi0787), .ZN(new_n30292_));
  NOR3_X1    g27036(.A1(new_n30264_), .A2(new_n12776_), .A3(new_n30257_), .ZN(new_n30293_));
  XOR2_X1    g27037(.A1(new_n30293_), .A2(new_n30292_), .Z(new_n30294_));
  OAI21_X1   g27038(.A1(new_n30294_), .A2(new_n14204_), .B(new_n15385_), .ZN(new_n30295_));
  OAI21_X1   g27039(.A1(new_n30291_), .A2(new_n30295_), .B(new_n30283_), .ZN(new_n30296_));
  AOI21_X1   g27040(.A1(new_n30296_), .A2(pi0644), .B(new_n12775_), .ZN(new_n30297_));
  NAND3_X1   g27041(.A1(new_n30287_), .A2(pi0644), .A3(new_n30284_), .ZN(new_n30298_));
  NAND2_X1   g27042(.A1(new_n30298_), .A2(new_n14205_), .ZN(new_n30299_));
  NAND4_X1   g27043(.A1(new_n30287_), .A2(pi0644), .A3(new_n14200_), .A4(new_n30284_), .ZN(new_n30300_));
  AOI21_X1   g27044(.A1(new_n30299_), .A2(new_n30300_), .B(new_n29811_), .ZN(new_n30301_));
  OAI21_X1   g27045(.A1(new_n30294_), .A2(pi0644), .B(new_n14243_), .ZN(new_n30302_));
  OAI21_X1   g27046(.A1(new_n30301_), .A2(new_n30302_), .B(new_n14204_), .ZN(new_n30303_));
  NOR2_X1    g27047(.A1(new_n30283_), .A2(new_n12775_), .ZN(new_n30304_));
  NAND2_X1   g27048(.A1(new_n30303_), .A2(new_n30304_), .ZN(new_n30305_));
  XOR2_X1    g27049(.A1(new_n30297_), .A2(new_n30305_), .Z(new_n30306_));
  NAND2_X1   g27050(.A1(po1038), .A2(pi0224), .ZN(new_n30307_));
  OAI21_X1   g27051(.A1(new_n30306_), .A2(po1038), .B(new_n30307_), .ZN(po0381));
  OAI21_X1   g27052(.A1(new_n2921_), .A2(new_n2752_), .B(pi0137), .ZN(new_n30309_));
  NAND2_X1   g27053(.A1(new_n30309_), .A2(pi0332), .ZN(new_n30310_));
  INV_X1     g27054(.I(new_n2969_), .ZN(new_n30311_));
  AOI21_X1   g27055(.A1(new_n2734_), .A2(new_n9239_), .B(new_n2961_), .ZN(new_n30312_));
  NOR2_X1    g27056(.A1(new_n30312_), .A2(new_n2968_), .ZN(new_n30313_));
  NOR3_X1    g27057(.A1(new_n2484_), .A2(new_n2806_), .A3(new_n9239_), .ZN(new_n30314_));
  OAI21_X1   g27058(.A1(new_n2886_), .A2(new_n30314_), .B(new_n2503_), .ZN(new_n30315_));
  AOI21_X1   g27059(.A1(new_n30315_), .A2(new_n3041_), .B(new_n2920_), .ZN(new_n30316_));
  NAND4_X1   g27060(.A1(new_n30313_), .A2(new_n30311_), .A3(new_n2776_), .A4(pi0332), .ZN(new_n30317_));
  XOR2_X1    g27061(.A1(new_n30310_), .A2(new_n30317_), .Z(new_n30318_));
  NOR2_X1    g27062(.A1(new_n2968_), .A2(new_n6427_), .ZN(new_n30319_));
  XOR2_X1    g27063(.A1(new_n30313_), .A2(new_n30319_), .Z(new_n30320_));
  NOR2_X1    g27064(.A1(new_n6382_), .A2(new_n2735_), .ZN(new_n30321_));
  NAND4_X1   g27065(.A1(new_n30320_), .A2(new_n2715_), .A3(new_n9237_), .A4(new_n30321_), .ZN(new_n30322_));
  NOR2_X1    g27066(.A1(new_n2729_), .A2(pi0137), .ZN(new_n30323_));
  INV_X1     g27067(.I(new_n30323_), .ZN(new_n30324_));
  AOI21_X1   g27068(.A1(new_n2908_), .A2(new_n30321_), .B(pi0032), .ZN(new_n30325_));
  INV_X1     g27069(.I(new_n30325_), .ZN(new_n30326_));
  AOI21_X1   g27070(.A1(new_n30326_), .A2(new_n30319_), .B(pi1093), .ZN(new_n30327_));
  AOI21_X1   g27071(.A1(new_n30327_), .A2(new_n30313_), .B(new_n30324_), .ZN(new_n30328_));
  OAI21_X1   g27072(.A1(new_n30322_), .A2(new_n2984_), .B(new_n30328_), .ZN(new_n30329_));
  INV_X1     g27073(.I(new_n30327_), .ZN(new_n30330_));
  AOI21_X1   g27074(.A1(new_n2969_), .A2(new_n6427_), .B(new_n30330_), .ZN(new_n30331_));
  AOI21_X1   g27075(.A1(new_n30319_), .A2(pi0032), .B(new_n30321_), .ZN(new_n30332_));
  OAI21_X1   g27076(.A1(new_n30332_), .A2(new_n2935_), .B(new_n2984_), .ZN(new_n30333_));
  NOR2_X1    g27077(.A1(new_n6427_), .A2(new_n30323_), .ZN(new_n30334_));
  NAND4_X1   g27078(.A1(new_n30331_), .A2(new_n2969_), .A3(new_n30333_), .A4(new_n30334_), .ZN(new_n30335_));
  OR2_X2     g27079(.A1(new_n30335_), .A2(new_n30322_), .Z(new_n30336_));
  NAND2_X1   g27080(.A1(new_n30335_), .A2(new_n30323_), .ZN(new_n30337_));
  OAI21_X1   g27081(.A1(new_n2969_), .A2(new_n2984_), .B(pi0332), .ZN(new_n30338_));
  NOR2_X1    g27082(.A1(new_n30331_), .A2(new_n30338_), .ZN(new_n30339_));
  AND4_X2    g27083(.A1(new_n30329_), .A2(new_n30336_), .A3(new_n30337_), .A4(new_n30339_), .Z(new_n30340_));
  OAI21_X1   g27084(.A1(new_n30316_), .A2(new_n2776_), .B(new_n30340_), .ZN(new_n30341_));
  XNOR2_X1   g27085(.A1(new_n30310_), .A2(new_n30341_), .ZN(new_n30342_));
  NAND2_X1   g27086(.A1(new_n30342_), .A2(new_n3030_), .ZN(new_n30343_));
  NAND2_X1   g27087(.A1(new_n3030_), .A2(pi0210), .ZN(new_n30344_));
  XOR2_X1    g27088(.A1(new_n30343_), .A2(new_n30344_), .Z(new_n30345_));
  NAND2_X1   g27089(.A1(new_n30345_), .A2(new_n30318_), .ZN(new_n30346_));
  NAND2_X1   g27090(.A1(new_n30315_), .A2(new_n3051_), .ZN(new_n30347_));
  AOI21_X1   g27091(.A1(new_n30347_), .A2(new_n2851_), .B(new_n2955_), .ZN(new_n30348_));
  INV_X1     g27092(.I(new_n30312_), .ZN(new_n30349_));
  AOI21_X1   g27093(.A1(pi0137), .A2(new_n2962_), .B(new_n2889_), .ZN(new_n30350_));
  NAND4_X1   g27094(.A1(new_n2752_), .A2(pi0095), .A3(pi0137), .A4(pi0332), .ZN(new_n30351_));
  NOR4_X1    g27095(.A1(new_n30350_), .A2(new_n2852_), .A3(new_n30349_), .A4(new_n30351_), .ZN(new_n30352_));
  XOR2_X1    g27096(.A1(new_n30352_), .A2(new_n30348_), .Z(new_n30353_));
  NAND2_X1   g27097(.A1(new_n30353_), .A2(pi0210), .ZN(new_n30354_));
  AOI21_X1   g27098(.A1(new_n30346_), .A2(new_n3098_), .B(new_n30354_), .ZN(new_n30355_));
  AOI21_X1   g27099(.A1(new_n3211_), .A2(new_n2776_), .B(new_n3183_), .ZN(new_n30356_));
  AOI21_X1   g27100(.A1(new_n3160_), .A2(new_n30356_), .B(new_n30355_), .ZN(new_n30357_));
  NAND2_X1   g27101(.A1(new_n30342_), .A2(new_n5500_), .ZN(new_n30358_));
  NAND2_X1   g27102(.A1(new_n5500_), .A2(pi0198), .ZN(new_n30359_));
  XOR2_X1    g27103(.A1(new_n30358_), .A2(new_n30359_), .Z(new_n30360_));
  NAND2_X1   g27104(.A1(new_n30360_), .A2(new_n30318_), .ZN(new_n30361_));
  NAND2_X1   g27105(.A1(new_n30361_), .A2(new_n3098_), .ZN(new_n30362_));
  NAND4_X1   g27106(.A1(new_n30362_), .A2(pi0198), .A3(new_n5507_), .A4(new_n30353_), .ZN(new_n30363_));
  OAI21_X1   g27107(.A1(new_n5502_), .A2(new_n5469_), .B(new_n2776_), .ZN(new_n30364_));
  AOI21_X1   g27108(.A1(new_n2776_), .A2(new_n5486_), .B(new_n30364_), .ZN(new_n30365_));
  AOI21_X1   g27109(.A1(new_n5492_), .A2(new_n30365_), .B(new_n3455_), .ZN(new_n30366_));
  OAI21_X1   g27110(.A1(new_n30357_), .A2(new_n30363_), .B(new_n30366_), .ZN(new_n30367_));
  XOR2_X1    g27111(.A1(new_n30367_), .A2(new_n3694_), .Z(new_n30368_));
  NOR2_X1    g27112(.A1(new_n6295_), .A2(new_n3208_), .ZN(new_n30369_));
  NOR3_X1    g27113(.A1(new_n3145_), .A2(new_n2776_), .A3(new_n3474_), .ZN(new_n30370_));
  INV_X1     g27114(.I(new_n30370_), .ZN(new_n30371_));
  NAND2_X1   g27115(.A1(new_n3205_), .A2(new_n9569_), .ZN(new_n30372_));
  OAI21_X1   g27116(.A1(new_n30371_), .A2(new_n30372_), .B(new_n3258_), .ZN(new_n30373_));
  NOR2_X1    g27117(.A1(new_n30369_), .A2(new_n30373_), .ZN(new_n30374_));
  AOI21_X1   g27118(.A1(new_n12112_), .A2(new_n3483_), .B(new_n30364_), .ZN(new_n30375_));
  NOR2_X1    g27119(.A1(new_n30370_), .A2(new_n9569_), .ZN(new_n30376_));
  NOR2_X1    g27120(.A1(new_n30370_), .A2(new_n6398_), .ZN(new_n30377_));
  NOR4_X1    g27121(.A1(new_n30376_), .A2(new_n30377_), .A3(pi0092), .A4(new_n3204_), .ZN(new_n30378_));
  OAI21_X1   g27122(.A1(new_n30375_), .A2(new_n30378_), .B(new_n30370_), .ZN(new_n30379_));
  OR3_X2     g27123(.A1(new_n30368_), .A2(new_n30374_), .A3(new_n30379_), .Z(new_n30380_));
  NOR2_X1    g27124(.A1(new_n3209_), .A2(pi0056), .ZN(new_n30381_));
  OAI21_X1   g27125(.A1(new_n8226_), .A2(new_n3426_), .B(new_n3201_), .ZN(new_n30383_));
  NAND2_X1   g27126(.A1(new_n30370_), .A2(new_n30383_), .ZN(new_n30384_));
  AOI21_X1   g27127(.A1(new_n30380_), .A2(new_n30381_), .B(new_n30384_), .ZN(po0382));
  INV_X1     g27128(.I(pi0231), .ZN(new_n30386_));
  NOR2_X1    g27129(.A1(new_n3005_), .A2(new_n30386_), .ZN(new_n30387_));
  INV_X1     g27130(.I(new_n30387_), .ZN(new_n30388_));
  NAND2_X1   g27131(.A1(new_n2694_), .A2(new_n2508_), .ZN(new_n30389_));
  OAI22_X1   g27132(.A1(new_n2858_), .A2(pi0070), .B1(new_n2692_), .B2(new_n2697_), .ZN(new_n30390_));
  NOR2_X1    g27133(.A1(new_n2807_), .A2(new_n30390_), .ZN(new_n30391_));
  NAND2_X1   g27134(.A1(new_n30389_), .A2(new_n30391_), .ZN(new_n30392_));
  NAND2_X1   g27135(.A1(new_n30392_), .A2(new_n3323_), .ZN(new_n30393_));
  NAND4_X1   g27136(.A1(new_n30393_), .A2(pi0038), .A3(pi0039), .A4(new_n5472_), .ZN(new_n30394_));
  NAND2_X1   g27137(.A1(new_n30393_), .A2(new_n5472_), .ZN(new_n30395_));
  NAND3_X1   g27138(.A1(new_n30395_), .A2(pi0039), .A3(new_n4368_), .ZN(new_n30396_));
  AOI21_X1   g27139(.A1(new_n30396_), .A2(new_n30394_), .B(new_n3145_), .ZN(new_n30397_));
  NAND3_X1   g27140(.A1(new_n30397_), .A2(pi0100), .A3(pi0228), .ZN(new_n30398_));
  INV_X1     g27141(.I(new_n30397_), .ZN(new_n30399_));
  NAND3_X1   g27142(.A1(new_n30399_), .A2(new_n3462_), .A3(pi0228), .ZN(new_n30400_));
  AOI21_X1   g27143(.A1(new_n6310_), .A2(new_n3171_), .B(new_n30388_), .ZN(new_n30401_));
  AOI21_X1   g27144(.A1(pi0100), .A2(new_n30387_), .B(new_n3411_), .ZN(new_n30402_));
  OAI21_X1   g27145(.A1(new_n30402_), .A2(new_n3212_), .B(new_n3455_), .ZN(new_n30403_));
  OAI21_X1   g27146(.A1(new_n30401_), .A2(new_n30403_), .B(pi0231), .ZN(new_n30404_));
  AOI21_X1   g27147(.A1(new_n30400_), .A2(new_n30398_), .B(new_n30404_), .ZN(new_n30405_));
  INV_X1     g27148(.I(new_n6312_), .ZN(new_n30406_));
  NOR2_X1    g27149(.A1(new_n30387_), .A2(new_n3303_), .ZN(new_n30407_));
  AOI21_X1   g27150(.A1(new_n30406_), .A2(new_n30407_), .B(pi0092), .ZN(new_n30408_));
  INV_X1     g27151(.I(new_n30408_), .ZN(new_n30409_));
  AOI21_X1   g27152(.A1(new_n10869_), .A2(new_n30388_), .B(new_n3235_), .ZN(new_n30410_));
  OAI21_X1   g27153(.A1(new_n30405_), .A2(new_n30409_), .B(new_n30410_), .ZN(new_n30411_));
  OR3_X2     g27154(.A1(new_n30411_), .A2(new_n3115_), .A3(new_n3175_), .Z(new_n30412_));
  NAND3_X1   g27155(.A1(new_n30411_), .A2(pi0054), .A3(new_n3175_), .ZN(new_n30413_));
  AOI21_X1   g27156(.A1(new_n30412_), .A2(new_n30413_), .B(new_n30388_), .ZN(new_n30414_));
  NAND2_X1   g27157(.A1(new_n3258_), .A2(pi0056), .ZN(new_n30415_));
  NAND2_X1   g27158(.A1(new_n30387_), .A2(pi0074), .ZN(new_n30416_));
  AOI21_X1   g27159(.A1(new_n3412_), .A2(new_n30416_), .B(new_n27651_), .ZN(new_n30417_));
  OAI21_X1   g27160(.A1(new_n30414_), .A2(new_n30415_), .B(new_n30417_), .ZN(new_n30418_));
  NAND2_X1   g27161(.A1(new_n30418_), .A2(new_n3201_), .ZN(new_n30419_));
  NOR3_X1    g27162(.A1(new_n6333_), .A2(new_n3219_), .A3(new_n30387_), .ZN(new_n30420_));
  NAND2_X1   g27163(.A1(new_n30388_), .A2(new_n3201_), .ZN(new_n30421_));
  AOI21_X1   g27164(.A1(new_n30419_), .A2(new_n30420_), .B(new_n30421_), .ZN(new_n30422_));
  NAND2_X1   g27165(.A1(new_n6331_), .A2(new_n3230_), .ZN(new_n30423_));
  OAI22_X1   g27166(.A1(new_n30422_), .A2(new_n30423_), .B1(new_n3230_), .B2(new_n30388_), .ZN(po0383));
  NOR2_X1    g27167(.A1(new_n5596_), .A2(new_n2481_), .ZN(new_n30425_));
  NAND2_X1   g27168(.A1(new_n8963_), .A2(new_n30425_), .ZN(new_n30426_));
  OAI21_X1   g27169(.A1(new_n2458_), .A2(new_n2490_), .B(new_n2672_), .ZN(new_n30427_));
  AOI21_X1   g27170(.A1(new_n30425_), .A2(new_n30427_), .B(pi0072), .ZN(new_n30428_));
  INV_X1     g27171(.I(new_n30428_), .ZN(new_n30429_));
  NAND3_X1   g27172(.A1(new_n8963_), .A2(pi1093), .A3(new_n30425_), .ZN(new_n30430_));
  NAND2_X1   g27173(.A1(new_n6402_), .A2(pi0829), .ZN(new_n30431_));
  AOI21_X1   g27174(.A1(new_n30430_), .A2(new_n30431_), .B(new_n30429_), .ZN(new_n30432_));
  AOI21_X1   g27175(.A1(new_n5561_), .A2(new_n2987_), .B(new_n30428_), .ZN(new_n30433_));
  NOR4_X1    g27176(.A1(new_n30432_), .A2(new_n5625_), .A3(new_n30426_), .A4(new_n30433_), .ZN(new_n30434_));
  AOI21_X1   g27177(.A1(new_n2480_), .A2(new_n6402_), .B(new_n5687_), .ZN(new_n30435_));
  AOI21_X1   g27178(.A1(new_n5625_), .A2(new_n30435_), .B(new_n10289_), .ZN(new_n30436_));
  OAI21_X1   g27179(.A1(new_n30434_), .A2(pi1093), .B(new_n30436_), .ZN(new_n30437_));
  AOI21_X1   g27180(.A1(new_n5561_), .A2(pi0072), .B(new_n30425_), .ZN(new_n30438_));
  INV_X1     g27181(.I(new_n30427_), .ZN(new_n30439_));
  NOR3_X1    g27182(.A1(new_n8970_), .A2(new_n2682_), .A3(new_n6403_), .ZN(new_n30440_));
  NOR2_X1    g27183(.A1(new_n8964_), .A2(new_n2981_), .ZN(new_n30441_));
  OAI21_X1   g27184(.A1(new_n30439_), .A2(new_n30440_), .B(new_n30441_), .ZN(new_n30442_));
  AOI21_X1   g27185(.A1(new_n2730_), .A2(pi1093), .B(new_n2721_), .ZN(new_n30443_));
  OAI21_X1   g27186(.A1(new_n30442_), .A2(new_n30438_), .B(new_n30443_), .ZN(new_n30444_));
  AOI21_X1   g27187(.A1(new_n30437_), .A2(new_n9273_), .B(new_n30444_), .ZN(po0384));
  NAND3_X1   g27188(.A1(new_n5461_), .A2(pi0039), .A3(new_n9241_), .ZN(new_n30446_));
  AOI21_X1   g27189(.A1(new_n30446_), .A2(new_n3384_), .B(new_n6272_), .ZN(new_n30447_));
  NOR2_X1    g27190(.A1(new_n5695_), .A2(new_n2726_), .ZN(new_n30448_));
  INV_X1     g27191(.I(new_n2893_), .ZN(new_n30449_));
  NAND3_X1   g27192(.A1(new_n2794_), .A2(new_n3183_), .A3(new_n2436_), .ZN(new_n30450_));
  NAND2_X1   g27193(.A1(new_n7293_), .A2(new_n2985_), .ZN(new_n30451_));
  AOI21_X1   g27194(.A1(new_n30449_), .A2(new_n30450_), .B(new_n30451_), .ZN(new_n30452_));
  AOI22_X1   g27195(.A1(new_n30452_), .A2(new_n30448_), .B1(new_n9291_), .B2(new_n30447_), .ZN(new_n30453_));
  OAI21_X1   g27196(.A1(new_n30453_), .A2(new_n3005_), .B(new_n9285_), .ZN(po0385));
  NOR2_X1    g27197(.A1(new_n13677_), .A2(new_n7611_), .ZN(new_n30455_));
  NAND3_X1   g27198(.A1(new_n12780_), .A2(pi1091), .A3(new_n5684_), .ZN(new_n30456_));
  NAND3_X1   g27199(.A1(new_n12782_), .A2(new_n2726_), .A3(new_n5684_), .ZN(new_n30457_));
  AOI21_X1   g27200(.A1(new_n30457_), .A2(new_n30456_), .B(new_n12801_), .ZN(new_n30458_));
  NOR2_X1    g27201(.A1(new_n30458_), .A2(new_n10925_), .ZN(new_n30459_));
  NAND2_X1   g27202(.A1(new_n12782_), .A2(pi1091), .ZN(new_n30460_));
  NOR3_X1    g27203(.A1(new_n6432_), .A2(new_n2726_), .A3(new_n5531_), .ZN(new_n30461_));
  XOR2_X1    g27204(.A1(new_n30460_), .A2(new_n30461_), .Z(new_n30462_));
  NOR4_X1    g27205(.A1(new_n30462_), .A2(new_n10925_), .A3(new_n3145_), .A4(new_n12801_), .ZN(new_n30463_));
  XNOR2_X1   g27206(.A1(new_n30463_), .A2(new_n30459_), .ZN(new_n30464_));
  AOI21_X1   g27207(.A1(new_n30464_), .A2(new_n7611_), .B(new_n30455_), .ZN(new_n30465_));
  NAND2_X1   g27208(.A1(new_n30465_), .A2(new_n5454_), .ZN(new_n30466_));
  XOR2_X1    g27209(.A1(new_n30466_), .A2(new_n13516_), .Z(new_n30467_));
  NOR2_X1    g27210(.A1(new_n5385_), .A2(pi0120), .ZN(new_n30468_));
  AOI21_X1   g27211(.A1(new_n13676_), .A2(new_n30468_), .B(new_n5438_), .ZN(new_n30469_));
  NAND2_X1   g27212(.A1(new_n5438_), .A2(new_n10925_), .ZN(new_n30470_));
  OAI21_X1   g27213(.A1(new_n13677_), .A2(new_n30470_), .B(new_n5434_), .ZN(new_n30471_));
  NAND2_X1   g27214(.A1(new_n30471_), .A2(pi0215), .ZN(new_n30472_));
  XOR2_X1    g27215(.A1(new_n30472_), .A2(new_n13309_), .Z(new_n30473_));
  NAND2_X1   g27216(.A1(new_n30473_), .A2(new_n30469_), .ZN(new_n30474_));
  NAND2_X1   g27217(.A1(new_n30474_), .A2(new_n3098_), .ZN(new_n30475_));
  NAND2_X1   g27218(.A1(new_n30464_), .A2(new_n5385_), .ZN(new_n30476_));
  OAI21_X1   g27219(.A1(new_n5385_), .A2(new_n13677_), .B(new_n30476_), .ZN(new_n30477_));
  NAND2_X1   g27220(.A1(new_n13677_), .A2(new_n3312_), .ZN(new_n30478_));
  NAND4_X1   g27221(.A1(new_n30477_), .A2(new_n3111_), .A3(new_n30475_), .A4(new_n30478_), .ZN(new_n30479_));
  NAND2_X1   g27222(.A1(new_n30471_), .A2(pi0223), .ZN(new_n30480_));
  XOR2_X1    g27223(.A1(new_n30480_), .A2(new_n13466_), .Z(new_n30481_));
  AOI21_X1   g27224(.A1(new_n30481_), .A2(new_n30469_), .B(pi0299), .ZN(new_n30482_));
  OAI21_X1   g27225(.A1(new_n30467_), .A2(new_n30479_), .B(new_n30482_), .ZN(new_n30483_));
  NAND2_X1   g27226(.A1(new_n30465_), .A2(new_n5398_), .ZN(new_n30484_));
  XOR2_X1    g27227(.A1(new_n30484_), .A2(new_n12982_), .Z(new_n30485_));
  NAND2_X1   g27228(.A1(new_n30485_), .A2(new_n30477_), .ZN(new_n30486_));
  NAND2_X1   g27229(.A1(new_n30486_), .A2(new_n3090_), .ZN(new_n30487_));
  OAI21_X1   g27230(.A1(new_n13013_), .A2(new_n5683_), .B(new_n2794_), .ZN(new_n30488_));
  NAND3_X1   g27231(.A1(new_n13128_), .A2(new_n13129_), .A3(new_n30488_), .ZN(new_n30489_));
  NOR2_X1    g27232(.A1(pi0829), .A2(pi1091), .ZN(new_n30490_));
  AND2_X2    g27233(.A1(new_n30489_), .A2(new_n30490_), .Z(new_n30491_));
  AND2_X2    g27234(.A1(new_n13034_), .A2(new_n13033_), .Z(new_n30492_));
  AOI21_X1   g27235(.A1(new_n5683_), .A2(new_n30490_), .B(new_n13013_), .ZN(new_n30493_));
  OAI21_X1   g27236(.A1(new_n30492_), .A2(pi0032), .B(new_n30493_), .ZN(new_n30494_));
  AOI21_X1   g27237(.A1(new_n5469_), .A2(new_n5691_), .B(new_n2980_), .ZN(new_n30495_));
  NOR3_X1    g27238(.A1(new_n30491_), .A2(new_n30494_), .A3(new_n30495_), .ZN(new_n30496_));
  OAI22_X1   g27239(.A1(new_n13041_), .A2(new_n6402_), .B1(new_n13006_), .B2(new_n13058_), .ZN(new_n30497_));
  AND3_X2    g27240(.A1(new_n30497_), .A2(new_n2984_), .A3(new_n5468_), .Z(new_n30498_));
  INV_X1     g27241(.I(new_n13028_), .ZN(new_n30499_));
  NAND3_X1   g27242(.A1(new_n12996_), .A2(new_n2486_), .A3(new_n5464_), .ZN(new_n30500_));
  AOI21_X1   g27243(.A1(new_n30499_), .A2(new_n30500_), .B(new_n8380_), .ZN(new_n30501_));
  NOR2_X1    g27244(.A1(new_n5532_), .A2(pi1093), .ZN(new_n30502_));
  OAI21_X1   g27245(.A1(new_n30501_), .A2(new_n3721_), .B(new_n30502_), .ZN(new_n30503_));
  NOR2_X1    g27246(.A1(new_n13033_), .A2(new_n3183_), .ZN(new_n30504_));
  AOI21_X1   g27247(.A1(new_n30503_), .A2(new_n30504_), .B(new_n13053_), .ZN(new_n30505_));
  NOR4_X1    g27248(.A1(new_n30498_), .A2(new_n5533_), .A3(new_n5692_), .A4(new_n30505_), .ZN(new_n30506_));
  NOR2_X1    g27249(.A1(new_n13053_), .A2(new_n5691_), .ZN(new_n30507_));
  AOI21_X1   g27250(.A1(new_n30494_), .A2(new_n30507_), .B(new_n30489_), .ZN(new_n30508_));
  OAI21_X1   g27251(.A1(new_n30506_), .A2(new_n30496_), .B(new_n30508_), .ZN(new_n30509_));
  NAND2_X1   g27252(.A1(new_n30509_), .A2(new_n3259_), .ZN(new_n30510_));
  NOR3_X1    g27253(.A1(new_n13676_), .A2(new_n3183_), .A3(new_n3092_), .ZN(new_n30511_));
  NAND4_X1   g27254(.A1(new_n30487_), .A2(new_n30483_), .A3(new_n30510_), .A4(new_n30511_), .ZN(new_n30512_));
  AOI21_X1   g27255(.A1(new_n30512_), .A2(new_n8345_), .B(new_n6281_), .ZN(po0387));
  NOR2_X1    g27256(.A1(new_n5507_), .A2(new_n3455_), .ZN(new_n30514_));
  INV_X1     g27257(.I(new_n2524_), .ZN(new_n30515_));
  NOR2_X1    g27258(.A1(new_n2647_), .A2(new_n2492_), .ZN(new_n30516_));
  XOR2_X1    g27259(.A1(new_n30516_), .A2(new_n2563_), .Z(new_n30517_));
  AOI21_X1   g27260(.A1(new_n2555_), .A2(new_n12074_), .B(new_n2513_), .ZN(new_n30518_));
  AOI21_X1   g27261(.A1(new_n2861_), .A2(new_n2859_), .B(new_n2552_), .ZN(new_n30519_));
  NOR4_X1    g27262(.A1(new_n30519_), .A2(new_n30518_), .A3(new_n2453_), .A4(new_n2862_), .ZN(new_n30520_));
  AOI21_X1   g27263(.A1(new_n30517_), .A2(new_n30520_), .B(new_n2528_), .ZN(new_n30521_));
  OR4_X2     g27264(.A1(new_n30515_), .A2(new_n30521_), .A3(new_n2689_), .A4(new_n2878_), .Z(new_n30522_));
  NOR2_X1    g27265(.A1(new_n30522_), .A2(new_n2692_), .ZN(new_n30523_));
  XOR2_X1    g27266(.A1(new_n30522_), .A2(new_n5606_), .Z(new_n30524_));
  NAND2_X1   g27267(.A1(new_n30524_), .A2(new_n2508_), .ZN(new_n30525_));
  OAI21_X1   g27268(.A1(new_n30525_), .A2(new_n30523_), .B(pi0070), .ZN(new_n30526_));
  AOI21_X1   g27269(.A1(new_n30523_), .A2(new_n30525_), .B(new_n30526_), .ZN(new_n30527_));
  XOR2_X1    g27270(.A1(new_n30527_), .A2(new_n9238_), .Z(new_n30528_));
  NOR3_X1    g27271(.A1(new_n2485_), .A2(pi0072), .A3(new_n2805_), .ZN(new_n30529_));
  OAI21_X1   g27272(.A1(new_n30529_), .A2(new_n2713_), .B(new_n2715_), .ZN(new_n30530_));
  OAI21_X1   g27273(.A1(new_n30528_), .A2(new_n30530_), .B(pi0032), .ZN(new_n30531_));
  NAND3_X1   g27274(.A1(new_n2502_), .A2(pi0032), .A3(new_n8320_), .ZN(new_n30532_));
  NOR2_X1    g27275(.A1(new_n2773_), .A2(new_n30532_), .ZN(new_n30533_));
  NOR2_X1    g27276(.A1(new_n30531_), .A2(new_n30533_), .ZN(new_n30534_));
  NAND2_X1   g27277(.A1(new_n30531_), .A2(new_n30533_), .ZN(new_n30535_));
  NAND2_X1   g27278(.A1(new_n30535_), .A2(new_n2436_), .ZN(new_n30536_));
  OAI21_X1   g27279(.A1(new_n30536_), .A2(new_n30534_), .B(new_n2793_), .ZN(new_n30537_));
  NAND2_X1   g27280(.A1(new_n30537_), .A2(pi0039), .ZN(new_n30538_));
  NOR2_X1    g27281(.A1(new_n6272_), .A2(pi0299), .ZN(new_n30539_));
  AOI21_X1   g27282(.A1(new_n5461_), .A2(pi0299), .B(new_n30539_), .ZN(new_n30540_));
  NOR2_X1    g27283(.A1(new_n5436_), .A2(new_n2981_), .ZN(new_n30541_));
  NAND4_X1   g27284(.A1(new_n9205_), .A2(pi0039), .A3(pi0287), .A4(pi0835), .ZN(new_n30542_));
  NOR4_X1    g27285(.A1(new_n30540_), .A2(new_n5408_), .A3(new_n30541_), .A4(new_n30542_), .ZN(new_n30543_));
  XNOR2_X1   g27286(.A1(new_n30538_), .A2(new_n30543_), .ZN(new_n30544_));
  NAND4_X1   g27287(.A1(new_n30544_), .A2(pi0038), .A3(pi0100), .A4(new_n3160_), .ZN(new_n30545_));
  NAND2_X1   g27288(.A1(new_n30544_), .A2(new_n3160_), .ZN(new_n30546_));
  NAND3_X1   g27289(.A1(new_n30546_), .A2(pi0038), .A3(new_n3462_), .ZN(new_n30547_));
  NAND2_X1   g27290(.A1(new_n30547_), .A2(new_n30545_), .ZN(new_n30548_));
  NAND4_X1   g27291(.A1(new_n30548_), .A2(pi0087), .A3(new_n5488_), .A4(new_n5492_), .ZN(new_n30549_));
  NAND2_X1   g27292(.A1(new_n30549_), .A2(new_n30514_), .ZN(new_n30550_));
  NOR2_X1    g27293(.A1(new_n30549_), .A2(new_n30514_), .ZN(new_n30551_));
  NOR2_X1    g27294(.A1(new_n30551_), .A2(new_n3189_), .ZN(new_n30552_));
  AOI21_X1   g27295(.A1(new_n30552_), .A2(new_n30550_), .B(new_n6291_), .ZN(new_n30553_));
  NOR3_X1    g27296(.A1(new_n5497_), .A2(new_n12144_), .A3(new_n6297_), .ZN(new_n30554_));
  OAI21_X1   g27297(.A1(new_n30553_), .A2(pi0054), .B(new_n30554_), .ZN(new_n30555_));
  AOI21_X1   g27298(.A1(new_n30555_), .A2(new_n12147_), .B(new_n5544_), .ZN(po0389));
  INV_X1     g27299(.I(pi0230), .ZN(new_n30557_));
  NOR2_X1    g27300(.A1(new_n8684_), .A2(pi1143), .ZN(new_n30558_));
  NOR2_X1    g27301(.A1(pi0211), .A2(pi1144), .ZN(new_n30559_));
  NOR2_X1    g27302(.A1(new_n30558_), .A2(new_n30559_), .ZN(new_n30560_));
  INV_X1     g27303(.I(new_n30560_), .ZN(new_n30561_));
  NOR2_X1    g27304(.A1(new_n30561_), .A2(new_n3098_), .ZN(new_n30562_));
  AOI21_X1   g27305(.A1(pi0199), .A2(pi1142), .B(pi0200), .ZN(new_n30563_));
  AOI21_X1   g27306(.A1(new_n8549_), .A2(pi1143), .B(new_n8555_), .ZN(new_n30564_));
  NAND2_X1   g27307(.A1(new_n30564_), .A2(new_n30563_), .ZN(new_n30565_));
  AOI21_X1   g27308(.A1(new_n30565_), .A2(new_n3057_), .B(new_n8549_), .ZN(new_n30566_));
  INV_X1     g27309(.I(new_n30566_), .ZN(new_n30567_));
  NOR2_X1    g27310(.A1(new_n8545_), .A2(pi0299), .ZN(new_n30568_));
  AOI21_X1   g27311(.A1(new_n30568_), .A2(pi0200), .B(pi1142), .ZN(new_n30569_));
  INV_X1     g27312(.I(new_n30569_), .ZN(new_n30570_));
  INV_X1     g27313(.I(new_n30563_), .ZN(new_n30571_));
  NOR2_X1    g27314(.A1(new_n30571_), .A2(new_n8549_), .ZN(new_n30572_));
  AOI21_X1   g27315(.A1(new_n30570_), .A2(new_n30572_), .B(pi1143), .ZN(new_n30573_));
  INV_X1     g27316(.I(new_n30573_), .ZN(new_n30574_));
  NOR2_X1    g27317(.A1(new_n8549_), .A2(new_n8545_), .ZN(new_n30575_));
  AOI21_X1   g27318(.A1(new_n30574_), .A2(new_n30575_), .B(pi0299), .ZN(new_n30576_));
  NOR4_X1    g27319(.A1(new_n30576_), .A2(new_n8545_), .A3(new_n8546_), .A4(new_n30567_), .ZN(new_n30577_));
  NAND2_X1   g27320(.A1(new_n30566_), .A2(new_n8547_), .ZN(new_n30578_));
  NOR2_X1    g27321(.A1(new_n30576_), .A2(new_n30578_), .ZN(new_n30579_));
  NOR3_X1    g27322(.A1(new_n30579_), .A2(new_n8546_), .A3(new_n30566_), .ZN(new_n30580_));
  NOR2_X1    g27323(.A1(new_n30580_), .A2(new_n30577_), .ZN(new_n30581_));
  NAND2_X1   g27324(.A1(new_n30581_), .A2(new_n3098_), .ZN(new_n30582_));
  OAI21_X1   g27325(.A1(new_n30582_), .A2(new_n8739_), .B(new_n8685_), .ZN(new_n30583_));
  AND2_X2    g27326(.A1(new_n30583_), .A2(new_n30562_), .Z(new_n30584_));
  INV_X1     g27327(.I(new_n30582_), .ZN(new_n30585_));
  NOR2_X1    g27328(.A1(pi0212), .A2(pi0214), .ZN(new_n30586_));
  NOR2_X1    g27329(.A1(new_n3098_), .A2(pi1142), .ZN(new_n30587_));
  NOR2_X1    g27330(.A1(new_n8684_), .A2(new_n3098_), .ZN(new_n30588_));
  XOR2_X1    g27331(.A1(new_n30588_), .A2(new_n30587_), .Z(new_n30589_));
  NAND2_X1   g27332(.A1(new_n30589_), .A2(pi1143), .ZN(new_n30590_));
  OAI21_X1   g27333(.A1(new_n30561_), .A2(new_n3098_), .B(new_n8685_), .ZN(new_n30591_));
  NOR4_X1    g27334(.A1(new_n30585_), .A2(new_n30586_), .A3(new_n30590_), .A4(new_n30591_), .ZN(new_n30592_));
  OAI21_X1   g27335(.A1(new_n30584_), .A2(pi0219), .B(new_n30592_), .ZN(new_n30593_));
  NOR2_X1    g27336(.A1(new_n30586_), .A2(pi0211), .ZN(new_n30594_));
  NOR2_X1    g27337(.A1(new_n30594_), .A2(new_n8683_), .ZN(new_n30595_));
  NOR2_X1    g27338(.A1(new_n7240_), .A2(new_n30595_), .ZN(new_n30596_));
  INV_X1     g27339(.I(new_n8740_), .ZN(new_n30597_));
  NOR3_X1    g27340(.A1(new_n30597_), .A2(pi0211), .A3(new_n3650_), .ZN(new_n30599_));
  AOI21_X1   g27341(.A1(new_n30596_), .A2(new_n30599_), .B(pi1142), .ZN(new_n30600_));
  NOR2_X1    g27342(.A1(new_n30600_), .A2(new_n8688_), .ZN(new_n30601_));
  NOR2_X1    g27343(.A1(new_n30601_), .A2(po1038), .ZN(new_n30602_));
  NAND2_X1   g27344(.A1(new_n30581_), .A2(new_n30594_), .ZN(new_n30603_));
  INV_X1     g27345(.I(new_n30594_), .ZN(new_n30604_));
  NOR2_X1    g27346(.A1(new_n30604_), .A2(new_n3098_), .ZN(new_n30605_));
  XOR2_X1    g27347(.A1(new_n30603_), .A2(new_n30605_), .Z(new_n30606_));
  OAI21_X1   g27348(.A1(new_n30606_), .A2(new_n3814_), .B(new_n8683_), .ZN(new_n30607_));
  NAND3_X1   g27349(.A1(new_n30607_), .A2(new_n30585_), .A3(new_n30594_), .ZN(new_n30608_));
  AOI21_X1   g27350(.A1(new_n30593_), .A2(new_n30602_), .B(new_n30608_), .ZN(new_n30609_));
  NOR2_X1    g27351(.A1(new_n3098_), .A2(new_n13778_), .ZN(new_n30610_));
  INV_X1     g27352(.I(new_n30610_), .ZN(new_n30611_));
  NOR2_X1    g27353(.A1(new_n3098_), .A2(new_n13614_), .ZN(new_n30612_));
  NOR2_X1    g27354(.A1(new_n3098_), .A2(new_n13817_), .ZN(new_n30613_));
  INV_X1     g27355(.I(new_n30613_), .ZN(new_n30614_));
  NOR2_X1    g27356(.A1(new_n8683_), .A2(pi0211), .ZN(new_n30615_));
  INV_X1     g27357(.I(new_n30615_), .ZN(new_n30616_));
  NOR2_X1    g27358(.A1(new_n30614_), .A2(new_n30616_), .ZN(new_n30617_));
  NOR3_X1    g27359(.A1(new_n30611_), .A2(pi0212), .A3(new_n8685_), .ZN(new_n30618_));
  NOR2_X1    g27360(.A1(new_n3098_), .A2(pi0219), .ZN(new_n30619_));
  INV_X1     g27361(.I(new_n30619_), .ZN(new_n30620_));
  NOR2_X1    g27362(.A1(new_n8684_), .A2(new_n13969_), .ZN(new_n30621_));
  NOR2_X1    g27363(.A1(new_n14006_), .A2(pi0211), .ZN(new_n30622_));
  NOR2_X1    g27364(.A1(new_n30621_), .A2(new_n30622_), .ZN(new_n30623_));
  NOR2_X1    g27365(.A1(new_n30623_), .A2(new_n8685_), .ZN(new_n30624_));
  NOR2_X1    g27366(.A1(new_n13969_), .A2(pi0211), .ZN(new_n30625_));
  NOR2_X1    g27367(.A1(new_n30625_), .A2(new_n8685_), .ZN(new_n30626_));
  INV_X1     g27368(.I(new_n30626_), .ZN(new_n30627_));
  NOR4_X1    g27369(.A1(new_n8684_), .A2(new_n8685_), .A3(new_n13778_), .A4(pi1154), .ZN(new_n30628_));
  AOI21_X1   g27370(.A1(new_n30627_), .A2(new_n30628_), .B(new_n8739_), .ZN(new_n30629_));
  OAI21_X1   g27371(.A1(new_n30627_), .A2(new_n30628_), .B(new_n30629_), .ZN(new_n30630_));
  INV_X1     g27372(.I(new_n30630_), .ZN(new_n30631_));
  AOI21_X1   g27373(.A1(new_n8739_), .A2(new_n30624_), .B(new_n30631_), .ZN(new_n30632_));
  NOR2_X1    g27374(.A1(new_n30632_), .A2(new_n30620_), .ZN(new_n30633_));
  INV_X1     g27375(.I(new_n30632_), .ZN(new_n30634_));
  NOR2_X1    g27376(.A1(new_n13614_), .A2(pi0211), .ZN(new_n30635_));
  NOR2_X1    g27377(.A1(new_n30635_), .A2(new_n8685_), .ZN(new_n30636_));
  NOR2_X1    g27378(.A1(new_n13817_), .A2(pi0211), .ZN(new_n30637_));
  NAND2_X1   g27379(.A1(new_n8740_), .A2(new_n30637_), .ZN(new_n30638_));
  XNOR2_X1   g27380(.A1(new_n30638_), .A2(new_n30636_), .ZN(new_n30639_));
  NOR2_X1    g27381(.A1(new_n8685_), .A2(pi0211), .ZN(new_n30640_));
  NAND2_X1   g27382(.A1(new_n8739_), .A2(pi0213), .ZN(new_n30641_));
  AOI21_X1   g27383(.A1(pi1155), .A2(new_n30640_), .B(new_n30641_), .ZN(new_n30642_));
  OAI21_X1   g27384(.A1(new_n9213_), .A2(new_n30639_), .B(new_n30642_), .ZN(new_n30643_));
  NAND2_X1   g27385(.A1(new_n30643_), .A2(new_n8683_), .ZN(new_n30644_));
  NAND2_X1   g27386(.A1(new_n30634_), .A2(new_n30644_), .ZN(new_n30645_));
  OAI22_X1   g27387(.A1(new_n30645_), .A2(new_n7240_), .B1(new_n30618_), .B2(new_n30633_), .ZN(new_n30646_));
  NAND2_X1   g27388(.A1(new_n30585_), .A2(new_n30646_), .ZN(new_n30647_));
  AOI21_X1   g27389(.A1(new_n30647_), .A2(new_n28364_), .B(new_n28529_), .ZN(new_n30648_));
  AOI21_X1   g27390(.A1(new_n30609_), .A2(new_n30648_), .B(new_n30557_), .ZN(new_n30649_));
  NOR2_X1    g27391(.A1(new_n8555_), .A2(pi0199), .ZN(new_n30650_));
  NOR2_X1    g27392(.A1(new_n8549_), .A2(pi0200), .ZN(new_n30651_));
  NOR2_X1    g27393(.A1(new_n30650_), .A2(new_n30651_), .ZN(new_n30652_));
  NOR2_X1    g27394(.A1(new_n30652_), .A2(pi0299), .ZN(new_n30653_));
  INV_X1     g27395(.I(new_n30653_), .ZN(new_n30654_));
  NOR2_X1    g27396(.A1(new_n8549_), .A2(pi1153), .ZN(new_n30655_));
  NOR2_X1    g27397(.A1(new_n30654_), .A2(new_n30655_), .ZN(new_n30656_));
  NOR2_X1    g27398(.A1(new_n9214_), .A2(new_n13778_), .ZN(new_n30657_));
  NOR2_X1    g27399(.A1(new_n30656_), .A2(new_n30657_), .ZN(new_n30658_));
  NOR2_X1    g27400(.A1(pi0200), .A2(pi0299), .ZN(new_n30659_));
  OAI21_X1   g27401(.A1(new_n8549_), .A2(pi1153), .B(new_n30659_), .ZN(new_n30660_));
  NAND2_X1   g27402(.A1(pi0199), .A2(pi1155), .ZN(new_n30661_));
  AOI21_X1   g27403(.A1(new_n30660_), .A2(new_n13817_), .B(new_n30661_), .ZN(new_n30662_));
  AOI21_X1   g27404(.A1(pi1154), .A2(new_n30662_), .B(new_n30658_), .ZN(new_n30663_));
  NOR2_X1    g27405(.A1(new_n30663_), .A2(new_n3098_), .ZN(new_n30664_));
  INV_X1     g27406(.I(new_n30664_), .ZN(new_n30665_));
  NOR2_X1    g27407(.A1(new_n30651_), .A2(pi0299), .ZN(new_n30666_));
  NOR2_X1    g27408(.A1(new_n30666_), .A2(pi1155), .ZN(new_n30667_));
  INV_X1     g27409(.I(new_n30652_), .ZN(new_n30668_));
  NOR2_X1    g27410(.A1(new_n30668_), .A2(pi0299), .ZN(new_n30669_));
  INV_X1     g27411(.I(new_n30669_), .ZN(new_n30670_));
  AOI21_X1   g27412(.A1(new_n30670_), .A2(pi1155), .B(new_n30667_), .ZN(new_n30671_));
  NOR2_X1    g27413(.A1(new_n30671_), .A2(new_n13817_), .ZN(new_n30672_));
  NOR2_X1    g27414(.A1(new_n8555_), .A2(pi0299), .ZN(new_n30673_));
  INV_X1     g27415(.I(new_n30673_), .ZN(new_n30674_));
  NOR2_X1    g27416(.A1(new_n13778_), .A2(pi0199), .ZN(new_n30675_));
  INV_X1     g27417(.I(new_n30675_), .ZN(new_n30676_));
  NOR2_X1    g27418(.A1(new_n30674_), .A2(new_n30676_), .ZN(new_n30677_));
  NOR2_X1    g27419(.A1(new_n30677_), .A2(pi1154), .ZN(new_n30678_));
  INV_X1     g27420(.I(new_n30678_), .ZN(new_n30679_));
  NOR2_X1    g27421(.A1(new_n8555_), .A2(pi1155), .ZN(new_n30680_));
  NOR2_X1    g27422(.A1(new_n9209_), .A2(new_n30680_), .ZN(new_n30681_));
  INV_X1     g27423(.I(new_n30681_), .ZN(new_n30682_));
  NOR2_X1    g27424(.A1(new_n30682_), .A2(new_n13969_), .ZN(new_n30683_));
  INV_X1     g27425(.I(new_n30683_), .ZN(new_n30684_));
  NOR2_X1    g27426(.A1(new_n30675_), .A2(new_n8555_), .ZN(new_n30685_));
  NOR2_X1    g27427(.A1(new_n30685_), .A2(new_n8774_), .ZN(new_n30686_));
  AOI21_X1   g27428(.A1(new_n30684_), .A2(new_n30686_), .B(new_n30679_), .ZN(new_n30687_));
  INV_X1     g27429(.I(new_n30687_), .ZN(new_n30688_));
  OAI21_X1   g27430(.A1(new_n30688_), .A2(new_n30672_), .B(pi0208), .ZN(new_n30689_));
  XOR2_X1    g27431(.A1(new_n30689_), .A2(new_n8547_), .Z(new_n30690_));
  OR2_X2     g27432(.A1(new_n30690_), .A2(new_n30665_), .Z(new_n30691_));
  NOR2_X1    g27433(.A1(pi0207), .A2(pi0299), .ZN(new_n30692_));
  NOR2_X1    g27434(.A1(new_n30692_), .A2(pi0208), .ZN(new_n30693_));
  INV_X1     g27435(.I(new_n30693_), .ZN(new_n30694_));
  NOR2_X1    g27436(.A1(new_n8775_), .A2(pi1155), .ZN(new_n30695_));
  AOI21_X1   g27437(.A1(pi1155), .A2(new_n30673_), .B(new_n30695_), .ZN(new_n30696_));
  NOR2_X1    g27438(.A1(new_n30696_), .A2(pi1156), .ZN(new_n30697_));
  INV_X1     g27439(.I(new_n9214_), .ZN(new_n30698_));
  NOR2_X1    g27440(.A1(new_n13778_), .A2(pi0200), .ZN(new_n30699_));
  NOR2_X1    g27441(.A1(new_n30698_), .A2(new_n30699_), .ZN(new_n30700_));
  INV_X1     g27442(.I(new_n30700_), .ZN(new_n30701_));
  NOR2_X1    g27443(.A1(new_n30701_), .A2(new_n13969_), .ZN(new_n30702_));
  NOR2_X1    g27444(.A1(new_n30697_), .A2(new_n30702_), .ZN(new_n30703_));
  INV_X1     g27445(.I(new_n30703_), .ZN(new_n30704_));
  AOI21_X1   g27446(.A1(new_n30704_), .A2(pi0207), .B(new_n30694_), .ZN(new_n30705_));
  NAND2_X1   g27447(.A1(new_n13817_), .A2(pi0299), .ZN(new_n30706_));
  NAND3_X1   g27448(.A1(new_n30705_), .A2(pi1157), .A3(new_n30706_), .ZN(new_n30707_));
  INV_X1     g27449(.I(new_n30699_), .ZN(new_n30708_));
  NOR2_X1    g27450(.A1(new_n30708_), .A2(new_n8549_), .ZN(new_n30709_));
  AOI21_X1   g27451(.A1(new_n30709_), .A2(new_n3098_), .B(pi1156), .ZN(new_n30710_));
  INV_X1     g27452(.I(new_n30710_), .ZN(new_n30711_));
  NAND2_X1   g27453(.A1(pi0200), .A2(pi1155), .ZN(new_n30712_));
  AOI21_X1   g27454(.A1(new_n30711_), .A2(new_n30654_), .B(new_n30712_), .ZN(new_n30713_));
  NOR2_X1    g27455(.A1(new_n30614_), .A2(new_n8546_), .ZN(new_n30714_));
  OAI21_X1   g27456(.A1(pi0207), .A2(new_n30714_), .B(new_n30713_), .ZN(new_n30715_));
  OR2_X2     g27457(.A1(new_n30715_), .A2(new_n14006_), .Z(new_n30716_));
  AOI21_X1   g27458(.A1(new_n30691_), .A2(new_n30707_), .B(new_n30716_), .ZN(new_n30717_));
  INV_X1     g27459(.I(new_n8686_), .ZN(new_n30718_));
  AOI21_X1   g27460(.A1(new_n30668_), .A2(pi1154), .B(pi1153), .ZN(new_n30719_));
  OAI22_X1   g27461(.A1(new_n30719_), .A2(new_n30708_), .B1(new_n13614_), .B2(new_n9209_), .ZN(new_n30720_));
  INV_X1     g27462(.I(new_n30720_), .ZN(new_n30721_));
  NOR2_X1    g27463(.A1(new_n8549_), .A2(new_n8555_), .ZN(new_n30722_));
  NOR2_X1    g27464(.A1(new_n30722_), .A2(pi0299), .ZN(new_n30723_));
  NOR2_X1    g27465(.A1(new_n30723_), .A2(new_n13614_), .ZN(new_n30724_));
  NOR3_X1    g27466(.A1(new_n30724_), .A2(new_n30662_), .A3(pi1154), .ZN(new_n30725_));
  NOR2_X1    g27467(.A1(new_n30721_), .A2(new_n30725_), .ZN(new_n30726_));
  AOI21_X1   g27468(.A1(pi1155), .A2(new_n9214_), .B(new_n30695_), .ZN(new_n30727_));
  INV_X1     g27469(.I(new_n30727_), .ZN(new_n30728_));
  NOR2_X1    g27470(.A1(new_n30728_), .A2(new_n13969_), .ZN(new_n30729_));
  INV_X1     g27471(.I(new_n30729_), .ZN(new_n30730_));
  AOI21_X1   g27472(.A1(new_n30730_), .A2(new_n30686_), .B(new_n30679_), .ZN(new_n30731_));
  INV_X1     g27473(.I(new_n30731_), .ZN(new_n30732_));
  NOR2_X1    g27474(.A1(new_n3098_), .A2(new_n13969_), .ZN(new_n30733_));
  OAI21_X1   g27475(.A1(new_n30732_), .A2(new_n8546_), .B(new_n8545_), .ZN(new_n30734_));
  INV_X1     g27476(.I(new_n30659_), .ZN(new_n30735_));
  NOR2_X1    g27477(.A1(new_n8549_), .A2(pi1155), .ZN(new_n30736_));
  NAND3_X1   g27478(.A1(new_n30723_), .A2(pi1156), .A3(new_n30736_), .ZN(new_n30737_));
  INV_X1     g27479(.I(new_n30723_), .ZN(new_n30738_));
  INV_X1     g27480(.I(new_n30736_), .ZN(new_n30739_));
  NAND3_X1   g27481(.A1(new_n30738_), .A2(pi1156), .A3(new_n30739_), .ZN(new_n30740_));
  AOI21_X1   g27482(.A1(new_n30740_), .A2(new_n30737_), .B(new_n30735_), .ZN(new_n30741_));
  INV_X1     g27483(.I(new_n30741_), .ZN(new_n30742_));
  INV_X1     g27484(.I(new_n30733_), .ZN(new_n30743_));
  NOR2_X1    g27485(.A1(new_n14006_), .A2(pi0208), .ZN(new_n30744_));
  INV_X1     g27486(.I(new_n30744_), .ZN(new_n30745_));
  NOR2_X1    g27487(.A1(new_n30743_), .A2(new_n30745_), .ZN(new_n30746_));
  INV_X1     g27488(.I(new_n30746_), .ZN(new_n30747_));
  AOI21_X1   g27489(.A1(new_n8545_), .A2(new_n30747_), .B(new_n30742_), .ZN(new_n30748_));
  AOI21_X1   g27490(.A1(new_n30734_), .A2(new_n30726_), .B(new_n30748_), .ZN(new_n30749_));
  NOR2_X1    g27491(.A1(new_n30650_), .A2(pi0299), .ZN(new_n30750_));
  INV_X1     g27492(.I(new_n30750_), .ZN(new_n30751_));
  OAI21_X1   g27493(.A1(new_n30709_), .A2(new_n30750_), .B(pi0299), .ZN(new_n30752_));
  OAI21_X1   g27494(.A1(new_n13969_), .A2(new_n30751_), .B(new_n30752_), .ZN(new_n30753_));
  INV_X1     g27495(.I(new_n30753_), .ZN(new_n30754_));
  NOR2_X1    g27496(.A1(new_n8546_), .A2(new_n3098_), .ZN(new_n30755_));
  INV_X1     g27497(.I(new_n30755_), .ZN(new_n30756_));
  AOI21_X1   g27498(.A1(new_n30754_), .A2(new_n30756_), .B(new_n8545_), .ZN(new_n30757_));
  INV_X1     g27499(.I(new_n30757_), .ZN(new_n30758_));
  NOR3_X1    g27500(.A1(new_n30749_), .A2(new_n30711_), .A3(new_n30758_), .ZN(new_n30759_));
  NAND2_X1   g27501(.A1(new_n30759_), .A2(pi0211), .ZN(new_n30760_));
  NOR2_X1    g27502(.A1(new_n30610_), .A2(pi0207), .ZN(new_n30761_));
  NOR2_X1    g27503(.A1(new_n30761_), .A2(pi0208), .ZN(new_n30762_));
  AOI21_X1   g27504(.A1(new_n30687_), .A2(new_n30761_), .B(pi0208), .ZN(new_n30763_));
  NOR2_X1    g27505(.A1(new_n30674_), .A2(new_n13614_), .ZN(new_n30764_));
  AOI21_X1   g27506(.A1(new_n13614_), .A2(new_n8774_), .B(new_n30764_), .ZN(new_n30765_));
  AOI21_X1   g27507(.A1(new_n30765_), .A2(pi1155), .B(new_n13817_), .ZN(new_n30766_));
  NAND2_X1   g27508(.A1(pi0200), .A2(pi1153), .ZN(new_n30767_));
  NOR2_X1    g27509(.A1(new_n13817_), .A2(new_n13778_), .ZN(new_n30768_));
  INV_X1     g27510(.I(new_n30768_), .ZN(new_n30769_));
  NOR3_X1    g27511(.A1(new_n30769_), .A2(new_n30698_), .A3(new_n30767_), .ZN(new_n30770_));
  NAND2_X1   g27512(.A1(new_n30658_), .A2(new_n30770_), .ZN(new_n30771_));
  XOR2_X1    g27513(.A1(new_n30771_), .A2(new_n30766_), .Z(new_n30772_));
  INV_X1     g27514(.I(new_n30772_), .ZN(new_n30773_));
  NAND2_X1   g27515(.A1(new_n30773_), .A2(pi0207), .ZN(new_n30774_));
  NOR2_X1    g27516(.A1(new_n30667_), .A2(new_n13969_), .ZN(new_n30775_));
  NAND2_X1   g27517(.A1(new_n30674_), .A2(pi1155), .ZN(new_n30776_));
  NAND4_X1   g27518(.A1(new_n30776_), .A2(pi1156), .A3(new_n9209_), .A4(new_n30673_), .ZN(new_n30777_));
  XOR2_X1    g27519(.A1(new_n30777_), .A2(new_n30775_), .Z(new_n30778_));
  INV_X1     g27520(.I(new_n30778_), .ZN(new_n30779_));
  AOI21_X1   g27521(.A1(pi0208), .A2(new_n14006_), .B(new_n8545_), .ZN(new_n30780_));
  NAND2_X1   g27522(.A1(new_n30779_), .A2(new_n30780_), .ZN(new_n30781_));
  OAI21_X1   g27523(.A1(new_n30774_), .A2(new_n30763_), .B(new_n30781_), .ZN(new_n30782_));
  NOR2_X1    g27524(.A1(new_n9208_), .A2(pi1155), .ZN(new_n30783_));
  AOI21_X1   g27525(.A1(pi0299), .A2(new_n30783_), .B(new_n30668_), .ZN(new_n30784_));
  NOR2_X1    g27526(.A1(new_n30711_), .A2(new_n30784_), .ZN(new_n30785_));
  NAND3_X1   g27527(.A1(new_n30782_), .A2(new_n30762_), .A3(new_n30785_), .ZN(new_n30786_));
  XOR2_X1    g27528(.A1(new_n30759_), .A2(new_n30718_), .Z(new_n30787_));
  NOR2_X1    g27529(.A1(new_n30787_), .A2(new_n30786_), .ZN(new_n30788_));
  XOR2_X1    g27530(.A1(new_n30788_), .A2(new_n30760_), .Z(new_n30789_));
  OAI21_X1   g27531(.A1(new_n30789_), .A2(new_n8739_), .B(new_n30718_), .ZN(new_n30790_));
  NAND2_X1   g27532(.A1(new_n30790_), .A2(new_n30717_), .ZN(new_n30791_));
  NAND2_X1   g27533(.A1(new_n30713_), .A2(pi0207), .ZN(new_n30792_));
  NAND2_X1   g27534(.A1(new_n30792_), .A2(new_n8546_), .ZN(new_n30793_));
  NAND2_X1   g27535(.A1(new_n30793_), .A2(pi1157), .ZN(new_n30794_));
  NOR2_X1    g27536(.A1(new_n30726_), .A2(new_n8546_), .ZN(new_n30795_));
  XOR2_X1    g27537(.A1(new_n30795_), .A2(new_n8547_), .Z(new_n30796_));
  NAND2_X1   g27538(.A1(new_n30796_), .A2(new_n30687_), .ZN(new_n30797_));
  NOR2_X1    g27539(.A1(new_n30797_), .A2(new_n14006_), .ZN(new_n30798_));
  XNOR2_X1   g27540(.A1(new_n30798_), .A2(new_n30794_), .ZN(new_n30799_));
  AOI21_X1   g27541(.A1(new_n30742_), .A2(pi0207), .B(pi0208), .ZN(new_n30800_));
  NAND2_X1   g27542(.A1(new_n30799_), .A2(new_n30800_), .ZN(new_n30801_));
  AOI21_X1   g27543(.A1(new_n30801_), .A2(new_n8685_), .B(pi0212), .ZN(new_n30802_));
  AOI21_X1   g27544(.A1(new_n30797_), .A2(new_n30793_), .B(pi1157), .ZN(new_n30803_));
  NOR2_X1    g27545(.A1(new_n30672_), .A2(new_n30729_), .ZN(new_n30804_));
  NOR2_X1    g27546(.A1(new_n30750_), .A2(new_n13778_), .ZN(new_n30805_));
  NOR2_X1    g27547(.A1(new_n3098_), .A2(pi1155), .ZN(new_n30806_));
  NOR2_X1    g27548(.A1(new_n30805_), .A2(new_n30806_), .ZN(new_n30807_));
  NAND2_X1   g27549(.A1(new_n30804_), .A2(new_n30807_), .ZN(new_n30808_));
  NOR2_X1    g27550(.A1(new_n30808_), .A2(pi0207), .ZN(new_n30809_));
  NOR2_X1    g27551(.A1(new_n30705_), .A2(new_n14006_), .ZN(new_n30810_));
  INV_X1     g27552(.I(new_n30810_), .ZN(new_n30811_));
  INV_X1     g27553(.I(new_n30568_), .ZN(new_n30812_));
  INV_X1     g27554(.I(new_n30666_), .ZN(new_n30813_));
  AOI21_X1   g27555(.A1(pi1153), .A2(new_n30813_), .B(new_n30721_), .ZN(new_n30814_));
  INV_X1     g27556(.I(new_n30814_), .ZN(new_n30815_));
  NOR2_X1    g27557(.A1(new_n30815_), .A2(new_n30812_), .ZN(new_n30816_));
  NOR4_X1    g27558(.A1(new_n30811_), .A2(new_n8546_), .A3(new_n30809_), .A4(new_n30816_), .ZN(new_n30817_));
  OAI21_X1   g27559(.A1(new_n30803_), .A2(pi0211), .B(new_n30817_), .ZN(new_n30818_));
  AOI21_X1   g27560(.A1(new_n30818_), .A2(new_n8685_), .B(new_n30760_), .ZN(new_n30819_));
  NAND2_X1   g27561(.A1(new_n30802_), .A2(new_n30819_), .ZN(new_n30820_));
  AOI21_X1   g27562(.A1(new_n30791_), .A2(new_n8683_), .B(new_n30820_), .ZN(new_n30821_));
  INV_X1     g27563(.I(new_n30640_), .ZN(new_n30822_));
  NOR2_X1    g27564(.A1(new_n30786_), .A2(new_n30822_), .ZN(new_n30823_));
  NOR2_X1    g27565(.A1(new_n30801_), .A2(new_n30823_), .ZN(new_n30824_));
  NAND2_X1   g27566(.A1(new_n30802_), .A2(new_n30824_), .ZN(new_n30825_));
  AOI21_X1   g27567(.A1(new_n30804_), .A2(new_n30807_), .B(new_n8545_), .ZN(new_n30826_));
  INV_X1     g27568(.I(new_n30826_), .ZN(new_n30827_));
  NOR2_X1    g27569(.A1(new_n3098_), .A2(pi1153), .ZN(new_n30828_));
  INV_X1     g27570(.I(new_n30828_), .ZN(new_n30829_));
  NOR3_X1    g27571(.A1(new_n30815_), .A2(new_n8545_), .A3(new_n30829_), .ZN(new_n30830_));
  NOR2_X1    g27572(.A1(new_n30827_), .A2(new_n30830_), .ZN(new_n30831_));
  NOR4_X1    g27573(.A1(new_n30808_), .A2(new_n8545_), .A3(new_n30815_), .A4(new_n30829_), .ZN(new_n30832_));
  NOR3_X1    g27574(.A1(new_n30831_), .A2(new_n30832_), .A3(new_n8546_), .ZN(new_n30833_));
  NOR2_X1    g27575(.A1(new_n30757_), .A2(pi1157), .ZN(new_n30834_));
  NAND2_X1   g27576(.A1(new_n30822_), .A2(new_n30829_), .ZN(new_n30835_));
  OAI21_X1   g27577(.A1(new_n30810_), .A2(new_n30835_), .B(new_n30834_), .ZN(new_n30836_));
  OAI21_X1   g27578(.A1(new_n30833_), .A2(new_n30836_), .B(new_n8739_), .ZN(new_n30837_));
  NOR2_X1    g27579(.A1(pi0211), .A2(pi0214), .ZN(new_n30838_));
  NAND4_X1   g27580(.A1(new_n30717_), .A2(pi0211), .A3(new_n30837_), .A4(new_n30838_), .ZN(new_n30839_));
  AOI21_X1   g27581(.A1(new_n30825_), .A2(new_n30839_), .B(new_n8683_), .ZN(new_n30840_));
  OAI21_X1   g27582(.A1(new_n30821_), .A2(po1038), .B(new_n30840_), .ZN(new_n30841_));
  NAND3_X1   g27583(.A1(new_n30841_), .A2(new_n30634_), .A3(new_n30644_), .ZN(new_n30842_));
  INV_X1     g27584(.I(new_n30601_), .ZN(new_n30843_));
  INV_X1     g27585(.I(new_n30834_), .ZN(new_n30844_));
  NOR2_X1    g27586(.A1(new_n3098_), .A2(new_n3650_), .ZN(new_n30845_));
  NOR3_X1    g27587(.A1(new_n30721_), .A2(new_n8545_), .A3(new_n30725_), .ZN(new_n30846_));
  INV_X1     g27588(.I(new_n30845_), .ZN(new_n30847_));
  NAND2_X1   g27589(.A1(new_n30846_), .A2(new_n30847_), .ZN(new_n30848_));
  NAND2_X1   g27590(.A1(new_n30848_), .A2(new_n8546_), .ZN(new_n30849_));
  NOR2_X1    g27591(.A1(new_n30679_), .A2(new_n13969_), .ZN(new_n30850_));
  NAND2_X1   g27592(.A1(pi0299), .A2(pi1143), .ZN(new_n30851_));
  NOR2_X1    g27593(.A1(pi1154), .A2(pi1155), .ZN(new_n30852_));
  AOI21_X1   g27594(.A1(new_n30698_), .A2(new_n30852_), .B(new_n8555_), .ZN(new_n30853_));
  INV_X1     g27595(.I(new_n30685_), .ZN(new_n30855_));
  AOI21_X1   g27596(.A1(new_n30855_), .A2(new_n3098_), .B(new_n13817_), .ZN(new_n30856_));
  AND2_X2    g27597(.A1(new_n30856_), .A2(pi1156), .Z(new_n30857_));
  NAND2_X1   g27598(.A1(pi0299), .A2(pi1143), .ZN(new_n30858_));
  AOI21_X1   g27599(.A1(new_n30851_), .A2(new_n30858_), .B(new_n8545_), .ZN(new_n30859_));
  AOI22_X1   g27600(.A1(new_n30849_), .A2(new_n30859_), .B1(new_n30844_), .B2(new_n30845_), .ZN(new_n30860_));
  NOR2_X1    g27601(.A1(new_n30723_), .A2(pi1156), .ZN(new_n30861_));
  AOI21_X1   g27602(.A1(new_n30696_), .A2(new_n30861_), .B(new_n30739_), .ZN(new_n30862_));
  NOR2_X1    g27603(.A1(new_n30862_), .A2(new_n3098_), .ZN(new_n30863_));
  NAND2_X1   g27604(.A1(pi0207), .A2(pi0299), .ZN(new_n30864_));
  NOR2_X1    g27605(.A1(new_n30864_), .A2(new_n3650_), .ZN(new_n30865_));
  XNOR2_X1   g27606(.A1(new_n30863_), .A2(new_n30865_), .ZN(new_n30866_));
  NOR4_X1    g27607(.A1(new_n30860_), .A2(new_n8684_), .A3(new_n30745_), .A4(new_n30866_), .ZN(new_n30867_));
  XOR2_X1    g27608(.A1(new_n30867_), .A2(new_n30597_), .Z(new_n30868_));
  NOR2_X1    g27609(.A1(new_n3098_), .A2(pi1144), .ZN(new_n30869_));
  OR3_X2     g27610(.A1(new_n30758_), .A2(pi1157), .A3(new_n30869_), .Z(new_n30870_));
  OAI21_X1   g27611(.A1(new_n3057_), .A2(new_n30864_), .B(new_n30863_), .ZN(new_n30871_));
  NAND4_X1   g27612(.A1(new_n30862_), .A2(pi0207), .A3(pi0299), .A4(pi1144), .ZN(new_n30872_));
  NAND3_X1   g27613(.A1(new_n30871_), .A2(new_n30744_), .A3(new_n30872_), .ZN(new_n30873_));
  NOR2_X1    g27614(.A1(new_n8685_), .A2(pi0212), .ZN(new_n30874_));
  NOR2_X1    g27615(.A1(new_n8739_), .A2(pi0214), .ZN(new_n30875_));
  NOR2_X1    g27616(.A1(new_n30874_), .A2(new_n30875_), .ZN(new_n30876_));
  NOR2_X1    g27617(.A1(new_n30876_), .A2(new_n8684_), .ZN(new_n30877_));
  AOI21_X1   g27618(.A1(new_n30870_), .A2(new_n30873_), .B(new_n30877_), .ZN(new_n30878_));
  NAND2_X1   g27619(.A1(pi0299), .A2(pi1144), .ZN(new_n30879_));
  AOI21_X1   g27620(.A1(new_n30846_), .A2(new_n30879_), .B(pi0208), .ZN(new_n30880_));
  NOR3_X1    g27621(.A1(new_n30853_), .A2(pi0299), .A3(pi1144), .ZN(new_n30881_));
  NOR2_X1    g27622(.A1(new_n30881_), .A2(new_n13778_), .ZN(new_n30882_));
  OAI21_X1   g27623(.A1(new_n30857_), .A2(pi1144), .B(new_n30613_), .ZN(new_n30883_));
  NAND3_X1   g27624(.A1(new_n30850_), .A2(pi0299), .A3(new_n3057_), .ZN(new_n30884_));
  AOI21_X1   g27625(.A1(new_n30883_), .A2(new_n30727_), .B(new_n30884_), .ZN(new_n30885_));
  NOR4_X1    g27626(.A1(new_n30669_), .A2(new_n8545_), .A3(new_n13778_), .A4(new_n30869_), .ZN(new_n30886_));
  OAI21_X1   g27627(.A1(new_n30885_), .A2(new_n30882_), .B(new_n30886_), .ZN(new_n30887_));
  OR3_X2     g27628(.A1(new_n30878_), .A2(new_n30880_), .A3(new_n30887_), .Z(new_n30888_));
  NOR2_X1    g27629(.A1(new_n30597_), .A2(new_n8684_), .ZN(new_n30889_));
  NOR2_X1    g27630(.A1(new_n30889_), .A2(pi0219), .ZN(new_n30890_));
  OAI21_X1   g27631(.A1(new_n30868_), .A2(new_n30888_), .B(new_n30890_), .ZN(new_n30891_));
  NOR2_X1    g27632(.A1(new_n30586_), .A2(pi0219), .ZN(new_n30892_));
  NOR2_X1    g27633(.A1(new_n30594_), .A2(new_n30892_), .ZN(new_n30893_));
  INV_X1     g27634(.I(new_n30893_), .ZN(new_n30894_));
  NAND2_X1   g27635(.A1(new_n30772_), .A2(pi0207), .ZN(new_n30895_));
  XOR2_X1    g27636(.A1(new_n30895_), .A2(new_n30864_), .Z(new_n30896_));
  NAND2_X1   g27637(.A1(new_n30896_), .A2(pi1142), .ZN(new_n30897_));
  NOR2_X1    g27638(.A1(new_n30810_), .A2(new_n30834_), .ZN(new_n30898_));
  INV_X1     g27639(.I(new_n30677_), .ZN(new_n30899_));
  NAND3_X1   g27640(.A1(new_n8545_), .A2(new_n13817_), .A3(new_n13969_), .ZN(new_n30900_));
  NOR2_X1    g27641(.A1(new_n3098_), .A2(new_n3814_), .ZN(new_n30901_));
  INV_X1     g27642(.I(new_n30901_), .ZN(new_n30902_));
  NAND4_X1   g27643(.A1(new_n30804_), .A2(new_n30899_), .A3(new_n30900_), .A4(new_n30902_), .ZN(new_n30903_));
  AOI21_X1   g27644(.A1(new_n30903_), .A2(new_n3098_), .B(new_n3814_), .ZN(new_n30904_));
  NAND4_X1   g27645(.A1(new_n8689_), .A2(pi0208), .A3(new_n30893_), .A4(new_n30901_), .ZN(new_n30905_));
  NOR3_X1    g27646(.A1(new_n30898_), .A2(new_n30904_), .A3(new_n30905_), .ZN(new_n30906_));
  AOI21_X1   g27647(.A1(new_n30897_), .A2(new_n30906_), .B(po1038), .ZN(new_n30907_));
  NOR3_X1    g27648(.A1(new_n30801_), .A2(new_n30894_), .A3(new_n30907_), .ZN(new_n30908_));
  NOR2_X1    g27649(.A1(pi0209), .A2(pi0213), .ZN(new_n30909_));
  INV_X1     g27650(.I(new_n30909_), .ZN(new_n30910_));
  AOI21_X1   g27651(.A1(new_n30908_), .A2(new_n30891_), .B(new_n30910_), .ZN(new_n30911_));
  NOR4_X1    g27652(.A1(new_n30911_), .A2(new_n30557_), .A3(new_n27639_), .A4(new_n30843_), .ZN(new_n30912_));
  NAND2_X1   g27653(.A1(new_n30842_), .A2(new_n30912_), .ZN(new_n30913_));
  XNOR2_X1   g27654(.A1(new_n30913_), .A2(new_n30649_), .ZN(po0390));
  NOR2_X1    g27655(.A1(new_n8739_), .A2(new_n8683_), .ZN(new_n30915_));
  INV_X1     g27656(.I(new_n30915_), .ZN(new_n30916_));
  XOR2_X1    g27657(.A1(new_n30630_), .A2(new_n30916_), .Z(new_n30917_));
  INV_X1     g27658(.I(new_n30596_), .ZN(new_n30918_));
  NOR2_X1    g27659(.A1(new_n8684_), .A2(new_n13778_), .ZN(new_n30919_));
  NOR2_X1    g27660(.A1(new_n30919_), .A2(new_n30625_), .ZN(new_n30920_));
  NOR2_X1    g27661(.A1(new_n30920_), .A2(new_n8685_), .ZN(new_n30921_));
  INV_X1     g27662(.I(new_n30921_), .ZN(new_n30922_));
  NOR2_X1    g27663(.A1(new_n30637_), .A2(new_n8683_), .ZN(new_n30923_));
  INV_X1     g27664(.I(new_n30923_), .ZN(new_n30924_));
  NOR4_X1    g27665(.A1(new_n30918_), .A2(new_n28529_), .A3(new_n30922_), .A4(new_n30924_), .ZN(new_n30925_));
  AOI21_X1   g27666(.A1(new_n30917_), .A2(new_n30925_), .B(new_n30557_), .ZN(new_n30926_));
  NOR2_X1    g27667(.A1(new_n8774_), .A2(new_n13817_), .ZN(new_n30927_));
  NOR2_X1    g27668(.A1(new_n13614_), .A2(new_n13817_), .ZN(new_n30928_));
  XOR2_X1    g27669(.A1(new_n30927_), .A2(new_n30928_), .Z(new_n30929_));
  NAND2_X1   g27670(.A1(new_n30929_), .A2(new_n9214_), .ZN(new_n30930_));
  INV_X1     g27671(.I(new_n30650_), .ZN(new_n30931_));
  NOR2_X1    g27672(.A1(new_n30931_), .A2(new_n13614_), .ZN(new_n30932_));
  INV_X1     g27673(.I(new_n30932_), .ZN(new_n30933_));
  NOR2_X1    g27674(.A1(new_n30933_), .A2(pi0299), .ZN(new_n30934_));
  NOR2_X1    g27675(.A1(new_n30934_), .A2(pi0207), .ZN(new_n30935_));
  AOI21_X1   g27676(.A1(new_n30930_), .A2(new_n30935_), .B(new_n8546_), .ZN(new_n30936_));
  NOR2_X1    g27677(.A1(new_n30934_), .A2(new_n8545_), .ZN(new_n30937_));
  NOR3_X1    g27678(.A1(new_n30930_), .A2(new_n8545_), .A3(new_n30614_), .ZN(new_n30938_));
  XOR2_X1    g27679(.A1(new_n30938_), .A2(new_n30937_), .Z(new_n30939_));
  OAI21_X1   g27680(.A1(new_n8773_), .A2(new_n13614_), .B(new_n3098_), .ZN(new_n30940_));
  AOI21_X1   g27681(.A1(new_n30940_), .A2(new_n30706_), .B(new_n9090_), .ZN(new_n30941_));
  NAND2_X1   g27682(.A1(new_n30939_), .A2(new_n30941_), .ZN(new_n30942_));
  XOR2_X1    g27683(.A1(new_n30942_), .A2(new_n30936_), .Z(new_n30943_));
  INV_X1     g27684(.I(new_n30876_), .ZN(new_n30944_));
  NOR2_X1    g27685(.A1(new_n30612_), .A2(pi0207), .ZN(new_n30945_));
  INV_X1     g27686(.I(new_n30945_), .ZN(new_n30946_));
  NOR2_X1    g27687(.A1(new_n30659_), .A2(pi1153), .ZN(new_n30947_));
  NOR3_X1    g27688(.A1(new_n30947_), .A2(new_n13817_), .A3(new_n9214_), .ZN(new_n30948_));
  NOR2_X1    g27689(.A1(new_n13614_), .A2(pi1154), .ZN(new_n30949_));
  INV_X1     g27690(.I(new_n30949_), .ZN(new_n30950_));
  NOR2_X1    g27691(.A1(new_n30750_), .A2(new_n30950_), .ZN(new_n30951_));
  NOR2_X1    g27692(.A1(new_n30951_), .A2(new_n30948_), .ZN(new_n30952_));
  NAND2_X1   g27693(.A1(new_n30952_), .A2(pi0207), .ZN(new_n30953_));
  AOI21_X1   g27694(.A1(new_n30953_), .A2(new_n30946_), .B(pi0208), .ZN(new_n30954_));
  NAND2_X1   g27695(.A1(new_n8775_), .A2(pi0207), .ZN(new_n30955_));
  NAND3_X1   g27696(.A1(new_n30952_), .A2(pi0207), .A3(pi1153), .ZN(new_n30956_));
  XOR2_X1    g27697(.A1(new_n30956_), .A2(new_n30955_), .Z(new_n30957_));
  AOI21_X1   g27698(.A1(new_n30957_), .A2(pi0208), .B(new_n30954_), .ZN(new_n30958_));
  NAND2_X1   g27699(.A1(new_n30958_), .A2(new_n30944_), .ZN(new_n30959_));
  XOR2_X1    g27700(.A1(new_n30959_), .A2(new_n30877_), .Z(new_n30960_));
  NOR2_X1    g27701(.A1(new_n30943_), .A2(new_n30960_), .ZN(new_n30961_));
  NAND2_X1   g27702(.A1(new_n30958_), .A2(new_n30597_), .ZN(new_n30962_));
  NOR2_X1    g27703(.A1(new_n30812_), .A2(new_n8546_), .ZN(new_n30963_));
  NOR2_X1    g27704(.A1(new_n8546_), .A2(pi0207), .ZN(new_n30964_));
  NOR2_X1    g27705(.A1(new_n8545_), .A2(pi0208), .ZN(new_n30965_));
  NOR2_X1    g27706(.A1(new_n30964_), .A2(new_n30965_), .ZN(new_n30966_));
  INV_X1     g27707(.I(new_n30966_), .ZN(new_n30967_));
  NAND2_X1   g27708(.A1(new_n30967_), .A2(new_n30963_), .ZN(new_n30968_));
  NOR2_X1    g27709(.A1(new_n8774_), .A2(new_n13614_), .ZN(new_n30969_));
  AOI21_X1   g27710(.A1(pi0200), .A2(new_n13614_), .B(new_n9209_), .ZN(new_n30970_));
  NAND2_X1   g27711(.A1(new_n30970_), .A2(pi1154), .ZN(new_n30971_));
  INV_X1     g27712(.I(new_n30971_), .ZN(new_n30972_));
  AOI21_X1   g27713(.A1(new_n30934_), .A2(new_n13817_), .B(new_n30972_), .ZN(new_n30973_));
  INV_X1     g27714(.I(new_n30973_), .ZN(new_n30974_));
  NAND2_X1   g27715(.A1(new_n30974_), .A2(new_n30969_), .ZN(new_n30975_));
  NAND2_X1   g27716(.A1(new_n30975_), .A2(new_n30968_), .ZN(new_n30976_));
  INV_X1     g27717(.I(new_n30976_), .ZN(new_n30977_));
  NOR2_X1    g27718(.A1(new_n30977_), .A2(new_n7240_), .ZN(new_n30978_));
  INV_X1     g27719(.I(new_n30892_), .ZN(new_n30979_));
  NOR2_X1    g27720(.A1(new_n8684_), .A2(pi1153), .ZN(new_n30980_));
  NOR2_X1    g27721(.A1(pi0211), .A2(pi1154), .ZN(new_n30981_));
  NOR2_X1    g27722(.A1(new_n30980_), .A2(new_n30981_), .ZN(new_n30982_));
  INV_X1     g27723(.I(new_n30982_), .ZN(new_n30983_));
  AOI21_X1   g27724(.A1(new_n30983_), .A2(new_n30597_), .B(new_n30979_), .ZN(new_n30984_));
  OAI21_X1   g27725(.A1(new_n30597_), .A2(new_n30635_), .B(new_n30984_), .ZN(new_n30985_));
  INV_X1     g27726(.I(new_n30985_), .ZN(new_n30986_));
  AOI21_X1   g27727(.A1(new_n30986_), .A2(po1038), .B(pi1152), .ZN(new_n30987_));
  INV_X1     g27728(.I(new_n30987_), .ZN(new_n30988_));
  NAND2_X1   g27729(.A1(new_n30876_), .A2(new_n30822_), .ZN(new_n30989_));
  NOR2_X1    g27730(.A1(new_n30988_), .A2(new_n30989_), .ZN(new_n30990_));
  AOI21_X1   g27731(.A1(new_n30978_), .A2(new_n30990_), .B(pi0219), .ZN(new_n30991_));
  NOR2_X1    g27732(.A1(new_n30991_), .A2(new_n8684_), .ZN(new_n30992_));
  OAI21_X1   g27733(.A1(new_n30961_), .A2(new_n30962_), .B(new_n30992_), .ZN(new_n30993_));
  NOR2_X1    g27734(.A1(new_n8684_), .A2(new_n13817_), .ZN(new_n30994_));
  INV_X1     g27735(.I(new_n30994_), .ZN(new_n30995_));
  NAND2_X1   g27736(.A1(new_n8686_), .A2(new_n13817_), .ZN(new_n30996_));
  NAND2_X1   g27737(.A1(new_n30718_), .A2(pi1154), .ZN(new_n30997_));
  AOI21_X1   g27738(.A1(new_n30997_), .A2(new_n30996_), .B(new_n13614_), .ZN(new_n30998_));
  AOI21_X1   g27739(.A1(new_n30998_), .A2(new_n30995_), .B(new_n8739_), .ZN(new_n30999_));
  OAI21_X1   g27740(.A1(new_n30995_), .A2(new_n30998_), .B(new_n30999_), .ZN(new_n31000_));
  INV_X1     g27741(.I(new_n31000_), .ZN(new_n31001_));
  INV_X1     g27742(.I(pi1152), .ZN(new_n31002_));
  INV_X1     g27743(.I(new_n30874_), .ZN(new_n31003_));
  NOR2_X1    g27744(.A1(new_n30983_), .A2(new_n31003_), .ZN(new_n31004_));
  OAI22_X1   g27745(.A1(new_n30918_), .A2(new_n31002_), .B1(pi0219), .B2(new_n31004_), .ZN(new_n31005_));
  NAND2_X1   g27746(.A1(new_n31001_), .A2(new_n31005_), .ZN(new_n31006_));
  NOR2_X1    g27747(.A1(new_n8773_), .A2(pi1153), .ZN(new_n31007_));
  NOR2_X1    g27748(.A1(new_n30738_), .A2(new_n31007_), .ZN(new_n31008_));
  INV_X1     g27749(.I(new_n31008_), .ZN(new_n31009_));
  NOR2_X1    g27750(.A1(new_n31009_), .A2(new_n8545_), .ZN(new_n31010_));
  NOR2_X1    g27751(.A1(new_n8773_), .A2(pi0299), .ZN(new_n31011_));
  NAND3_X1   g27752(.A1(new_n31011_), .A2(pi1153), .A3(pi1154), .ZN(new_n31012_));
  INV_X1     g27753(.I(new_n31011_), .ZN(new_n31013_));
  NAND3_X1   g27754(.A1(new_n31013_), .A2(new_n13614_), .A3(pi1154), .ZN(new_n31014_));
  AOI21_X1   g27755(.A1(new_n31014_), .A2(new_n31012_), .B(new_n30738_), .ZN(new_n31015_));
  NOR2_X1    g27756(.A1(pi0199), .A2(pi1153), .ZN(new_n31016_));
  NOR2_X1    g27757(.A1(new_n30654_), .A2(new_n31016_), .ZN(new_n31017_));
  NOR2_X1    g27758(.A1(new_n31015_), .A2(new_n31017_), .ZN(new_n31018_));
  INV_X1     g27759(.I(new_n31018_), .ZN(new_n31019_));
  XOR2_X1    g27760(.A1(new_n31008_), .A2(new_n9090_), .Z(new_n31020_));
  NOR2_X1    g27761(.A1(new_n31019_), .A2(new_n31020_), .ZN(new_n31021_));
  XNOR2_X1   g27762(.A1(new_n31021_), .A2(new_n31010_), .ZN(new_n31022_));
  INV_X1     g27763(.I(new_n31022_), .ZN(new_n31023_));
  NOR2_X1    g27764(.A1(new_n31022_), .A2(new_n8684_), .ZN(new_n31024_));
  NOR2_X1    g27765(.A1(new_n8549_), .A2(new_n13614_), .ZN(new_n31025_));
  OAI21_X1   g27766(.A1(pi1154), .A2(new_n30673_), .B(new_n31025_), .ZN(new_n31026_));
  OAI21_X1   g27767(.A1(new_n30813_), .A2(new_n31026_), .B(new_n13817_), .ZN(new_n31027_));
  NAND2_X1   g27768(.A1(new_n31027_), .A2(new_n30934_), .ZN(new_n31028_));
  NOR2_X1    g27769(.A1(new_n8549_), .A2(new_n3098_), .ZN(new_n31029_));
  INV_X1     g27770(.I(new_n31029_), .ZN(new_n31030_));
  AOI21_X1   g27771(.A1(new_n31030_), .A2(new_n13614_), .B(new_n8555_), .ZN(new_n31031_));
  INV_X1     g27772(.I(new_n31031_), .ZN(new_n31032_));
  NOR2_X1    g27773(.A1(new_n31032_), .A2(new_n30651_), .ZN(new_n31033_));
  NAND2_X1   g27774(.A1(new_n31028_), .A2(pi0208), .ZN(new_n31034_));
  XOR2_X1    g27775(.A1(new_n31034_), .A2(new_n9090_), .Z(new_n31035_));
  NAND2_X1   g27776(.A1(new_n31035_), .A2(new_n31033_), .ZN(new_n31036_));
  INV_X1     g27777(.I(new_n31036_), .ZN(new_n31037_));
  AOI21_X1   g27778(.A1(new_n30693_), .A2(new_n31028_), .B(new_n31037_), .ZN(new_n31038_));
  NOR2_X1    g27779(.A1(new_n31038_), .A2(pi0211), .ZN(new_n31039_));
  NOR2_X1    g27780(.A1(new_n31039_), .A2(new_n31024_), .ZN(new_n31040_));
  NAND2_X1   g27781(.A1(new_n31040_), .A2(pi0219), .ZN(new_n31041_));
  NAND2_X1   g27782(.A1(new_n30586_), .A2(pi0219), .ZN(new_n31042_));
  XNOR2_X1   g27783(.A1(new_n31041_), .A2(new_n31042_), .ZN(new_n31043_));
  OAI21_X1   g27784(.A1(new_n31043_), .A2(new_n31022_), .B(new_n7240_), .ZN(new_n31044_));
  NOR2_X1    g27785(.A1(new_n30669_), .A2(new_n30947_), .ZN(new_n31045_));
  OR2_X2     g27786(.A1(new_n31045_), .A2(new_n30948_), .Z(new_n31046_));
  NOR2_X1    g27787(.A1(new_n31046_), .A2(new_n8545_), .ZN(new_n31047_));
  NOR2_X1    g27788(.A1(new_n31047_), .A2(new_n30945_), .ZN(new_n31048_));
  NOR2_X1    g27789(.A1(new_n31048_), .A2(pi0208), .ZN(new_n31049_));
  NOR2_X1    g27790(.A1(new_n8774_), .A2(pi1153), .ZN(new_n31050_));
  NOR2_X1    g27791(.A1(new_n31050_), .A2(new_n8545_), .ZN(new_n31051_));
  NOR2_X1    g27792(.A1(new_n30674_), .A2(new_n8549_), .ZN(new_n31052_));
  INV_X1     g27793(.I(new_n31052_), .ZN(new_n31053_));
  NOR3_X1    g27794(.A1(new_n31046_), .A2(new_n8545_), .A3(new_n31053_), .ZN(new_n31054_));
  XOR2_X1    g27795(.A1(new_n31054_), .A2(new_n31051_), .Z(new_n31055_));
  AOI21_X1   g27796(.A1(new_n31055_), .A2(pi0208), .B(new_n31049_), .ZN(new_n31056_));
  NAND2_X1   g27797(.A1(new_n31056_), .A2(pi0214), .ZN(new_n31057_));
  XOR2_X1    g27798(.A1(new_n31057_), .A2(new_n30718_), .Z(new_n31058_));
  AOI21_X1   g27799(.A1(new_n31058_), .A2(new_n31038_), .B(pi0212), .ZN(new_n31059_));
  NOR2_X1    g27800(.A1(new_n31018_), .A2(new_n8545_), .ZN(new_n31060_));
  NOR2_X1    g27801(.A1(new_n31060_), .A2(new_n8546_), .ZN(new_n31061_));
  INV_X1     g27802(.I(new_n31033_), .ZN(new_n31062_));
  NAND2_X1   g27803(.A1(new_n31062_), .A2(pi0207), .ZN(new_n31063_));
  NOR2_X1    g27804(.A1(new_n31015_), .A2(new_n30927_), .ZN(new_n31064_));
  NOR3_X1    g27805(.A1(new_n8545_), .A2(new_n3098_), .A3(pi1154), .ZN(new_n31065_));
  NAND2_X1   g27806(.A1(new_n31064_), .A2(new_n31065_), .ZN(new_n31066_));
  XOR2_X1    g27807(.A1(new_n31066_), .A2(new_n31063_), .Z(new_n31067_));
  NAND2_X1   g27808(.A1(new_n31067_), .A2(new_n30714_), .ZN(new_n31068_));
  XNOR2_X1   g27809(.A1(new_n31068_), .A2(new_n31061_), .ZN(new_n31069_));
  NOR2_X1    g27810(.A1(new_n31056_), .A2(new_n8684_), .ZN(new_n31070_));
  AOI21_X1   g27811(.A1(new_n31069_), .A2(new_n8684_), .B(new_n31070_), .ZN(new_n31071_));
  OR3_X2     g27812(.A1(new_n31059_), .A2(new_n8685_), .A3(new_n31071_), .Z(new_n31072_));
  NAND3_X1   g27813(.A1(new_n31044_), .A2(new_n8683_), .A3(new_n31072_), .ZN(new_n31073_));
  NAND2_X1   g27814(.A1(new_n31071_), .A2(pi0214), .ZN(new_n31074_));
  XOR2_X1    g27815(.A1(new_n31074_), .A2(new_n30597_), .Z(new_n31075_));
  AND3_X2    g27816(.A1(new_n31073_), .A2(new_n31023_), .A3(new_n31075_), .Z(new_n31076_));
  OAI21_X1   g27817(.A1(new_n31076_), .A2(new_n31006_), .B(new_n30993_), .ZN(new_n31077_));
  NAND2_X1   g27818(.A1(new_n31077_), .A2(pi0213), .ZN(new_n31078_));
  NOR2_X1    g27819(.A1(new_n28364_), .A2(new_n28529_), .ZN(new_n31079_));
  INV_X1     g27820(.I(new_n31079_), .ZN(new_n31080_));
  XOR2_X1    g27821(.A1(new_n31078_), .A2(new_n31080_), .Z(new_n31081_));
  INV_X1     g27822(.I(new_n30762_), .ZN(new_n31082_));
  NOR2_X1    g27823(.A1(new_n3098_), .A2(pi0207), .ZN(new_n31083_));
  NOR2_X1    g27824(.A1(new_n8773_), .A2(pi1154), .ZN(new_n31084_));
  NAND2_X1   g27825(.A1(new_n31084_), .A2(new_n30610_), .ZN(new_n31085_));
  XOR2_X1    g27826(.A1(new_n31085_), .A2(new_n31083_), .Z(new_n31086_));
  OR2_X2     g27827(.A1(new_n31036_), .A2(new_n31086_), .Z(new_n31087_));
  AOI21_X1   g27828(.A1(new_n31087_), .A2(new_n31082_), .B(new_n31028_), .ZN(new_n31088_));
  INV_X1     g27829(.I(new_n31088_), .ZN(new_n31089_));
  NOR2_X1    g27830(.A1(new_n8740_), .A2(new_n30586_), .ZN(new_n31090_));
  INV_X1     g27831(.I(new_n31090_), .ZN(new_n31091_));
  NAND2_X1   g27832(.A1(new_n8546_), .A2(new_n8684_), .ZN(new_n31092_));
  OAI21_X1   g27833(.A1(new_n31060_), .A2(new_n31092_), .B(new_n30733_), .ZN(new_n31093_));
  NAND2_X1   g27834(.A1(new_n31062_), .A2(new_n8545_), .ZN(new_n31094_));
  AOI21_X1   g27835(.A1(new_n31094_), .A2(new_n30733_), .B(pi0208), .ZN(new_n31095_));
  OAI21_X1   g27836(.A1(new_n31019_), .A2(new_n30733_), .B(new_n8545_), .ZN(new_n31096_));
  AOI21_X1   g27837(.A1(new_n31093_), .A2(new_n31095_), .B(new_n31096_), .ZN(new_n31097_));
  OAI21_X1   g27838(.A1(new_n31097_), .A2(new_n31091_), .B(pi0211), .ZN(new_n31098_));
  OAI21_X1   g27839(.A1(new_n31089_), .A2(new_n31098_), .B(new_n8683_), .ZN(new_n31099_));
  INV_X1     g27840(.I(new_n30875_), .ZN(new_n31100_));
  NAND2_X1   g27841(.A1(new_n30586_), .A2(pi0211), .ZN(new_n31101_));
  NOR4_X1    g27842(.A1(new_n31069_), .A2(new_n31100_), .A3(new_n31023_), .A4(new_n31101_), .ZN(new_n31102_));
  NAND2_X1   g27843(.A1(new_n31099_), .A2(new_n31102_), .ZN(new_n31103_));
  NOR2_X1    g27844(.A1(new_n31069_), .A2(new_n30597_), .ZN(new_n31104_));
  XOR2_X1    g27845(.A1(new_n31104_), .A2(new_n30889_), .Z(new_n31105_));
  NAND3_X1   g27846(.A1(new_n31105_), .A2(pi0219), .A3(new_n31088_), .ZN(new_n31106_));
  NAND3_X1   g27847(.A1(new_n31106_), .A2(pi1152), .A3(new_n31103_), .ZN(new_n31107_));
  NOR2_X1    g27848(.A1(new_n7240_), .A2(new_n31002_), .ZN(new_n31108_));
  XOR2_X1    g27849(.A1(new_n31107_), .A2(new_n31108_), .Z(new_n31109_));
  OR2_X2     g27850(.A1(new_n30943_), .A2(new_n8684_), .Z(new_n31110_));
  OAI21_X1   g27851(.A1(new_n3098_), .A2(pi1155), .B(new_n30940_), .ZN(new_n31111_));
  NAND2_X1   g27852(.A1(new_n31111_), .A2(pi0207), .ZN(new_n31112_));
  AOI21_X1   g27853(.A1(new_n30933_), .A2(pi0299), .B(new_n30614_), .ZN(new_n31113_));
  NOR3_X1    g27854(.A1(new_n30932_), .A2(new_n3098_), .A3(pi1154), .ZN(new_n31114_));
  NOR2_X1    g27855(.A1(new_n31113_), .A2(new_n31114_), .ZN(new_n31115_));
  OAI22_X1   g27856(.A1(new_n30783_), .A2(new_n30930_), .B1(new_n31115_), .B2(new_n13778_), .ZN(new_n31116_));
  INV_X1     g27857(.I(new_n31116_), .ZN(new_n31117_));
  AOI22_X1   g27858(.A1(new_n31117_), .A2(new_n8545_), .B1(pi0208), .B2(new_n31112_), .ZN(new_n31118_));
  AOI21_X1   g27859(.A1(new_n31117_), .A2(new_n8545_), .B(new_n30762_), .ZN(new_n31119_));
  NOR3_X1    g27860(.A1(new_n31118_), .A2(new_n31119_), .A3(pi0211), .ZN(new_n31120_));
  AOI22_X1   g27861(.A1(new_n31110_), .A2(new_n8740_), .B1(new_n8684_), .B2(new_n31120_), .ZN(new_n31121_));
  NOR2_X1    g27862(.A1(new_n31091_), .A2(pi0211), .ZN(new_n31122_));
  AOI21_X1   g27863(.A1(new_n30977_), .A2(new_n31122_), .B(new_n30743_), .ZN(new_n31123_));
  NOR2_X1    g27864(.A1(new_n31120_), .A2(new_n31123_), .ZN(new_n31124_));
  OAI21_X1   g27865(.A1(new_n31121_), .A2(new_n31124_), .B(new_n8683_), .ZN(new_n31125_));
  NOR2_X1    g27866(.A1(new_n30586_), .A2(new_n8683_), .ZN(new_n31126_));
  NAND2_X1   g27867(.A1(new_n30943_), .A2(new_n31126_), .ZN(new_n31127_));
  NAND2_X1   g27868(.A1(new_n31126_), .A2(pi0211), .ZN(new_n31128_));
  XOR2_X1    g27869(.A1(new_n31127_), .A2(new_n31128_), .Z(new_n31129_));
  NAND2_X1   g27870(.A1(new_n31129_), .A2(new_n30976_), .ZN(new_n31130_));
  NAND2_X1   g27871(.A1(new_n30977_), .A2(new_n30586_), .ZN(new_n31131_));
  NAND3_X1   g27872(.A1(new_n31130_), .A2(new_n31125_), .A3(new_n31131_), .ZN(new_n31132_));
  NOR2_X1    g27873(.A1(new_n31109_), .A2(new_n31132_), .ZN(new_n31133_));
  OAI21_X1   g27874(.A1(new_n8555_), .A2(pi0299), .B(pi0199), .ZN(new_n31134_));
  AOI21_X1   g27875(.A1(new_n30699_), .A2(new_n9208_), .B(pi1154), .ZN(new_n31135_));
  NOR3_X1    g27876(.A1(new_n31135_), .A2(new_n13778_), .A3(new_n31134_), .ZN(new_n31136_));
  NAND2_X1   g27877(.A1(new_n31136_), .A2(pi0207), .ZN(new_n31137_));
  XOR2_X1    g27878(.A1(new_n31136_), .A2(new_n8547_), .Z(new_n31138_));
  NAND2_X1   g27879(.A1(new_n30687_), .A2(new_n31138_), .ZN(new_n31139_));
  XNOR2_X1   g27880(.A1(new_n31139_), .A2(new_n31137_), .ZN(new_n31140_));
  INV_X1     g27881(.I(new_n31140_), .ZN(new_n31141_));
  AOI21_X1   g27882(.A1(new_n30734_), .A2(new_n31136_), .B(new_n8684_), .ZN(new_n31142_));
  OAI21_X1   g27883(.A1(new_n30731_), .A2(new_n8545_), .B(new_n30743_), .ZN(new_n31143_));
  NAND2_X1   g27884(.A1(new_n31143_), .A2(new_n8546_), .ZN(new_n31144_));
  NAND4_X1   g27885(.A1(new_n30687_), .A2(new_n8545_), .A3(pi0208), .A4(new_n30611_), .ZN(new_n31145_));
  NOR3_X1    g27886(.A1(new_n31144_), .A2(new_n8684_), .A3(new_n31145_), .ZN(new_n31146_));
  XNOR2_X1   g27887(.A1(new_n31146_), .A2(new_n31142_), .ZN(new_n31147_));
  NAND2_X1   g27888(.A1(new_n31147_), .A2(pi0214), .ZN(new_n31148_));
  XOR2_X1    g27889(.A1(new_n31148_), .A2(new_n30597_), .Z(new_n31149_));
  NOR2_X1    g27890(.A1(new_n30688_), .A2(new_n30672_), .ZN(new_n31150_));
  NOR2_X1    g27891(.A1(new_n31150_), .A2(new_n8545_), .ZN(new_n31151_));
  XOR2_X1    g27892(.A1(new_n31151_), .A2(new_n9090_), .Z(new_n31152_));
  AOI21_X1   g27893(.A1(new_n13778_), .A2(new_n8772_), .B(new_n30722_), .ZN(new_n31153_));
  NOR2_X1    g27894(.A1(new_n31153_), .A2(pi0299), .ZN(new_n31154_));
  NOR2_X1    g27895(.A1(new_n31154_), .A2(new_n31135_), .ZN(new_n31155_));
  INV_X1     g27896(.I(new_n31155_), .ZN(new_n31156_));
  OAI22_X1   g27897(.A1(new_n31152_), .A2(new_n30614_), .B1(new_n30690_), .B2(new_n31156_), .ZN(new_n31157_));
  NOR2_X1    g27898(.A1(new_n30604_), .A2(pi0219), .ZN(new_n31158_));
  NOR2_X1    g27899(.A1(new_n31157_), .A2(new_n31158_), .ZN(new_n31159_));
  NAND2_X1   g27900(.A1(new_n7240_), .A2(pi0213), .ZN(new_n31160_));
  OAI21_X1   g27901(.A1(new_n31159_), .A2(new_n31160_), .B(new_n8683_), .ZN(new_n31161_));
  AOI21_X1   g27902(.A1(new_n31149_), .A2(new_n31141_), .B(new_n31161_), .ZN(new_n31162_));
  NAND2_X1   g27903(.A1(new_n31157_), .A2(pi0214), .ZN(new_n31163_));
  XOR2_X1    g27904(.A1(new_n31163_), .A2(new_n8686_), .Z(new_n31164_));
  OAI21_X1   g27905(.A1(new_n31164_), .A2(new_n31145_), .B(new_n8739_), .ZN(new_n31165_));
  NOR2_X1    g27906(.A1(new_n31147_), .A2(new_n8685_), .ZN(new_n31166_));
  NAND2_X1   g27907(.A1(new_n31165_), .A2(new_n31166_), .ZN(new_n31167_));
  OAI21_X1   g27908(.A1(new_n31162_), .A2(new_n31167_), .B(new_n28364_), .ZN(new_n31168_));
  AOI21_X1   g27909(.A1(new_n31081_), .A2(new_n31133_), .B(new_n31168_), .ZN(new_n31169_));
  NOR2_X1    g27910(.A1(new_n31157_), .A2(pi0211), .ZN(new_n31170_));
  NOR2_X1    g27911(.A1(new_n30808_), .A2(new_n8545_), .ZN(new_n31171_));
  INV_X1     g27912(.I(new_n31171_), .ZN(new_n31172_));
  NAND2_X1   g27913(.A1(new_n31156_), .A2(new_n30568_), .ZN(new_n31173_));
  NAND4_X1   g27914(.A1(new_n31172_), .A2(pi0208), .A3(new_n30693_), .A4(new_n31173_), .ZN(new_n31174_));
  AOI21_X1   g27915(.A1(new_n31174_), .A2(new_n30808_), .B(new_n8545_), .ZN(new_n31175_));
  NOR2_X1    g27916(.A1(new_n31175_), .A2(new_n30828_), .ZN(new_n31176_));
  NOR2_X1    g27917(.A1(new_n31176_), .A2(new_n8684_), .ZN(new_n31177_));
  NOR2_X1    g27918(.A1(new_n31177_), .A2(new_n31170_), .ZN(new_n31178_));
  NOR2_X1    g27919(.A1(new_n31175_), .A2(pi0214), .ZN(new_n31179_));
  NAND2_X1   g27920(.A1(new_n30828_), .A2(pi0211), .ZN(new_n31180_));
  NAND2_X1   g27921(.A1(new_n31178_), .A2(pi0214), .ZN(new_n31181_));
  XOR2_X1    g27922(.A1(new_n31181_), .A2(new_n8740_), .Z(new_n31182_));
  OAI21_X1   g27923(.A1(new_n31182_), .A2(new_n31140_), .B(new_n8683_), .ZN(new_n31183_));
  OAI22_X1   g27924(.A1(new_n31183_), .A2(new_n8739_), .B1(new_n31179_), .B2(new_n31180_), .ZN(new_n31184_));
  NAND3_X1   g27925(.A1(new_n31184_), .A2(new_n8685_), .A3(new_n31178_), .ZN(new_n31185_));
  INV_X1     g27926(.I(new_n31006_), .ZN(new_n31186_));
  NOR2_X1    g27927(.A1(new_n31186_), .A2(po1038), .ZN(new_n31187_));
  AOI21_X1   g27928(.A1(new_n31141_), .A2(new_n30604_), .B(new_n8683_), .ZN(new_n31188_));
  OAI21_X1   g27929(.A1(new_n31175_), .A2(new_n30604_), .B(new_n31188_), .ZN(new_n31189_));
  AOI21_X1   g27930(.A1(new_n31185_), .A2(new_n31187_), .B(new_n31189_), .ZN(new_n31190_));
  NOR2_X1    g27931(.A1(new_n31141_), .A2(new_n8683_), .ZN(new_n31191_));
  OR3_X2     g27932(.A1(new_n31183_), .A2(po1038), .A3(new_n31191_), .Z(new_n31192_));
  NAND2_X1   g27933(.A1(new_n31178_), .A2(new_n8685_), .ZN(new_n31193_));
  NOR2_X1    g27934(.A1(new_n31176_), .A2(new_n8685_), .ZN(new_n31194_));
  XOR2_X1    g27935(.A1(new_n31194_), .A2(new_n8686_), .Z(new_n31195_));
  NAND2_X1   g27936(.A1(new_n31195_), .A2(new_n31141_), .ZN(new_n31196_));
  NOR2_X1    g27937(.A1(new_n30557_), .A2(new_n2768_), .ZN(new_n31197_));
  NAND4_X1   g27938(.A1(new_n31196_), .A2(new_n30987_), .A3(new_n31193_), .A4(new_n31197_), .ZN(new_n31198_));
  AOI21_X1   g27939(.A1(new_n31192_), .A2(new_n8739_), .B(new_n31198_), .ZN(new_n31199_));
  OAI21_X1   g27940(.A1(new_n31190_), .A2(pi0213), .B(new_n31199_), .ZN(new_n31200_));
  NOR2_X1    g27941(.A1(new_n31169_), .A2(new_n31200_), .ZN(new_n31201_));
  XOR2_X1    g27942(.A1(new_n31201_), .A2(new_n30926_), .Z(po0391));
  INV_X1     g27943(.I(new_n30612_), .ZN(new_n31203_));
  INV_X1     g27944(.I(new_n30952_), .ZN(new_n31204_));
  NOR2_X1    g27945(.A1(new_n30814_), .A2(new_n8545_), .ZN(new_n31205_));
  XOR2_X1    g27946(.A1(new_n31205_), .A2(new_n9090_), .Z(new_n31206_));
  NOR2_X1    g27947(.A1(new_n30814_), .A2(new_n8546_), .ZN(new_n31207_));
  XOR2_X1    g27948(.A1(new_n31207_), .A2(new_n9090_), .Z(new_n31208_));
  OAI22_X1   g27949(.A1(new_n31203_), .A2(new_n31206_), .B1(new_n31208_), .B2(new_n31204_), .ZN(new_n31209_));
  NOR2_X1    g27950(.A1(new_n31209_), .A2(pi0211), .ZN(new_n31210_));
  NOR2_X1    g27951(.A1(pi0207), .A2(pi0208), .ZN(new_n31211_));
  AOI21_X1   g27952(.A1(new_n30726_), .A2(new_n9090_), .B(new_n31211_), .ZN(new_n31212_));
  INV_X1     g27953(.I(new_n31212_), .ZN(new_n31213_));
  AOI21_X1   g27954(.A1(new_n8547_), .A2(new_n30973_), .B(new_n31213_), .ZN(new_n31214_));
  INV_X1     g27955(.I(new_n31214_), .ZN(new_n31215_));
  AOI21_X1   g27956(.A1(new_n31215_), .A2(pi0211), .B(new_n31091_), .ZN(new_n31216_));
  NAND2_X1   g27957(.A1(new_n31216_), .A2(pi0219), .ZN(new_n31217_));
  NOR2_X1    g27958(.A1(new_n31210_), .A2(new_n31217_), .ZN(new_n31218_));
  NAND2_X1   g27959(.A1(new_n31117_), .A2(pi0207), .ZN(new_n31219_));
  NOR2_X1    g27960(.A1(new_n31082_), .A2(new_n8546_), .ZN(new_n31220_));
  NOR2_X1    g27961(.A1(new_n30773_), .A2(new_n30762_), .ZN(new_n31221_));
  INV_X1     g27962(.I(new_n31221_), .ZN(new_n31222_));
  AOI22_X1   g27963(.A1(new_n31222_), .A2(pi0207), .B1(new_n31219_), .B2(new_n31220_), .ZN(new_n31223_));
  NOR2_X1    g27964(.A1(new_n30664_), .A2(new_n8545_), .ZN(new_n31224_));
  XOR2_X1    g27965(.A1(new_n31224_), .A2(new_n8547_), .Z(new_n31225_));
  NAND2_X1   g27966(.A1(new_n31225_), .A2(new_n30613_), .ZN(new_n31226_));
  NAND2_X1   g27967(.A1(new_n30930_), .A2(pi0207), .ZN(new_n31227_));
  NOR4_X1    g27968(.A1(new_n30665_), .A2(new_n8545_), .A3(pi0299), .A4(new_n30933_), .ZN(new_n31228_));
  AOI21_X1   g27969(.A1(new_n31228_), .A2(new_n31227_), .B(new_n8546_), .ZN(new_n31229_));
  OAI21_X1   g27970(.A1(new_n31227_), .A2(new_n31228_), .B(new_n31229_), .ZN(new_n31230_));
  NAND2_X1   g27971(.A1(new_n31230_), .A2(new_n31226_), .ZN(new_n31231_));
  NAND2_X1   g27972(.A1(new_n31231_), .A2(pi0211), .ZN(new_n31232_));
  NOR2_X1    g27973(.A1(new_n31090_), .A2(new_n8684_), .ZN(new_n31233_));
  XOR2_X1    g27974(.A1(new_n31232_), .A2(new_n31233_), .Z(new_n31234_));
  NAND2_X1   g27975(.A1(new_n31231_), .A2(new_n8740_), .ZN(new_n31235_));
  XOR2_X1    g27976(.A1(new_n31235_), .A2(new_n30889_), .Z(new_n31236_));
  OAI22_X1   g27977(.A1(new_n31236_), .A2(new_n31209_), .B1(new_n31234_), .B2(new_n31223_), .ZN(new_n31237_));
  INV_X1     g27978(.I(new_n30586_), .ZN(new_n31238_));
  NOR4_X1    g27979(.A1(new_n31215_), .A2(new_n8683_), .A3(new_n31238_), .A4(new_n31091_), .ZN(new_n31239_));
  AOI21_X1   g27980(.A1(new_n31237_), .A2(new_n31239_), .B(new_n31218_), .ZN(new_n31240_));
  AOI21_X1   g27981(.A1(new_n30704_), .A2(new_n8545_), .B(new_n8546_), .ZN(new_n31241_));
  INV_X1     g27982(.I(new_n31241_), .ZN(new_n31242_));
  NOR2_X1    g27983(.A1(new_n30807_), .A2(pi0207), .ZN(new_n31243_));
  NAND2_X1   g27984(.A1(new_n31242_), .A2(new_n31243_), .ZN(new_n31244_));
  AOI21_X1   g27985(.A1(new_n31244_), .A2(new_n30729_), .B(new_n30705_), .ZN(new_n31245_));
  NOR2_X1    g27986(.A1(new_n31245_), .A2(new_n14006_), .ZN(new_n31246_));
  NAND3_X1   g27987(.A1(new_n30728_), .A2(pi0207), .A3(pi1156), .ZN(new_n31247_));
  NAND3_X1   g27988(.A1(new_n30727_), .A2(pi0207), .A3(new_n13969_), .ZN(new_n31248_));
  AOI21_X1   g27989(.A1(new_n31247_), .A2(new_n31248_), .B(new_n30899_), .ZN(new_n31249_));
  NAND2_X1   g27990(.A1(new_n31249_), .A2(pi0208), .ZN(new_n31250_));
  NAND2_X1   g27991(.A1(new_n31250_), .A2(new_n30754_), .ZN(new_n31251_));
  NAND3_X1   g27992(.A1(new_n31251_), .A2(pi0207), .A3(pi1157), .ZN(new_n31252_));
  AOI21_X1   g27993(.A1(new_n31252_), .A2(new_n30758_), .B(new_n30711_), .ZN(new_n31253_));
  NAND2_X1   g27994(.A1(new_n31253_), .A2(pi1157), .ZN(new_n31254_));
  XOR2_X1    g27995(.A1(new_n31254_), .A2(new_n31246_), .Z(new_n31255_));
  OAI21_X1   g27996(.A1(new_n31255_), .A2(new_n3098_), .B(new_n30829_), .ZN(new_n31256_));
  NAND2_X1   g27997(.A1(new_n31256_), .A2(new_n8740_), .ZN(new_n31257_));
  XOR2_X1    g27998(.A1(new_n31257_), .A2(new_n30889_), .Z(new_n31258_));
  AOI21_X1   g27999(.A1(new_n30683_), .A2(pi0207), .B(new_n30807_), .ZN(new_n31259_));
  OAI22_X1   g28000(.A1(new_n30715_), .A2(new_n8546_), .B1(new_n30679_), .B2(new_n31259_), .ZN(new_n31260_));
  NAND4_X1   g28001(.A1(new_n8555_), .A2(new_n3098_), .A3(pi0199), .A4(pi1155), .ZN(new_n31262_));
  AOI21_X1   g28002(.A1(new_n31262_), .A2(new_n13778_), .B(new_n8555_), .ZN(new_n31263_));
  NOR2_X1    g28003(.A1(new_n3098_), .A2(pi1156), .ZN(new_n31264_));
  OAI21_X1   g28004(.A1(new_n31263_), .A2(pi0207), .B(new_n31264_), .ZN(new_n31265_));
  NOR3_X1    g28005(.A1(new_n31265_), .A2(new_n14006_), .A3(new_n30706_), .ZN(new_n31266_));
  NAND2_X1   g28006(.A1(new_n31260_), .A2(new_n31266_), .ZN(new_n31267_));
  XOR2_X1    g28007(.A1(new_n31246_), .A2(new_n31267_), .Z(new_n31268_));
  INV_X1     g28008(.I(new_n31268_), .ZN(new_n31269_));
  INV_X1     g28009(.I(new_n30713_), .ZN(new_n31270_));
  NAND3_X1   g28010(.A1(new_n30677_), .A2(pi1156), .A3(new_n8547_), .ZN(new_n31271_));
  NAND3_X1   g28011(.A1(new_n30899_), .A2(new_n13969_), .A3(new_n8547_), .ZN(new_n31272_));
  AOI21_X1   g28012(.A1(new_n31272_), .A2(new_n31271_), .B(new_n30682_), .ZN(new_n31273_));
  AOI21_X1   g28013(.A1(new_n31273_), .A2(pi0208), .B(pi0207), .ZN(new_n31274_));
  NOR2_X1    g28014(.A1(new_n31273_), .A2(pi0208), .ZN(new_n31275_));
  NOR3_X1    g28015(.A1(new_n31274_), .A2(new_n31275_), .A3(new_n31270_), .ZN(new_n31276_));
  NOR4_X1    g28016(.A1(new_n31274_), .A2(new_n31275_), .A3(new_n14006_), .A4(new_n30742_), .ZN(new_n31277_));
  AOI21_X1   g28017(.A1(new_n31276_), .A2(new_n14006_), .B(new_n31277_), .ZN(new_n31278_));
  AND2_X2    g28018(.A1(new_n31278_), .A2(new_n30586_), .Z(new_n31279_));
  NAND2_X1   g28019(.A1(new_n31268_), .A2(pi0211), .ZN(new_n31280_));
  INV_X1     g28020(.I(new_n30805_), .ZN(new_n31281_));
  AOI21_X1   g28021(.A1(new_n30684_), .A2(new_n31281_), .B(new_n8545_), .ZN(new_n31282_));
  NOR2_X1    g28022(.A1(new_n8546_), .A2(new_n14006_), .ZN(new_n31283_));
  INV_X1     g28023(.I(new_n31283_), .ZN(new_n31284_));
  NOR2_X1    g28024(.A1(new_n30781_), .A2(new_n31284_), .ZN(new_n31285_));
  NOR2_X1    g28025(.A1(new_n31285_), .A2(new_n31282_), .ZN(new_n31286_));
  NOR2_X1    g28026(.A1(new_n30779_), .A2(pi0207), .ZN(new_n31287_));
  INV_X1     g28027(.I(new_n31287_), .ZN(new_n31288_));
  INV_X1     g28028(.I(new_n30785_), .ZN(new_n31289_));
  NOR3_X1    g28029(.A1(new_n31289_), .A2(new_n8545_), .A3(new_n31282_), .ZN(new_n31290_));
  NOR3_X1    g28030(.A1(new_n31290_), .A2(pi1157), .A3(new_n31220_), .ZN(new_n31291_));
  NOR3_X1    g28031(.A1(new_n31286_), .A2(new_n31288_), .A3(new_n31291_), .ZN(new_n31292_));
  INV_X1     g28032(.I(new_n31292_), .ZN(new_n31293_));
  AOI21_X1   g28033(.A1(new_n31293_), .A2(new_n8684_), .B(new_n30876_), .ZN(new_n31294_));
  AOI21_X1   g28034(.A1(new_n31280_), .A2(new_n31294_), .B(new_n31279_), .ZN(new_n31295_));
  OAI21_X1   g28035(.A1(new_n31090_), .A2(pi0211), .B(pi0219), .ZN(new_n31296_));
  NOR2_X1    g28036(.A1(new_n31256_), .A2(new_n31296_), .ZN(new_n31297_));
  OAI21_X1   g28037(.A1(new_n31297_), .A2(new_n31295_), .B(new_n31269_), .ZN(new_n31298_));
  OAI21_X1   g28038(.A1(new_n31258_), .A2(new_n31298_), .B(pi0209), .ZN(new_n31299_));
  NOR2_X1    g28039(.A1(new_n7240_), .A2(new_n28364_), .ZN(new_n31300_));
  XOR2_X1    g28040(.A1(new_n31299_), .A2(new_n31300_), .Z(new_n31301_));
  OAI21_X1   g28041(.A1(new_n31301_), .A2(new_n31240_), .B(new_n28529_), .ZN(new_n31302_));
  OAI21_X1   g28042(.A1(new_n13614_), .A2(pi0211), .B(pi0219), .ZN(new_n31303_));
  NOR2_X1    g28043(.A1(new_n13778_), .A2(pi0211), .ZN(new_n31304_));
  NOR2_X1    g28044(.A1(new_n30994_), .A2(new_n31304_), .ZN(new_n31305_));
  INV_X1     g28045(.I(new_n31305_), .ZN(new_n31306_));
  OAI21_X1   g28046(.A1(new_n30983_), .A2(new_n30597_), .B(new_n8683_), .ZN(new_n31307_));
  AOI21_X1   g28047(.A1(new_n31306_), .A2(new_n30944_), .B(new_n31307_), .ZN(new_n31308_));
  AOI21_X1   g28048(.A1(pi0219), .A2(new_n30876_), .B(new_n31308_), .ZN(new_n31309_));
  NAND4_X1   g28049(.A1(new_n31302_), .A2(po1038), .A3(new_n31303_), .A4(new_n31309_), .ZN(new_n31310_));
  NAND2_X1   g28050(.A1(new_n31310_), .A2(pi0230), .ZN(new_n31311_));
  INV_X1     g28051(.I(new_n31223_), .ZN(new_n31312_));
  NOR2_X1    g28052(.A1(new_n31214_), .A2(new_n30733_), .ZN(new_n31313_));
  NOR2_X1    g28053(.A1(new_n8684_), .A2(new_n14006_), .ZN(new_n31314_));
  NOR4_X1    g28054(.A1(new_n8555_), .A2(new_n3098_), .A3(new_n13614_), .A4(pi0199), .ZN(new_n31315_));
  NOR2_X1    g28055(.A1(new_n8545_), .A2(new_n8546_), .ZN(new_n31316_));
  AND2_X2    g28056(.A1(new_n31315_), .A2(new_n31316_), .Z(new_n31317_));
  NOR2_X1    g28057(.A1(new_n30816_), .A2(new_n30694_), .ZN(new_n31318_));
  OAI21_X1   g28058(.A1(new_n31318_), .A2(new_n31317_), .B(pi1157), .ZN(new_n31319_));
  XOR2_X1    g28059(.A1(new_n31319_), .A2(new_n31314_), .Z(new_n31320_));
  NAND2_X1   g28060(.A1(new_n31214_), .A2(new_n30944_), .ZN(new_n31321_));
  OAI21_X1   g28061(.A1(new_n31320_), .A2(new_n31321_), .B(new_n8684_), .ZN(new_n31322_));
  NOR2_X1    g28062(.A1(new_n31313_), .A2(new_n30597_), .ZN(new_n31323_));
  XOR2_X1    g28063(.A1(new_n31323_), .A2(new_n30889_), .Z(new_n31324_));
  AOI22_X1   g28064(.A1(new_n31322_), .A2(new_n31313_), .B1(new_n31324_), .B2(new_n31312_), .ZN(new_n31325_));
  AOI21_X1   g28065(.A1(new_n31214_), .A2(new_n31091_), .B(new_n8683_), .ZN(new_n31326_));
  NAND2_X1   g28066(.A1(new_n31216_), .A2(new_n31326_), .ZN(new_n31327_));
  AOI21_X1   g28067(.A1(new_n31327_), .A2(new_n31223_), .B(new_n8684_), .ZN(new_n31328_));
  NOR3_X1    g28068(.A1(new_n31215_), .A2(new_n8683_), .A3(new_n31238_), .ZN(new_n31329_));
  OAI21_X1   g28069(.A1(new_n31328_), .A2(pi0209), .B(new_n31329_), .ZN(new_n31330_));
  NOR2_X1    g28070(.A1(new_n31278_), .A2(new_n31090_), .ZN(new_n31331_));
  NAND2_X1   g28071(.A1(new_n31278_), .A2(pi0211), .ZN(new_n31332_));
  NAND3_X1   g28072(.A1(new_n31332_), .A2(pi0219), .A3(new_n31090_), .ZN(new_n31333_));
  OAI21_X1   g28073(.A1(new_n31331_), .A2(new_n31333_), .B(new_n31293_), .ZN(new_n31334_));
  AOI21_X1   g28074(.A1(new_n31334_), .A2(pi0211), .B(pi0209), .ZN(new_n31335_));
  OAI21_X1   g28075(.A1(new_n31325_), .A2(new_n31330_), .B(new_n31335_), .ZN(new_n31336_));
  XOR2_X1    g28076(.A1(new_n31246_), .A2(new_n31314_), .Z(new_n31337_));
  NAND2_X1   g28077(.A1(new_n31337_), .A2(new_n31276_), .ZN(new_n31338_));
  NAND2_X1   g28078(.A1(new_n31338_), .A2(new_n30876_), .ZN(new_n31339_));
  INV_X1     g28079(.I(new_n31249_), .ZN(new_n31340_));
  NOR4_X1    g28080(.A1(new_n30735_), .A2(new_n30736_), .A3(new_n8545_), .A4(pi1156), .ZN(new_n31341_));
  OAI21_X1   g28081(.A1(new_n31341_), .A2(pi1156), .B(new_n30700_), .ZN(new_n31342_));
  AOI21_X1   g28082(.A1(new_n31340_), .A2(new_n31342_), .B(new_n31284_), .ZN(new_n31343_));
  NOR3_X1    g28083(.A1(new_n31253_), .A2(new_n30748_), .A3(new_n31343_), .ZN(new_n31344_));
  NAND3_X1   g28084(.A1(new_n31339_), .A2(pi0211), .A3(new_n31344_), .ZN(new_n31345_));
  NOR2_X1    g28085(.A1(new_n31279_), .A2(pi0219), .ZN(new_n31346_));
  NOR2_X1    g28086(.A1(new_n31292_), .A2(new_n30597_), .ZN(new_n31347_));
  XOR2_X1    g28087(.A1(new_n31347_), .A2(new_n30889_), .Z(new_n31348_));
  INV_X1     g28088(.I(new_n9213_), .ZN(new_n31349_));
  NOR3_X1    g28089(.A1(new_n30623_), .A2(new_n30916_), .A3(pi0214), .ZN(new_n31350_));
  NAND2_X1   g28090(.A1(new_n31350_), .A2(new_n31304_), .ZN(new_n31351_));
  AOI21_X1   g28091(.A1(new_n31349_), .A2(new_n30876_), .B(new_n31351_), .ZN(new_n31352_));
  OAI21_X1   g28092(.A1(new_n31352_), .A2(new_n30624_), .B(pi0212), .ZN(new_n31353_));
  NAND2_X1   g28093(.A1(new_n31353_), .A2(new_n28529_), .ZN(new_n31354_));
  NOR3_X1    g28094(.A1(new_n7240_), .A2(new_n30557_), .A3(new_n3611_), .ZN(new_n31355_));
  NAND4_X1   g28095(.A1(new_n31348_), .A2(new_n31344_), .A3(new_n31354_), .A4(new_n31355_), .ZN(new_n31356_));
  AOI21_X1   g28096(.A1(new_n31345_), .A2(new_n31346_), .B(new_n31356_), .ZN(new_n31357_));
  NAND2_X1   g28097(.A1(new_n31357_), .A2(new_n31336_), .ZN(new_n31358_));
  XOR2_X1    g28098(.A1(new_n31311_), .A2(new_n31358_), .Z(po0392));
  NOR2_X1    g28099(.A1(new_n3235_), .A2(new_n3462_), .ZN(new_n31360_));
  OAI21_X1   g28100(.A1(new_n5507_), .A2(pi0087), .B(new_n31360_), .ZN(new_n31361_));
  OAI21_X1   g28101(.A1(new_n30399_), .A2(new_n31361_), .B(new_n3455_), .ZN(new_n31362_));
  AOI22_X1   g28102(.A1(new_n31362_), .A2(new_n5488_), .B1(pi0092), .B2(new_n10621_), .ZN(new_n31363_));
  INV_X1     g28103(.I(new_n6287_), .ZN(new_n31364_));
  NOR4_X1    g28104(.A1(new_n5544_), .A2(new_n3175_), .A3(new_n8226_), .A4(new_n31364_), .ZN(new_n31365_));
  NAND3_X1   g28105(.A1(new_n31365_), .A2(new_n5491_), .A3(new_n5496_), .ZN(new_n31366_));
  NOR2_X1    g28106(.A1(new_n31363_), .A2(new_n31366_), .ZN(po0393));
  NOR2_X1    g28107(.A1(new_n30966_), .A2(new_n8555_), .ZN(new_n31368_));
  NOR2_X1    g28108(.A1(new_n31368_), .A2(pi1144), .ZN(new_n31369_));
  NOR2_X1    g28109(.A1(new_n8549_), .A2(pi1143), .ZN(new_n31370_));
  XNOR2_X1   g28110(.A1(new_n30722_), .A2(new_n31370_), .ZN(new_n31371_));
  NOR2_X1    g28111(.A1(new_n31371_), .A2(new_n3057_), .ZN(new_n31372_));
  INV_X1     g28112(.I(new_n30963_), .ZN(new_n31373_));
  OR3_X2     g28113(.A1(new_n31373_), .A2(new_n3098_), .A3(new_n30564_), .Z(new_n31374_));
  OAI22_X1   g28114(.A1(new_n31372_), .A2(new_n31374_), .B1(new_n8549_), .B2(new_n31369_), .ZN(new_n31375_));
  NOR2_X1    g28115(.A1(new_n31371_), .A2(new_n3518_), .ZN(new_n31376_));
  AND2_X2    g28116(.A1(new_n31375_), .A2(new_n31376_), .Z(new_n31377_));
  INV_X1     g28117(.I(new_n31377_), .ZN(new_n31378_));
  INV_X1     g28118(.I(new_n31126_), .ZN(new_n31379_));
  NOR2_X1    g28119(.A1(new_n3650_), .A2(pi0211), .ZN(new_n31380_));
  NAND2_X1   g28120(.A1(new_n31380_), .A2(pi0299), .ZN(new_n31381_));
  NOR2_X1    g28121(.A1(new_n30560_), .A2(new_n8739_), .ZN(new_n31382_));
  NOR2_X1    g28122(.A1(new_n8684_), .A2(pi1144), .ZN(new_n31383_));
  INV_X1     g28123(.I(new_n31383_), .ZN(new_n31384_));
  OAI21_X1   g28124(.A1(pi0211), .A2(pi1145), .B(new_n31384_), .ZN(new_n31385_));
  XOR2_X1    g28125(.A1(new_n30560_), .A2(new_n30597_), .Z(new_n31386_));
  NAND2_X1   g28126(.A1(new_n31386_), .A2(new_n31385_), .ZN(new_n31387_));
  XOR2_X1    g28127(.A1(new_n31387_), .A2(new_n31382_), .Z(new_n31388_));
  OAI22_X1   g28128(.A1(new_n31388_), .A2(new_n30620_), .B1(new_n31379_), .B2(new_n31381_), .ZN(new_n31389_));
  NAND2_X1   g28129(.A1(new_n31388_), .A2(new_n30596_), .ZN(new_n31390_));
  NOR2_X1    g28130(.A1(new_n30918_), .A2(new_n8683_), .ZN(new_n31391_));
  XOR2_X1    g28131(.A1(new_n31390_), .A2(new_n31391_), .Z(new_n31392_));
  NOR3_X1    g28132(.A1(new_n31392_), .A2(pi0211), .A3(new_n3650_), .ZN(new_n31393_));
  NAND2_X1   g28133(.A1(new_n31393_), .A2(po1038), .ZN(new_n31394_));
  AOI21_X1   g28134(.A1(new_n31394_), .A2(new_n31389_), .B(new_n31378_), .ZN(new_n31395_));
  NAND2_X1   g28135(.A1(new_n31395_), .A2(pi0213), .ZN(new_n31396_));
  NOR3_X1    g28136(.A1(new_n31003_), .A2(new_n8684_), .A3(new_n14006_), .ZN(new_n31397_));
  NOR3_X1    g28137(.A1(new_n31003_), .A2(pi0211), .A3(pi1157), .ZN(new_n31398_));
  OAI21_X1   g28138(.A1(new_n31397_), .A2(new_n31398_), .B(pi1158), .ZN(new_n31399_));
  NAND2_X1   g28139(.A1(new_n31399_), .A2(new_n31350_), .ZN(new_n31400_));
  INV_X1     g28140(.I(new_n30625_), .ZN(new_n31401_));
  AOI21_X1   g28141(.A1(new_n31349_), .A2(new_n31401_), .B(new_n31003_), .ZN(new_n31402_));
  INV_X1     g28142(.I(new_n31402_), .ZN(new_n31403_));
  NOR2_X1    g28143(.A1(po1038), .A2(pi0212), .ZN(new_n31404_));
  NOR3_X1    g28144(.A1(new_n8684_), .A2(new_n8685_), .A3(new_n13817_), .ZN(new_n31405_));
  NOR3_X1    g28145(.A1(new_n8685_), .A2(pi0211), .A3(pi1154), .ZN(new_n31406_));
  OAI21_X1   g28146(.A1(new_n31405_), .A2(new_n31406_), .B(pi1155), .ZN(new_n31407_));
  AOI21_X1   g28147(.A1(new_n31403_), .A2(new_n31404_), .B(new_n31407_), .ZN(new_n31408_));
  INV_X1     g28148(.I(new_n31408_), .ZN(new_n31409_));
  AOI21_X1   g28149(.A1(new_n31409_), .A2(new_n31400_), .B(pi0213), .ZN(new_n31410_));
  AND2_X2    g28150(.A1(new_n31410_), .A2(pi0209), .Z(new_n31411_));
  AOI21_X1   g28151(.A1(new_n31396_), .A2(new_n31411_), .B(po1038), .ZN(new_n31412_));
  NOR3_X1    g28152(.A1(new_n30611_), .A2(new_n8739_), .A3(new_n8685_), .ZN(new_n31413_));
  NOR3_X1    g28153(.A1(new_n30610_), .A2(new_n8739_), .A3(pi0214), .ZN(new_n31414_));
  OAI21_X1   g28154(.A1(new_n31413_), .A2(new_n31414_), .B(new_n30617_), .ZN(new_n31415_));
  AOI21_X1   g28155(.A1(new_n31415_), .A2(new_n30743_), .B(new_n31003_), .ZN(new_n31416_));
  NOR2_X1    g28156(.A1(new_n31400_), .A2(new_n30620_), .ZN(new_n31417_));
  OAI21_X1   g28157(.A1(new_n31377_), .A2(new_n31416_), .B(new_n31417_), .ZN(new_n31418_));
  OAI21_X1   g28158(.A1(new_n31412_), .A2(new_n31418_), .B(pi0230), .ZN(new_n31419_));
  INV_X1     g28159(.I(new_n30651_), .ZN(new_n31420_));
  NOR2_X1    g28160(.A1(new_n8555_), .A2(new_n13969_), .ZN(new_n31421_));
  NOR3_X1    g28161(.A1(new_n31420_), .A2(pi1158), .A3(new_n31421_), .ZN(new_n31422_));
  NAND3_X1   g28162(.A1(new_n31420_), .A2(new_n13929_), .A3(new_n31421_), .ZN(new_n31423_));
  INV_X1     g28163(.I(new_n31423_), .ZN(new_n31424_));
  NOR2_X1    g28164(.A1(new_n31424_), .A2(new_n31422_), .ZN(new_n31425_));
  NOR2_X1    g28165(.A1(new_n31425_), .A2(pi0299), .ZN(new_n31426_));
  NOR4_X1    g28166(.A1(new_n31171_), .A2(new_n30694_), .A3(new_n31242_), .A4(new_n31426_), .ZN(new_n31427_));
  NAND2_X1   g28167(.A1(new_n31427_), .A2(pi0211), .ZN(new_n31428_));
  INV_X1     g28168(.I(new_n31425_), .ZN(new_n31429_));
  OAI21_X1   g28169(.A1(new_n30731_), .A2(new_n8545_), .B(new_n31342_), .ZN(new_n31430_));
  NAND2_X1   g28170(.A1(new_n30747_), .A2(new_n30812_), .ZN(new_n31431_));
  AOI22_X1   g28171(.A1(new_n31430_), .A2(new_n31283_), .B1(new_n31429_), .B2(new_n31431_), .ZN(new_n31432_));
  NOR2_X1    g28172(.A1(new_n30731_), .A2(new_n8546_), .ZN(new_n31433_));
  XOR2_X1    g28173(.A1(new_n31433_), .A2(new_n9090_), .Z(new_n31434_));
  NAND2_X1   g28174(.A1(new_n8549_), .A2(new_n13969_), .ZN(new_n31435_));
  AOI22_X1   g28175(.A1(new_n31011_), .A2(new_n31435_), .B1(pi0199), .B2(pi1158), .ZN(new_n31436_));
  INV_X1     g28176(.I(new_n31436_), .ZN(new_n31437_));
  NOR3_X1    g28177(.A1(new_n31437_), .A2(pi0200), .A3(new_n8545_), .ZN(new_n31438_));
  NOR3_X1    g28178(.A1(new_n31438_), .A2(pi0208), .A3(pi1157), .ZN(new_n31439_));
  NAND2_X1   g28179(.A1(new_n30753_), .A2(new_n30733_), .ZN(new_n31440_));
  NOR4_X1    g28180(.A1(new_n31434_), .A2(new_n31432_), .A3(new_n31439_), .A4(new_n31440_), .ZN(new_n31441_));
  XOR2_X1    g28181(.A1(new_n31427_), .A2(new_n8686_), .Z(new_n31442_));
  NAND2_X1   g28182(.A1(new_n31442_), .A2(new_n31441_), .ZN(new_n31443_));
  XNOR2_X1   g28183(.A1(new_n31443_), .A2(new_n31428_), .ZN(new_n31444_));
  OAI21_X1   g28184(.A1(new_n31444_), .A2(new_n8739_), .B(new_n30718_), .ZN(new_n31445_));
  NOR2_X1    g28185(.A1(new_n31289_), .A2(pi0207), .ZN(new_n31446_));
  NOR2_X1    g28186(.A1(new_n30688_), .A2(new_n30610_), .ZN(new_n31447_));
  NOR2_X1    g28187(.A1(new_n31447_), .A2(new_n8545_), .ZN(new_n31448_));
  OAI21_X1   g28188(.A1(new_n31448_), .A2(new_n31446_), .B(pi0208), .ZN(new_n31449_));
  INV_X1     g28189(.I(new_n30965_), .ZN(new_n31450_));
  NOR3_X1    g28190(.A1(new_n31437_), .A2(new_n30735_), .A3(new_n31450_), .ZN(new_n31451_));
  NAND2_X1   g28191(.A1(new_n31451_), .A2(pi0208), .ZN(new_n31452_));
  XNOR2_X1   g28192(.A1(new_n31449_), .A2(new_n31452_), .ZN(new_n31453_));
  OAI21_X1   g28193(.A1(new_n31453_), .A2(new_n30611_), .B(new_n14006_), .ZN(new_n31454_));
  INV_X1     g28194(.I(new_n31448_), .ZN(new_n31455_));
  NAND2_X1   g28195(.A1(new_n31053_), .A2(new_n13969_), .ZN(new_n31456_));
  NOR3_X1    g28196(.A1(new_n30654_), .A2(new_n8549_), .A3(new_n13929_), .ZN(new_n31457_));
  AOI21_X1   g28197(.A1(new_n31457_), .A2(new_n31456_), .B(pi1158), .ZN(new_n31458_));
  OAI21_X1   g28198(.A1(new_n31458_), .A2(new_n8555_), .B(new_n30568_), .ZN(new_n31459_));
  NAND2_X1   g28199(.A1(new_n31459_), .A2(new_n30611_), .ZN(new_n31460_));
  NAND3_X1   g28200(.A1(new_n31460_), .A2(new_n30744_), .A3(new_n31283_), .ZN(new_n31461_));
  NAND2_X1   g28201(.A1(new_n31455_), .A2(new_n31461_), .ZN(new_n31462_));
  AND3_X2    g28202(.A1(new_n31454_), .A2(new_n31287_), .A3(new_n31462_), .Z(new_n31463_));
  NOR2_X1    g28203(.A1(new_n30687_), .A2(new_n8546_), .ZN(new_n31464_));
  XOR2_X1    g28204(.A1(new_n31464_), .A2(new_n8547_), .Z(new_n31465_));
  NOR3_X1    g28205(.A1(new_n31429_), .A2(pi0208), .A3(new_n30812_), .ZN(new_n31466_));
  INV_X1     g28206(.I(new_n31466_), .ZN(new_n31467_));
  NOR2_X1    g28207(.A1(new_n31467_), .A2(new_n30742_), .ZN(new_n31468_));
  NAND3_X1   g28208(.A1(new_n31465_), .A2(new_n8685_), .A3(new_n31468_), .ZN(new_n31469_));
  NAND2_X1   g28209(.A1(new_n31469_), .A2(new_n8739_), .ZN(new_n31470_));
  INV_X1     g28210(.I(new_n31470_), .ZN(new_n31471_));
  NAND3_X1   g28211(.A1(new_n30827_), .A2(pi0207), .A3(pi1158), .ZN(new_n31472_));
  NAND3_X1   g28212(.A1(new_n30808_), .A2(pi0207), .A3(new_n13929_), .ZN(new_n31473_));
  AOI21_X1   g28213(.A1(new_n31472_), .A2(new_n31473_), .B(new_n30688_), .ZN(new_n31474_));
  INV_X1     g28214(.I(new_n31474_), .ZN(new_n31475_));
  NOR2_X1    g28215(.A1(new_n30745_), .A2(new_n8684_), .ZN(new_n31476_));
  NOR2_X1    g28216(.A1(new_n3098_), .A2(new_n13929_), .ZN(new_n31477_));
  INV_X1     g28217(.I(new_n31477_), .ZN(new_n31478_));
  AOI21_X1   g28218(.A1(new_n31478_), .A2(new_n8773_), .B(new_n8545_), .ZN(new_n31479_));
  AOI21_X1   g28219(.A1(new_n13969_), .A2(new_n30674_), .B(new_n30654_), .ZN(new_n31480_));
  INV_X1     g28220(.I(new_n31480_), .ZN(new_n31481_));
  AOI21_X1   g28221(.A1(new_n31011_), .A2(pi1158), .B(pi1157), .ZN(new_n31482_));
  AOI21_X1   g28222(.A1(new_n8545_), .A2(new_n31482_), .B(new_n31481_), .ZN(new_n31483_));
  OAI21_X1   g28223(.A1(new_n31483_), .A2(new_n31476_), .B(new_n31479_), .ZN(new_n31484_));
  OR2_X2     g28224(.A1(new_n31484_), .A2(new_n31284_), .Z(new_n31485_));
  AOI21_X1   g28225(.A1(new_n30703_), .A2(new_n8545_), .B(new_n31478_), .ZN(new_n31486_));
  NAND2_X1   g28226(.A1(new_n31427_), .A2(new_n31486_), .ZN(new_n31487_));
  AOI21_X1   g28227(.A1(new_n31475_), .A2(new_n31485_), .B(new_n31487_), .ZN(new_n31488_));
  AOI21_X1   g28228(.A1(new_n30754_), .A2(pi0299), .B(new_n30864_), .ZN(new_n31489_));
  NOR3_X1    g28229(.A1(new_n30753_), .A2(pi0207), .A3(new_n3098_), .ZN(new_n31490_));
  OAI21_X1   g28230(.A1(new_n31489_), .A2(new_n31490_), .B(pi1158), .ZN(new_n31491_));
  NAND2_X1   g28231(.A1(new_n30651_), .A2(pi1156), .ZN(new_n31492_));
  NOR2_X1    g28232(.A1(new_n31492_), .A2(new_n30812_), .ZN(new_n31493_));
  OAI21_X1   g28233(.A1(new_n31479_), .A2(pi0208), .B(new_n31493_), .ZN(new_n31494_));
  NAND2_X1   g28234(.A1(new_n31494_), .A2(new_n14006_), .ZN(new_n31495_));
  NAND4_X1   g28235(.A1(new_n31491_), .A2(pi0208), .A3(pi0211), .A4(new_n31495_), .ZN(new_n31496_));
  OAI21_X1   g28236(.A1(new_n31475_), .A2(new_n31496_), .B(pi0214), .ZN(new_n31497_));
  OAI21_X1   g28237(.A1(new_n31488_), .A2(new_n31497_), .B(new_n31471_), .ZN(new_n31498_));
  NAND3_X1   g28238(.A1(new_n31498_), .A2(new_n8683_), .A3(new_n7240_), .ZN(new_n31499_));
  NAND3_X1   g28239(.A1(new_n31445_), .A2(new_n31463_), .A3(new_n31499_), .ZN(new_n31500_));
  NOR2_X1    g28240(.A1(new_n3098_), .A2(pi1145), .ZN(new_n31501_));
  INV_X1     g28241(.I(new_n30671_), .ZN(new_n31502_));
  NOR2_X1    g28242(.A1(new_n3098_), .A2(new_n3518_), .ZN(new_n31503_));
  OAI21_X1   g28243(.A1(new_n13817_), .A2(pi1156), .B(new_n31502_), .ZN(new_n31504_));
  AOI21_X1   g28244(.A1(new_n8772_), .A2(pi1157), .B(pi0299), .ZN(new_n31505_));
  AOI21_X1   g28245(.A1(new_n30754_), .A2(new_n31505_), .B(pi0207), .ZN(new_n31506_));
  NAND2_X1   g28246(.A1(new_n31506_), .A2(new_n8546_), .ZN(new_n31507_));
  INV_X1     g28247(.I(new_n31501_), .ZN(new_n31508_));
  NOR2_X1    g28248(.A1(new_n31508_), .A2(new_n8545_), .ZN(new_n31509_));
  AOI22_X1   g28249(.A1(new_n31507_), .A2(new_n31509_), .B1(new_n31504_), .B2(new_n31501_), .ZN(new_n31510_));
  INV_X1     g28250(.I(new_n31503_), .ZN(new_n31511_));
  NAND2_X1   g28251(.A1(pi1154), .A2(pi1156), .ZN(new_n31512_));
  AOI21_X1   g28252(.A1(new_n30856_), .A2(new_n31511_), .B(new_n31512_), .ZN(new_n31513_));
  OAI21_X1   g28253(.A1(new_n30728_), .A2(new_n31513_), .B(new_n31501_), .ZN(new_n31514_));
  OAI21_X1   g28254(.A1(new_n31510_), .A2(new_n31514_), .B(pi0211), .ZN(new_n31515_));
  NAND2_X1   g28255(.A1(new_n31438_), .A2(pi1157), .ZN(new_n31516_));
  AOI21_X1   g28256(.A1(new_n31459_), .A2(new_n8546_), .B(new_n31516_), .ZN(new_n31517_));
  NAND2_X1   g28257(.A1(new_n30754_), .A2(new_n31505_), .ZN(new_n31518_));
  NOR2_X1    g28258(.A1(new_n30869_), .A2(pi0207), .ZN(new_n31519_));
  NAND2_X1   g28259(.A1(new_n31518_), .A2(new_n31519_), .ZN(new_n31520_));
  NOR4_X1    g28260(.A1(new_n31517_), .A2(pi0208), .A3(new_n30887_), .A4(new_n31520_), .ZN(new_n31521_));
  OAI21_X1   g28261(.A1(new_n31521_), .A2(pi1144), .B(pi0299), .ZN(new_n31522_));
  INV_X1     g28262(.I(new_n30588_), .ZN(new_n31523_));
  NOR2_X1    g28263(.A1(new_n31503_), .A2(pi0208), .ZN(new_n31524_));
  NOR4_X1    g28264(.A1(new_n31482_), .A2(new_n31523_), .A3(new_n31492_), .A4(new_n31524_), .ZN(new_n31525_));
  NAND2_X1   g28265(.A1(new_n31483_), .A2(new_n31525_), .ZN(new_n31526_));
  NOR2_X1    g28266(.A1(new_n31522_), .A2(new_n31526_), .ZN(new_n31527_));
  XNOR2_X1   g28267(.A1(new_n31527_), .A2(new_n31515_), .ZN(new_n31528_));
  OAI21_X1   g28268(.A1(new_n31528_), .A2(new_n8685_), .B(new_n31471_), .ZN(new_n31529_));
  INV_X1     g28269(.I(new_n31517_), .ZN(new_n31530_));
  NOR2_X1    g28270(.A1(new_n31506_), .A2(new_n30847_), .ZN(new_n31531_));
  NAND4_X1   g28271(.A1(new_n31530_), .A2(new_n8546_), .A3(new_n30859_), .A4(new_n31531_), .ZN(new_n31532_));
  AOI21_X1   g28272(.A1(new_n31532_), .A2(new_n3650_), .B(new_n3098_), .ZN(new_n31533_));
  NAND4_X1   g28273(.A1(new_n31465_), .A2(new_n9213_), .A3(new_n30604_), .A4(new_n31468_), .ZN(new_n31534_));
  NAND3_X1   g28274(.A1(new_n31529_), .A2(new_n8683_), .A3(new_n31534_), .ZN(new_n31535_));
  NAND2_X1   g28275(.A1(new_n31522_), .A2(pi0214), .ZN(new_n31536_));
  XOR2_X1    g28276(.A1(new_n31536_), .A2(new_n30718_), .Z(new_n31537_));
  AOI21_X1   g28277(.A1(new_n31537_), .A2(new_n31533_), .B(pi0212), .ZN(new_n31538_));
  NAND2_X1   g28278(.A1(new_n31528_), .A2(pi0214), .ZN(new_n31539_));
  NOR2_X1    g28279(.A1(new_n31538_), .A2(new_n31539_), .ZN(new_n31540_));
  AOI21_X1   g28280(.A1(new_n31535_), .A2(new_n31540_), .B(new_n30910_), .ZN(new_n31541_));
  NAND2_X1   g28281(.A1(new_n31393_), .A2(new_n31410_), .ZN(new_n31542_));
  OAI21_X1   g28282(.A1(new_n31541_), .A2(new_n31542_), .B(new_n31500_), .ZN(new_n31543_));
  NAND2_X1   g28283(.A1(new_n31265_), .A2(pi1157), .ZN(new_n31544_));
  NAND4_X1   g28284(.A1(new_n31451_), .A2(new_n8545_), .A3(pi1157), .A4(new_n30706_), .ZN(new_n31545_));
  NOR2_X1    g28285(.A1(new_n30704_), .A2(new_n31545_), .ZN(new_n31546_));
  OR2_X2     g28286(.A1(new_n31546_), .A2(new_n31544_), .Z(new_n31547_));
  AOI21_X1   g28287(.A1(new_n31546_), .A2(new_n31544_), .B(pi0208), .ZN(new_n31548_));
  NAND2_X1   g28288(.A1(new_n31150_), .A2(pi0207), .ZN(new_n31549_));
  AOI21_X1   g28289(.A1(new_n31547_), .A2(new_n31548_), .B(new_n31549_), .ZN(new_n31550_));
  NOR2_X1    g28290(.A1(new_n31451_), .A2(pi1157), .ZN(new_n31551_));
  OAI21_X1   g28291(.A1(pi0208), .A2(new_n30613_), .B(new_n31551_), .ZN(new_n31552_));
  OAI21_X1   g28292(.A1(new_n31552_), .A2(new_n31459_), .B(pi0214), .ZN(new_n31553_));
  OAI21_X1   g28293(.A1(new_n31550_), .A2(new_n31553_), .B(new_n8739_), .ZN(new_n31554_));
  NAND3_X1   g28294(.A1(new_n31463_), .A2(pi0214), .A3(new_n31554_), .ZN(new_n31555_));
  NAND4_X1   g28295(.A1(new_n31465_), .A2(pi0219), .A3(new_n30604_), .A4(new_n31468_), .ZN(new_n31556_));
  NAND2_X1   g28296(.A1(new_n31556_), .A2(new_n8684_), .ZN(new_n31557_));
  NAND3_X1   g28297(.A1(new_n31557_), .A2(pi0230), .A3(pi0237), .ZN(new_n31558_));
  AOI21_X1   g28298(.A1(new_n31441_), .A2(new_n30874_), .B(new_n31558_), .ZN(new_n31559_));
  NAND3_X1   g28299(.A1(new_n31543_), .A2(new_n31555_), .A3(new_n31559_), .ZN(new_n31560_));
  XOR2_X1    g28300(.A1(new_n31560_), .A2(new_n31419_), .Z(po0394));
  NOR2_X1    g28301(.A1(new_n30654_), .A2(new_n30950_), .ZN(new_n31562_));
  NOR2_X1    g28302(.A1(new_n31562_), .A2(new_n8545_), .ZN(new_n31563_));
  NAND3_X1   g28303(.A1(new_n30664_), .A2(pi0207), .A3(new_n31064_), .ZN(new_n31564_));
  NAND2_X1   g28304(.A1(new_n31564_), .A2(new_n31563_), .ZN(new_n31565_));
  NAND4_X1   g28305(.A1(new_n30664_), .A2(pi0207), .A3(new_n31064_), .A4(new_n31562_), .ZN(new_n31566_));
  NAND3_X1   g28306(.A1(new_n31565_), .A2(pi0208), .A3(new_n31566_), .ZN(new_n31567_));
  NAND2_X1   g28307(.A1(new_n31226_), .A2(new_n31567_), .ZN(new_n31568_));
  INV_X1     g28308(.I(new_n31211_), .ZN(new_n31569_));
  AOI21_X1   g28309(.A1(new_n13614_), .A2(new_n30614_), .B(new_n30652_), .ZN(new_n31570_));
  OAI21_X1   g28310(.A1(new_n31064_), .A2(new_n31569_), .B(new_n31570_), .ZN(new_n31571_));
  NOR2_X1    g28311(.A1(new_n30723_), .A2(pi0207), .ZN(new_n31572_));
  AOI21_X1   g28312(.A1(new_n31571_), .A2(new_n31572_), .B(new_n31111_), .ZN(new_n31573_));
  OAI21_X1   g28313(.A1(new_n31573_), .A2(pi0207), .B(new_n30762_), .ZN(new_n31574_));
  NAND2_X1   g28314(.A1(new_n30774_), .A2(new_n31574_), .ZN(new_n31575_));
  NOR3_X1    g28315(.A1(new_n31575_), .A2(pi0211), .A3(pi0214), .ZN(new_n31576_));
  NOR2_X1    g28316(.A1(new_n31206_), .A2(new_n31203_), .ZN(new_n31577_));
  NOR2_X1    g28317(.A1(new_n30669_), .A2(new_n13614_), .ZN(new_n31578_));
  INV_X1     g28318(.I(new_n31578_), .ZN(new_n31579_));
  NOR3_X1    g28319(.A1(new_n30815_), .A2(new_n8545_), .A3(new_n31579_), .ZN(new_n31580_));
  NOR3_X1    g28320(.A1(new_n31580_), .A2(new_n8545_), .A3(new_n31015_), .ZN(new_n31581_));
  INV_X1     g28321(.I(new_n31015_), .ZN(new_n31582_));
  NOR4_X1    g28322(.A1(new_n30815_), .A2(new_n8545_), .A3(new_n31582_), .A4(new_n31579_), .ZN(new_n31583_));
  NOR3_X1    g28323(.A1(new_n31581_), .A2(new_n8546_), .A3(new_n31583_), .ZN(new_n31584_));
  NOR2_X1    g28324(.A1(new_n31577_), .A2(new_n31584_), .ZN(new_n31585_));
  OAI21_X1   g28325(.A1(new_n31585_), .A2(new_n30718_), .B(pi0212), .ZN(new_n31586_));
  NOR2_X1    g28326(.A1(new_n31003_), .A2(new_n8684_), .ZN(new_n31587_));
  NAND2_X1   g28327(.A1(new_n31568_), .A2(new_n30874_), .ZN(new_n31588_));
  XOR2_X1    g28328(.A1(new_n31588_), .A2(new_n31587_), .Z(new_n31589_));
  NAND2_X1   g28329(.A1(new_n31575_), .A2(pi0219), .ZN(new_n31590_));
  OAI22_X1   g28330(.A1(new_n31589_), .A2(new_n31590_), .B1(new_n31576_), .B2(new_n31586_), .ZN(new_n31591_));
  NOR2_X1    g28331(.A1(new_n8684_), .A2(pi0214), .ZN(new_n31592_));
  NOR2_X1    g28332(.A1(new_n30640_), .A2(new_n31592_), .ZN(new_n31593_));
  INV_X1     g28333(.I(new_n31593_), .ZN(new_n31594_));
  NAND3_X1   g28334(.A1(new_n31591_), .A2(new_n31568_), .A3(new_n31594_), .ZN(new_n31595_));
  NOR3_X1    g28335(.A1(new_n31213_), .A2(new_n8547_), .A3(new_n31562_), .ZN(new_n31596_));
  NOR2_X1    g28336(.A1(new_n31596_), .A2(new_n31582_), .ZN(new_n31597_));
  OAI21_X1   g28337(.A1(po1038), .A2(new_n31238_), .B(new_n31597_), .ZN(new_n31598_));
  NAND3_X1   g28338(.A1(new_n31595_), .A2(new_n28364_), .A3(new_n31598_), .ZN(new_n31599_));
  NOR2_X1    g28339(.A1(new_n30966_), .A2(new_n8773_), .ZN(new_n31600_));
  NOR2_X1    g28340(.A1(new_n31600_), .A2(pi0299), .ZN(new_n31601_));
  NOR2_X1    g28341(.A1(new_n31601_), .A2(new_n30588_), .ZN(new_n31602_));
  NOR2_X1    g28342(.A1(new_n31013_), .A2(new_n30966_), .ZN(new_n31603_));
  NOR2_X1    g28343(.A1(new_n31603_), .A2(pi0214), .ZN(new_n31604_));
  NAND2_X1   g28344(.A1(new_n31604_), .A2(pi0212), .ZN(new_n31605_));
  NOR2_X1    g28345(.A1(new_n31605_), .A2(new_n31602_), .ZN(new_n31606_));
  INV_X1     g28346(.I(new_n31606_), .ZN(new_n31607_));
  NOR2_X1    g28347(.A1(new_n31607_), .A2(new_n13614_), .ZN(new_n31608_));
  NOR2_X1    g28348(.A1(new_n31608_), .A2(new_n30892_), .ZN(new_n31609_));
  NOR2_X1    g28349(.A1(po1038), .A2(pi1151), .ZN(new_n31610_));
  NAND2_X1   g28350(.A1(new_n31610_), .A2(pi1152), .ZN(new_n31611_));
  OAI21_X1   g28351(.A1(new_n31609_), .A2(new_n31611_), .B(new_n8683_), .ZN(new_n31612_));
  INV_X1     g28352(.I(new_n31603_), .ZN(new_n31613_));
  NOR2_X1    g28353(.A1(new_n31613_), .A2(new_n13614_), .ZN(new_n31614_));
  NOR2_X1    g28354(.A1(new_n31306_), .A2(new_n3098_), .ZN(new_n31615_));
  OAI21_X1   g28355(.A1(new_n31614_), .A2(new_n31091_), .B(new_n31615_), .ZN(new_n31616_));
  NOR3_X1    g28356(.A1(new_n31601_), .A2(new_n8684_), .A3(new_n13614_), .ZN(new_n31617_));
  NOR2_X1    g28357(.A1(new_n31617_), .A2(new_n8740_), .ZN(new_n31618_));
  NAND2_X1   g28358(.A1(new_n31616_), .A2(new_n31618_), .ZN(new_n31619_));
  INV_X1     g28359(.I(new_n31614_), .ZN(new_n31620_));
  NAND2_X1   g28360(.A1(new_n31620_), .A2(new_n30614_), .ZN(new_n31621_));
  NAND4_X1   g28361(.A1(new_n31612_), .A2(new_n8684_), .A3(new_n31619_), .A4(new_n31621_), .ZN(new_n31622_));
  NAND2_X1   g28362(.A1(new_n30706_), .A2(pi0211), .ZN(new_n31623_));
  NOR2_X1    g28363(.A1(new_n31062_), .A2(new_n8546_), .ZN(new_n31624_));
  NOR2_X1    g28364(.A1(new_n31053_), .A2(new_n30694_), .ZN(new_n31625_));
  AOI21_X1   g28365(.A1(new_n31624_), .A2(new_n31625_), .B(pi0207), .ZN(new_n31626_));
  NOR2_X1    g28366(.A1(new_n31626_), .A2(new_n31062_), .ZN(new_n31627_));
  NAND2_X1   g28367(.A1(new_n31627_), .A2(pi0211), .ZN(new_n31628_));
  XOR2_X1    g28368(.A1(new_n31628_), .A2(new_n31623_), .Z(new_n31629_));
  AOI21_X1   g28369(.A1(new_n31629_), .A2(new_n30806_), .B(new_n31091_), .ZN(new_n31630_));
  NAND2_X1   g28370(.A1(new_n31031_), .A2(pi0208), .ZN(new_n31631_));
  NOR2_X1    g28371(.A1(new_n31032_), .A2(pi0207), .ZN(new_n31632_));
  NOR2_X1    g28372(.A1(new_n8775_), .A2(new_n8545_), .ZN(new_n31633_));
  OAI21_X1   g28373(.A1(new_n31632_), .A2(new_n31633_), .B(new_n30693_), .ZN(new_n31634_));
  NAND4_X1   g28374(.A1(new_n31634_), .A2(new_n8684_), .A3(new_n30706_), .A4(new_n31631_), .ZN(new_n31635_));
  OAI21_X1   g28375(.A1(new_n31635_), .A2(new_n30597_), .B(new_n8684_), .ZN(new_n31636_));
  NAND2_X1   g28376(.A1(new_n31634_), .A2(new_n31631_), .ZN(new_n31637_));
  NOR2_X1    g28377(.A1(new_n31637_), .A2(new_n31091_), .ZN(new_n31638_));
  AOI21_X1   g28378(.A1(new_n8773_), .A2(new_n31203_), .B(new_n9090_), .ZN(new_n31639_));
  NAND2_X1   g28379(.A1(pi0200), .A2(pi0207), .ZN(new_n31640_));
  NAND2_X1   g28380(.A1(new_n31640_), .A2(new_n8549_), .ZN(new_n31641_));
  AOI21_X1   g28381(.A1(new_n31641_), .A2(new_n3098_), .B(new_n8546_), .ZN(new_n31642_));
  INV_X1     g28382(.I(new_n31642_), .ZN(new_n31643_));
  NOR2_X1    g28383(.A1(new_n9214_), .A2(new_n13614_), .ZN(new_n31644_));
  NOR3_X1    g28384(.A1(new_n9258_), .A2(new_n31644_), .A3(new_n8545_), .ZN(new_n31645_));
  AOI21_X1   g28385(.A1(new_n8545_), .A2(new_n31203_), .B(new_n31645_), .ZN(new_n31646_));
  NOR2_X1    g28386(.A1(new_n31646_), .A2(new_n31643_), .ZN(new_n31647_));
  NOR2_X1    g28387(.A1(new_n31647_), .A2(new_n31639_), .ZN(new_n31648_));
  INV_X1     g28388(.I(new_n31648_), .ZN(new_n31649_));
  NAND3_X1   g28389(.A1(new_n31636_), .A2(new_n31638_), .A3(new_n31649_), .ZN(new_n31650_));
  INV_X1     g28390(.I(new_n31610_), .ZN(new_n31651_));
  OAI21_X1   g28391(.A1(new_n9209_), .A2(pi0208), .B(pi0207), .ZN(new_n31652_));
  AOI21_X1   g28392(.A1(new_n8555_), .A2(new_n13614_), .B(new_n9090_), .ZN(new_n31653_));
  NOR2_X1    g28393(.A1(new_n31203_), .A2(pi0211), .ZN(new_n31654_));
  NAND2_X1   g28394(.A1(new_n31238_), .A2(pi0219), .ZN(new_n31655_));
  NOR4_X1    g28395(.A1(new_n31651_), .A2(new_n31653_), .A3(new_n31654_), .A4(new_n31655_), .ZN(new_n31656_));
  OAI21_X1   g28396(.A1(new_n31656_), .A2(pi0219), .B(new_n31305_), .ZN(new_n31657_));
  AOI21_X1   g28397(.A1(new_n31650_), .A2(new_n3098_), .B(new_n31657_), .ZN(new_n31658_));
  NOR2_X1    g28398(.A1(new_n8773_), .A2(new_n8545_), .ZN(new_n31659_));
  INV_X1     g28399(.I(new_n31659_), .ZN(new_n31660_));
  AOI21_X1   g28400(.A1(new_n8546_), .A2(new_n30738_), .B(new_n31660_), .ZN(new_n31661_));
  NOR2_X1    g28401(.A1(new_n30652_), .A2(new_n30812_), .ZN(new_n31662_));
  NOR2_X1    g28402(.A1(new_n31661_), .A2(new_n31662_), .ZN(new_n31663_));
  INV_X1     g28403(.I(new_n31663_), .ZN(new_n31664_));
  NAND3_X1   g28404(.A1(new_n31635_), .A2(new_n30597_), .A3(new_n31664_), .ZN(new_n31665_));
  AOI21_X1   g28405(.A1(new_n31665_), .A2(new_n31617_), .B(pi0219), .ZN(new_n31666_));
  NOR2_X1    g28406(.A1(new_n31664_), .A2(pi0214), .ZN(new_n31667_));
  AOI21_X1   g28407(.A1(new_n31667_), .A2(new_n31620_), .B(pi0212), .ZN(new_n31668_));
  INV_X1     g28408(.I(new_n31668_), .ZN(new_n31669_));
  INV_X1     g28409(.I(pi1151), .ZN(new_n31670_));
  NOR2_X1    g28410(.A1(po1038), .A2(new_n31670_), .ZN(new_n31671_));
  NOR3_X1    g28411(.A1(new_n31663_), .A2(pi0219), .A3(new_n31671_), .ZN(new_n31672_));
  NAND3_X1   g28412(.A1(new_n31608_), .A2(pi0209), .A3(pi0214), .ZN(new_n31673_));
  NOR4_X1    g28413(.A1(new_n31673_), .A2(new_n31666_), .A3(new_n31669_), .A4(new_n31672_), .ZN(new_n31674_));
  OAI21_X1   g28414(.A1(pi1152), .A2(new_n31658_), .B(new_n31674_), .ZN(new_n31675_));
  OAI21_X1   g28415(.A1(new_n31630_), .A2(new_n31675_), .B(new_n31622_), .ZN(new_n31676_));
  NOR2_X1    g28416(.A1(pi0207), .A2(pi0208), .ZN(new_n31677_));
  NOR2_X1    g28417(.A1(new_n30735_), .A2(new_n31677_), .ZN(new_n31678_));
  NOR2_X1    g28418(.A1(new_n31007_), .A2(new_n31678_), .ZN(new_n31679_));
  INV_X1     g28419(.I(new_n31679_), .ZN(new_n31680_));
  AOI21_X1   g28420(.A1(new_n31680_), .A2(new_n8685_), .B(pi0212), .ZN(new_n31681_));
  INV_X1     g28421(.I(new_n31681_), .ZN(new_n31682_));
  INV_X1     g28422(.I(new_n31050_), .ZN(new_n31683_));
  NOR3_X1    g28423(.A1(new_n31679_), .A2(pi0212), .A3(new_n31594_), .ZN(new_n31684_));
  NAND2_X1   g28424(.A1(new_n8686_), .A2(new_n30613_), .ZN(new_n31685_));
  OAI21_X1   g28425(.A1(new_n31684_), .A2(new_n31685_), .B(new_n31683_), .ZN(new_n31686_));
  AOI21_X1   g28426(.A1(new_n30652_), .A2(new_n30568_), .B(new_n8546_), .ZN(new_n31687_));
  OAI21_X1   g28427(.A1(new_n31687_), .A2(new_n30735_), .B(pi0207), .ZN(new_n31688_));
  AOI21_X1   g28428(.A1(new_n30756_), .A2(new_n8545_), .B(new_n8555_), .ZN(new_n31689_));
  INV_X1     g28429(.I(new_n31689_), .ZN(new_n31690_));
  AND2_X2    g28430(.A1(new_n31688_), .A2(new_n31690_), .Z(new_n31691_));
  INV_X1     g28431(.I(new_n31691_), .ZN(new_n31692_));
  NOR2_X1    g28432(.A1(new_n31692_), .A2(new_n8683_), .ZN(new_n31693_));
  AOI21_X1   g28433(.A1(new_n31693_), .A2(new_n31686_), .B(new_n30838_), .ZN(new_n31694_));
  INV_X1     g28434(.I(new_n31678_), .ZN(new_n31695_));
  NOR2_X1    g28435(.A1(new_n31695_), .A2(new_n8684_), .ZN(new_n31696_));
  AOI21_X1   g28436(.A1(new_n31691_), .A2(new_n8684_), .B(new_n31696_), .ZN(new_n31697_));
  AND2_X2    g28437(.A1(new_n31697_), .A2(new_n31683_), .Z(new_n31698_));
  NOR2_X1    g28438(.A1(new_n31680_), .A2(new_n31238_), .ZN(new_n31699_));
  INV_X1     g28439(.I(new_n31699_), .ZN(new_n31700_));
  NOR2_X1    g28440(.A1(new_n31698_), .A2(new_n31700_), .ZN(new_n31701_));
  INV_X1     g28441(.I(new_n31701_), .ZN(new_n31702_));
  NAND2_X1   g28442(.A1(new_n31702_), .A2(pi0219), .ZN(new_n31703_));
  INV_X1     g28443(.I(new_n31016_), .ZN(new_n31704_));
  AOI21_X1   g28444(.A1(new_n13614_), .A2(new_n30666_), .B(new_n30764_), .ZN(new_n31706_));
  AOI21_X1   g28445(.A1(new_n30652_), .A2(new_n30568_), .B(new_n8546_), .ZN(new_n31708_));
  NAND4_X1   g28446(.A1(new_n31703_), .A2(new_n30762_), .A3(new_n31671_), .A4(new_n31708_), .ZN(new_n31709_));
  OAI21_X1   g28447(.A1(new_n31709_), .A2(new_n31694_), .B(new_n31682_), .ZN(new_n31710_));
  AOI21_X1   g28448(.A1(new_n31708_), .A2(new_n30762_), .B(new_n8685_), .ZN(new_n31711_));
  NOR2_X1    g28449(.A1(new_n8685_), .A2(new_n3098_), .ZN(new_n31712_));
  XOR2_X1    g28450(.A1(new_n31711_), .A2(new_n31712_), .Z(new_n31713_));
  NAND4_X1   g28451(.A1(new_n31676_), .A2(new_n31710_), .A3(new_n31305_), .A4(new_n31713_), .ZN(new_n31714_));
  NOR4_X1    g28452(.A1(new_n28529_), .A2(new_n8683_), .A3(pi0211), .A4(pi1153), .ZN(new_n31715_));
  OAI21_X1   g28453(.A1(new_n31308_), .A2(new_n30596_), .B(new_n31715_), .ZN(new_n31716_));
  NAND2_X1   g28454(.A1(new_n31585_), .A2(new_n8684_), .ZN(new_n31717_));
  OAI21_X1   g28455(.A1(new_n8684_), .A2(new_n31597_), .B(new_n31717_), .ZN(new_n31718_));
  NAND2_X1   g28456(.A1(new_n31718_), .A2(new_n31126_), .ZN(new_n31719_));
  AOI21_X1   g28457(.A1(new_n31714_), .A2(new_n31716_), .B(new_n31719_), .ZN(new_n31720_));
  AOI21_X1   g28458(.A1(new_n31599_), .A2(new_n31720_), .B(new_n30557_), .ZN(new_n31721_));
  NOR2_X1    g28459(.A1(new_n30876_), .A2(pi0211), .ZN(new_n31722_));
  INV_X1     g28460(.I(new_n31722_), .ZN(new_n31723_));
  NOR2_X1    g28461(.A1(new_n31723_), .A2(new_n13614_), .ZN(new_n31724_));
  INV_X1     g28462(.I(new_n31724_), .ZN(new_n31725_));
  NAND2_X1   g28463(.A1(new_n30596_), .A2(pi1151), .ZN(new_n31726_));
  AOI21_X1   g28464(.A1(new_n31726_), .A2(new_n8688_), .B(new_n31725_), .ZN(new_n31727_));
  INV_X1     g28465(.I(new_n31727_), .ZN(new_n31728_));
  INV_X1     g28466(.I(new_n31597_), .ZN(new_n31729_));
  AOI21_X1   g28467(.A1(new_n30814_), .A2(new_n30692_), .B(new_n31571_), .ZN(new_n31730_));
  NOR2_X1    g28468(.A1(new_n31318_), .A2(new_n31730_), .ZN(new_n31731_));
  INV_X1     g28469(.I(new_n31731_), .ZN(new_n31732_));
  NOR2_X1    g28470(.A1(new_n31732_), .A2(new_n8684_), .ZN(new_n31733_));
  INV_X1     g28471(.I(new_n31733_), .ZN(new_n31734_));
  NAND2_X1   g28472(.A1(new_n31717_), .A2(new_n31734_), .ZN(new_n31735_));
  NOR2_X1    g28473(.A1(new_n31735_), .A2(new_n8685_), .ZN(new_n31736_));
  XOR2_X1    g28474(.A1(new_n31736_), .A2(new_n30597_), .Z(new_n31737_));
  OAI21_X1   g28475(.A1(new_n31737_), .A2(new_n31729_), .B(new_n8683_), .ZN(new_n31738_));
  AOI21_X1   g28476(.A1(new_n9077_), .A2(new_n13614_), .B(new_n30889_), .ZN(new_n31739_));
  NAND2_X1   g28477(.A1(new_n8687_), .A2(new_n30892_), .ZN(new_n31740_));
  INV_X1     g28478(.I(new_n31740_), .ZN(new_n31741_));
  NOR2_X1    g28479(.A1(po1038), .A2(pi1151), .ZN(new_n31742_));
  OAI21_X1   g28480(.A1(new_n31597_), .A2(new_n8683_), .B(new_n31742_), .ZN(new_n31743_));
  NAND2_X1   g28481(.A1(new_n31738_), .A2(new_n31743_), .ZN(new_n31744_));
  NOR2_X1    g28482(.A1(new_n31597_), .A2(new_n8684_), .ZN(new_n31745_));
  AOI21_X1   g28483(.A1(new_n8684_), .A2(new_n31731_), .B(new_n31745_), .ZN(new_n31746_));
  NAND2_X1   g28484(.A1(new_n31746_), .A2(pi0212), .ZN(new_n31747_));
  XOR2_X1    g28485(.A1(new_n31747_), .A2(new_n8740_), .Z(new_n31748_));
  AOI21_X1   g28486(.A1(new_n31717_), .A2(new_n31734_), .B(new_n31748_), .ZN(new_n31749_));
  NAND2_X1   g28487(.A1(new_n28364_), .A2(new_n31002_), .ZN(new_n31750_));
  AOI21_X1   g28488(.A1(new_n31744_), .A2(new_n31749_), .B(new_n31750_), .ZN(new_n31751_));
  NAND3_X1   g28489(.A1(new_n31746_), .A2(new_n8740_), .A3(new_n31729_), .ZN(new_n31752_));
  NOR3_X1    g28490(.A1(new_n31746_), .A2(new_n30597_), .A3(new_n31729_), .ZN(new_n31753_));
  NOR2_X1    g28491(.A1(new_n31753_), .A2(new_n8683_), .ZN(new_n31754_));
  AOI21_X1   g28492(.A1(new_n31754_), .A2(new_n31752_), .B(po1038), .ZN(new_n31755_));
  NOR2_X1    g28493(.A1(new_n7240_), .A2(new_n31740_), .ZN(new_n31756_));
  INV_X1     g28494(.I(new_n31756_), .ZN(new_n31757_));
  NOR2_X1    g28495(.A1(new_n30918_), .A2(new_n8689_), .ZN(new_n31758_));
  NOR2_X1    g28496(.A1(new_n31758_), .A2(pi1151), .ZN(new_n31759_));
  NOR3_X1    g28497(.A1(new_n31759_), .A2(new_n31739_), .A3(new_n31757_), .ZN(new_n31760_));
  NAND2_X1   g28498(.A1(new_n31755_), .A2(new_n31760_), .ZN(new_n31761_));
  NAND2_X1   g28499(.A1(new_n31738_), .A2(new_n31761_), .ZN(new_n31762_));
  NOR2_X1    g28500(.A1(new_n7240_), .A2(pi0219), .ZN(new_n31763_));
  AOI21_X1   g28501(.A1(new_n31763_), .A2(new_n31724_), .B(pi1151), .ZN(new_n31764_));
  NOR2_X1    g28502(.A1(new_n30876_), .A2(pi0219), .ZN(new_n31765_));
  INV_X1     g28503(.I(new_n31765_), .ZN(new_n31766_));
  NOR2_X1    g28504(.A1(new_n31718_), .A2(new_n31766_), .ZN(new_n31767_));
  NAND2_X1   g28505(.A1(po1038), .A2(new_n31765_), .ZN(new_n31768_));
  XOR2_X1    g28506(.A1(new_n31767_), .A2(new_n31768_), .Z(new_n31769_));
  OAI21_X1   g28507(.A1(new_n31769_), .A2(new_n31729_), .B(new_n31764_), .ZN(new_n31770_));
  NOR2_X1    g28508(.A1(new_n31735_), .A2(new_n8739_), .ZN(new_n31771_));
  XOR2_X1    g28509(.A1(new_n31771_), .A2(new_n8740_), .Z(new_n31772_));
  NOR2_X1    g28510(.A1(new_n31732_), .A2(pi1152), .ZN(new_n31773_));
  NAND4_X1   g28511(.A1(new_n31762_), .A2(new_n31770_), .A3(new_n31772_), .A4(new_n31773_), .ZN(new_n31774_));
  OAI21_X1   g28512(.A1(new_n31774_), .A2(new_n31751_), .B(new_n31728_), .ZN(new_n31775_));
  OAI21_X1   g28513(.A1(pi0211), .A2(new_n31597_), .B(new_n31734_), .ZN(new_n31776_));
  NOR2_X1    g28514(.A1(new_n31718_), .A2(new_n8739_), .ZN(new_n31777_));
  XOR2_X1    g28515(.A1(new_n31777_), .A2(new_n8740_), .Z(new_n31778_));
  AOI22_X1   g28516(.A1(new_n31778_), .A2(new_n31776_), .B1(pi0219), .B2(new_n31755_), .ZN(new_n31779_));
  NOR2_X1    g28517(.A1(new_n31718_), .A2(new_n8685_), .ZN(new_n31780_));
  XOR2_X1    g28518(.A1(new_n31780_), .A2(new_n30597_), .Z(new_n31781_));
  NOR3_X1    g28519(.A1(new_n31779_), .A2(new_n31729_), .A3(new_n31781_), .ZN(new_n31782_));
  NAND2_X1   g28520(.A1(new_n31775_), .A2(new_n31782_), .ZN(new_n31783_));
  NOR2_X1    g28521(.A1(new_n31614_), .A2(new_n30588_), .ZN(new_n31784_));
  INV_X1     g28522(.I(new_n31784_), .ZN(new_n31785_));
  AOI21_X1   g28523(.A1(new_n31785_), .A2(new_n30597_), .B(new_n31680_), .ZN(new_n31786_));
  INV_X1     g28524(.I(new_n31786_), .ZN(new_n31787_));
  AOI21_X1   g28525(.A1(new_n31698_), .A2(new_n30875_), .B(new_n8683_), .ZN(new_n31788_));
  OAI21_X1   g28526(.A1(new_n31702_), .A2(new_n31787_), .B(new_n31788_), .ZN(new_n31789_));
  XOR2_X1    g28527(.A1(new_n31789_), .A2(new_n31349_), .Z(new_n31790_));
  AOI21_X1   g28528(.A1(new_n31756_), .A2(new_n31739_), .B(pi1151), .ZN(new_n31791_));
  NAND2_X1   g28529(.A1(new_n31653_), .A2(new_n30876_), .ZN(new_n31792_));
  NOR2_X1    g28530(.A1(pi0219), .A2(pi0299), .ZN(new_n31793_));
  NAND2_X1   g28531(.A1(new_n30597_), .A2(new_n31793_), .ZN(new_n31794_));
  NAND4_X1   g28532(.A1(new_n31638_), .A2(pi0211), .A3(new_n31792_), .A4(new_n31794_), .ZN(new_n31795_));
  AOI21_X1   g28533(.A1(new_n31795_), .A2(new_n31648_), .B(new_n8684_), .ZN(new_n31796_));
  INV_X1     g28534(.I(new_n31653_), .ZN(new_n31797_));
  NOR2_X1    g28535(.A1(new_n31797_), .A2(new_n8683_), .ZN(new_n31798_));
  OAI21_X1   g28536(.A1(new_n31796_), .A2(po1038), .B(new_n31798_), .ZN(new_n31799_));
  INV_X1     g28537(.I(new_n10253_), .ZN(new_n31800_));
  AOI21_X1   g28538(.A1(new_n31700_), .A2(new_n31800_), .B(new_n31620_), .ZN(new_n31801_));
  INV_X1     g28539(.I(new_n31604_), .ZN(new_n31802_));
  NOR2_X1    g28540(.A1(pi0212), .A2(pi0219), .ZN(new_n31803_));
  AOI21_X1   g28541(.A1(new_n31785_), .A2(new_n31803_), .B(new_n31802_), .ZN(new_n31804_));
  INV_X1     g28542(.I(new_n31804_), .ZN(new_n31805_));
  INV_X1     g28543(.I(new_n31654_), .ZN(new_n31806_));
  OAI21_X1   g28544(.A1(new_n31003_), .A2(new_n31806_), .B(new_n31613_), .ZN(new_n31807_));
  NAND2_X1   g28545(.A1(new_n31608_), .A2(new_n31604_), .ZN(new_n31808_));
  AOI21_X1   g28546(.A1(new_n31805_), .A2(new_n31807_), .B(new_n31808_), .ZN(new_n31809_));
  AOI21_X1   g28547(.A1(new_n31613_), .A2(pi0219), .B(po1038), .ZN(new_n31810_));
  NAND3_X1   g28548(.A1(new_n31801_), .A2(pi1152), .A3(new_n31727_), .ZN(new_n31812_));
  AOI21_X1   g28549(.A1(new_n31799_), .A2(new_n31791_), .B(new_n31812_), .ZN(new_n31813_));
  AOI21_X1   g28550(.A1(new_n31790_), .A2(new_n31813_), .B(new_n31760_), .ZN(new_n31814_));
  AOI22_X1   g28551(.A1(new_n31627_), .A2(pi1153), .B1(pi0211), .B2(new_n31601_), .ZN(new_n31815_));
  INV_X1     g28552(.I(new_n31627_), .ZN(new_n31816_));
  NOR2_X1    g28553(.A1(new_n31664_), .A2(new_n31614_), .ZN(new_n31817_));
  INV_X1     g28554(.I(new_n31817_), .ZN(new_n31818_));
  AOI21_X1   g28555(.A1(new_n31816_), .A2(new_n8684_), .B(new_n31818_), .ZN(new_n31819_));
  NAND2_X1   g28556(.A1(new_n31620_), .A2(pi0214), .ZN(new_n31820_));
  NAND3_X1   g28557(.A1(new_n31819_), .A2(pi0214), .A3(new_n31663_), .ZN(new_n31821_));
  XNOR2_X1   g28558(.A1(new_n31821_), .A2(new_n31820_), .ZN(new_n31822_));
  AND2_X2    g28559(.A1(new_n31822_), .A2(new_n8739_), .Z(new_n31823_));
  OAI21_X1   g28560(.A1(new_n31823_), .A2(new_n9213_), .B(new_n31819_), .ZN(new_n31824_));
  INV_X1     g28561(.I(new_n31824_), .ZN(new_n31825_));
  INV_X1     g28562(.I(new_n31667_), .ZN(new_n31826_));
  NOR2_X1    g28563(.A1(new_n31815_), .A2(new_n31826_), .ZN(new_n31827_));
  OAI21_X1   g28564(.A1(new_n31816_), .A2(new_n8685_), .B(pi0212), .ZN(new_n31828_));
  OAI21_X1   g28565(.A1(new_n31827_), .A2(new_n31828_), .B(new_n8683_), .ZN(new_n31829_));
  NOR2_X1    g28566(.A1(new_n31825_), .A2(new_n31829_), .ZN(new_n31830_));
  NOR2_X1    g28567(.A1(new_n31663_), .A2(pi0214), .ZN(new_n31831_));
  INV_X1     g28568(.I(new_n31831_), .ZN(new_n31832_));
  NOR2_X1    g28569(.A1(new_n31668_), .A2(new_n31832_), .ZN(new_n31833_));
  NOR4_X1    g28570(.A1(new_n31830_), .A2(new_n31814_), .A3(new_n31815_), .A4(new_n31833_), .ZN(new_n31834_));
  NAND4_X1   g28571(.A1(new_n31834_), .A2(pi0209), .A3(pi0230), .A4(pi0238), .ZN(new_n31835_));
  AOI21_X1   g28572(.A1(new_n31783_), .A2(new_n28529_), .B(new_n31835_), .ZN(new_n31836_));
  XOR2_X1    g28573(.A1(new_n31836_), .A2(new_n31721_), .Z(po0395));
  NOR2_X1    g28574(.A1(new_n31803_), .A2(new_n8685_), .ZN(new_n31838_));
  INV_X1     g28575(.I(new_n31838_), .ZN(new_n31839_));
  NOR2_X1    g28576(.A1(new_n30687_), .A2(new_n31450_), .ZN(new_n31840_));
  INV_X1     g28577(.I(new_n31840_), .ZN(new_n31841_));
  NOR2_X1    g28578(.A1(new_n31841_), .A2(new_n31839_), .ZN(new_n31842_));
  NAND3_X1   g28579(.A1(new_n31144_), .A2(new_n8684_), .A3(new_n30743_), .ZN(new_n31843_));
  NOR2_X1    g28580(.A1(new_n30610_), .A2(new_n8684_), .ZN(new_n31844_));
  OAI21_X1   g28581(.A1(new_n31447_), .A2(new_n31082_), .B(new_n31844_), .ZN(new_n31845_));
  INV_X1     g28582(.I(new_n31842_), .ZN(new_n31846_));
  AND3_X2    g28583(.A1(new_n31846_), .A2(new_n8685_), .A3(new_n31845_), .Z(new_n31847_));
  AOI21_X1   g28584(.A1(new_n31841_), .A2(pi0212), .B(po1038), .ZN(new_n31848_));
  INV_X1     g28585(.I(new_n31848_), .ZN(new_n31849_));
  OAI21_X1   g28586(.A1(new_n31843_), .A2(new_n31847_), .B(new_n31849_), .ZN(new_n31850_));
  NOR2_X1    g28587(.A1(new_n3098_), .A2(new_n13817_), .ZN(new_n31851_));
  AOI21_X1   g28588(.A1(new_n31841_), .A2(pi0211), .B(new_n8685_), .ZN(new_n31852_));
  NAND4_X1   g28589(.A1(new_n31850_), .A2(new_n31842_), .A3(new_n31851_), .A4(new_n31852_), .ZN(new_n31853_));
  NOR2_X1    g28590(.A1(new_n7240_), .A2(new_n30923_), .ZN(new_n31854_));
  NOR2_X1    g28591(.A1(new_n30922_), .A2(new_n31379_), .ZN(new_n31855_));
  AOI21_X1   g28592(.A1(new_n31854_), .A2(new_n31855_), .B(pi0213), .ZN(new_n31856_));
  NAND2_X1   g28593(.A1(new_n31853_), .A2(new_n31856_), .ZN(new_n31857_));
  NAND2_X1   g28594(.A1(new_n31856_), .A2(pi0209), .ZN(new_n31858_));
  XNOR2_X1   g28595(.A1(new_n31857_), .A2(new_n31858_), .ZN(new_n31859_));
  NOR2_X1    g28596(.A1(new_n31467_), .A2(new_n31551_), .ZN(new_n31860_));
  INV_X1     g28597(.I(new_n31860_), .ZN(new_n31861_));
  AOI21_X1   g28598(.A1(new_n31861_), .A2(new_n30838_), .B(new_n30743_), .ZN(new_n31862_));
  NOR2_X1    g28599(.A1(new_n31861_), .A2(new_n31839_), .ZN(new_n31863_));
  AOI21_X1   g28600(.A1(new_n31862_), .A2(new_n31863_), .B(new_n31844_), .ZN(new_n31864_));
  NOR2_X1    g28601(.A1(new_n31864_), .A2(new_n31530_), .ZN(new_n31865_));
  AOI21_X1   g28602(.A1(new_n31861_), .A2(pi0212), .B(po1038), .ZN(new_n31866_));
  NOR4_X1    g28603(.A1(new_n31861_), .A2(new_n8684_), .A3(new_n8685_), .A4(new_n31803_), .ZN(new_n31868_));
  OAI21_X1   g28604(.A1(new_n31865_), .A2(new_n31866_), .B(new_n31868_), .ZN(new_n31869_));
  OAI21_X1   g28605(.A1(new_n31859_), .A2(new_n31869_), .B(pi0230), .ZN(new_n31870_));
  INV_X1     g28606(.I(new_n31863_), .ZN(new_n31871_));
  NOR2_X1    g28607(.A1(new_n31866_), .A2(pi0209), .ZN(new_n31872_));
  NAND2_X1   g28608(.A1(new_n31861_), .A2(pi0211), .ZN(new_n31873_));
  NOR2_X1    g28609(.A1(new_n31871_), .A2(new_n31399_), .ZN(new_n31874_));
  OAI21_X1   g28610(.A1(new_n31403_), .A2(new_n28529_), .B(new_n8683_), .ZN(new_n31875_));
  NAND4_X1   g28611(.A1(new_n31874_), .A2(new_n31862_), .A3(new_n31873_), .A4(new_n31875_), .ZN(new_n31876_));
  OAI21_X1   g28612(.A1(new_n31876_), .A2(new_n31872_), .B(new_n31871_), .ZN(new_n31877_));
  NAND2_X1   g28613(.A1(new_n31843_), .A2(new_n31852_), .ZN(new_n31878_));
  NOR3_X1    g28614(.A1(new_n8546_), .A2(new_n3098_), .A3(new_n14006_), .ZN(new_n31879_));
  OAI21_X1   g28615(.A1(new_n31551_), .A2(new_n31879_), .B(pi0211), .ZN(new_n31880_));
  NAND2_X1   g28616(.A1(new_n31880_), .A2(new_n8685_), .ZN(new_n31881_));
  NOR3_X1    g28617(.A1(new_n31484_), .A2(pi0209), .A3(new_n14006_), .ZN(new_n31882_));
  NOR2_X1    g28618(.A1(new_n31477_), .A2(new_n8546_), .ZN(new_n31883_));
  NOR2_X1    g28619(.A1(new_n31494_), .A2(new_n8546_), .ZN(new_n31884_));
  XOR2_X1    g28620(.A1(new_n31884_), .A2(new_n31883_), .Z(new_n31885_));
  NAND4_X1   g28621(.A1(new_n31882_), .A2(new_n31848_), .A3(new_n31881_), .A4(new_n31885_), .ZN(new_n31886_));
  AOI21_X1   g28622(.A1(new_n31878_), .A2(new_n31842_), .B(new_n31886_), .ZN(new_n31887_));
  NAND2_X1   g28623(.A1(new_n31877_), .A2(new_n31887_), .ZN(new_n31888_));
  NAND2_X1   g28624(.A1(new_n31888_), .A2(new_n31846_), .ZN(new_n31889_));
  NAND3_X1   g28625(.A1(pi0208), .A2(pi0299), .A3(pi1157), .ZN(new_n31890_));
  NAND3_X1   g28626(.A1(new_n31840_), .A2(pi0214), .A3(pi1157), .ZN(new_n31891_));
  OAI21_X1   g28627(.A1(new_n31891_), .A2(new_n31890_), .B(new_n8684_), .ZN(new_n31892_));
  NAND4_X1   g28628(.A1(new_n31883_), .A2(new_n8545_), .A3(pi0230), .A4(pi0239), .ZN(new_n31893_));
  AOI21_X1   g28629(.A1(new_n31474_), .A2(pi0208), .B(new_n31893_), .ZN(new_n31894_));
  NAND3_X1   g28630(.A1(new_n31889_), .A2(new_n31892_), .A3(new_n31894_), .ZN(new_n31895_));
  XOR2_X1    g28631(.A1(new_n31870_), .A2(new_n31895_), .Z(po0396));
  NOR2_X1    g28632(.A1(new_n8549_), .A2(new_n3518_), .ZN(new_n31897_));
  NOR2_X1    g28633(.A1(new_n31897_), .A2(pi0200), .ZN(new_n31898_));
  INV_X1     g28634(.I(new_n31898_), .ZN(new_n31899_));
  NOR2_X1    g28635(.A1(new_n3350_), .A2(pi0199), .ZN(new_n31900_));
  INV_X1     g28636(.I(new_n31900_), .ZN(new_n31901_));
  AOI21_X1   g28637(.A1(new_n31901_), .A2(pi0200), .B(pi0299), .ZN(new_n31902_));
  NOR2_X1    g28638(.A1(new_n3518_), .A2(pi0199), .ZN(new_n31903_));
  NOR4_X1    g28639(.A1(new_n30812_), .A2(new_n31901_), .A3(pi0200), .A4(new_n31897_), .ZN(new_n31904_));
  NOR2_X1    g28640(.A1(new_n31904_), .A2(new_n30967_), .ZN(new_n31905_));
  AOI21_X1   g28641(.A1(new_n31905_), .A2(new_n8547_), .B(new_n31902_), .ZN(new_n31906_));
  NOR2_X1    g28642(.A1(new_n31906_), .A2(new_n31899_), .ZN(new_n31907_));
  INV_X1     g28643(.I(new_n31902_), .ZN(new_n31908_));
  NOR2_X1    g28644(.A1(pi0199), .A2(pi1145), .ZN(new_n31909_));
  AOI21_X1   g28645(.A1(new_n31908_), .A2(new_n31909_), .B(new_n8555_), .ZN(new_n31910_));
  INV_X1     g28646(.I(new_n31910_), .ZN(new_n31911_));
  NOR2_X1    g28647(.A1(new_n3098_), .A2(new_n3350_), .ZN(new_n31912_));
  NOR2_X1    g28648(.A1(new_n31912_), .A2(new_n8546_), .ZN(new_n31913_));
  INV_X1     g28649(.I(new_n31913_), .ZN(new_n31914_));
  OAI21_X1   g28650(.A1(new_n31904_), .A2(new_n31914_), .B(new_n31911_), .ZN(new_n31915_));
  NAND2_X1   g28651(.A1(new_n31911_), .A2(new_n31899_), .ZN(new_n31916_));
  OAI21_X1   g28652(.A1(new_n31915_), .A2(new_n31916_), .B(pi0207), .ZN(new_n31917_));
  NAND3_X1   g28653(.A1(new_n31917_), .A2(new_n31450_), .A3(new_n31908_), .ZN(new_n31918_));
  NAND2_X1   g28654(.A1(new_n31918_), .A2(new_n31898_), .ZN(new_n31919_));
  NOR2_X1    g28655(.A1(new_n31919_), .A2(pi0299), .ZN(new_n31920_));
  NOR2_X1    g28656(.A1(new_n31920_), .A2(new_n8685_), .ZN(new_n31921_));
  XOR2_X1    g28657(.A1(new_n31921_), .A2(new_n8740_), .Z(new_n31922_));
  NAND2_X1   g28658(.A1(new_n31922_), .A2(new_n31907_), .ZN(new_n31923_));
  NAND2_X1   g28659(.A1(new_n31915_), .A2(pi0207), .ZN(new_n31924_));
  OAI21_X1   g28660(.A1(new_n31450_), .A2(new_n31911_), .B(new_n31924_), .ZN(new_n31925_));
  NOR2_X1    g28661(.A1(new_n31925_), .A2(pi0299), .ZN(new_n31926_));
  NOR2_X1    g28662(.A1(new_n31926_), .A2(pi0211), .ZN(new_n31927_));
  INV_X1     g28663(.I(new_n31927_), .ZN(new_n31928_));
  AOI21_X1   g28664(.A1(new_n31911_), .A2(new_n9090_), .B(new_n31905_), .ZN(new_n31929_));
  NOR3_X1    g28665(.A1(new_n31920_), .A2(pi0214), .A3(new_n31929_), .ZN(new_n31930_));
  OAI21_X1   g28666(.A1(new_n31930_), .A2(new_n31928_), .B(pi0212), .ZN(new_n31931_));
  AOI21_X1   g28667(.A1(new_n31923_), .A2(new_n31931_), .B(new_n8683_), .ZN(new_n31932_));
  XOR2_X1    g28668(.A1(new_n31932_), .A2(new_n9213_), .Z(new_n31933_));
  NAND2_X1   g28669(.A1(new_n31933_), .A2(new_n31907_), .ZN(new_n31934_));
  INV_X1     g28670(.I(new_n31934_), .ZN(new_n31935_));
  NOR2_X1    g28671(.A1(new_n8684_), .A2(new_n8683_), .ZN(new_n31936_));
  INV_X1     g28672(.I(new_n31936_), .ZN(new_n31937_));
  AOI21_X1   g28673(.A1(new_n7240_), .A2(new_n31238_), .B(new_n31937_), .ZN(new_n31938_));
  INV_X1     g28674(.I(new_n31938_), .ZN(new_n31939_));
  INV_X1     g28675(.I(pi1147), .ZN(new_n31940_));
  INV_X1     g28676(.I(pi1149), .ZN(new_n31941_));
  NAND2_X1   g28677(.A1(new_n31940_), .A2(new_n31941_), .ZN(new_n31942_));
  AOI21_X1   g28678(.A1(new_n31929_), .A2(new_n30604_), .B(new_n8683_), .ZN(new_n31943_));
  NAND2_X1   g28679(.A1(new_n31943_), .A2(po1038), .ZN(new_n31944_));
  AOI21_X1   g28680(.A1(new_n31928_), .A2(new_n31944_), .B(new_n31238_), .ZN(new_n31945_));
  INV_X1     g28681(.I(new_n31945_), .ZN(new_n31946_));
  NOR2_X1    g28682(.A1(new_n30586_), .A2(new_n3098_), .ZN(new_n31947_));
  INV_X1     g28683(.I(new_n31947_), .ZN(new_n31948_));
  NAND3_X1   g28684(.A1(new_n31946_), .A2(new_n8683_), .A3(new_n31948_), .ZN(new_n31949_));
  AOI21_X1   g28685(.A1(new_n31949_), .A2(new_n31929_), .B(new_n31942_), .ZN(new_n31950_));
  NOR2_X1    g28686(.A1(new_n31756_), .A2(pi1147), .ZN(new_n31951_));
  OAI21_X1   g28687(.A1(new_n31950_), .A2(new_n31939_), .B(new_n31951_), .ZN(new_n31952_));
  INV_X1     g28688(.I(pi1148), .ZN(new_n31953_));
  NOR2_X1    g28689(.A1(po1038), .A2(new_n31940_), .ZN(new_n31954_));
  INV_X1     g28690(.I(new_n31758_), .ZN(new_n31955_));
  INV_X1     g28691(.I(new_n31920_), .ZN(new_n31956_));
  NOR2_X1    g28692(.A1(new_n31926_), .A2(new_n8684_), .ZN(new_n31957_));
  AOI21_X1   g28693(.A1(new_n31957_), .A2(pi0212), .B(pi0214), .ZN(new_n31958_));
  INV_X1     g28694(.I(new_n31926_), .ZN(new_n31959_));
  NAND2_X1   g28695(.A1(new_n31959_), .A2(new_n8686_), .ZN(new_n31960_));
  NAND2_X1   g28696(.A1(new_n31929_), .A2(pi0219), .ZN(new_n31961_));
  NOR4_X1    g28697(.A1(new_n31958_), .A2(new_n31956_), .A3(new_n31960_), .A4(new_n31961_), .ZN(new_n31962_));
  NOR2_X1    g28698(.A1(new_n31946_), .A2(new_n31962_), .ZN(new_n31963_));
  OAI21_X1   g28699(.A1(pi0214), .A2(new_n31929_), .B(new_n31957_), .ZN(new_n31965_));
  NAND2_X1   g28700(.A1(new_n31929_), .A2(pi0212), .ZN(new_n31966_));
  NAND2_X1   g28701(.A1(new_n31966_), .A2(new_n8685_), .ZN(new_n31967_));
  NAND2_X1   g28702(.A1(new_n31927_), .A2(new_n31967_), .ZN(new_n31968_));
  NAND3_X1   g28703(.A1(new_n31965_), .A2(new_n8683_), .A3(new_n31968_), .ZN(new_n31969_));
  NAND2_X1   g28704(.A1(new_n31963_), .A2(new_n31969_), .ZN(new_n31970_));
  NAND4_X1   g28705(.A1(new_n31970_), .A2(pi1147), .A3(new_n31955_), .A4(new_n31907_), .ZN(new_n31971_));
  XOR2_X1    g28706(.A1(new_n31971_), .A2(new_n31954_), .Z(new_n31972_));
  AOI21_X1   g28707(.A1(new_n8689_), .A2(new_n31723_), .B(new_n30918_), .ZN(new_n31973_));
  AOI21_X1   g28708(.A1(pi1147), .A2(new_n31973_), .B(new_n31945_), .ZN(new_n31974_));
  NOR2_X1    g28709(.A1(new_n31953_), .A2(new_n31941_), .ZN(new_n31975_));
  INV_X1     g28710(.I(new_n31975_), .ZN(new_n31976_));
  OAI21_X1   g28711(.A1(new_n31974_), .A2(new_n31969_), .B(new_n31976_), .ZN(new_n31977_));
  NOR2_X1    g28712(.A1(new_n9078_), .A2(new_n30979_), .ZN(new_n31978_));
  INV_X1     g28713(.I(new_n31907_), .ZN(new_n31979_));
  INV_X1     g28714(.I(new_n31978_), .ZN(new_n31980_));
  OAI21_X1   g28715(.A1(new_n31940_), .A2(new_n31980_), .B(new_n31979_), .ZN(new_n31981_));
  AOI21_X1   g28716(.A1(new_n31981_), .A2(po1038), .B(new_n31978_), .ZN(new_n31982_));
  NAND2_X1   g28717(.A1(new_n12654_), .A2(pi0213), .ZN(new_n31983_));
  AOI21_X1   g28718(.A1(new_n31919_), .A2(new_n31982_), .B(new_n31983_), .ZN(new_n31984_));
  AOI21_X1   g28719(.A1(new_n31977_), .A2(new_n31984_), .B(pi1149), .ZN(new_n31985_));
  OAI21_X1   g28720(.A1(new_n31972_), .A2(new_n31985_), .B(new_n31953_), .ZN(new_n31986_));
  AOI21_X1   g28721(.A1(new_n31935_), .A2(new_n31952_), .B(new_n31986_), .ZN(new_n31987_));
  NAND2_X1   g28722(.A1(new_n31935_), .A2(new_n31962_), .ZN(new_n31988_));
  NAND2_X1   g28723(.A1(new_n31988_), .A2(new_n31238_), .ZN(new_n31989_));
  AOI21_X1   g28724(.A1(pi0214), .A2(pi0219), .B(pi0212), .ZN(new_n31990_));
  NOR2_X1    g28725(.A1(pi0214), .A2(pi0219), .ZN(new_n31991_));
  NOR3_X1    g28726(.A1(new_n31990_), .A2(new_n8684_), .A3(new_n31991_), .ZN(new_n31992_));
  NOR2_X1    g28727(.A1(new_n30918_), .A2(new_n31992_), .ZN(new_n31993_));
  OAI21_X1   g28728(.A1(new_n31963_), .A2(new_n31942_), .B(new_n31993_), .ZN(new_n31994_));
  NOR2_X1    g28729(.A1(new_n31763_), .A2(pi0214), .ZN(new_n31995_));
  INV_X1     g28730(.I(new_n31995_), .ZN(new_n31996_));
  NOR2_X1    g28731(.A1(new_n31996_), .A2(pi1147), .ZN(new_n31997_));
  AOI21_X1   g28732(.A1(new_n31994_), .A2(new_n31997_), .B(new_n31979_), .ZN(new_n31998_));
  NAND2_X1   g28733(.A1(new_n31989_), .A2(new_n31998_), .ZN(new_n31999_));
  OAI21_X1   g28734(.A1(new_n31999_), .A2(new_n31987_), .B(new_n28364_), .ZN(new_n32000_));
  NAND2_X1   g28735(.A1(new_n31919_), .A2(new_n3098_), .ZN(new_n32001_));
  NOR2_X1    g28736(.A1(new_n8684_), .A2(pi1145), .ZN(new_n32002_));
  AOI21_X1   g28737(.A1(new_n8684_), .A2(new_n3350_), .B(new_n32002_), .ZN(new_n32003_));
  NAND2_X1   g28738(.A1(new_n32003_), .A2(pi0299), .ZN(new_n32004_));
  INV_X1     g28739(.I(new_n32004_), .ZN(new_n32005_));
  NOR2_X1    g28740(.A1(new_n32005_), .A2(new_n8685_), .ZN(new_n32006_));
  INV_X1     g28741(.I(new_n32006_), .ZN(new_n32007_));
  INV_X1     g28742(.I(new_n31912_), .ZN(new_n32008_));
  NOR2_X1    g28743(.A1(new_n32008_), .A2(new_n8684_), .ZN(new_n32009_));
  NOR2_X1    g28744(.A1(new_n31907_), .A2(pi0214), .ZN(new_n32010_));
  NOR2_X1    g28745(.A1(new_n32010_), .A2(pi0212), .ZN(new_n32011_));
  AOI21_X1   g28746(.A1(new_n32011_), .A2(pi0219), .B(new_n32009_), .ZN(new_n32012_));
  INV_X1     g28747(.I(new_n32012_), .ZN(new_n32013_));
  NAND2_X1   g28748(.A1(new_n32010_), .A2(new_n8739_), .ZN(new_n32014_));
  NAND4_X1   g28749(.A1(new_n32013_), .A2(new_n31907_), .A3(new_n32009_), .A4(new_n32014_), .ZN(new_n32015_));
  AOI21_X1   g28750(.A1(new_n32015_), .A2(new_n32007_), .B(new_n32001_), .ZN(new_n32016_));
  NOR3_X1    g28751(.A1(new_n31503_), .A2(pi0211), .A3(new_n30586_), .ZN(new_n32017_));
  AOI21_X1   g28752(.A1(new_n31907_), .A2(new_n30586_), .B(new_n8683_), .ZN(new_n32018_));
  INV_X1     g28753(.I(new_n32018_), .ZN(new_n32019_));
  AOI21_X1   g28754(.A1(new_n31349_), .A2(new_n3518_), .B(new_n8684_), .ZN(new_n32020_));
  NOR2_X1    g28755(.A1(new_n32003_), .A2(new_n8739_), .ZN(new_n32021_));
  NOR2_X1    g28756(.A1(new_n8684_), .A2(new_n3350_), .ZN(new_n32022_));
  XOR2_X1    g28757(.A1(new_n32003_), .A2(new_n30597_), .Z(new_n32023_));
  NAND2_X1   g28758(.A1(new_n32023_), .A2(new_n32022_), .ZN(new_n32024_));
  XOR2_X1    g28759(.A1(new_n32024_), .A2(new_n32021_), .Z(new_n32025_));
  INV_X1     g28760(.I(new_n32025_), .ZN(new_n32026_));
  AOI21_X1   g28761(.A1(new_n32026_), .A2(new_n31379_), .B(new_n32020_), .ZN(new_n32027_));
  NOR2_X1    g28762(.A1(new_n31980_), .A2(new_n7240_), .ZN(new_n32028_));
  NOR3_X1    g28763(.A1(new_n32027_), .A2(new_n31940_), .A3(new_n32028_), .ZN(new_n32029_));
  INV_X1     g28764(.I(new_n32029_), .ZN(new_n32030_));
  NOR4_X1    g28765(.A1(new_n32030_), .A2(new_n32001_), .A3(new_n32017_), .A4(new_n32019_), .ZN(new_n32031_));
  OAI21_X1   g28766(.A1(po1038), .A2(new_n32016_), .B(new_n32031_), .ZN(new_n32032_));
  INV_X1     g28767(.I(new_n32032_), .ZN(new_n32033_));
  OAI21_X1   g28768(.A1(new_n31979_), .A2(new_n32012_), .B(new_n31968_), .ZN(new_n32034_));
  NAND2_X1   g28769(.A1(new_n31957_), .A2(new_n31508_), .ZN(new_n32035_));
  OAI21_X1   g28770(.A1(new_n31925_), .A2(new_n32007_), .B(new_n31960_), .ZN(new_n32036_));
  NOR2_X1    g28771(.A1(new_n32009_), .A2(new_n10253_), .ZN(new_n32037_));
  NOR2_X1    g28772(.A1(new_n32037_), .A2(pi0212), .ZN(new_n32038_));
  AOI21_X1   g28773(.A1(new_n31925_), .A2(new_n32038_), .B(new_n8685_), .ZN(new_n32039_));
  NAND4_X1   g28774(.A1(new_n32034_), .A2(new_n32036_), .A3(new_n32035_), .A4(new_n32039_), .ZN(new_n32040_));
  NOR2_X1    g28775(.A1(new_n32027_), .A2(pi1147), .ZN(new_n32041_));
  AND3_X2    g28776(.A1(new_n31943_), .A2(new_n31238_), .A3(new_n31508_), .Z(new_n32042_));
  NAND3_X1   g28777(.A1(new_n31927_), .A2(new_n32041_), .A3(new_n32042_), .ZN(new_n32043_));
  AOI21_X1   g28778(.A1(new_n32040_), .A2(new_n7240_), .B(new_n32043_), .ZN(new_n32044_));
  NOR2_X1    g28779(.A1(new_n32044_), .A2(new_n32033_), .ZN(new_n32045_));
  NOR2_X1    g28780(.A1(new_n32045_), .A2(new_n28529_), .ZN(new_n32046_));
  AOI21_X1   g28781(.A1(new_n32000_), .A2(new_n32046_), .B(new_n30557_), .ZN(new_n32047_));
  NOR2_X1    g28782(.A1(po1038), .A2(new_n30595_), .ZN(new_n32048_));
  INV_X1     g28783(.I(new_n32048_), .ZN(new_n32049_));
  NOR2_X1    g28784(.A1(new_n32049_), .A2(new_n31948_), .ZN(new_n32050_));
  INV_X1     g28785(.I(new_n32050_), .ZN(new_n32051_));
  NOR2_X1    g28786(.A1(new_n31663_), .A2(po1038), .ZN(new_n32052_));
  NAND2_X1   g28787(.A1(new_n32052_), .A2(new_n31992_), .ZN(new_n32053_));
  AOI21_X1   g28788(.A1(new_n32053_), .A2(new_n32051_), .B(new_n30918_), .ZN(new_n32054_));
  INV_X1     g28789(.I(new_n32054_), .ZN(new_n32055_));
  INV_X1     g28790(.I(new_n31633_), .ZN(new_n32056_));
  NAND2_X1   g28791(.A1(new_n8775_), .A2(new_n8547_), .ZN(new_n32057_));
  NAND2_X1   g28792(.A1(new_n9090_), .A2(new_n8774_), .ZN(new_n32058_));
  AOI21_X1   g28793(.A1(new_n32057_), .A2(new_n32058_), .B(new_n30751_), .ZN(new_n32059_));
  AOI21_X1   g28794(.A1(new_n32059_), .A2(new_n32056_), .B(pi0299), .ZN(new_n32060_));
  OAI21_X1   g28795(.A1(new_n32056_), .A2(new_n32059_), .B(new_n32060_), .ZN(new_n32061_));
  INV_X1     g28796(.I(new_n32061_), .ZN(new_n32062_));
  NOR2_X1    g28797(.A1(new_n32062_), .A2(new_n31660_), .ZN(new_n32063_));
  NOR2_X1    g28798(.A1(new_n30718_), .A2(new_n3098_), .ZN(new_n32064_));
  NOR2_X1    g28799(.A1(new_n32063_), .A2(new_n32064_), .ZN(new_n32065_));
  INV_X1     g28800(.I(new_n32065_), .ZN(new_n32066_));
  AOI21_X1   g28801(.A1(new_n32066_), .A2(new_n8739_), .B(pi0219), .ZN(new_n32067_));
  INV_X1     g28802(.I(new_n32063_), .ZN(new_n32068_));
  NAND3_X1   g28803(.A1(new_n32068_), .A2(pi0212), .A3(new_n31523_), .ZN(new_n32069_));
  AOI21_X1   g28804(.A1(new_n32069_), .A2(new_n8685_), .B(new_n32061_), .ZN(new_n32070_));
  NOR2_X1    g28805(.A1(new_n32062_), .A2(pi0211), .ZN(new_n32071_));
  NOR2_X1    g28806(.A1(new_n32071_), .A2(new_n8740_), .ZN(new_n32072_));
  NOR2_X1    g28807(.A1(new_n32072_), .A2(new_n32068_), .ZN(new_n32073_));
  AOI21_X1   g28808(.A1(new_n32063_), .A2(new_n8685_), .B(pi0212), .ZN(new_n32074_));
  AOI22_X1   g28809(.A1(new_n32073_), .A2(new_n32074_), .B1(pi0214), .B2(new_n32061_), .ZN(new_n32075_));
  INV_X1     g28810(.I(new_n32075_), .ZN(new_n32076_));
  NAND2_X1   g28811(.A1(new_n32076_), .A2(new_n32070_), .ZN(new_n32077_));
  AND2_X2    g28812(.A1(new_n32077_), .A2(new_n32067_), .Z(new_n32078_));
  AOI21_X1   g28813(.A1(new_n32068_), .A2(pi0219), .B(po1038), .ZN(new_n32079_));
  INV_X1     g28814(.I(new_n32079_), .ZN(new_n32080_));
  NOR2_X1    g28815(.A1(new_n32078_), .A2(new_n32080_), .ZN(new_n32081_));
  NOR2_X1    g28816(.A1(new_n32081_), .A2(new_n31996_), .ZN(new_n32082_));
  NOR2_X1    g28817(.A1(new_n32082_), .A2(new_n31940_), .ZN(new_n32083_));
  NAND2_X1   g28818(.A1(pi1147), .A2(pi1149), .ZN(new_n32084_));
  XOR2_X1    g28819(.A1(new_n32083_), .A2(new_n32084_), .Z(new_n32085_));
  OAI21_X1   g28820(.A1(new_n32085_), .A2(new_n32055_), .B(pi1148), .ZN(new_n32086_));
  NAND2_X1   g28821(.A1(new_n12654_), .A2(new_n31600_), .ZN(new_n32087_));
  INV_X1     g28822(.I(new_n32087_), .ZN(new_n32088_));
  NOR2_X1    g28823(.A1(new_n12654_), .A2(pi0219), .ZN(new_n32089_));
  INV_X1     g28824(.I(new_n32089_), .ZN(new_n32090_));
  NOR2_X1    g28825(.A1(new_n32090_), .A2(new_n31723_), .ZN(new_n32091_));
  NOR2_X1    g28826(.A1(new_n32091_), .A2(new_n32088_), .ZN(new_n32092_));
  NOR2_X1    g28827(.A1(new_n31695_), .A2(pi0214), .ZN(new_n32093_));
  NOR2_X1    g28828(.A1(new_n32093_), .A2(pi0212), .ZN(new_n32094_));
  NOR2_X1    g28829(.A1(new_n31697_), .A2(new_n8685_), .ZN(new_n32095_));
  INV_X1     g28830(.I(new_n32095_), .ZN(new_n32096_));
  AOI21_X1   g28831(.A1(new_n32096_), .A2(new_n32094_), .B(pi0219), .ZN(new_n32097_));
  NOR2_X1    g28832(.A1(new_n31678_), .A2(new_n8685_), .ZN(new_n32098_));
  XOR2_X1    g28833(.A1(new_n32098_), .A2(new_n30718_), .Z(new_n32099_));
  NOR2_X1    g28834(.A1(new_n31692_), .A2(new_n32099_), .ZN(new_n32100_));
  NOR3_X1    g28835(.A1(new_n32097_), .A2(pi0212), .A3(new_n32100_), .ZN(new_n32101_));
  NOR2_X1    g28836(.A1(new_n32101_), .A2(new_n31697_), .ZN(new_n32102_));
  INV_X1     g28837(.I(new_n32102_), .ZN(new_n32103_));
  NOR2_X1    g28838(.A1(new_n32100_), .A2(new_n30597_), .ZN(new_n32104_));
  NOR2_X1    g28839(.A1(new_n32103_), .A2(new_n32104_), .ZN(new_n32105_));
  NOR3_X1    g28840(.A1(new_n31697_), .A2(new_n8739_), .A3(new_n8683_), .ZN(new_n32106_));
  NOR2_X1    g28841(.A1(new_n32106_), .A2(po1038), .ZN(new_n32107_));
  INV_X1     g28842(.I(new_n32107_), .ZN(new_n32108_));
  NOR2_X1    g28843(.A1(new_n32105_), .A2(new_n32108_), .ZN(new_n32109_));
  NAND2_X1   g28844(.A1(new_n31940_), .A2(new_n31941_), .ZN(new_n32110_));
  NOR2_X1    g28845(.A1(new_n31450_), .A2(new_n9209_), .ZN(new_n32111_));
  NOR2_X1    g28846(.A1(new_n32111_), .A2(pi0299), .ZN(new_n32112_));
  NAND2_X1   g28847(.A1(new_n32112_), .A2(new_n31643_), .ZN(new_n32113_));
  NOR2_X1    g28848(.A1(new_n31652_), .A2(new_n8555_), .ZN(new_n32114_));
  NAND2_X1   g28849(.A1(new_n32113_), .A2(pi0214), .ZN(new_n32115_));
  XOR2_X1    g28850(.A1(new_n32115_), .A2(new_n30718_), .Z(new_n32116_));
  NAND2_X1   g28851(.A1(new_n32116_), .A2(new_n32114_), .ZN(new_n32117_));
  NAND2_X1   g28852(.A1(new_n32117_), .A2(pi0212), .ZN(new_n32118_));
  NOR2_X1    g28853(.A1(new_n32114_), .A2(pi0214), .ZN(new_n32119_));
  NOR2_X1    g28854(.A1(new_n32119_), .A2(pi0212), .ZN(new_n32120_));
  NAND2_X1   g28855(.A1(new_n32120_), .A2(pi0219), .ZN(new_n32121_));
  AOI21_X1   g28856(.A1(new_n32121_), .A2(new_n8685_), .B(new_n32113_), .ZN(new_n32122_));
  INV_X1     g28857(.I(new_n32114_), .ZN(new_n32123_));
  NOR2_X1    g28858(.A1(new_n32123_), .A2(po1038), .ZN(new_n32124_));
  NOR2_X1    g28859(.A1(new_n31810_), .A2(new_n32124_), .ZN(new_n32125_));
  NAND2_X1   g28860(.A1(new_n32122_), .A2(new_n32125_), .ZN(new_n32126_));
  AOI21_X1   g28861(.A1(new_n32118_), .A2(new_n32126_), .B(new_n32113_), .ZN(new_n32127_));
  NOR2_X1    g28862(.A1(new_n32127_), .A2(new_n31756_), .ZN(new_n32128_));
  NOR2_X1    g28863(.A1(new_n32128_), .A2(new_n31941_), .ZN(new_n32129_));
  XNOR2_X1   g28864(.A1(new_n32129_), .A2(new_n32084_), .ZN(new_n32130_));
  NAND2_X1   g28865(.A1(new_n30666_), .A2(new_n31640_), .ZN(new_n32131_));
  AOI21_X1   g28866(.A1(new_n32131_), .A2(pi0208), .B(pi0199), .ZN(new_n32132_));
  NOR2_X1    g28867(.A1(new_n31663_), .A2(new_n32132_), .ZN(new_n32133_));
  NOR2_X1    g28868(.A1(new_n32133_), .A2(pi0299), .ZN(new_n32134_));
  INV_X1     g28869(.I(new_n32052_), .ZN(new_n32135_));
  NOR2_X1    g28870(.A1(new_n31832_), .A2(pi0212), .ZN(new_n32136_));
  NOR3_X1    g28871(.A1(new_n31831_), .A2(new_n8684_), .A3(new_n3098_), .ZN(new_n32137_));
  AOI21_X1   g28872(.A1(pi0214), .A2(new_n10253_), .B(new_n31664_), .ZN(new_n32138_));
  NOR2_X1    g28873(.A1(new_n32138_), .A2(pi0212), .ZN(new_n32139_));
  NOR3_X1    g28874(.A1(new_n32139_), .A2(pi0219), .A3(new_n32137_), .ZN(new_n32140_));
  AOI21_X1   g28875(.A1(pi0219), .A2(new_n31800_), .B(new_n32049_), .ZN(new_n32141_));
  INV_X1     g28876(.I(new_n32141_), .ZN(new_n32142_));
  AOI21_X1   g28877(.A1(new_n32135_), .A2(new_n32142_), .B(new_n32140_), .ZN(new_n32143_));
  INV_X1     g28878(.I(new_n32143_), .ZN(new_n32144_));
  NOR2_X1    g28879(.A1(new_n32144_), .A2(new_n32134_), .ZN(new_n32145_));
  INV_X1     g28880(.I(new_n32145_), .ZN(new_n32146_));
  INV_X1     g28881(.I(new_n32134_), .ZN(new_n32147_));
  NOR2_X1    g28882(.A1(new_n32138_), .A2(new_n31664_), .ZN(new_n32148_));
  AOI21_X1   g28883(.A1(new_n32148_), .A2(new_n32147_), .B(pi0219), .ZN(new_n32149_));
  AOI21_X1   g28884(.A1(new_n8684_), .A2(new_n32149_), .B(new_n32146_), .ZN(new_n32150_));
  NOR2_X1    g28885(.A1(new_n32150_), .A2(new_n31758_), .ZN(new_n32151_));
  NOR2_X1    g28886(.A1(new_n30738_), .A2(new_n31211_), .ZN(new_n32152_));
  INV_X1     g28887(.I(new_n32152_), .ZN(new_n32153_));
  NOR2_X1    g28888(.A1(new_n32153_), .A2(new_n7240_), .ZN(new_n32154_));
  INV_X1     g28889(.I(new_n32154_), .ZN(new_n32155_));
  AOI21_X1   g28890(.A1(new_n32051_), .A2(new_n31939_), .B(new_n32155_), .ZN(new_n32156_));
  AND2_X2    g28891(.A1(new_n32156_), .A2(pi1148), .Z(new_n32157_));
  NAND4_X1   g28892(.A1(new_n32151_), .A2(new_n32110_), .A3(new_n32130_), .A4(new_n32157_), .ZN(new_n32158_));
  XOR2_X1    g28893(.A1(new_n32086_), .A2(new_n32158_), .Z(new_n32159_));
  NOR2_X1    g28894(.A1(new_n32159_), .A2(new_n28364_), .ZN(new_n32160_));
  XOR2_X1    g28895(.A1(new_n32160_), .A2(new_n31079_), .Z(new_n32161_));
  NAND2_X1   g28896(.A1(new_n32048_), .A2(pi0219), .ZN(new_n32162_));
  AOI21_X1   g28897(.A1(new_n32162_), .A2(new_n31511_), .B(new_n8684_), .ZN(new_n32163_));
  INV_X1     g28898(.I(new_n32163_), .ZN(new_n32164_));
  AOI21_X1   g28899(.A1(pi0219), .A2(new_n31678_), .B(po1038), .ZN(new_n32165_));
  OAI21_X1   g28900(.A1(new_n8546_), .A2(pi0299), .B(pi0207), .ZN(new_n32166_));
  NOR2_X1    g28901(.A1(new_n32166_), .A2(new_n8555_), .ZN(new_n32167_));
  AOI21_X1   g28902(.A1(new_n32167_), .A2(new_n32008_), .B(new_n8684_), .ZN(new_n32168_));
  AOI21_X1   g28903(.A1(new_n31692_), .A2(new_n8684_), .B(new_n32168_), .ZN(new_n32169_));
  NAND2_X1   g28904(.A1(new_n32169_), .A2(pi0214), .ZN(new_n32170_));
  NAND2_X1   g28905(.A1(new_n32170_), .A2(new_n32094_), .ZN(new_n32171_));
  AOI21_X1   g28906(.A1(new_n32006_), .A2(new_n32167_), .B(new_n30916_), .ZN(new_n32172_));
  NOR2_X1    g28907(.A1(new_n32169_), .A2(new_n32172_), .ZN(new_n32173_));
  NOR3_X1    g28908(.A1(new_n32030_), .A2(new_n8685_), .A3(new_n32173_), .ZN(new_n32174_));
  AOI21_X1   g28909(.A1(new_n32174_), .A2(new_n32171_), .B(new_n32165_), .ZN(new_n32175_));
  OAI21_X1   g28910(.A1(new_n32175_), .A2(new_n32164_), .B(new_n31953_), .ZN(new_n32176_));
  INV_X1     g28911(.I(new_n32041_), .ZN(new_n32177_));
  NOR3_X1    g28912(.A1(new_n32025_), .A2(new_n3098_), .A3(new_n31349_), .ZN(new_n32178_));
  AOI21_X1   g28913(.A1(pi0219), .A2(new_n32163_), .B(new_n32178_), .ZN(new_n32179_));
  INV_X1     g28914(.I(new_n32179_), .ZN(new_n32180_));
  NOR3_X1    g28915(.A1(new_n32177_), .A2(new_n32087_), .A3(new_n32180_), .ZN(new_n32181_));
  AOI21_X1   g28916(.A1(new_n32176_), .A2(new_n32181_), .B(new_n31941_), .ZN(new_n32182_));
  AOI21_X1   g28917(.A1(new_n31663_), .A2(new_n32004_), .B(new_n30597_), .ZN(new_n32183_));
  AOI21_X1   g28918(.A1(new_n31664_), .A2(new_n30586_), .B(pi0219), .ZN(new_n32184_));
  NOR4_X1    g28919(.A1(new_n31664_), .A2(new_n10253_), .A3(new_n30876_), .A4(new_n32009_), .ZN(new_n32185_));
  OAI21_X1   g28920(.A1(new_n32183_), .A2(new_n32184_), .B(new_n32185_), .ZN(new_n32186_));
  OAI21_X1   g28921(.A1(new_n32030_), .A2(new_n32186_), .B(new_n32135_), .ZN(new_n32187_));
  AOI21_X1   g28922(.A1(new_n32187_), .A2(new_n32163_), .B(pi1148), .ZN(new_n32188_));
  NOR2_X1    g28923(.A1(new_n32177_), .A2(new_n32180_), .ZN(new_n32189_));
  NOR2_X1    g28924(.A1(new_n32068_), .A2(po1038), .ZN(new_n32190_));
  NAND2_X1   g28925(.A1(new_n32189_), .A2(new_n32190_), .ZN(new_n32191_));
  INV_X1     g28926(.I(new_n32133_), .ZN(new_n32192_));
  NAND3_X1   g28927(.A1(new_n31126_), .A2(new_n30588_), .A3(pi1145), .ZN(new_n32193_));
  OAI21_X1   g28928(.A1(new_n32192_), .A2(new_n30892_), .B(new_n32193_), .ZN(new_n32194_));
  OAI21_X1   g28929(.A1(new_n32030_), .A2(new_n7240_), .B(new_n32194_), .ZN(new_n32195_));
  INV_X1     g28930(.I(new_n32183_), .ZN(new_n32196_));
  NOR2_X1    g28931(.A1(new_n32134_), .A2(pi0219), .ZN(new_n32197_));
  NOR2_X1    g28932(.A1(new_n31523_), .A2(pi1146), .ZN(new_n32198_));
  NOR4_X1    g28933(.A1(new_n32197_), .A2(new_n30876_), .A3(new_n32196_), .A4(new_n32198_), .ZN(new_n32199_));
  AOI21_X1   g28934(.A1(new_n32195_), .A2(new_n32199_), .B(pi1148), .ZN(new_n32200_));
  OAI21_X1   g28935(.A1(new_n32188_), .A2(new_n32191_), .B(new_n32200_), .ZN(new_n32201_));
  INV_X1     g28936(.I(new_n32113_), .ZN(new_n32202_));
  NOR2_X1    g28937(.A1(new_n32202_), .A2(new_n8739_), .ZN(new_n32203_));
  INV_X1     g28938(.I(new_n32022_), .ZN(new_n32204_));
  NAND2_X1   g28939(.A1(new_n32204_), .A2(new_n8685_), .ZN(new_n32205_));
  OAI21_X1   g28940(.A1(new_n32003_), .A2(new_n8685_), .B(new_n32205_), .ZN(new_n32206_));
  AOI21_X1   g28941(.A1(new_n32203_), .A2(pi0219), .B(new_n32206_), .ZN(new_n32207_));
  NAND2_X1   g28942(.A1(new_n32120_), .A2(new_n32114_), .ZN(new_n32208_));
  NOR2_X1    g28943(.A1(new_n32207_), .A2(new_n32208_), .ZN(new_n32209_));
  OAI21_X1   g28944(.A1(new_n32209_), .A2(new_n32009_), .B(new_n32114_), .ZN(new_n32210_));
  NAND3_X1   g28945(.A1(new_n32030_), .A2(new_n31953_), .A3(new_n32180_), .ZN(new_n32211_));
  NOR2_X1    g28946(.A1(new_n8739_), .A2(new_n3098_), .ZN(new_n32212_));
  INV_X1     g28947(.I(new_n32212_), .ZN(new_n32213_));
  NOR2_X1    g28948(.A1(new_n32213_), .A2(new_n30838_), .ZN(new_n32214_));
  INV_X1     g28949(.I(new_n32214_), .ZN(new_n32215_));
  AOI21_X1   g28950(.A1(new_n32153_), .A2(new_n3098_), .B(new_n8739_), .ZN(new_n32216_));
  NOR2_X1    g28951(.A1(new_n7240_), .A2(pi0219), .ZN(new_n32217_));
  INV_X1     g28952(.I(new_n32217_), .ZN(new_n32218_));
  AOI21_X1   g28953(.A1(new_n32215_), .A2(new_n32216_), .B(new_n32218_), .ZN(new_n32219_));
  INV_X1     g28954(.I(new_n31712_), .ZN(new_n32220_));
  AOI21_X1   g28955(.A1(new_n32153_), .A2(new_n32220_), .B(pi0212), .ZN(new_n32221_));
  INV_X1     g28956(.I(new_n32221_), .ZN(new_n32222_));
  NOR2_X1    g28957(.A1(new_n32152_), .A2(new_n8684_), .ZN(new_n32223_));
  NOR3_X1    g28958(.A1(new_n32219_), .A2(new_n32222_), .A3(new_n32223_), .ZN(new_n32224_));
  NAND3_X1   g28959(.A1(new_n32211_), .A2(new_n32041_), .A3(new_n32224_), .ZN(new_n32225_));
  NOR2_X1    g28960(.A1(new_n30604_), .A2(pi0219), .ZN(new_n32226_));
  NOR2_X1    g28961(.A1(new_n32113_), .A2(new_n32226_), .ZN(new_n32227_));
  NOR2_X1    g28962(.A1(new_n32227_), .A2(po1038), .ZN(new_n32228_));
  INV_X1     g28963(.I(new_n32228_), .ZN(new_n32229_));
  NOR2_X1    g28964(.A1(new_n32229_), .A2(new_n9209_), .ZN(new_n32230_));
  INV_X1     g28965(.I(new_n32230_), .ZN(new_n32231_));
  NAND4_X1   g28966(.A1(new_n32189_), .A2(pi1149), .A3(new_n32164_), .A4(new_n32231_), .ZN(new_n32232_));
  AOI21_X1   g28967(.A1(new_n32225_), .A2(new_n32210_), .B(new_n32232_), .ZN(new_n32233_));
  NAND2_X1   g28968(.A1(new_n32201_), .A2(new_n32233_), .ZN(new_n32234_));
  XNOR2_X1   g28969(.A1(new_n32234_), .A2(new_n32182_), .ZN(new_n32235_));
  NAND4_X1   g28970(.A1(new_n32161_), .A2(pi0230), .A3(pi0240), .A4(new_n32235_), .ZN(new_n32236_));
  XNOR2_X1   g28971(.A1(new_n32236_), .A2(new_n32047_), .ZN(po0397));
  NAND2_X1   g28972(.A1(new_n32082_), .A2(new_n31670_), .ZN(new_n32238_));
  NOR2_X1    g28973(.A1(new_n31756_), .A2(new_n31670_), .ZN(new_n32239_));
  INV_X1     g28974(.I(new_n32239_), .ZN(new_n32240_));
  NOR2_X1    g28975(.A1(new_n32127_), .A2(new_n32240_), .ZN(new_n32241_));
  INV_X1     g28976(.I(pi1150), .ZN(new_n32242_));
  INV_X1     g28977(.I(new_n32092_), .ZN(new_n32243_));
  NOR2_X1    g28978(.A1(pi1149), .A2(pi1150), .ZN(new_n32244_));
  INV_X1     g28979(.I(new_n32244_), .ZN(new_n32245_));
  NOR2_X1    g28980(.A1(new_n32245_), .A2(pi1151), .ZN(new_n32246_));
  OAI21_X1   g28981(.A1(new_n32243_), .A2(new_n32246_), .B(new_n32242_), .ZN(new_n32247_));
  NOR2_X1    g28982(.A1(new_n32241_), .A2(new_n32247_), .ZN(new_n32248_));
  NOR2_X1    g28983(.A1(new_n31938_), .A2(new_n31670_), .ZN(new_n32249_));
  INV_X1     g28984(.I(new_n32249_), .ZN(new_n32250_));
  AOI21_X1   g28985(.A1(new_n32250_), .A2(new_n32051_), .B(new_n32155_), .ZN(new_n32251_));
  OR2_X2     g28986(.A1(new_n32251_), .A2(pi1150), .Z(new_n32252_));
  NOR2_X1    g28987(.A1(new_n32055_), .A2(new_n31670_), .ZN(new_n32253_));
  AOI21_X1   g28988(.A1(new_n32253_), .A2(new_n32252_), .B(pi1149), .ZN(new_n32254_));
  OAI21_X1   g28989(.A1(new_n32238_), .A2(new_n32248_), .B(new_n32254_), .ZN(new_n32255_));
  NOR2_X1    g28990(.A1(new_n31973_), .A2(new_n31670_), .ZN(new_n32256_));
  INV_X1     g28991(.I(new_n32256_), .ZN(new_n32257_));
  NOR2_X1    g28992(.A1(new_n32109_), .A2(new_n32257_), .ZN(new_n32258_));
  INV_X1     g28993(.I(new_n31759_), .ZN(new_n32259_));
  NOR2_X1    g28994(.A1(new_n32150_), .A2(new_n32259_), .ZN(new_n32260_));
  NOR3_X1    g28995(.A1(new_n32258_), .A2(new_n32260_), .A3(pi1150), .ZN(new_n32261_));
  NAND2_X1   g28996(.A1(new_n32255_), .A2(new_n32261_), .ZN(new_n32262_));
  NAND2_X1   g28997(.A1(new_n32262_), .A2(pi0213), .ZN(new_n32263_));
  XOR2_X1    g28998(.A1(new_n32263_), .A2(new_n31080_), .Z(new_n32264_));
  OAI21_X1   g28999(.A1(new_n31728_), .A2(new_n31002_), .B(new_n32229_), .ZN(new_n32265_));
  OAI21_X1   g29000(.A1(new_n30694_), .A2(new_n9214_), .B(new_n31643_), .ZN(new_n32266_));
  NAND3_X1   g29001(.A1(new_n32266_), .A2(new_n8684_), .A3(new_n30829_), .ZN(new_n32267_));
  INV_X1     g29002(.I(new_n32267_), .ZN(new_n32268_));
  AOI21_X1   g29003(.A1(new_n32268_), .A2(new_n32120_), .B(pi0211), .ZN(new_n32269_));
  OAI21_X1   g29004(.A1(new_n32269_), .A2(new_n32123_), .B(new_n8683_), .ZN(new_n32270_));
  NAND2_X1   g29005(.A1(new_n32113_), .A2(new_n8684_), .ZN(new_n32271_));
  AOI21_X1   g29006(.A1(new_n32271_), .A2(new_n32119_), .B(pi0212), .ZN(new_n32272_));
  NOR2_X1    g29007(.A1(new_n32202_), .A2(new_n8684_), .ZN(new_n32273_));
  NOR2_X1    g29008(.A1(new_n32273_), .A2(new_n32114_), .ZN(new_n32274_));
  INV_X1     g29009(.I(new_n32274_), .ZN(new_n32275_));
  NOR3_X1    g29010(.A1(new_n32275_), .A2(new_n8685_), .A3(new_n32272_), .ZN(new_n32276_));
  NOR2_X1    g29011(.A1(new_n32268_), .A2(new_n32273_), .ZN(new_n32277_));
  INV_X1     g29012(.I(new_n32277_), .ZN(new_n32278_));
  NOR2_X1    g29013(.A1(new_n32278_), .A2(new_n32242_), .ZN(new_n32279_));
  AND4_X2    g29014(.A1(new_n32265_), .A2(new_n32276_), .A3(new_n32279_), .A4(new_n32270_), .Z(new_n32280_));
  AOI21_X1   g29015(.A1(new_n32061_), .A2(new_n30829_), .B(pi0211), .ZN(new_n32281_));
  INV_X1     g29016(.I(new_n32281_), .ZN(new_n32282_));
  OAI21_X1   g29017(.A1(new_n32063_), .A2(new_n32071_), .B(new_n31765_), .ZN(new_n32283_));
  NAND3_X1   g29018(.A1(new_n32063_), .A2(po1038), .A3(new_n31766_), .ZN(new_n32284_));
  AOI21_X1   g29019(.A1(new_n32283_), .A2(new_n32284_), .B(new_n32282_), .ZN(new_n32285_));
  OAI21_X1   g29020(.A1(new_n32280_), .A2(new_n31764_), .B(new_n32285_), .ZN(new_n32286_));
  AOI21_X1   g29021(.A1(new_n32107_), .A2(new_n31727_), .B(pi0219), .ZN(new_n32287_));
  NOR2_X1    g29022(.A1(new_n31691_), .A2(new_n8684_), .ZN(new_n32288_));
  NOR2_X1    g29023(.A1(new_n31695_), .A2(new_n31180_), .ZN(new_n32289_));
  XOR2_X1    g29024(.A1(new_n32288_), .A2(new_n32289_), .Z(new_n32290_));
  NAND2_X1   g29025(.A1(new_n32290_), .A2(new_n32094_), .ZN(new_n32291_));
  OAI21_X1   g29026(.A1(new_n32291_), .A2(new_n32104_), .B(new_n8739_), .ZN(new_n32292_));
  NAND2_X1   g29027(.A1(new_n32292_), .A2(new_n32100_), .ZN(new_n32293_));
  OAI21_X1   g29028(.A1(new_n32293_), .A2(new_n32287_), .B(new_n31002_), .ZN(new_n32294_));
  NAND2_X1   g29029(.A1(new_n31791_), .A2(pi1152), .ZN(new_n32295_));
  AOI21_X1   g29030(.A1(new_n32192_), .A2(pi0219), .B(po1038), .ZN(new_n32296_));
  INV_X1     g29031(.I(new_n32296_), .ZN(new_n32297_));
  NAND2_X1   g29032(.A1(new_n32297_), .A2(new_n32295_), .ZN(new_n32298_));
  NOR3_X1    g29033(.A1(new_n32133_), .A2(new_n8683_), .A3(new_n31947_), .ZN(new_n32299_));
  NOR4_X1    g29034(.A1(new_n31759_), .A2(new_n30654_), .A3(new_n31739_), .A4(new_n31757_), .ZN(new_n32300_));
  NAND2_X1   g29035(.A1(new_n32298_), .A2(new_n32300_), .ZN(new_n32301_));
  NAND2_X1   g29036(.A1(new_n32301_), .A2(new_n32108_), .ZN(new_n32302_));
  NOR2_X1    g29037(.A1(new_n32100_), .A2(new_n32093_), .ZN(new_n32303_));
  INV_X1     g29038(.I(new_n32303_), .ZN(new_n32304_));
  NOR4_X1    g29039(.A1(new_n31702_), .A2(new_n8683_), .A3(new_n32215_), .A4(new_n32304_), .ZN(new_n32305_));
  NAND2_X1   g29040(.A1(new_n32305_), .A2(new_n32302_), .ZN(new_n32306_));
  AOI21_X1   g29041(.A1(new_n30718_), .A2(new_n31793_), .B(new_n8739_), .ZN(new_n32307_));
  NOR2_X1    g29042(.A1(new_n32142_), .A2(new_n32307_), .ZN(new_n32308_));
  NOR2_X1    g29043(.A1(new_n32224_), .A2(new_n32308_), .ZN(new_n32309_));
  NAND2_X1   g29044(.A1(new_n32153_), .A2(new_n8683_), .ZN(new_n32310_));
  NAND2_X1   g29045(.A1(new_n32310_), .A2(new_n13614_), .ZN(new_n32311_));
  OAI21_X1   g29046(.A1(new_n32309_), .A2(new_n32311_), .B(new_n32214_), .ZN(new_n32312_));
  OAI21_X1   g29047(.A1(new_n32052_), .A2(pi1151), .B(new_n31002_), .ZN(new_n32313_));
  NOR2_X1    g29048(.A1(new_n31723_), .A2(new_n30620_), .ZN(new_n32314_));
  INV_X1     g29049(.I(new_n32314_), .ZN(new_n32315_));
  AOI21_X1   g29050(.A1(new_n31670_), .A2(pi1152), .B(pi1153), .ZN(new_n32316_));
  NOR2_X1    g29051(.A1(new_n32315_), .A2(new_n32316_), .ZN(new_n32317_));
  AOI21_X1   g29052(.A1(new_n31727_), .A2(new_n32317_), .B(new_n32245_), .ZN(new_n32318_));
  OAI21_X1   g29053(.A1(new_n32312_), .A2(new_n32313_), .B(new_n32318_), .ZN(new_n32319_));
  NOR3_X1    g29054(.A1(new_n32310_), .A2(pi0211), .A3(new_n32214_), .ZN(new_n32320_));
  INV_X1     g29055(.I(new_n32320_), .ZN(new_n32321_));
  NOR2_X1    g29056(.A1(new_n32321_), .A2(new_n32051_), .ZN(new_n32322_));
  OAI21_X1   g29057(.A1(new_n32322_), .A2(new_n32152_), .B(po1038), .ZN(new_n32323_));
  INV_X1     g29058(.I(new_n32323_), .ZN(new_n32324_));
  INV_X1     g29059(.I(new_n31760_), .ZN(new_n32325_));
  NOR2_X1    g29060(.A1(new_n31664_), .A2(new_n8683_), .ZN(new_n32326_));
  NOR2_X1    g29061(.A1(new_n32326_), .A2(po1038), .ZN(new_n32327_));
  INV_X1     g29062(.I(new_n32327_), .ZN(new_n32328_));
  NAND2_X1   g29063(.A1(new_n32328_), .A2(new_n32295_), .ZN(new_n32329_));
  NOR2_X1    g29064(.A1(pi0211), .A2(pi1153), .ZN(new_n32330_));
  NOR3_X1    g29065(.A1(new_n31664_), .A2(new_n3098_), .A3(new_n31090_), .ZN(new_n32331_));
  NOR3_X1    g29066(.A1(new_n31663_), .A2(new_n3098_), .A3(new_n31091_), .ZN(new_n32332_));
  OAI21_X1   g29067(.A1(new_n32331_), .A2(new_n32332_), .B(new_n32330_), .ZN(new_n32333_));
  NAND2_X1   g29068(.A1(new_n31663_), .A2(new_n31800_), .ZN(new_n32334_));
  NAND2_X1   g29069(.A1(new_n32334_), .A2(new_n8740_), .ZN(new_n32335_));
  NAND4_X1   g29070(.A1(new_n32329_), .A2(new_n32184_), .A3(new_n32333_), .A4(new_n32335_), .ZN(new_n32336_));
  NAND3_X1   g29071(.A1(new_n32336_), .A2(new_n32325_), .A3(new_n32312_), .ZN(new_n32337_));
  NAND3_X1   g29072(.A1(new_n32337_), .A2(new_n32319_), .A3(new_n32324_), .ZN(new_n32338_));
  NAND3_X1   g29073(.A1(new_n32338_), .A2(new_n32306_), .A3(new_n32242_), .ZN(new_n32339_));
  AOI21_X1   g29074(.A1(new_n31607_), .A2(pi0219), .B(po1038), .ZN(new_n32340_));
  NOR2_X1    g29075(.A1(new_n31601_), .A2(pi0212), .ZN(new_n32341_));
  NOR3_X1    g29076(.A1(new_n31802_), .A2(new_n8684_), .A3(new_n32341_), .ZN(new_n32342_));
  INV_X1     g29077(.I(new_n32342_), .ZN(new_n32343_));
  NAND2_X1   g29078(.A1(new_n31802_), .A2(new_n32341_), .ZN(new_n32344_));
  NOR2_X1    g29079(.A1(new_n32344_), .A2(new_n10253_), .ZN(new_n32345_));
  NOR2_X1    g29080(.A1(new_n32345_), .A2(pi0219), .ZN(new_n32346_));
  NAND2_X1   g29081(.A1(new_n32346_), .A2(new_n32343_), .ZN(new_n32347_));
  NAND2_X1   g29082(.A1(new_n32347_), .A2(new_n32340_), .ZN(new_n32348_));
  INV_X1     g29083(.I(new_n32348_), .ZN(new_n32349_));
  NAND2_X1   g29084(.A1(new_n31741_), .A2(pi0299), .ZN(new_n32350_));
  AOI21_X1   g29085(.A1(new_n32295_), .A2(new_n32350_), .B(new_n31739_), .ZN(new_n32351_));
  INV_X1     g29086(.I(new_n32340_), .ZN(new_n32352_));
  OR2_X2     g29087(.A1(new_n31809_), .A2(new_n32352_), .Z(new_n32353_));
  NAND2_X1   g29088(.A1(new_n32353_), .A2(new_n32325_), .ZN(new_n32354_));
  OAI21_X1   g29089(.A1(new_n32354_), .A2(new_n32351_), .B(new_n32349_), .ZN(new_n32355_));
  AOI21_X1   g29090(.A1(pi1150), .A2(new_n32317_), .B(new_n31727_), .ZN(new_n32356_));
  NOR2_X1    g29091(.A1(new_n32353_), .A2(new_n32356_), .ZN(new_n32357_));
  AOI21_X1   g29092(.A1(new_n32192_), .A2(new_n32315_), .B(po1038), .ZN(new_n32358_));
  NAND2_X1   g29093(.A1(new_n32330_), .A2(pi0299), .ZN(new_n32359_));
  NAND4_X1   g29094(.A1(new_n32358_), .A2(new_n31941_), .A3(new_n31764_), .A4(new_n32359_), .ZN(new_n32360_));
  AOI21_X1   g29095(.A1(new_n32355_), .A2(new_n32357_), .B(new_n32360_), .ZN(new_n32361_));
  NAND3_X1   g29096(.A1(new_n32361_), .A2(new_n32294_), .A3(new_n32339_), .ZN(new_n32362_));
  AOI21_X1   g29097(.A1(new_n31791_), .A2(new_n7240_), .B(pi0219), .ZN(new_n32363_));
  NAND2_X1   g29098(.A1(new_n32359_), .A2(new_n8685_), .ZN(new_n32364_));
  NOR2_X1    g29099(.A1(new_n32062_), .A2(new_n32364_), .ZN(new_n32365_));
  AOI21_X1   g29100(.A1(new_n8685_), .A2(new_n32365_), .B(new_n32073_), .ZN(new_n32366_));
  NOR2_X1    g29101(.A1(new_n32074_), .A2(new_n32365_), .ZN(new_n32367_));
  NOR3_X1    g29102(.A1(new_n32366_), .A2(new_n32363_), .A3(new_n32367_), .ZN(new_n32368_));
  INV_X1     g29103(.I(new_n32120_), .ZN(new_n32369_));
  INV_X1     g29104(.I(new_n32203_), .ZN(new_n32370_));
  OAI21_X1   g29105(.A1(new_n8683_), .A2(new_n32370_), .B(new_n32278_), .ZN(new_n32371_));
  NAND3_X1   g29106(.A1(new_n32371_), .A2(pi0214), .A3(new_n32228_), .ZN(new_n32372_));
  NOR2_X1    g29107(.A1(new_n32278_), .A2(new_n8685_), .ZN(new_n32373_));
  NAND2_X1   g29108(.A1(new_n32373_), .A2(new_n31760_), .ZN(new_n32374_));
  AOI21_X1   g29109(.A1(new_n32372_), .A2(new_n32369_), .B(new_n32374_), .ZN(new_n32375_));
  OAI21_X1   g29110(.A1(new_n32368_), .A2(pi1152), .B(new_n32375_), .ZN(new_n32376_));
  AOI21_X1   g29111(.A1(new_n32362_), .A2(new_n32286_), .B(new_n32376_), .ZN(new_n32377_));
  AOI21_X1   g29112(.A1(new_n32264_), .A2(new_n32377_), .B(new_n30557_), .ZN(new_n32378_));
  NAND2_X1   g29113(.A1(new_n31668_), .A2(pi0219), .ZN(new_n32379_));
  AOI21_X1   g29114(.A1(new_n32379_), .A2(new_n8685_), .B(new_n31816_), .ZN(new_n32380_));
  AOI21_X1   g29115(.A1(new_n32380_), .A2(pi1152), .B(pi0212), .ZN(new_n32381_));
  NAND2_X1   g29116(.A1(new_n31604_), .A2(new_n8739_), .ZN(new_n32382_));
  AOI21_X1   g29117(.A1(new_n31785_), .A2(new_n32382_), .B(new_n30597_), .ZN(new_n32383_));
  NAND3_X1   g29118(.A1(new_n31637_), .A2(new_n31653_), .A3(new_n8740_), .ZN(new_n32384_));
  XNOR2_X1   g29119(.A1(new_n32383_), .A2(new_n32384_), .ZN(new_n32385_));
  NAND2_X1   g29120(.A1(new_n7240_), .A2(new_n8683_), .ZN(new_n32386_));
  NAND2_X1   g29121(.A1(new_n32386_), .A2(new_n31653_), .ZN(new_n32387_));
  OAI21_X1   g29122(.A1(new_n32387_), .A2(new_n31002_), .B(new_n8683_), .ZN(new_n32388_));
  AOI21_X1   g29123(.A1(new_n31620_), .A2(pi0219), .B(po1038), .ZN(new_n32389_));
  INV_X1     g29124(.I(new_n32389_), .ZN(new_n32390_));
  AOI22_X1   g29125(.A1(new_n31804_), .A2(new_n31620_), .B1(new_n32390_), .B2(new_n32142_), .ZN(new_n32391_));
  INV_X1     g29126(.I(new_n32391_), .ZN(new_n32392_));
  OAI21_X1   g29127(.A1(new_n32343_), .A2(new_n8685_), .B(new_n31523_), .ZN(new_n32393_));
  NAND2_X1   g29128(.A1(new_n32393_), .A2(new_n31601_), .ZN(new_n32394_));
  NAND2_X1   g29129(.A1(new_n32394_), .A2(new_n32346_), .ZN(new_n32395_));
  NOR2_X1    g29130(.A1(new_n31804_), .A2(pi0299), .ZN(new_n32396_));
  AOI21_X1   g29131(.A1(new_n32395_), .A2(new_n32396_), .B(new_n31620_), .ZN(new_n32397_));
  AOI21_X1   g29132(.A1(new_n32397_), .A2(new_n32389_), .B(pi1152), .ZN(new_n32398_));
  AOI22_X1   g29133(.A1(new_n32398_), .A2(new_n32392_), .B1(new_n32385_), .B2(new_n32388_), .ZN(new_n32399_));
  NOR3_X1    g29134(.A1(new_n32399_), .A2(pi1150), .A3(pi1151), .ZN(new_n32400_));
  AOI21_X1   g29135(.A1(new_n31692_), .A2(new_n31683_), .B(pi0299), .ZN(new_n32401_));
  NAND2_X1   g29136(.A1(new_n32401_), .A2(pi0219), .ZN(new_n32402_));
  AOI21_X1   g29137(.A1(new_n32402_), .A2(new_n31238_), .B(new_n31680_), .ZN(new_n32403_));
  AOI21_X1   g29138(.A1(new_n7240_), .A2(new_n31002_), .B(new_n8683_), .ZN(new_n32404_));
  NAND2_X1   g29139(.A1(new_n31801_), .A2(new_n32404_), .ZN(new_n32405_));
  INV_X1     g29140(.I(new_n31993_), .ZN(new_n32406_));
  NOR2_X1    g29141(.A1(new_n32406_), .A2(new_n32250_), .ZN(new_n32407_));
  OAI21_X1   g29142(.A1(new_n32403_), .A2(new_n32405_), .B(new_n32407_), .ZN(new_n32408_));
  OAI22_X1   g29143(.A1(new_n32400_), .A2(new_n32408_), .B1(new_n31816_), .B2(new_n32381_), .ZN(new_n32409_));
  AOI21_X1   g29144(.A1(new_n31825_), .A2(new_n32409_), .B(new_n31941_), .ZN(new_n32410_));
  AOI21_X1   g29145(.A1(new_n31691_), .A2(new_n8685_), .B(new_n8739_), .ZN(new_n32411_));
  NAND2_X1   g29146(.A1(new_n32096_), .A2(new_n32411_), .ZN(new_n32412_));
  AOI21_X1   g29147(.A1(new_n32412_), .A2(new_n31682_), .B(new_n32401_), .ZN(new_n32413_));
  AND4_X2    g29148(.A1(pi0219), .A2(new_n32413_), .A3(pi1152), .A4(new_n31678_), .Z(new_n32414_));
  NOR2_X1    g29149(.A1(new_n31819_), .A2(new_n8739_), .ZN(new_n32415_));
  XOR2_X1    g29150(.A1(new_n32415_), .A2(new_n30597_), .Z(new_n32416_));
  NOR3_X1    g29151(.A1(new_n32416_), .A2(new_n31816_), .A3(new_n32240_), .ZN(new_n32417_));
  OAI21_X1   g29152(.A1(new_n32380_), .A2(new_n32414_), .B(new_n32417_), .ZN(new_n32418_));
  NAND2_X1   g29153(.A1(new_n32418_), .A2(new_n32390_), .ZN(new_n32419_));
  AOI21_X1   g29154(.A1(new_n32419_), .A2(new_n32052_), .B(new_n32242_), .ZN(new_n32420_));
  INV_X1     g29155(.I(new_n32398_), .ZN(new_n32421_));
  AOI21_X1   g29156(.A1(po1038), .A2(new_n31653_), .B(new_n32397_), .ZN(new_n32422_));
  OAI21_X1   g29157(.A1(new_n32422_), .A2(new_n8683_), .B(pi1152), .ZN(new_n32423_));
  NOR2_X1    g29158(.A1(new_n31611_), .A2(new_n31797_), .ZN(new_n32424_));
  OAI21_X1   g29159(.A1(new_n7240_), .A2(new_n31978_), .B(pi1151), .ZN(new_n32425_));
  OAI21_X1   g29160(.A1(new_n31818_), .A2(new_n31002_), .B(new_n31980_), .ZN(new_n32426_));
  NAND2_X1   g29161(.A1(new_n32426_), .A2(new_n31627_), .ZN(new_n32427_));
  AOI21_X1   g29162(.A1(new_n32427_), .A2(new_n7240_), .B(new_n32425_), .ZN(new_n32428_));
  AOI21_X1   g29163(.A1(new_n32315_), .A2(new_n31680_), .B(new_n32425_), .ZN(new_n32429_));
  NOR2_X1    g29164(.A1(new_n31620_), .A2(new_n31651_), .ZN(new_n32430_));
  NAND3_X1   g29165(.A1(new_n31670_), .A2(pi1150), .A3(pi1152), .ZN(new_n32431_));
  NOR4_X1    g29166(.A1(new_n32430_), .A2(new_n31996_), .A3(new_n32429_), .A4(new_n32431_), .ZN(new_n32432_));
  OAI21_X1   g29167(.A1(new_n32428_), .A2(new_n32424_), .B(new_n32432_), .ZN(new_n32433_));
  AOI21_X1   g29168(.A1(new_n32423_), .A2(new_n32421_), .B(new_n32433_), .ZN(new_n32434_));
  XOR2_X1    g29169(.A1(new_n32420_), .A2(new_n32434_), .Z(new_n32435_));
  NAND2_X1   g29170(.A1(new_n31824_), .A2(new_n31002_), .ZN(new_n32436_));
  AOI21_X1   g29171(.A1(new_n31816_), .A2(new_n31593_), .B(new_n8739_), .ZN(new_n32437_));
  NOR3_X1    g29172(.A1(new_n31822_), .A2(new_n8739_), .A3(new_n31818_), .ZN(new_n32438_));
  XOR2_X1    g29173(.A1(new_n32438_), .A2(new_n32437_), .Z(new_n32439_));
  NAND2_X1   g29174(.A1(new_n32387_), .A2(new_n31002_), .ZN(new_n32440_));
  NAND3_X1   g29175(.A1(new_n31804_), .A2(new_n31653_), .A3(new_n32440_), .ZN(new_n32441_));
  NAND2_X1   g29176(.A1(new_n32441_), .A2(new_n32259_), .ZN(new_n32442_));
  NAND3_X1   g29177(.A1(new_n32442_), .A2(pi1152), .A3(new_n32391_), .ZN(new_n32443_));
  OAI21_X1   g29178(.A1(new_n32257_), .A2(new_n32405_), .B(new_n8683_), .ZN(new_n32444_));
  INV_X1     g29179(.I(new_n31801_), .ZN(new_n32445_));
  NOR3_X1    g29180(.A1(new_n31679_), .A2(pi0214), .A3(new_n10253_), .ZN(new_n32446_));
  NAND2_X1   g29181(.A1(new_n31614_), .A2(pi0212), .ZN(new_n32447_));
  OAI22_X1   g29182(.A1(new_n31787_), .A2(new_n32445_), .B1(new_n32446_), .B2(new_n32447_), .ZN(new_n32448_));
  NAND4_X1   g29183(.A1(new_n32448_), .A2(pi0219), .A3(pi1149), .A4(new_n32444_), .ZN(new_n32449_));
  AOI21_X1   g29184(.A1(new_n32443_), .A2(new_n32242_), .B(new_n32449_), .ZN(new_n32450_));
  NAND4_X1   g29185(.A1(new_n32435_), .A2(new_n32436_), .A3(new_n32439_), .A4(new_n32450_), .ZN(new_n32451_));
  OAI21_X1   g29186(.A1(new_n32451_), .A2(new_n32410_), .B(pi0209), .ZN(new_n32452_));
  AOI21_X1   g29187(.A1(new_n32410_), .A2(new_n32451_), .B(new_n32452_), .ZN(new_n32453_));
  XOR2_X1    g29188(.A1(new_n32453_), .A2(new_n31079_), .Z(new_n32454_));
  NAND4_X1   g29189(.A1(new_n32454_), .A2(pi0230), .A3(pi0241), .A4(new_n31834_), .ZN(new_n32455_));
  XNOR2_X1   g29190(.A1(new_n32455_), .A2(new_n32378_), .ZN(po0398));
  NOR2_X1    g29191(.A1(new_n31903_), .A2(new_n8555_), .ZN(new_n32457_));
  NOR2_X1    g29192(.A1(new_n32457_), .A2(pi0299), .ZN(new_n32458_));
  AOI21_X1   g29193(.A1(pi0199), .A2(pi1144), .B(pi0200), .ZN(new_n32459_));
  NAND2_X1   g29194(.A1(new_n31900_), .A2(new_n32459_), .ZN(new_n32460_));
  NOR2_X1    g29195(.A1(new_n32458_), .A2(new_n32460_), .ZN(new_n32461_));
  NOR2_X1    g29196(.A1(new_n32461_), .A2(new_n8546_), .ZN(new_n32462_));
  XOR2_X1    g29197(.A1(new_n32462_), .A2(new_n8547_), .Z(new_n32463_));
  NAND4_X1   g29198(.A1(new_n27298_), .A2(pi0199), .A3(new_n8555_), .A4(new_n3057_), .ZN(new_n32464_));
  AOI21_X1   g29199(.A1(new_n32464_), .A2(new_n3518_), .B(new_n8549_), .ZN(new_n32465_));
  NAND2_X1   g29200(.A1(new_n32463_), .A2(new_n32465_), .ZN(new_n32466_));
  INV_X1     g29201(.I(new_n32466_), .ZN(new_n32467_));
  INV_X1     g29202(.I(new_n32461_), .ZN(new_n32468_));
  NOR2_X1    g29203(.A1(new_n32468_), .A2(new_n31450_), .ZN(new_n32469_));
  NOR2_X1    g29204(.A1(new_n32467_), .A2(new_n32469_), .ZN(new_n32470_));
  INV_X1     g29205(.I(new_n32470_), .ZN(new_n32471_));
  NOR2_X1    g29206(.A1(new_n32471_), .A2(new_n31912_), .ZN(new_n32472_));
  INV_X1     g29207(.I(new_n32472_), .ZN(new_n32473_));
  NOR2_X1    g29208(.A1(new_n32473_), .A2(pi0211), .ZN(new_n32474_));
  NOR2_X1    g29209(.A1(new_n32471_), .A2(new_n31503_), .ZN(new_n32475_));
  AOI21_X1   g29210(.A1(pi0211), .A2(new_n32475_), .B(new_n32474_), .ZN(new_n32476_));
  NOR2_X1    g29211(.A1(new_n32468_), .A2(new_n30966_), .ZN(new_n32477_));
  NOR2_X1    g29212(.A1(new_n32467_), .A2(new_n32477_), .ZN(new_n32478_));
  AOI21_X1   g29213(.A1(new_n32478_), .A2(new_n8685_), .B(pi0212), .ZN(new_n32479_));
  NAND2_X1   g29214(.A1(new_n32479_), .A2(pi0219), .ZN(new_n32480_));
  AOI21_X1   g29215(.A1(new_n8685_), .A2(new_n32480_), .B(new_n32476_), .ZN(new_n32481_));
  INV_X1     g29216(.I(new_n32478_), .ZN(new_n32482_));
  AOI21_X1   g29217(.A1(new_n32482_), .A2(new_n30604_), .B(new_n8683_), .ZN(new_n32483_));
  AOI21_X1   g29218(.A1(new_n32483_), .A2(po1038), .B(new_n30594_), .ZN(new_n32484_));
  NOR2_X1    g29219(.A1(new_n32003_), .A2(pi0214), .ZN(new_n32485_));
  AOI21_X1   g29220(.A1(pi0214), .A2(new_n31385_), .B(new_n32485_), .ZN(new_n32486_));
  AOI21_X1   g29221(.A1(new_n32003_), .A2(pi0214), .B(new_n8739_), .ZN(new_n32487_));
  XOR2_X1    g29222(.A1(new_n32487_), .A2(new_n30916_), .Z(new_n32488_));
  NOR2_X1    g29223(.A1(new_n32488_), .A2(new_n32486_), .ZN(new_n32489_));
  AOI21_X1   g29224(.A1(new_n8684_), .A2(pi1144), .B(new_n8683_), .ZN(new_n32490_));
  NOR3_X1    g29225(.A1(new_n32489_), .A2(new_n30918_), .A3(new_n32490_), .ZN(new_n32491_));
  INV_X1     g29226(.I(new_n32491_), .ZN(new_n32492_));
  NOR4_X1    g29227(.A1(new_n32484_), .A2(new_n30879_), .A3(new_n32470_), .A4(new_n32492_), .ZN(new_n32493_));
  NOR2_X1    g29228(.A1(new_n32481_), .A2(new_n32493_), .ZN(new_n32494_));
  NOR2_X1    g29229(.A1(new_n32475_), .A2(new_n8685_), .ZN(new_n32495_));
  XOR2_X1    g29230(.A1(new_n32495_), .A2(new_n8686_), .Z(new_n32496_));
  NAND4_X1   g29231(.A1(new_n32496_), .A2(pi0299), .A3(pi1144), .A4(new_n32471_), .ZN(new_n32497_));
  NAND2_X1   g29232(.A1(new_n32497_), .A2(new_n8739_), .ZN(new_n32498_));
  NOR2_X1    g29233(.A1(new_n32476_), .A2(new_n8685_), .ZN(new_n32499_));
  NAND2_X1   g29234(.A1(new_n32498_), .A2(new_n32499_), .ZN(new_n32500_));
  NOR2_X1    g29235(.A1(new_n32500_), .A2(new_n32494_), .ZN(new_n32501_));
  INV_X1     g29236(.I(new_n32501_), .ZN(new_n32502_));
  NOR2_X1    g29237(.A1(new_n30590_), .A2(new_n8739_), .ZN(new_n32503_));
  XOR2_X1    g29238(.A1(new_n30590_), .A2(new_n30597_), .Z(new_n32504_));
  NAND2_X1   g29239(.A1(new_n32504_), .A2(new_n30562_), .ZN(new_n32505_));
  NOR2_X1    g29240(.A1(new_n32469_), .A2(pi0219), .ZN(new_n32506_));
  OAI21_X1   g29241(.A1(new_n32505_), .A2(new_n32503_), .B(new_n32506_), .ZN(new_n32507_));
  AOI21_X1   g29242(.A1(new_n32503_), .A2(new_n32505_), .B(new_n32507_), .ZN(new_n32508_));
  OAI21_X1   g29243(.A1(new_n31238_), .A2(new_n32477_), .B(new_n32467_), .ZN(new_n32509_));
  OAI21_X1   g29244(.A1(new_n32508_), .A2(new_n32509_), .B(new_n8683_), .ZN(new_n32510_));
  NOR4_X1    g29245(.A1(new_n32468_), .A2(new_n30604_), .A3(new_n30901_), .A4(new_n30966_), .ZN(new_n32511_));
  NOR3_X1    g29246(.A1(new_n32468_), .A2(new_n8684_), .A3(new_n31450_), .ZN(new_n32512_));
  OAI21_X1   g29247(.A1(new_n32511_), .A2(new_n32512_), .B(new_n31300_), .ZN(new_n32513_));
  AOI21_X1   g29248(.A1(new_n30843_), .A2(new_n28529_), .B(new_n32513_), .ZN(new_n32514_));
  AOI21_X1   g29249(.A1(new_n32510_), .A2(new_n32514_), .B(pi0213), .ZN(new_n32515_));
  OAI21_X1   g29250(.A1(new_n32502_), .A2(new_n32515_), .B(pi0230), .ZN(new_n32516_));
  NOR2_X1    g29251(.A1(new_n30609_), .A2(new_n28529_), .ZN(new_n32517_));
  XOR2_X1    g29252(.A1(new_n32517_), .A2(new_n31079_), .Z(new_n32518_));
  INV_X1     g29253(.I(new_n32490_), .ZN(new_n32520_));
  NAND2_X1   g29254(.A1(po1038), .A2(pi0299), .ZN(new_n32521_));
  INV_X1     g29255(.I(new_n32521_), .ZN(new_n32522_));
  NOR2_X1    g29256(.A1(new_n30580_), .A2(new_n30577_), .ZN(new_n32524_));
  NOR4_X1    g29257(.A1(new_n32524_), .A2(new_n30557_), .A3(new_n5364_), .A4(new_n3098_), .ZN(new_n32525_));
  NAND2_X1   g29258(.A1(new_n32518_), .A2(new_n32525_), .ZN(new_n32526_));
  XOR2_X1    g29259(.A1(new_n32516_), .A2(new_n32526_), .Z(po0399));
  NOR3_X1    g29260(.A1(pi0081), .A2(pi0085), .A3(pi0314), .ZN(new_n32528_));
  NOR2_X1    g29261(.A1(new_n32528_), .A2(new_n2630_), .ZN(new_n32529_));
  INV_X1     g29262(.I(new_n32529_), .ZN(new_n32530_));
  NAND2_X1   g29263(.A1(pi0276), .A2(pi0802), .ZN(new_n32531_));
  NOR2_X1    g29264(.A1(new_n32530_), .A2(new_n32531_), .ZN(new_n32532_));
  INV_X1     g29265(.I(new_n32532_), .ZN(new_n32533_));
  NOR2_X1    g29266(.A1(new_n32533_), .A2(pi1091), .ZN(new_n32534_));
  INV_X1     g29267(.I(new_n32534_), .ZN(new_n32535_));
  AND2_X2    g29268(.A1(pi0271), .A2(pi0273), .Z(new_n32536_));
  INV_X1     g29269(.I(new_n32536_), .ZN(new_n32537_));
  NOR2_X1    g29270(.A1(new_n32535_), .A2(new_n32537_), .ZN(new_n32538_));
  NOR2_X1    g29271(.A1(new_n32538_), .A2(new_n3098_), .ZN(new_n32539_));
  AOI21_X1   g29272(.A1(new_n2630_), .A2(new_n2575_), .B(new_n9231_), .ZN(new_n32540_));
  INV_X1     g29273(.I(new_n32540_), .ZN(new_n32541_));
  NOR2_X1    g29274(.A1(new_n32541_), .A2(new_n32531_), .ZN(new_n32542_));
  INV_X1     g29275(.I(new_n32542_), .ZN(new_n32543_));
  NAND2_X1   g29276(.A1(pi0273), .A2(pi1091), .ZN(new_n32544_));
  NAND2_X1   g29277(.A1(new_n32543_), .A2(new_n32544_), .ZN(new_n32545_));
  NAND2_X1   g29278(.A1(new_n32545_), .A2(pi0271), .ZN(new_n32546_));
  INV_X1     g29279(.I(new_n32546_), .ZN(new_n32547_));
  NOR2_X1    g29280(.A1(new_n32547_), .A2(pi1091), .ZN(new_n32548_));
  NOR2_X1    g29281(.A1(new_n32548_), .A2(new_n8549_), .ZN(new_n32549_));
  NOR2_X1    g29282(.A1(new_n32538_), .A2(new_n32547_), .ZN(new_n32550_));
  NAND2_X1   g29283(.A1(new_n32550_), .A2(new_n2726_), .ZN(new_n32551_));
  INV_X1     g29284(.I(new_n32551_), .ZN(new_n32552_));
  NOR2_X1    g29285(.A1(new_n32552_), .A2(pi0199), .ZN(new_n32553_));
  NOR2_X1    g29286(.A1(new_n32553_), .A2(new_n32549_), .ZN(new_n32554_));
  INV_X1     g29287(.I(new_n32554_), .ZN(new_n32555_));
  AOI21_X1   g29288(.A1(new_n32555_), .A2(new_n32534_), .B(pi0299), .ZN(new_n32556_));
  INV_X1     g29289(.I(new_n32556_), .ZN(new_n32557_));
  NOR2_X1    g29290(.A1(new_n32548_), .A2(pi0200), .ZN(new_n32558_));
  NOR2_X1    g29291(.A1(new_n32557_), .A2(new_n32558_), .ZN(new_n32559_));
  NOR2_X1    g29292(.A1(new_n32559_), .A2(new_n32539_), .ZN(new_n32560_));
  NAND3_X1   g29293(.A1(new_n32560_), .A2(new_n13778_), .A3(new_n32535_), .ZN(new_n32561_));
  NAND2_X1   g29294(.A1(new_n32561_), .A2(pi0243), .ZN(new_n32562_));
  NOR2_X1    g29295(.A1(new_n32543_), .A2(pi1091), .ZN(new_n32563_));
  INV_X1     g29296(.I(new_n32563_), .ZN(new_n32564_));
  NOR2_X1    g29297(.A1(new_n32564_), .A2(new_n32537_), .ZN(new_n32565_));
  NOR2_X1    g29298(.A1(new_n32565_), .A2(new_n3098_), .ZN(new_n32566_));
  NOR2_X1    g29299(.A1(new_n32557_), .A2(new_n32553_), .ZN(new_n32567_));
  NOR2_X1    g29300(.A1(new_n32567_), .A2(new_n32566_), .ZN(new_n32568_));
  AOI21_X1   g29301(.A1(new_n32554_), .A2(pi0299), .B(pi0200), .ZN(new_n32569_));
  NOR2_X1    g29302(.A1(new_n32569_), .A2(new_n32535_), .ZN(new_n32570_));
  INV_X1     g29303(.I(new_n32570_), .ZN(new_n32571_));
  OAI21_X1   g29304(.A1(pi1155), .A2(new_n32571_), .B(new_n32568_), .ZN(new_n32572_));
  NOR2_X1    g29305(.A1(new_n32557_), .A2(new_n32549_), .ZN(new_n32573_));
  INV_X1     g29306(.I(new_n32548_), .ZN(new_n32574_));
  NOR2_X1    g29307(.A1(new_n32574_), .A2(new_n3098_), .ZN(new_n32575_));
  NOR2_X1    g29308(.A1(new_n32573_), .A2(new_n32575_), .ZN(new_n32576_));
  NAND3_X1   g29309(.A1(new_n32572_), .A2(pi0243), .A3(new_n32576_), .ZN(new_n32577_));
  XOR2_X1    g29310(.A1(new_n32577_), .A2(new_n32562_), .Z(new_n32578_));
  INV_X1     g29311(.I(pi0243), .ZN(new_n32579_));
  NOR2_X1    g29312(.A1(new_n32571_), .A2(new_n32549_), .ZN(new_n32580_));
  INV_X1     g29313(.I(new_n32559_), .ZN(new_n32581_));
  NOR2_X1    g29314(.A1(new_n32581_), .A2(new_n32553_), .ZN(new_n32582_));
  NOR2_X1    g29315(.A1(new_n32582_), .A2(new_n32566_), .ZN(new_n32583_));
  INV_X1     g29316(.I(new_n32583_), .ZN(new_n32584_));
  NOR2_X1    g29317(.A1(new_n32584_), .A2(new_n32580_), .ZN(new_n32585_));
  INV_X1     g29318(.I(new_n32585_), .ZN(new_n32586_));
  INV_X1     g29319(.I(new_n32573_), .ZN(new_n32587_));
  NOR2_X1    g29320(.A1(new_n32587_), .A2(new_n32558_), .ZN(new_n32588_));
  NOR2_X1    g29321(.A1(new_n32588_), .A2(new_n32575_), .ZN(new_n32589_));
  INV_X1     g29322(.I(new_n32589_), .ZN(new_n32590_));
  NAND2_X1   g29323(.A1(new_n32590_), .A2(new_n32579_), .ZN(new_n32591_));
  OAI21_X1   g29324(.A1(new_n32586_), .A2(new_n32579_), .B(new_n32591_), .ZN(new_n32592_));
  NOR2_X1    g29325(.A1(new_n32559_), .A2(new_n32566_), .ZN(new_n32593_));
  INV_X1     g29326(.I(new_n32593_), .ZN(new_n32594_));
  NOR2_X1    g29327(.A1(new_n32594_), .A2(new_n32573_), .ZN(new_n32595_));
  NOR2_X1    g29328(.A1(new_n32595_), .A2(new_n32579_), .ZN(new_n32596_));
  INV_X1     g29329(.I(new_n32539_), .ZN(new_n32597_));
  NOR2_X1    g29330(.A1(new_n32597_), .A2(new_n32574_), .ZN(new_n32598_));
  NOR2_X1    g29331(.A1(new_n32570_), .A2(new_n32598_), .ZN(new_n32599_));
  INV_X1     g29332(.I(new_n32599_), .ZN(new_n32600_));
  NOR4_X1    g29333(.A1(new_n32594_), .A2(new_n32600_), .A3(new_n32579_), .A4(new_n13778_), .ZN(new_n32601_));
  XOR2_X1    g29334(.A1(new_n32596_), .A2(new_n32601_), .Z(new_n32602_));
  NOR2_X1    g29335(.A1(new_n32571_), .A2(new_n32553_), .ZN(new_n32603_));
  NOR2_X1    g29336(.A1(new_n32603_), .A2(new_n32575_), .ZN(new_n32604_));
  INV_X1     g29337(.I(new_n32604_), .ZN(new_n32605_));
  NOR2_X1    g29338(.A1(pi0211), .A2(pi1157), .ZN(new_n32606_));
  NOR3_X1    g29339(.A1(new_n32605_), .A2(new_n13969_), .A3(new_n32606_), .ZN(new_n32607_));
  AOI21_X1   g29340(.A1(new_n32602_), .A2(new_n32607_), .B(new_n32592_), .ZN(new_n32608_));
  NAND2_X1   g29341(.A1(pi0243), .A2(pi1155), .ZN(new_n32609_));
  NOR2_X1    g29342(.A1(new_n32583_), .A2(new_n13778_), .ZN(new_n32610_));
  XOR2_X1    g29343(.A1(new_n32610_), .A2(new_n32609_), .Z(new_n32611_));
  NOR3_X1    g29344(.A1(new_n32611_), .A2(new_n13778_), .A3(new_n32600_), .ZN(new_n32612_));
  INV_X1     g29345(.I(new_n32567_), .ZN(new_n32613_));
  NAND3_X1   g29346(.A1(new_n32593_), .A2(new_n32613_), .A3(pi0243), .ZN(new_n32614_));
  NAND2_X1   g29347(.A1(new_n32614_), .A2(new_n13778_), .ZN(new_n32615_));
  NOR2_X1    g29348(.A1(new_n32580_), .A2(new_n32575_), .ZN(new_n32616_));
  NAND3_X1   g29349(.A1(new_n32615_), .A2(pi0243), .A3(new_n32616_), .ZN(new_n32617_));
  NOR2_X1    g29350(.A1(pi1156), .A2(pi1157), .ZN(new_n32618_));
  NOR2_X1    g29351(.A1(new_n32556_), .A2(new_n32566_), .ZN(new_n32619_));
  NAND2_X1   g29352(.A1(new_n13778_), .A2(pi0243), .ZN(new_n32620_));
  NAND4_X1   g29353(.A1(new_n32604_), .A2(pi1091), .A3(new_n32619_), .A4(new_n32620_), .ZN(new_n32621_));
  AOI21_X1   g29354(.A1(new_n32617_), .A2(new_n32618_), .B(new_n32621_), .ZN(new_n32622_));
  OAI21_X1   g29355(.A1(new_n32612_), .A2(pi0243), .B(new_n32622_), .ZN(new_n32623_));
  OAI21_X1   g29356(.A1(new_n32623_), .A2(new_n32608_), .B(new_n13969_), .ZN(new_n32624_));
  INV_X1     g29357(.I(pi0267), .ZN(new_n32625_));
  INV_X1     g29358(.I(pi0253), .ZN(new_n32626_));
  INV_X1     g29359(.I(pi0254), .ZN(new_n32627_));
  NOR2_X1    g29360(.A1(new_n32626_), .A2(new_n32627_), .ZN(new_n32628_));
  INV_X1     g29361(.I(new_n32628_), .ZN(new_n32629_));
  NOR2_X1    g29362(.A1(new_n32629_), .A2(new_n32625_), .ZN(new_n32630_));
  INV_X1     g29363(.I(new_n32630_), .ZN(new_n32631_));
  NOR2_X1    g29364(.A1(new_n32631_), .A2(pi0263), .ZN(new_n32632_));
  AOI22_X1   g29365(.A1(new_n32624_), .A2(new_n32578_), .B1(pi0219), .B2(new_n32632_), .ZN(new_n32633_));
  NOR2_X1    g29366(.A1(new_n32603_), .A2(new_n32566_), .ZN(new_n32634_));
  NAND3_X1   g29367(.A1(new_n32634_), .A2(pi0243), .A3(pi1155), .ZN(new_n32635_));
  INV_X1     g29368(.I(new_n32634_), .ZN(new_n32636_));
  NAND3_X1   g29369(.A1(new_n32636_), .A2(pi0243), .A3(new_n13778_), .ZN(new_n32637_));
  NAND2_X1   g29370(.A1(new_n32637_), .A2(new_n32635_), .ZN(new_n32638_));
  NOR2_X1    g29371(.A1(new_n32570_), .A2(new_n32566_), .ZN(new_n32639_));
  INV_X1     g29372(.I(new_n32639_), .ZN(new_n32640_));
  NOR2_X1    g29373(.A1(pi1155), .A2(pi1156), .ZN(new_n32641_));
  NAND2_X1   g29374(.A1(new_n32640_), .A2(new_n32641_), .ZN(new_n32642_));
  AOI22_X1   g29375(.A1(new_n32638_), .A2(new_n32573_), .B1(pi0243), .B2(new_n32642_), .ZN(new_n32643_));
  NOR2_X1    g29376(.A1(new_n32559_), .A2(new_n32575_), .ZN(new_n32644_));
  NAND2_X1   g29377(.A1(new_n32644_), .A2(pi0243), .ZN(new_n32645_));
  OAI22_X1   g29378(.A1(new_n32643_), .A2(new_n32645_), .B1(pi0211), .B2(new_n14006_), .ZN(new_n32646_));
  INV_X1     g29379(.I(new_n32644_), .ZN(new_n32647_));
  NOR2_X1    g29380(.A1(pi0243), .A2(pi1155), .ZN(new_n32648_));
  AOI21_X1   g29381(.A1(new_n32586_), .A2(new_n32648_), .B(new_n32647_), .ZN(new_n32649_));
  NOR3_X1    g29382(.A1(new_n32649_), .A2(new_n32589_), .A3(new_n32639_), .ZN(new_n32650_));
  NOR2_X1    g29383(.A1(new_n32579_), .A2(new_n2726_), .ZN(new_n32651_));
  NOR2_X1    g29384(.A1(new_n32588_), .A2(new_n32539_), .ZN(new_n32652_));
  INV_X1     g29385(.I(new_n32652_), .ZN(new_n32653_));
  NAND2_X1   g29386(.A1(new_n32653_), .A2(new_n2726_), .ZN(new_n32654_));
  AOI21_X1   g29387(.A1(new_n32654_), .A2(new_n32604_), .B(new_n32651_), .ZN(new_n32655_));
  OAI21_X1   g29388(.A1(new_n32650_), .A2(new_n32609_), .B(new_n32655_), .ZN(new_n32656_));
  NAND4_X1   g29389(.A1(new_n32656_), .A2(new_n32646_), .A3(pi1156), .A4(new_n32592_), .ZN(new_n32657_));
  NOR2_X1    g29390(.A1(new_n32633_), .A2(new_n32657_), .ZN(new_n32658_));
  NOR2_X1    g29391(.A1(new_n32582_), .A2(new_n32598_), .ZN(new_n32659_));
  INV_X1     g29392(.I(new_n32649_), .ZN(new_n32660_));
  NOR2_X1    g29393(.A1(new_n32570_), .A2(new_n32539_), .ZN(new_n32661_));
  INV_X1     g29394(.I(new_n32661_), .ZN(new_n32662_));
  NOR4_X1    g29395(.A1(new_n32660_), .A2(pi0243), .A3(new_n32588_), .A4(new_n32662_), .ZN(new_n32663_));
  OAI21_X1   g29396(.A1(new_n32663_), .A2(pi1155), .B(new_n32659_), .ZN(new_n32664_));
  NOR2_X1    g29397(.A1(new_n32582_), .A2(new_n32579_), .ZN(new_n32665_));
  INV_X1     g29398(.I(new_n32665_), .ZN(new_n32666_));
  NOR2_X1    g29399(.A1(new_n32588_), .A2(new_n32603_), .ZN(new_n32667_));
  INV_X1     g29400(.I(new_n32667_), .ZN(new_n32668_));
  NOR2_X1    g29401(.A1(new_n32580_), .A2(new_n32539_), .ZN(new_n32669_));
  INV_X1     g29402(.I(new_n32669_), .ZN(new_n32670_));
  NOR4_X1    g29403(.A1(new_n32668_), .A2(new_n32579_), .A3(new_n32598_), .A4(new_n32670_), .ZN(new_n32671_));
  AOI21_X1   g29404(.A1(new_n32671_), .A2(new_n32666_), .B(pi1155), .ZN(new_n32672_));
  OAI21_X1   g29405(.A1(new_n32666_), .A2(new_n32671_), .B(new_n32672_), .ZN(new_n32673_));
  NAND2_X1   g29406(.A1(new_n32664_), .A2(new_n32673_), .ZN(new_n32674_));
  NOR2_X1    g29407(.A1(new_n32559_), .A2(new_n32598_), .ZN(new_n32675_));
  NOR2_X1    g29408(.A1(new_n32661_), .A2(pi0243), .ZN(new_n32676_));
  AOI21_X1   g29409(.A1(new_n32675_), .A2(pi0243), .B(new_n32676_), .ZN(new_n32677_));
  NOR2_X1    g29410(.A1(new_n32556_), .A2(new_n32539_), .ZN(new_n32678_));
  NOR2_X1    g29411(.A1(pi0243), .A2(pi1091), .ZN(new_n32679_));
  INV_X1     g29412(.I(new_n32679_), .ZN(new_n32680_));
  OAI21_X1   g29413(.A1(new_n32619_), .A2(new_n32680_), .B(new_n32678_), .ZN(new_n32681_));
  NAND2_X1   g29414(.A1(new_n32678_), .A2(pi1155), .ZN(new_n32682_));
  XNOR2_X1   g29415(.A1(new_n32681_), .A2(new_n32682_), .ZN(new_n32683_));
  OAI21_X1   g29416(.A1(new_n32683_), .A2(new_n32579_), .B(new_n13969_), .ZN(new_n32684_));
  OAI21_X1   g29417(.A1(new_n32684_), .A2(new_n13778_), .B(new_n32677_), .ZN(new_n32685_));
  NOR2_X1    g29418(.A1(new_n32567_), .A2(new_n32598_), .ZN(new_n32686_));
  NOR2_X1    g29419(.A1(new_n32573_), .A2(new_n32539_), .ZN(new_n32687_));
  NOR2_X1    g29420(.A1(new_n32687_), .A2(pi0243), .ZN(new_n32688_));
  AOI21_X1   g29421(.A1(pi0243), .A2(new_n32686_), .B(new_n32688_), .ZN(new_n32689_));
  INV_X1     g29422(.I(new_n32606_), .ZN(new_n32690_));
  INV_X1     g29423(.I(new_n32675_), .ZN(new_n32691_));
  INV_X1     g29424(.I(new_n32689_), .ZN(new_n32692_));
  NAND3_X1   g29425(.A1(new_n32692_), .A2(pi1156), .A3(new_n32561_), .ZN(new_n32693_));
  NAND3_X1   g29426(.A1(new_n32693_), .A2(new_n13778_), .A3(new_n32691_), .ZN(new_n32694_));
  AOI21_X1   g29427(.A1(new_n32694_), .A2(new_n32661_), .B(new_n32690_), .ZN(new_n32695_));
  INV_X1     g29428(.I(new_n32560_), .ZN(new_n32696_));
  NOR3_X1    g29429(.A1(new_n32696_), .A2(new_n32579_), .A3(new_n32573_), .ZN(new_n32697_));
  INV_X1     g29430(.I(new_n32678_), .ZN(new_n32698_));
  AOI21_X1   g29431(.A1(new_n32605_), .A2(new_n32648_), .B(new_n32698_), .ZN(new_n32699_));
  OAI21_X1   g29432(.A1(new_n32699_), .A2(new_n32697_), .B(new_n13969_), .ZN(new_n32700_));
  NOR2_X1    g29433(.A1(new_n32700_), .A2(new_n32677_), .ZN(new_n32701_));
  NOR4_X1    g29434(.A1(new_n32695_), .A2(new_n14006_), .A3(new_n32689_), .A4(new_n32701_), .ZN(new_n32702_));
  AOI21_X1   g29435(.A1(new_n32702_), .A2(new_n32685_), .B(pi1156), .ZN(new_n32703_));
  OAI21_X1   g29436(.A1(new_n32674_), .A2(new_n32703_), .B(new_n8683_), .ZN(new_n32704_));
  NOR2_X1    g29437(.A1(new_n32579_), .A2(pi1091), .ZN(new_n32705_));
  INV_X1     g29438(.I(new_n32705_), .ZN(new_n32706_));
  OAI21_X1   g29439(.A1(new_n32674_), .A2(new_n13969_), .B(new_n32706_), .ZN(new_n32707_));
  NAND2_X1   g29440(.A1(new_n32707_), .A2(new_n32652_), .ZN(new_n32708_));
  NAND2_X1   g29441(.A1(new_n32708_), .A2(new_n14006_), .ZN(new_n32709_));
  AOI21_X1   g29442(.A1(new_n32696_), .A2(pi1155), .B(new_n32609_), .ZN(new_n32710_));
  NOR3_X1    g29443(.A1(new_n32560_), .A2(pi0243), .A3(new_n13778_), .ZN(new_n32711_));
  OAI21_X1   g29444(.A1(new_n32710_), .A2(new_n32711_), .B(new_n32599_), .ZN(new_n32712_));
  NOR2_X1    g29445(.A1(new_n32700_), .A2(new_n32712_), .ZN(new_n32713_));
  NOR2_X1    g29446(.A1(new_n32549_), .A2(pi1155), .ZN(new_n32714_));
  NAND2_X1   g29447(.A1(new_n32712_), .A2(new_n32714_), .ZN(new_n32715_));
  NAND2_X1   g29448(.A1(new_n32693_), .A2(new_n14006_), .ZN(new_n32716_));
  NAND3_X1   g29449(.A1(new_n32716_), .A2(new_n32705_), .A3(new_n32715_), .ZN(new_n32717_));
  INV_X1     g29450(.I(new_n32632_), .ZN(new_n32718_));
  NOR2_X1    g29451(.A1(new_n2726_), .A2(pi0299), .ZN(new_n32719_));
  NAND2_X1   g29452(.A1(new_n31153_), .A2(new_n32651_), .ZN(new_n32720_));
  XOR2_X1    g29453(.A1(new_n32720_), .A2(new_n32719_), .Z(new_n32721_));
  NOR2_X1    g29454(.A1(new_n32721_), .A2(new_n13969_), .ZN(new_n32722_));
  NOR2_X1    g29455(.A1(new_n31420_), .A2(pi0299), .ZN(new_n32723_));
  NOR2_X1    g29456(.A1(new_n32723_), .A2(new_n2726_), .ZN(new_n32724_));
  INV_X1     g29457(.I(new_n32724_), .ZN(new_n32725_));
  OAI21_X1   g29458(.A1(new_n2726_), .A2(new_n13778_), .B(new_n32680_), .ZN(new_n32726_));
  NAND3_X1   g29459(.A1(new_n32726_), .A2(pi1156), .A3(new_n30659_), .ZN(new_n32727_));
  AOI21_X1   g29460(.A1(new_n32727_), .A2(new_n32706_), .B(new_n32725_), .ZN(new_n32728_));
  NOR2_X1    g29461(.A1(new_n32728_), .A2(new_n32606_), .ZN(new_n32729_));
  AOI21_X1   g29462(.A1(new_n32722_), .A2(new_n32729_), .B(new_n8683_), .ZN(new_n32730_));
  NOR2_X1    g29463(.A1(new_n31011_), .A2(new_n2726_), .ZN(new_n32731_));
  OAI21_X1   g29464(.A1(new_n32722_), .A2(new_n32731_), .B(new_n31052_), .ZN(new_n32732_));
  INV_X1     g29465(.I(new_n32731_), .ZN(new_n32733_));
  NAND2_X1   g29466(.A1(new_n30931_), .A2(new_n32719_), .ZN(new_n32734_));
  NOR2_X1    g29467(.A1(new_n32705_), .A2(pi1155), .ZN(new_n32735_));
  INV_X1     g29468(.I(new_n32735_), .ZN(new_n32736_));
  NOR2_X1    g29469(.A1(new_n30698_), .A2(new_n2726_), .ZN(new_n32737_));
  OAI21_X1   g29470(.A1(pi1156), .A2(new_n32736_), .B(new_n32737_), .ZN(new_n32738_));
  NAND4_X1   g29471(.A1(new_n32733_), .A2(pi1156), .A3(pi1157), .A4(new_n32726_), .ZN(new_n32740_));
  NAND2_X1   g29472(.A1(new_n32732_), .A2(new_n32740_), .ZN(new_n32741_));
  AOI21_X1   g29473(.A1(new_n32741_), .A2(new_n32728_), .B(new_n8684_), .ZN(new_n32742_));
  NOR2_X1    g29474(.A1(new_n9258_), .A2(new_n2726_), .ZN(new_n32743_));
  INV_X1     g29475(.I(new_n32743_), .ZN(new_n32744_));
  NOR3_X1    g29476(.A1(new_n32744_), .A2(new_n13778_), .A3(new_n32706_), .ZN(new_n32745_));
  NOR3_X1    g29477(.A1(new_n32743_), .A2(new_n13778_), .A3(new_n32705_), .ZN(new_n32746_));
  OAI21_X1   g29478(.A1(new_n32745_), .A2(new_n32746_), .B(new_n32737_), .ZN(new_n32747_));
  NOR2_X1    g29479(.A1(new_n32719_), .A2(pi0200), .ZN(new_n32748_));
  AOI21_X1   g29480(.A1(new_n32747_), .A2(new_n32748_), .B(new_n13969_), .ZN(new_n32749_));
  NAND2_X1   g29481(.A1(new_n32749_), .A2(pi1157), .ZN(new_n32750_));
  AOI21_X1   g29482(.A1(new_n32750_), .A2(new_n2726_), .B(new_n3098_), .ZN(new_n32751_));
  INV_X1     g29483(.I(new_n32749_), .ZN(new_n32752_));
  NOR3_X1    g29484(.A1(new_n32721_), .A2(new_n32724_), .A3(new_n32736_), .ZN(new_n32753_));
  NOR2_X1    g29485(.A1(new_n30674_), .A2(new_n2726_), .ZN(new_n32754_));
  OAI21_X1   g29486(.A1(pi1156), .A2(new_n32736_), .B(new_n32754_), .ZN(new_n32755_));
  OAI21_X1   g29487(.A1(new_n32738_), .A2(new_n32755_), .B(pi1157), .ZN(new_n32756_));
  NOR2_X1    g29488(.A1(new_n32753_), .A2(new_n32756_), .ZN(new_n32757_));
  XNOR2_X1   g29489(.A1(new_n32757_), .A2(new_n31314_), .ZN(new_n32758_));
  NOR2_X1    g29490(.A1(new_n32758_), .A2(new_n32752_), .ZN(new_n32759_));
  INV_X1     g29491(.I(new_n32754_), .ZN(new_n32760_));
  NAND4_X1   g29492(.A1(new_n30666_), .A2(pi1091), .A3(pi1155), .A4(new_n32705_), .ZN(new_n32761_));
  NAND2_X1   g29493(.A1(new_n30666_), .A2(pi1091), .ZN(new_n32762_));
  NAND3_X1   g29494(.A1(new_n32762_), .A2(pi1155), .A3(new_n32706_), .ZN(new_n32763_));
  AOI21_X1   g29495(.A1(new_n32763_), .A2(new_n32761_), .B(new_n32760_), .ZN(new_n32764_));
  OAI21_X1   g29496(.A1(new_n32764_), .A2(pi1156), .B(new_n30622_), .ZN(new_n32765_));
  OAI21_X1   g29497(.A1(new_n32732_), .A2(new_n32765_), .B(pi0219), .ZN(new_n32766_));
  NOR4_X1    g29498(.A1(new_n32759_), .A2(new_n32742_), .A3(new_n32751_), .A4(new_n32766_), .ZN(new_n32767_));
  XNOR2_X1   g29499(.A1(new_n32767_), .A2(new_n32730_), .ZN(new_n32768_));
  INV_X1     g29500(.I(pi0272), .ZN(new_n32769_));
  INV_X1     g29501(.I(pi0275), .ZN(new_n32770_));
  INV_X1     g29502(.I(pi0283), .ZN(new_n32771_));
  NOR3_X1    g29503(.A1(new_n32769_), .A2(new_n32770_), .A3(new_n32771_), .ZN(new_n32772_));
  NAND2_X1   g29504(.A1(new_n32772_), .A2(pi0268), .ZN(new_n32773_));
  INV_X1     g29505(.I(new_n30621_), .ZN(new_n32774_));
  OAI21_X1   g29506(.A1(pi0211), .A2(new_n13778_), .B(new_n32774_), .ZN(new_n32775_));
  NOR3_X1    g29507(.A1(new_n32775_), .A2(new_n8683_), .A3(new_n14006_), .ZN(new_n32776_));
  XOR2_X1    g29508(.A1(new_n32776_), .A2(new_n30615_), .Z(new_n32777_));
  AOI21_X1   g29509(.A1(new_n32777_), .A2(pi1091), .B(new_n32705_), .ZN(new_n32778_));
  NAND2_X1   g29510(.A1(new_n32550_), .A2(new_n32705_), .ZN(new_n32779_));
  OAI21_X1   g29511(.A1(new_n32775_), .A2(new_n2726_), .B(new_n8683_), .ZN(new_n32780_));
  NAND4_X1   g29512(.A1(new_n32779_), .A2(pi0243), .A3(new_n32538_), .A4(new_n32780_), .ZN(new_n32781_));
  NOR4_X1    g29513(.A1(new_n32548_), .A2(new_n32579_), .A3(new_n32537_), .A4(new_n32564_), .ZN(new_n32783_));
  OAI21_X1   g29514(.A1(new_n8683_), .A2(new_n32783_), .B(new_n32781_), .ZN(new_n32784_));
  NAND2_X1   g29515(.A1(new_n32784_), .A2(po1038), .ZN(new_n32785_));
  NOR2_X1    g29516(.A1(new_n32718_), .A2(new_n7240_), .ZN(new_n32786_));
  XOR2_X1    g29517(.A1(new_n32785_), .A2(new_n32786_), .Z(new_n32787_));
  OAI21_X1   g29518(.A1(new_n32787_), .A2(new_n32778_), .B(new_n32773_), .ZN(new_n32788_));
  NAND3_X1   g29519(.A1(new_n32788_), .A2(pi0211), .A3(new_n7240_), .ZN(new_n32789_));
  AOI21_X1   g29520(.A1(new_n32718_), .A2(new_n32768_), .B(new_n32789_), .ZN(new_n32790_));
  OAI21_X1   g29521(.A1(new_n32717_), .A2(new_n32684_), .B(new_n32790_), .ZN(new_n32791_));
  AOI21_X1   g29522(.A1(new_n32709_), .A2(new_n32713_), .B(new_n32791_), .ZN(new_n32792_));
  OAI21_X1   g29523(.A1(new_n32658_), .A2(new_n32704_), .B(new_n32792_), .ZN(new_n32793_));
  NAND4_X1   g29524(.A1(pi0199), .A2(pi0200), .A3(pi1155), .A4(pi1156), .ZN(new_n32794_));
  INV_X1     g29525(.I(new_n30722_), .ZN(new_n32795_));
  OAI21_X1   g29526(.A1(new_n32795_), .A2(new_n13969_), .B(new_n30680_), .ZN(new_n32796_));
  AOI21_X1   g29527(.A1(new_n32796_), .A2(new_n32794_), .B(new_n8549_), .ZN(new_n32797_));
  OAI21_X1   g29528(.A1(new_n32797_), .A2(pi1157), .B(pi0200), .ZN(new_n32798_));
  NAND2_X1   g29529(.A1(new_n32798_), .A2(pi0230), .ZN(new_n32799_));
  NOR2_X1    g29530(.A1(new_n12655_), .A2(new_n30557_), .ZN(new_n32800_));
  XNOR2_X1   g29531(.A1(new_n32799_), .A2(new_n32800_), .ZN(new_n32801_));
  AOI21_X1   g29532(.A1(new_n32801_), .A2(new_n32777_), .B(pi0230), .ZN(new_n32802_));
  INV_X1     g29533(.I(new_n32778_), .ZN(new_n32803_));
  NAND2_X1   g29534(.A1(new_n32768_), .A2(po1038), .ZN(new_n32804_));
  NOR2_X1    g29535(.A1(new_n7240_), .A2(new_n32773_), .ZN(new_n32805_));
  XNOR2_X1   g29536(.A1(new_n32804_), .A2(new_n32805_), .ZN(new_n32806_));
  NAND2_X1   g29537(.A1(new_n32806_), .A2(new_n32803_), .ZN(new_n32807_));
  AOI21_X1   g29538(.A1(new_n32793_), .A2(new_n32802_), .B(new_n32807_), .ZN(po0400));
  INV_X1     g29539(.I(new_n32178_), .ZN(new_n32809_));
  NOR4_X1    g29540(.A1(new_n32009_), .A2(new_n30597_), .A3(new_n10253_), .A4(new_n30979_), .ZN(new_n32810_));
  NOR3_X1    g29541(.A1(new_n32037_), .A2(new_n30979_), .A3(new_n8740_), .ZN(new_n32811_));
  OAI21_X1   g29542(.A1(new_n32811_), .A2(new_n32810_), .B(new_n32005_), .ZN(new_n32812_));
  OAI21_X1   g29543(.A1(new_n32177_), .A2(new_n32812_), .B(new_n3098_), .ZN(new_n32813_));
  NAND3_X1   g29544(.A1(new_n31378_), .A2(new_n7240_), .A3(new_n32193_), .ZN(new_n32814_));
  AND3_X2    g29545(.A1(new_n32029_), .A2(new_n32026_), .A3(new_n32814_), .Z(new_n32815_));
  AOI21_X1   g29546(.A1(new_n32815_), .A2(new_n32813_), .B(new_n32041_), .ZN(new_n32816_));
  OAI21_X1   g29547(.A1(new_n32816_), .A2(new_n32809_), .B(pi0213), .ZN(new_n32817_));
  XOR2_X1    g29548(.A1(new_n32817_), .A2(new_n31080_), .Z(new_n32818_));
  AOI21_X1   g29549(.A1(new_n32818_), .A2(new_n31395_), .B(new_n30557_), .ZN(new_n32819_));
  INV_X1     g29550(.I(new_n32045_), .ZN(new_n32820_));
  NOR4_X1    g29551(.A1(new_n8684_), .A2(new_n3098_), .A3(new_n3057_), .A4(pi1145), .ZN(new_n32822_));
  OAI21_X1   g29552(.A1(new_n30560_), .A2(new_n32220_), .B(pi0212), .ZN(new_n32823_));
  AOI21_X1   g29553(.A1(new_n8685_), .A2(new_n32822_), .B(new_n32823_), .ZN(new_n32824_));
  NOR2_X1    g29554(.A1(new_n32822_), .A2(new_n8685_), .ZN(new_n32825_));
  XOR2_X1    g29555(.A1(new_n32825_), .A2(new_n8740_), .Z(new_n32826_));
  NAND2_X1   g29556(.A1(new_n31929_), .A2(new_n32826_), .ZN(new_n32827_));
  NOR2_X1    g29557(.A1(new_n31380_), .A2(new_n8683_), .ZN(new_n32828_));
  NAND2_X1   g29558(.A1(new_n32828_), .A2(new_n30619_), .ZN(new_n32829_));
  AOI21_X1   g29559(.A1(new_n31946_), .A2(new_n31940_), .B(new_n32829_), .ZN(new_n32830_));
  AOI21_X1   g29560(.A1(new_n32830_), .A2(new_n32827_), .B(new_n32824_), .ZN(new_n32831_));
  NAND2_X1   g29561(.A1(new_n8739_), .A2(pi0214), .ZN(new_n32832_));
  NAND2_X1   g29562(.A1(new_n31956_), .A2(new_n32832_), .ZN(new_n32833_));
  AOI21_X1   g29563(.A1(new_n32833_), .A2(new_n32822_), .B(pi0219), .ZN(new_n32834_));
  NAND2_X1   g29564(.A1(new_n31920_), .A2(new_n32824_), .ZN(new_n32835_));
  NOR2_X1    g29565(.A1(po1038), .A2(pi1147), .ZN(new_n32836_));
  INV_X1     g29566(.I(new_n32836_), .ZN(new_n32837_));
  OAI21_X1   g29567(.A1(new_n32834_), .A2(new_n32835_), .B(new_n32837_), .ZN(new_n32838_));
  NAND2_X1   g29568(.A1(new_n31919_), .A2(pi0299), .ZN(new_n32839_));
  XOR2_X1    g29569(.A1(new_n32839_), .A2(new_n31523_), .Z(new_n32840_));
  NAND2_X1   g29570(.A1(new_n32840_), .A2(pi1143), .ZN(new_n32841_));
  OAI21_X1   g29571(.A1(new_n31907_), .A2(new_n8684_), .B(new_n31238_), .ZN(new_n32842_));
  NOR4_X1    g29572(.A1(new_n31959_), .A2(new_n31080_), .A3(new_n32842_), .A4(new_n32019_), .ZN(new_n32843_));
  NAND4_X1   g29573(.A1(new_n32838_), .A2(new_n31393_), .A3(new_n32841_), .A4(new_n32843_), .ZN(new_n32844_));
  OAI21_X1   g29574(.A1(new_n32844_), .A2(new_n32831_), .B(new_n28529_), .ZN(new_n32845_));
  NAND4_X1   g29575(.A1(new_n32820_), .A2(new_n32845_), .A3(pi0230), .A4(pi0244), .ZN(new_n32846_));
  XNOR2_X1   g29576(.A1(new_n32846_), .A2(new_n32819_), .ZN(po0401));
  NOR2_X1    g29577(.A1(new_n31955_), .A2(new_n3350_), .ZN(new_n32848_));
  INV_X1     g29578(.I(new_n32848_), .ZN(new_n32849_));
  NOR2_X1    g29579(.A1(new_n32849_), .A2(new_n31951_), .ZN(new_n32850_));
  AOI21_X1   g29580(.A1(pi1147), .A2(new_n32406_), .B(new_n32850_), .ZN(new_n32851_));
  NOR2_X1    g29581(.A1(new_n30588_), .A2(new_n8685_), .ZN(new_n32852_));
  NAND2_X1   g29582(.A1(new_n32475_), .A2(new_n3098_), .ZN(new_n32853_));
  INV_X1     g29583(.I(new_n32853_), .ZN(new_n32854_));
  NOR2_X1    g29584(.A1(new_n32473_), .A2(new_n8684_), .ZN(new_n32855_));
  AOI21_X1   g29585(.A1(new_n8684_), .A2(new_n32854_), .B(new_n32855_), .ZN(new_n32856_));
  NOR3_X1    g29586(.A1(new_n32856_), .A2(new_n8685_), .A3(new_n32482_), .ZN(new_n32857_));
  XOR2_X1    g29587(.A1(new_n32857_), .A2(new_n32852_), .Z(new_n32858_));
  NAND2_X1   g29588(.A1(new_n32473_), .A2(new_n30594_), .ZN(new_n32859_));
  AOI21_X1   g29589(.A1(new_n32859_), .A2(new_n32483_), .B(po1038), .ZN(new_n32860_));
  NAND2_X1   g29590(.A1(new_n32480_), .A2(new_n32482_), .ZN(new_n32861_));
  AND3_X2    g29591(.A1(new_n32860_), .A2(new_n30588_), .A3(new_n32861_), .Z(new_n32862_));
  OAI21_X1   g29592(.A1(pi0212), .A2(new_n32862_), .B(new_n32858_), .ZN(new_n32863_));
  OAI21_X1   g29593(.A1(new_n32854_), .A2(pi0211), .B(new_n32478_), .ZN(new_n32864_));
  NAND2_X1   g29594(.A1(new_n32864_), .A2(new_n32479_), .ZN(new_n32865_));
  NOR2_X1    g29595(.A1(new_n32848_), .A2(pi1147), .ZN(new_n32866_));
  INV_X1     g29596(.I(new_n32866_), .ZN(new_n32867_));
  NOR2_X1    g29597(.A1(new_n32867_), .A2(new_n31757_), .ZN(new_n32868_));
  OAI21_X1   g29598(.A1(new_n32868_), .A2(new_n8689_), .B(new_n31722_), .ZN(new_n32869_));
  INV_X1     g29599(.I(new_n32869_), .ZN(new_n32870_));
  AOI22_X1   g29600(.A1(new_n32865_), .A2(new_n8683_), .B1(new_n32860_), .B2(new_n32870_), .ZN(new_n32871_));
  NOR2_X1    g29601(.A1(new_n32009_), .A2(new_n8685_), .ZN(new_n32872_));
  AOI21_X1   g29602(.A1(new_n32872_), .A2(pi0212), .B(pi0299), .ZN(new_n32873_));
  NOR2_X1    g29603(.A1(new_n32476_), .A2(new_n32873_), .ZN(new_n32874_));
  OAI21_X1   g29604(.A1(pi0214), .A2(new_n32864_), .B(new_n32874_), .ZN(new_n32875_));
  OAI21_X1   g29605(.A1(new_n32875_), .A2(new_n32871_), .B(new_n31953_), .ZN(new_n32876_));
  AOI21_X1   g29606(.A1(new_n32482_), .A2(new_n8739_), .B(pi0219), .ZN(new_n32877_));
  AOI21_X1   g29607(.A1(new_n32874_), .A2(new_n32877_), .B(new_n32478_), .ZN(new_n32878_));
  NOR2_X1    g29608(.A1(new_n32867_), .A2(new_n31953_), .ZN(new_n32879_));
  INV_X1     g29609(.I(new_n32850_), .ZN(new_n32880_));
  NOR2_X1    g29610(.A1(new_n32880_), .A2(new_n8685_), .ZN(new_n32881_));
  OAI21_X1   g29611(.A1(new_n32860_), .A2(new_n32879_), .B(new_n32881_), .ZN(new_n32882_));
  NOR2_X1    g29612(.A1(new_n32856_), .A2(new_n8685_), .ZN(new_n32883_));
  AOI21_X1   g29613(.A1(new_n8685_), .A2(new_n32854_), .B(new_n32883_), .ZN(new_n32884_));
  AOI21_X1   g29614(.A1(new_n32853_), .A2(new_n32479_), .B(pi0219), .ZN(new_n32885_));
  AOI21_X1   g29615(.A1(new_n32860_), .A2(new_n32885_), .B(pi0212), .ZN(new_n32886_));
  NOR4_X1    g29616(.A1(new_n32884_), .A2(new_n32878_), .A3(new_n32882_), .A4(new_n32886_), .ZN(new_n32887_));
  NAND2_X1   g29617(.A1(new_n32887_), .A2(new_n32876_), .ZN(new_n32888_));
  NAND2_X1   g29618(.A1(new_n32863_), .A2(new_n32888_), .ZN(new_n32889_));
  AOI21_X1   g29619(.A1(new_n32889_), .A2(new_n32851_), .B(new_n28529_), .ZN(new_n32890_));
  XOR2_X1    g29620(.A1(new_n32890_), .A2(new_n31079_), .Z(new_n32891_));
  AOI21_X1   g29621(.A1(new_n32891_), .A2(new_n32501_), .B(new_n30557_), .ZN(new_n32892_));
  INV_X1     g29622(.I(new_n32872_), .ZN(new_n32893_));
  XNOR2_X1   g29623(.A1(pi0200), .A2(pi1146), .ZN(new_n32894_));
  NOR2_X1    g29624(.A1(new_n32894_), .A2(new_n31030_), .ZN(new_n32895_));
  AOI21_X1   g29625(.A1(new_n32895_), .A2(pi0208), .B(pi0207), .ZN(new_n32896_));
  INV_X1     g29626(.I(new_n32895_), .ZN(new_n32897_));
  AOI21_X1   g29627(.A1(new_n32897_), .A2(new_n8546_), .B(new_n30735_), .ZN(new_n32898_));
  INV_X1     g29628(.I(new_n32898_), .ZN(new_n32899_));
  NOR2_X1    g29629(.A1(new_n32899_), .A2(new_n32896_), .ZN(new_n32900_));
  AOI22_X1   g29630(.A1(new_n32895_), .A2(new_n30666_), .B1(pi0207), .B2(pi1146), .ZN(new_n32901_));
  NAND2_X1   g29631(.A1(new_n32901_), .A2(pi0208), .ZN(new_n32902_));
  NOR2_X1    g29632(.A1(new_n31420_), .A2(pi1146), .ZN(new_n32903_));
  NOR3_X1    g29633(.A1(new_n31908_), .A2(new_n8546_), .A3(new_n32903_), .ZN(new_n32905_));
  XNOR2_X1   g29634(.A1(new_n32902_), .A2(new_n32905_), .ZN(new_n32906_));
  NAND2_X1   g29635(.A1(new_n32906_), .A2(new_n31912_), .ZN(new_n32907_));
  INV_X1     g29636(.I(new_n32907_), .ZN(new_n32908_));
  AOI21_X1   g29637(.A1(new_n3098_), .A2(new_n32897_), .B(new_n32908_), .ZN(new_n32909_));
  NOR2_X1    g29638(.A1(new_n32909_), .A2(pi0299), .ZN(new_n32910_));
  INV_X1     g29639(.I(new_n32910_), .ZN(new_n32911_));
  NOR2_X1    g29640(.A1(new_n32908_), .A2(pi0299), .ZN(new_n32912_));
  INV_X1     g29641(.I(new_n32912_), .ZN(new_n32913_));
  NOR3_X1    g29642(.A1(new_n32911_), .A2(new_n8684_), .A3(new_n32913_), .ZN(new_n32914_));
  NOR2_X1    g29643(.A1(new_n8684_), .A2(new_n3098_), .ZN(new_n32915_));
  OAI21_X1   g29644(.A1(new_n32914_), .A2(new_n32915_), .B(new_n32900_), .ZN(new_n32916_));
  OAI21_X1   g29645(.A1(new_n32916_), .A2(pi0214), .B(pi0212), .ZN(new_n32917_));
  NAND2_X1   g29646(.A1(new_n32916_), .A2(new_n8739_), .ZN(new_n32918_));
  NOR2_X1    g29647(.A1(new_n32913_), .A2(new_n8685_), .ZN(new_n32919_));
  AOI21_X1   g29648(.A1(new_n32918_), .A2(new_n32919_), .B(pi0219), .ZN(new_n32920_));
  INV_X1     g29649(.I(new_n32920_), .ZN(new_n32921_));
  OAI21_X1   g29650(.A1(new_n32921_), .A2(new_n32917_), .B(new_n32893_), .ZN(new_n32922_));
  NOR2_X1    g29651(.A1(new_n31908_), .A2(new_n32903_), .ZN(new_n32923_));
  INV_X1     g29652(.I(new_n32923_), .ZN(new_n32924_));
  NOR2_X1    g29653(.A1(new_n32924_), .A2(new_n8545_), .ZN(new_n32925_));
  AOI21_X1   g29654(.A1(pi1146), .A2(new_n30735_), .B(new_n30652_), .ZN(new_n32926_));
  XOR2_X1    g29655(.A1(new_n32923_), .A2(new_n8547_), .Z(new_n32927_));
  NAND2_X1   g29656(.A1(new_n32927_), .A2(new_n32926_), .ZN(new_n32928_));
  NOR2_X1    g29657(.A1(new_n32928_), .A2(new_n32925_), .ZN(new_n32929_));
  NAND2_X1   g29658(.A1(new_n32928_), .A2(new_n32925_), .ZN(new_n32930_));
  INV_X1     g29659(.I(new_n32930_), .ZN(new_n32931_));
  NOR2_X1    g29660(.A1(new_n32931_), .A2(new_n32929_), .ZN(new_n32932_));
  AOI21_X1   g29661(.A1(new_n32932_), .A2(pi0211), .B(new_n30586_), .ZN(new_n32933_));
  INV_X1     g29662(.I(new_n32926_), .ZN(new_n32934_));
  AOI21_X1   g29663(.A1(new_n32934_), .A2(new_n31913_), .B(pi0207), .ZN(new_n32935_));
  NOR2_X1    g29664(.A1(new_n32935_), .A2(new_n32924_), .ZN(new_n32936_));
  INV_X1     g29665(.I(new_n32936_), .ZN(new_n32937_));
  AOI21_X1   g29666(.A1(new_n31912_), .A2(pi0208), .B(pi0207), .ZN(new_n32938_));
  NOR2_X1    g29667(.A1(new_n32934_), .A2(new_n32938_), .ZN(new_n32939_));
  NAND2_X1   g29668(.A1(new_n32932_), .A2(new_n31991_), .ZN(new_n32940_));
  NAND2_X1   g29669(.A1(new_n32940_), .A2(pi0212), .ZN(new_n32941_));
  NOR2_X1    g29670(.A1(new_n32941_), .A2(new_n7240_), .ZN(new_n32942_));
  AOI21_X1   g29671(.A1(new_n32937_), .A2(new_n32939_), .B(new_n32942_), .ZN(new_n32943_));
  NOR2_X1    g29672(.A1(new_n8686_), .A2(new_n3098_), .ZN(new_n32944_));
  NOR2_X1    g29673(.A1(new_n32907_), .A2(new_n32213_), .ZN(new_n32945_));
  XOR2_X1    g29674(.A1(new_n32945_), .A2(new_n32944_), .Z(new_n32946_));
  INV_X1     g29675(.I(new_n32900_), .ZN(new_n32947_));
  AOI21_X1   g29676(.A1(new_n32947_), .A2(pi0211), .B(new_n30586_), .ZN(new_n32948_));
  OAI21_X1   g29677(.A1(new_n32947_), .A2(new_n31238_), .B(pi0219), .ZN(new_n32949_));
  AOI21_X1   g29678(.A1(po1038), .A2(new_n32949_), .B(new_n32948_), .ZN(new_n32950_));
  NAND2_X1   g29679(.A1(new_n32909_), .A2(pi0219), .ZN(new_n32951_));
  OAI21_X1   g29680(.A1(new_n32951_), .A2(new_n32950_), .B(new_n32901_), .ZN(new_n32952_));
  AOI21_X1   g29681(.A1(new_n32952_), .A2(new_n32946_), .B(new_n32867_), .ZN(new_n32953_));
  NAND2_X1   g29682(.A1(new_n32851_), .A2(new_n31953_), .ZN(new_n32954_));
  OAI22_X1   g29683(.A1(new_n32943_), .A2(new_n32933_), .B1(new_n32953_), .B2(new_n32954_), .ZN(new_n32955_));
  NAND2_X1   g29684(.A1(new_n32937_), .A2(new_n32939_), .ZN(new_n32956_));
  NOR2_X1    g29685(.A1(new_n32956_), .A2(pi0299), .ZN(new_n32957_));
  NOR2_X1    g29686(.A1(new_n32957_), .A2(new_n8685_), .ZN(new_n32958_));
  NOR2_X1    g29687(.A1(new_n30738_), .A2(new_n32903_), .ZN(new_n32959_));
  NAND2_X1   g29688(.A1(new_n32927_), .A2(new_n32959_), .ZN(new_n32960_));
  XOR2_X1    g29689(.A1(new_n32960_), .A2(new_n32925_), .Z(new_n32961_));
  INV_X1     g29690(.I(new_n32961_), .ZN(new_n32962_));
  NOR2_X1    g29691(.A1(new_n32959_), .A2(new_n8546_), .ZN(new_n32963_));
  NAND2_X1   g29692(.A1(new_n32925_), .A2(pi0208), .ZN(new_n32964_));
  XOR2_X1    g29693(.A1(new_n32964_), .A2(new_n32963_), .Z(new_n32965_));
  NOR2_X1    g29694(.A1(new_n32937_), .A2(pi0299), .ZN(new_n32966_));
  NOR2_X1    g29695(.A1(new_n32965_), .A2(new_n32966_), .ZN(new_n32967_));
  INV_X1     g29696(.I(new_n32967_), .ZN(new_n32968_));
  NOR2_X1    g29697(.A1(new_n32968_), .A2(pi0299), .ZN(new_n32969_));
  INV_X1     g29698(.I(new_n32969_), .ZN(new_n32970_));
  AOI21_X1   g29699(.A1(new_n32970_), .A2(new_n8684_), .B(new_n32962_), .ZN(new_n32971_));
  INV_X1     g29700(.I(new_n32971_), .ZN(new_n32972_));
  AOI21_X1   g29701(.A1(new_n32972_), .A2(new_n32958_), .B(new_n8739_), .ZN(new_n32973_));
  NAND2_X1   g29702(.A1(new_n32932_), .A2(new_n31523_), .ZN(new_n32974_));
  INV_X1     g29703(.I(new_n32932_), .ZN(new_n32975_));
  AOI21_X1   g29704(.A1(new_n32975_), .A2(new_n8685_), .B(pi0212), .ZN(new_n32976_));
  AOI22_X1   g29705(.A1(new_n32973_), .A2(new_n32976_), .B1(pi0214), .B2(new_n32974_), .ZN(new_n32977_));
  OAI21_X1   g29706(.A1(new_n31594_), .A2(pi1146), .B(new_n32214_), .ZN(new_n32978_));
  NAND4_X1   g29707(.A1(new_n32977_), .A2(new_n8683_), .A3(new_n32955_), .A4(new_n32978_), .ZN(new_n32979_));
  AOI21_X1   g29708(.A1(new_n32961_), .A2(new_n8685_), .B(pi0212), .ZN(new_n32980_));
  AOI21_X1   g29709(.A1(new_n32970_), .A2(new_n32980_), .B(pi0219), .ZN(new_n32981_));
  NOR2_X1    g29710(.A1(new_n32961_), .A2(new_n30594_), .ZN(new_n32982_));
  NOR2_X1    g29711(.A1(new_n32982_), .A2(new_n8683_), .ZN(new_n32983_));
  AOI21_X1   g29712(.A1(new_n32983_), .A2(po1038), .B(new_n30594_), .ZN(new_n32984_));
  NOR4_X1    g29713(.A1(new_n32984_), .A2(new_n31912_), .A3(new_n32880_), .A4(new_n32968_), .ZN(new_n32985_));
  NOR2_X1    g29714(.A1(new_n32969_), .A2(pi0212), .ZN(new_n32986_));
  NOR4_X1    g29715(.A1(new_n32986_), .A2(new_n30718_), .A3(new_n31912_), .A4(new_n32968_), .ZN(new_n32987_));
  OAI21_X1   g29716(.A1(new_n32985_), .A2(new_n32981_), .B(new_n32987_), .ZN(new_n32988_));
  NAND3_X1   g29717(.A1(new_n32979_), .A2(new_n31953_), .A3(new_n32988_), .ZN(new_n32989_));
  AOI21_X1   g29718(.A1(new_n32912_), .A2(new_n30604_), .B(new_n8683_), .ZN(new_n32990_));
  INV_X1     g29719(.I(new_n32990_), .ZN(new_n32991_));
  AOI21_X1   g29720(.A1(new_n30594_), .A2(new_n32907_), .B(new_n32991_), .ZN(new_n32992_));
  NOR3_X1    g29721(.A1(new_n32992_), .A2(po1038), .A3(new_n32870_), .ZN(new_n32993_));
  NOR3_X1    g29722(.A1(new_n32993_), .A2(new_n28529_), .A3(new_n32913_), .ZN(new_n32994_));
  NAND3_X1   g29723(.A1(new_n32989_), .A2(new_n32922_), .A3(new_n32994_), .ZN(new_n32995_));
  AOI21_X1   g29724(.A1(new_n32908_), .A2(new_n3098_), .B(new_n30604_), .ZN(new_n32996_));
  INV_X1     g29725(.I(new_n32996_), .ZN(new_n32997_));
  OAI21_X1   g29726(.A1(new_n32991_), .A2(new_n32837_), .B(new_n32997_), .ZN(new_n32998_));
  AOI21_X1   g29727(.A1(new_n32912_), .A2(pi0212), .B(pi0214), .ZN(new_n32999_));
  OAI21_X1   g29728(.A1(new_n32999_), .A2(new_n32004_), .B(new_n8683_), .ZN(new_n33000_));
  AOI21_X1   g29729(.A1(new_n32998_), .A2(new_n30869_), .B(new_n33000_), .ZN(new_n33001_));
  NAND2_X1   g29730(.A1(new_n32967_), .A2(new_n30879_), .ZN(new_n33002_));
  NAND2_X1   g29731(.A1(new_n32983_), .A2(new_n31954_), .ZN(new_n33003_));
  AOI21_X1   g29732(.A1(new_n33003_), .A2(new_n30604_), .B(new_n33002_), .ZN(new_n33004_));
  NOR3_X1    g29733(.A1(new_n32980_), .A2(pi0214), .A3(new_n32967_), .ZN(new_n33005_));
  OAI21_X1   g29734(.A1(new_n33005_), .A2(new_n32004_), .B(new_n8683_), .ZN(new_n33006_));
  AND2_X2    g29735(.A1(new_n32486_), .A2(pi0299), .Z(new_n33007_));
  OAI21_X1   g29736(.A1(new_n32912_), .A2(new_n33007_), .B(pi0212), .ZN(new_n33008_));
  OAI21_X1   g29737(.A1(new_n32968_), .A2(new_n33007_), .B(pi0212), .ZN(new_n33009_));
  NOR4_X1    g29738(.A1(new_n33009_), .A2(new_n33008_), .A3(new_n31953_), .A4(new_n32492_), .ZN(new_n33010_));
  OAI21_X1   g29739(.A1(new_n33004_), .A2(new_n33006_), .B(new_n33010_), .ZN(new_n33011_));
  OAI21_X1   g29740(.A1(new_n33011_), .A2(new_n33001_), .B(new_n28529_), .ZN(new_n33012_));
  NAND2_X1   g29741(.A1(new_n32911_), .A2(new_n8685_), .ZN(new_n33013_));
  NOR3_X1    g29742(.A1(new_n32913_), .A2(new_n8739_), .A3(new_n32004_), .ZN(new_n33014_));
  AOI21_X1   g29743(.A1(new_n33013_), .A2(new_n33014_), .B(new_n32900_), .ZN(new_n33015_));
  OAI21_X1   g29744(.A1(new_n33008_), .A2(new_n8683_), .B(new_n3098_), .ZN(new_n33016_));
  INV_X1     g29745(.I(new_n32957_), .ZN(new_n33017_));
  NAND2_X1   g29746(.A1(new_n32492_), .A2(new_n31953_), .ZN(new_n33018_));
  NAND4_X1   g29747(.A1(new_n33018_), .A2(pi0214), .A3(new_n31954_), .A4(new_n32895_), .ZN(new_n33019_));
  NOR3_X1    g29748(.A1(new_n33009_), .A2(new_n33017_), .A3(new_n33019_), .ZN(new_n33020_));
  NAND2_X1   g29749(.A1(new_n33020_), .A2(new_n33016_), .ZN(new_n33021_));
  NOR2_X1    g29750(.A1(new_n32968_), .A2(new_n32005_), .ZN(new_n33022_));
  NAND2_X1   g29751(.A1(new_n32958_), .A2(pi0212), .ZN(new_n33023_));
  OAI21_X1   g29752(.A1(new_n33022_), .A2(new_n33023_), .B(new_n32932_), .ZN(new_n33024_));
  AOI21_X1   g29753(.A1(new_n33024_), .A2(pi0214), .B(pi0219), .ZN(new_n33025_));
  NAND2_X1   g29754(.A1(new_n32948_), .A2(pi0211), .ZN(new_n33026_));
  NAND2_X1   g29755(.A1(new_n32911_), .A2(new_n33026_), .ZN(new_n33027_));
  AOI21_X1   g29756(.A1(new_n33027_), .A2(new_n30869_), .B(new_n32949_), .ZN(new_n33028_));
  OAI21_X1   g29757(.A1(new_n32932_), .A2(new_n30586_), .B(pi0211), .ZN(new_n33029_));
  AOI21_X1   g29758(.A1(new_n33029_), .A2(new_n33017_), .B(new_n33002_), .ZN(new_n33030_));
  OAI22_X1   g29759(.A1(new_n33028_), .A2(new_n32836_), .B1(new_n32941_), .B2(new_n33030_), .ZN(new_n33031_));
  NOR4_X1    g29760(.A1(new_n33031_), .A2(new_n33015_), .A3(new_n33021_), .A4(new_n33025_), .ZN(new_n33032_));
  AOI21_X1   g29761(.A1(new_n33032_), .A2(new_n33012_), .B(pi0209), .ZN(new_n33033_));
  NOR4_X1    g29762(.A1(new_n32995_), .A2(new_n30557_), .A3(new_n4955_), .A4(new_n33033_), .ZN(new_n33034_));
  XOR2_X1    g29763(.A1(new_n32892_), .A2(new_n33034_), .Z(po0402));
  AOI21_X1   g29764(.A1(new_n32048_), .A2(new_n32061_), .B(new_n32079_), .ZN(new_n33036_));
  AOI21_X1   g29765(.A1(new_n33036_), .A2(pi0219), .B(new_n32341_), .ZN(new_n33037_));
  NAND2_X1   g29766(.A1(new_n32063_), .A2(pi1146), .ZN(new_n33038_));
  NAND2_X1   g29767(.A1(new_n33038_), .A2(new_n32242_), .ZN(new_n33039_));
  INV_X1     g29768(.I(new_n32078_), .ZN(new_n33040_));
  OR3_X2     g29769(.A1(new_n33036_), .A2(pi0219), .A3(pi1146), .Z(new_n33041_));
  AOI22_X1   g29770(.A1(new_n33041_), .A2(new_n32063_), .B1(new_n31712_), .B2(new_n32022_), .ZN(new_n33042_));
  NAND2_X1   g29771(.A1(new_n32851_), .A2(new_n32063_), .ZN(new_n33043_));
  AOI21_X1   g29772(.A1(new_n33040_), .A2(new_n33042_), .B(new_n33043_), .ZN(new_n33044_));
  AOI21_X1   g29773(.A1(new_n33044_), .A2(new_n33039_), .B(pi1148), .ZN(new_n33045_));
  AOI21_X1   g29774(.A1(new_n8685_), .A2(new_n32120_), .B(new_n32275_), .ZN(new_n33047_));
  INV_X1     g29775(.I(new_n33047_), .ZN(new_n33048_));
  NOR3_X1    g29776(.A1(new_n32273_), .A2(new_n8685_), .A3(new_n32114_), .ZN(new_n33049_));
  AOI21_X1   g29777(.A1(pi0219), .A2(new_n32008_), .B(new_n32049_), .ZN(new_n33050_));
  INV_X1     g29778(.I(new_n33050_), .ZN(new_n33051_));
  AOI21_X1   g29779(.A1(new_n32231_), .A2(new_n33051_), .B(new_n33049_), .ZN(new_n33052_));
  NOR4_X1    g29780(.A1(new_n31643_), .A2(new_n3098_), .A3(new_n9209_), .A4(new_n31450_), .ZN(new_n33053_));
  NOR3_X1    g29781(.A1(new_n32111_), .A2(new_n31642_), .A3(new_n3098_), .ZN(new_n33054_));
  NOR2_X1    g29782(.A1(new_n33053_), .A2(new_n33054_), .ZN(new_n33055_));
  NOR4_X1    g29783(.A1(new_n33048_), .A2(new_n33052_), .A3(new_n3350_), .A4(new_n33055_), .ZN(new_n33056_));
  OR2_X2     g29784(.A1(new_n33056_), .A2(new_n32851_), .Z(new_n33057_));
  NOR2_X1    g29785(.A1(new_n32276_), .A2(pi0219), .ZN(new_n33058_));
  NOR3_X1    g29786(.A1(new_n33058_), .A2(new_n32117_), .A3(new_n32369_), .ZN(new_n33059_));
  INV_X1     g29787(.I(new_n33059_), .ZN(new_n33060_));
  NAND2_X1   g29788(.A1(new_n33060_), .A2(new_n32228_), .ZN(new_n33061_));
  OAI22_X1   g29789(.A1(new_n33061_), .A2(new_n32867_), .B1(po1038), .B2(new_n32123_), .ZN(new_n33062_));
  NAND4_X1   g29790(.A1(new_n33062_), .A2(pi1150), .A3(new_n33056_), .A4(new_n33057_), .ZN(new_n33063_));
  OAI21_X1   g29791(.A1(new_n33045_), .A2(new_n33063_), .B(pi1149), .ZN(new_n33064_));
  NAND2_X1   g29792(.A1(new_n32851_), .A2(new_n32866_), .ZN(new_n33065_));
  NOR2_X1    g29793(.A1(new_n32204_), .A2(new_n8683_), .ZN(new_n33066_));
  OAI21_X1   g29794(.A1(new_n33050_), .A2(new_n32307_), .B(new_n33066_), .ZN(new_n33067_));
  NOR2_X1    g29795(.A1(new_n33067_), .A2(new_n33051_), .ZN(new_n33068_));
  AOI21_X1   g29796(.A1(pi1150), .A2(new_n32088_), .B(new_n33068_), .ZN(new_n33069_));
  AOI21_X1   g29797(.A1(new_n33065_), .A2(new_n33069_), .B(new_n31953_), .ZN(new_n33070_));
  NAND2_X1   g29798(.A1(new_n32170_), .A2(new_n32411_), .ZN(new_n33071_));
  NOR2_X1    g29799(.A1(new_n31695_), .A2(new_n8739_), .ZN(new_n33072_));
  INV_X1     g29800(.I(new_n33072_), .ZN(new_n33073_));
  AOI21_X1   g29801(.A1(new_n32344_), .A2(new_n8683_), .B(new_n33073_), .ZN(new_n33074_));
  INV_X1     g29802(.I(new_n33074_), .ZN(new_n33075_));
  NOR2_X1    g29803(.A1(new_n32880_), .A2(new_n33075_), .ZN(new_n33076_));
  AOI21_X1   g29804(.A1(new_n33076_), .A2(new_n33071_), .B(new_n32165_), .ZN(new_n33077_));
  OAI21_X1   g29805(.A1(new_n33077_), .A2(new_n33051_), .B(new_n32242_), .ZN(new_n33078_));
  NAND2_X1   g29806(.A1(new_n32097_), .A2(new_n33050_), .ZN(new_n33079_));
  OAI21_X1   g29807(.A1(new_n32168_), .A2(pi0214), .B(new_n31696_), .ZN(new_n33080_));
  NAND2_X1   g29808(.A1(new_n33080_), .A2(new_n8739_), .ZN(new_n33081_));
  NAND3_X1   g29809(.A1(new_n32095_), .A2(new_n32165_), .A3(new_n33081_), .ZN(new_n33082_));
  AOI21_X1   g29810(.A1(new_n33079_), .A2(new_n33082_), .B(new_n32869_), .ZN(new_n33083_));
  NAND2_X1   g29811(.A1(new_n32134_), .A2(pi0219), .ZN(new_n33084_));
  NAND2_X1   g29812(.A1(new_n33084_), .A2(new_n32242_), .ZN(new_n33085_));
  AOI21_X1   g29813(.A1(new_n33078_), .A2(new_n33083_), .B(new_n33085_), .ZN(new_n33086_));
  NOR2_X1    g29814(.A1(new_n32135_), .A2(new_n32132_), .ZN(new_n33087_));
  NOR2_X1    g29815(.A1(new_n32870_), .A2(new_n32850_), .ZN(new_n33088_));
  NOR2_X1    g29816(.A1(new_n32299_), .A2(new_n31091_), .ZN(new_n33089_));
  NOR3_X1    g29817(.A1(new_n33089_), .A2(new_n32134_), .A3(new_n32198_), .ZN(new_n33090_));
  AOI21_X1   g29818(.A1(new_n33088_), .A2(new_n33090_), .B(new_n33087_), .ZN(new_n33091_));
  AOI21_X1   g29819(.A1(new_n31003_), .A2(new_n31793_), .B(new_n8684_), .ZN(new_n33092_));
  AOI21_X1   g29820(.A1(new_n32978_), .A2(new_n33092_), .B(new_n32851_), .ZN(new_n33093_));
  NAND4_X1   g29821(.A1(new_n33050_), .A2(pi1148), .A3(pi1150), .A4(new_n31603_), .ZN(new_n33094_));
  NOR4_X1    g29822(.A1(new_n33086_), .A2(new_n33091_), .A3(new_n33093_), .A4(new_n33094_), .ZN(new_n33095_));
  XOR2_X1    g29823(.A1(new_n33095_), .A2(new_n33070_), .Z(new_n33096_));
  NOR2_X1    g29824(.A1(new_n32136_), .A2(new_n31800_), .ZN(new_n33097_));
  NOR2_X1    g29825(.A1(new_n32139_), .A2(pi0219), .ZN(new_n33098_));
  NAND2_X1   g29826(.A1(new_n33098_), .A2(new_n33097_), .ZN(new_n33099_));
  AOI21_X1   g29827(.A1(new_n33099_), .A2(new_n32893_), .B(new_n31664_), .ZN(new_n33100_));
  AOI21_X1   g29828(.A1(new_n32870_), .A2(new_n33100_), .B(new_n32148_), .ZN(new_n33101_));
  NAND3_X1   g29829(.A1(new_n33088_), .A2(new_n32137_), .A3(new_n32334_), .ZN(new_n33102_));
  OAI21_X1   g29830(.A1(new_n33102_), .A2(new_n33101_), .B(new_n32135_), .ZN(new_n33103_));
  AOI21_X1   g29831(.A1(new_n32153_), .A2(pi0219), .B(po1038), .ZN(new_n33104_));
  NAND2_X1   g29832(.A1(new_n32222_), .A2(new_n8683_), .ZN(new_n33105_));
  NAND4_X1   g29833(.A1(new_n33105_), .A2(new_n32216_), .A3(pi0214), .A4(new_n32223_), .ZN(new_n33106_));
  NAND2_X1   g29834(.A1(new_n33106_), .A2(new_n33104_), .ZN(new_n33107_));
  NOR2_X1    g29835(.A1(new_n32850_), .A2(pi1150), .ZN(new_n33108_));
  NAND2_X1   g29836(.A1(new_n32050_), .A2(pi1146), .ZN(new_n33109_));
  AOI21_X1   g29837(.A1(new_n33108_), .A2(new_n33107_), .B(new_n33109_), .ZN(new_n33110_));
  NOR3_X1    g29838(.A1(new_n32870_), .A2(new_n32224_), .A3(new_n33110_), .ZN(new_n33111_));
  OAI21_X1   g29839(.A1(new_n33111_), .A2(new_n33067_), .B(new_n31953_), .ZN(new_n33112_));
  NAND2_X1   g29840(.A1(pi1149), .A2(pi1150), .ZN(new_n33113_));
  NOR2_X1    g29841(.A1(new_n33051_), .A2(new_n33113_), .ZN(new_n33114_));
  NAND4_X1   g29842(.A1(new_n33096_), .A2(new_n33103_), .A3(new_n33112_), .A4(new_n33114_), .ZN(new_n33115_));
  XOR2_X1    g29843(.A1(new_n33115_), .A2(new_n33064_), .Z(new_n33116_));
  OAI21_X1   g29844(.A1(new_n32109_), .A2(new_n31973_), .B(pi1150), .ZN(new_n33117_));
  XOR2_X1    g29845(.A1(new_n33117_), .A2(new_n33113_), .Z(new_n33118_));
  AOI21_X1   g29846(.A1(new_n33118_), .A2(new_n32151_), .B(new_n31953_), .ZN(new_n33119_));
  NOR2_X1    g29847(.A1(pi1149), .A2(pi1150), .ZN(new_n33120_));
  NOR2_X1    g29848(.A1(new_n32156_), .A2(new_n31941_), .ZN(new_n33121_));
  XOR2_X1    g29849(.A1(new_n33121_), .A2(new_n33113_), .Z(new_n33122_));
  NAND2_X1   g29850(.A1(new_n32092_), .A2(pi1148), .ZN(new_n33123_));
  NOR4_X1    g29851(.A1(new_n33122_), .A2(new_n32055_), .A3(new_n33120_), .A4(new_n33123_), .ZN(new_n33124_));
  XNOR2_X1   g29852(.A1(new_n33119_), .A2(new_n33124_), .ZN(new_n33125_));
  NAND2_X1   g29853(.A1(new_n33125_), .A2(pi0209), .ZN(new_n33126_));
  XOR2_X1    g29854(.A1(new_n33126_), .A2(new_n31080_), .Z(new_n33127_));
  AOI21_X1   g29855(.A1(new_n33127_), .A2(new_n33116_), .B(new_n30557_), .ZN(new_n33128_));
  NAND2_X1   g29856(.A1(new_n32909_), .A2(new_n31940_), .ZN(new_n33129_));
  NAND2_X1   g29857(.A1(new_n33129_), .A2(new_n12654_), .ZN(new_n33130_));
  NOR2_X1    g29858(.A1(new_n31980_), .A2(new_n32242_), .ZN(new_n33131_));
  AOI21_X1   g29859(.A1(new_n33130_), .A2(new_n33131_), .B(new_n31941_), .ZN(new_n33132_));
  NOR2_X1    g29860(.A1(new_n32910_), .A2(new_n8685_), .ZN(new_n33133_));
  NOR2_X1    g29861(.A1(new_n33133_), .A2(new_n30718_), .ZN(new_n33134_));
  INV_X1     g29862(.I(new_n33133_), .ZN(new_n33135_));
  NOR2_X1    g29863(.A1(new_n33135_), .A2(new_n8686_), .ZN(new_n33136_));
  OAI21_X1   g29864(.A1(new_n33136_), .A2(new_n33134_), .B(new_n32900_), .ZN(new_n33137_));
  NAND2_X1   g29865(.A1(new_n33137_), .A2(pi0212), .ZN(new_n33138_));
  NOR2_X1    g29866(.A1(new_n32900_), .A2(new_n30588_), .ZN(new_n33139_));
  OAI21_X1   g29867(.A1(new_n32947_), .A2(pi0214), .B(new_n8739_), .ZN(new_n33140_));
  OAI22_X1   g29868(.A1(new_n33138_), .A2(new_n33140_), .B1(new_n8685_), .B2(new_n33139_), .ZN(new_n33141_));
  NOR2_X1    g29869(.A1(new_n33141_), .A2(new_n32837_), .ZN(new_n33142_));
  NOR2_X1    g29870(.A1(new_n32837_), .A2(new_n8683_), .ZN(new_n33143_));
  XOR2_X1    g29871(.A1(new_n33142_), .A2(new_n33143_), .Z(new_n33144_));
  NAND2_X1   g29872(.A1(new_n32977_), .A2(new_n31954_), .ZN(new_n33145_));
  INV_X1     g29873(.I(new_n31954_), .ZN(new_n33146_));
  NOR2_X1    g29874(.A1(new_n33146_), .A2(new_n8683_), .ZN(new_n33147_));
  XOR2_X1    g29875(.A1(new_n33145_), .A2(new_n33147_), .Z(new_n33148_));
  NAND4_X1   g29876(.A1(new_n32975_), .A2(pi1150), .A3(new_n31996_), .A4(new_n32900_), .ZN(new_n33149_));
  NOR2_X1    g29877(.A1(new_n33148_), .A2(new_n33149_), .ZN(new_n33150_));
  NAND2_X1   g29878(.A1(new_n31757_), .A2(new_n32242_), .ZN(new_n33151_));
  AOI21_X1   g29879(.A1(new_n33150_), .A2(new_n33144_), .B(new_n33151_), .ZN(new_n33152_));
  NAND2_X1   g29880(.A1(po1038), .A2(pi1147), .ZN(new_n33153_));
  OAI21_X1   g29881(.A1(new_n8685_), .A2(new_n32910_), .B(new_n33138_), .ZN(new_n33154_));
  AOI21_X1   g29882(.A1(new_n33135_), .A2(new_n33140_), .B(pi0219), .ZN(new_n33155_));
  NAND2_X1   g29883(.A1(new_n33154_), .A2(new_n33155_), .ZN(new_n33156_));
  AOI21_X1   g29884(.A1(new_n32900_), .A2(pi0219), .B(new_n31940_), .ZN(new_n33157_));
  NAND2_X1   g29885(.A1(new_n33156_), .A2(new_n33157_), .ZN(new_n33158_));
  XOR2_X1    g29886(.A1(new_n33158_), .A2(new_n33153_), .Z(new_n33159_));
  AOI21_X1   g29887(.A1(new_n33017_), .A2(pi0214), .B(pi0212), .ZN(new_n33160_));
  OAI21_X1   g29888(.A1(new_n32976_), .A2(new_n32958_), .B(new_n8683_), .ZN(new_n33161_));
  OAI22_X1   g29889(.A1(new_n33161_), .A2(new_n33160_), .B1(new_n8683_), .B2(new_n32932_), .ZN(new_n33162_));
  NAND2_X1   g29890(.A1(new_n32932_), .A2(pi1147), .ZN(new_n33163_));
  XOR2_X1    g29891(.A1(new_n33163_), .A2(new_n33153_), .Z(new_n33164_));
  NOR3_X1    g29892(.A1(new_n32947_), .A2(new_n31941_), .A3(new_n33131_), .ZN(new_n33165_));
  NAND4_X1   g29893(.A1(new_n33159_), .A2(new_n33162_), .A3(new_n33164_), .A4(new_n33165_), .ZN(new_n33166_));
  NOR2_X1    g29894(.A1(new_n33166_), .A2(new_n33152_), .ZN(new_n33167_));
  XNOR2_X1   g29895(.A1(new_n33167_), .A2(new_n33132_), .ZN(new_n33168_));
  AOI21_X1   g29896(.A1(new_n32990_), .A2(new_n32997_), .B(new_n32837_), .ZN(new_n33169_));
  INV_X1     g29897(.I(new_n33169_), .ZN(new_n33170_));
  NOR3_X1    g29898(.A1(new_n32970_), .A2(pi0219), .A3(new_n30594_), .ZN(new_n33171_));
  OAI21_X1   g29899(.A1(new_n33171_), .A2(pi0212), .B(new_n32969_), .ZN(new_n33172_));
  NAND2_X1   g29900(.A1(new_n32321_), .A2(new_n31954_), .ZN(new_n33173_));
  NOR3_X1    g29901(.A1(new_n31993_), .A2(new_n31941_), .A3(pi1150), .ZN(new_n33174_));
  OAI21_X1   g29902(.A1(new_n33172_), .A2(new_n33173_), .B(new_n33174_), .ZN(new_n33175_));
  INV_X1     g29903(.I(new_n33139_), .ZN(new_n33176_));
  OAI21_X1   g29904(.A1(new_n32999_), .A2(new_n33176_), .B(new_n8683_), .ZN(new_n33177_));
  NAND2_X1   g29905(.A1(new_n32913_), .A2(new_n33176_), .ZN(new_n33178_));
  NOR2_X1    g29906(.A1(new_n30597_), .A2(new_n31953_), .ZN(new_n33179_));
  NAND4_X1   g29907(.A1(new_n33177_), .A2(new_n32910_), .A3(new_n33178_), .A4(new_n33179_), .ZN(new_n33180_));
  AOI21_X1   g29908(.A1(new_n33175_), .A2(new_n33170_), .B(new_n33180_), .ZN(new_n33181_));
  NAND2_X1   g29909(.A1(new_n9163_), .A2(new_n3229_), .ZN(new_n33188_));
  NOR2_X1    g29910(.A1(new_n33172_), .A2(new_n33188_), .ZN(new_n33189_));
  OAI21_X1   g29911(.A1(new_n33181_), .A2(pi1150), .B(new_n33189_), .ZN(new_n33190_));
  NAND2_X1   g29912(.A1(new_n30594_), .A2(new_n8683_), .ZN(new_n33191_));
  AOI21_X1   g29913(.A1(new_n32969_), .A2(new_n33191_), .B(new_n33146_), .ZN(new_n33192_));
  NOR2_X1    g29914(.A1(new_n32967_), .A2(pi0214), .ZN(new_n33193_));
  AOI21_X1   g29915(.A1(new_n33193_), .A2(new_n8739_), .B(new_n31523_), .ZN(new_n33194_));
  AOI21_X1   g29916(.A1(new_n32962_), .A2(new_n8739_), .B(pi0219), .ZN(new_n33195_));
  AOI21_X1   g29917(.A1(new_n33194_), .A2(new_n33195_), .B(pi0214), .ZN(new_n33196_));
  OAI21_X1   g29918(.A1(new_n33196_), .A2(new_n32961_), .B(new_n33192_), .ZN(new_n33197_));
  AOI21_X1   g29919(.A1(new_n8683_), .A2(new_n32946_), .B(new_n33170_), .ZN(new_n33198_));
  NOR3_X1    g29920(.A1(new_n33198_), .A2(pi1150), .A3(new_n31758_), .ZN(new_n33199_));
  AOI21_X1   g29921(.A1(new_n33199_), .A2(new_n33197_), .B(pi1149), .ZN(new_n33200_));
  NAND2_X1   g29922(.A1(new_n33194_), .A2(new_n8683_), .ZN(new_n33201_));
  OAI21_X1   g29923(.A1(new_n33201_), .A2(new_n32980_), .B(new_n32972_), .ZN(new_n33202_));
  INV_X1     g29924(.I(new_n31973_), .ZN(new_n33203_));
  AOI21_X1   g29925(.A1(new_n33203_), .A2(new_n32242_), .B(new_n8685_), .ZN(new_n33204_));
  NAND4_X1   g29926(.A1(new_n33202_), .A2(new_n33169_), .A3(new_n33192_), .A4(new_n33204_), .ZN(new_n33205_));
  NAND2_X1   g29927(.A1(new_n32921_), .A2(new_n33205_), .ZN(new_n33206_));
  NOR2_X1    g29928(.A1(new_n33139_), .A2(pi0214), .ZN(new_n33207_));
  AOI21_X1   g29929(.A1(new_n32917_), .A2(new_n33207_), .B(new_n32913_), .ZN(new_n33208_));
  NAND2_X1   g29930(.A1(new_n33206_), .A2(new_n33208_), .ZN(new_n33209_));
  AOI21_X1   g29931(.A1(new_n33190_), .A2(new_n33200_), .B(new_n33209_), .ZN(new_n33210_));
  OAI21_X1   g29932(.A1(new_n33210_), .A2(pi0213), .B(pi1148), .ZN(new_n33211_));
  OAI21_X1   g29933(.A1(new_n33168_), .A2(new_n33211_), .B(new_n28364_), .ZN(new_n33212_));
  NOR3_X1    g29934(.A1(new_n32995_), .A2(new_n30557_), .A3(new_n4549_), .ZN(new_n33213_));
  NAND2_X1   g29935(.A1(new_n33212_), .A2(new_n33213_), .ZN(new_n33214_));
  XNOR2_X1   g29936(.A1(new_n33214_), .A2(new_n33128_), .ZN(po0403));
  OAI21_X1   g29937(.A1(new_n32075_), .A2(new_n32080_), .B(new_n32239_), .ZN(new_n33216_));
  NAND2_X1   g29938(.A1(new_n32238_), .A2(new_n31940_), .ZN(new_n33217_));
  NAND2_X1   g29939(.A1(new_n32137_), .A2(new_n32334_), .ZN(new_n33218_));
  AOI21_X1   g29940(.A1(new_n33098_), .A2(new_n33218_), .B(new_n32328_), .ZN(new_n33219_));
  NOR2_X1    g29941(.A1(new_n33219_), .A2(new_n32028_), .ZN(new_n33220_));
  AOI21_X1   g29942(.A1(new_n33220_), .A2(pi1151), .B(pi1147), .ZN(new_n33221_));
  NAND2_X1   g29943(.A1(new_n32052_), .A2(pi1151), .ZN(new_n33222_));
  OAI21_X1   g29944(.A1(new_n33221_), .A2(new_n33222_), .B(new_n32242_), .ZN(new_n33223_));
  OAI21_X1   g29945(.A1(new_n32148_), .A2(pi0219), .B(new_n32327_), .ZN(new_n33224_));
  INV_X1     g29946(.I(new_n33224_), .ZN(new_n33225_));
  NOR2_X1    g29947(.A1(new_n33219_), .A2(new_n33225_), .ZN(new_n33226_));
  NAND2_X1   g29948(.A1(new_n33226_), .A2(new_n32239_), .ZN(new_n33227_));
  NAND3_X1   g29949(.A1(new_n31995_), .A2(new_n31940_), .A3(new_n31670_), .ZN(new_n33228_));
  NAND3_X1   g29950(.A1(new_n33227_), .A2(new_n33225_), .A3(new_n33228_), .ZN(new_n33229_));
  AOI21_X1   g29951(.A1(new_n32063_), .A2(new_n31766_), .B(new_n7240_), .ZN(new_n33230_));
  INV_X1     g29952(.I(new_n32028_), .ZN(new_n33231_));
  NOR2_X1    g29953(.A1(new_n32283_), .A2(new_n33231_), .ZN(new_n33232_));
  XOR2_X1    g29954(.A1(new_n33232_), .A2(new_n33230_), .Z(new_n33233_));
  NOR2_X1    g29955(.A1(new_n32190_), .A2(pi1151), .ZN(new_n33234_));
  NOR3_X1    g29956(.A1(new_n33234_), .A2(pi1147), .A3(new_n32242_), .ZN(new_n33235_));
  NAND4_X1   g29957(.A1(new_n33223_), .A2(new_n33229_), .A3(new_n33233_), .A4(new_n33235_), .ZN(new_n33236_));
  AOI21_X1   g29958(.A1(new_n33217_), .A2(new_n33236_), .B(new_n33216_), .ZN(new_n33237_));
  NOR2_X1    g29959(.A1(new_n33237_), .A2(new_n31953_), .ZN(new_n33238_));
  XOR2_X1    g29960(.A1(new_n33238_), .A2(new_n31975_), .Z(new_n33239_));
  INV_X1     g29961(.I(new_n32358_), .ZN(new_n33240_));
  NOR2_X1    g29962(.A1(new_n33049_), .A2(new_n32229_), .ZN(new_n33241_));
  NOR2_X1    g29963(.A1(new_n33241_), .A2(new_n31993_), .ZN(new_n33242_));
  NAND2_X1   g29964(.A1(new_n33242_), .A2(new_n31670_), .ZN(new_n33243_));
  AOI21_X1   g29965(.A1(new_n32228_), .A2(new_n32249_), .B(new_n32122_), .ZN(new_n33244_));
  NOR2_X1    g29966(.A1(new_n33244_), .A2(new_n32370_), .ZN(new_n33245_));
  NOR2_X1    g29967(.A1(new_n32259_), .A2(new_n32308_), .ZN(new_n33246_));
  INV_X1     g29968(.I(new_n33246_), .ZN(new_n33247_));
  AOI21_X1   g29969(.A1(new_n7240_), .A2(new_n32152_), .B(new_n33247_), .ZN(new_n33248_));
  NOR3_X1    g29970(.A1(new_n32257_), .A2(new_n32224_), .A3(new_n32308_), .ZN(new_n33249_));
  NOR3_X1    g29971(.A1(new_n33245_), .A2(pi1147), .A3(pi1150), .ZN(new_n33250_));
  NAND2_X1   g29972(.A1(new_n33060_), .A2(new_n33241_), .ZN(new_n33251_));
  INV_X1     g29973(.I(new_n33251_), .ZN(new_n33252_));
  OAI21_X1   g29974(.A1(new_n33252_), .A2(new_n32259_), .B(new_n31940_), .ZN(new_n33253_));
  NAND2_X1   g29975(.A1(new_n33061_), .A2(new_n32256_), .ZN(new_n33254_));
  NOR2_X1    g29976(.A1(new_n32251_), .A2(pi1147), .ZN(new_n33255_));
  NOR3_X1    g29977(.A1(new_n32324_), .A2(new_n31670_), .A3(new_n31993_), .ZN(new_n33256_));
  INV_X1     g29978(.I(new_n33256_), .ZN(new_n33257_));
  OAI21_X1   g29979(.A1(new_n33257_), .A2(new_n33255_), .B(pi1150), .ZN(new_n33258_));
  NOR2_X1    g29980(.A1(new_n33254_), .A2(new_n33258_), .ZN(new_n33259_));
  AOI22_X1   g29981(.A1(new_n33253_), .A2(new_n33259_), .B1(new_n33243_), .B2(new_n33250_), .ZN(new_n33260_));
  NOR2_X1    g29982(.A1(new_n32138_), .A2(new_n31090_), .ZN(new_n33261_));
  OAI21_X1   g29983(.A1(new_n32134_), .A2(new_n32296_), .B(new_n33261_), .ZN(new_n33262_));
  INV_X1     g29984(.I(new_n33262_), .ZN(new_n33263_));
  NOR2_X1    g29985(.A1(new_n33263_), .A2(new_n32240_), .ZN(new_n33264_));
  NOR2_X1    g29986(.A1(new_n33264_), .A2(pi1147), .ZN(new_n33265_));
  OAI21_X1   g29987(.A1(new_n32149_), .A2(new_n32297_), .B(new_n31995_), .ZN(new_n33266_));
  OR2_X2     g29988(.A1(new_n33266_), .A2(new_n31670_), .Z(new_n33267_));
  OAI21_X1   g29989(.A1(new_n33265_), .A2(new_n33267_), .B(new_n32242_), .ZN(new_n33268_));
  NOR2_X1    g29990(.A1(new_n12654_), .A2(new_n31740_), .ZN(new_n33269_));
  NOR2_X1    g29991(.A1(new_n32089_), .A2(pi0214), .ZN(new_n33270_));
  NOR3_X1    g29992(.A1(new_n33269_), .A2(pi1147), .A3(new_n31670_), .ZN(new_n33271_));
  AOI21_X1   g29993(.A1(new_n33268_), .A2(new_n33271_), .B(new_n31975_), .ZN(new_n33272_));
  NAND3_X1   g29994(.A1(new_n32091_), .A2(new_n31940_), .A3(pi1151), .ZN(new_n33273_));
  NOR2_X1    g29995(.A1(new_n33087_), .A2(pi1151), .ZN(new_n33274_));
  NOR3_X1    g29996(.A1(new_n33274_), .A2(new_n31940_), .A3(pi1150), .ZN(new_n33275_));
  AOI21_X1   g29997(.A1(new_n33275_), .A2(new_n33273_), .B(new_n32028_), .ZN(new_n33276_));
  NOR4_X1    g29998(.A1(new_n33260_), .A2(new_n33240_), .A3(new_n33272_), .A4(new_n33276_), .ZN(new_n33277_));
  NAND2_X1   g29999(.A1(new_n33239_), .A2(new_n33277_), .ZN(new_n33278_));
  AOI21_X1   g30000(.A1(new_n31613_), .A2(new_n32307_), .B(new_n32352_), .ZN(new_n33279_));
  INV_X1     g30001(.I(new_n33279_), .ZN(new_n33280_));
  NOR2_X1    g30002(.A1(new_n31606_), .A2(new_n31810_), .ZN(new_n33281_));
  AOI21_X1   g30003(.A1(new_n33280_), .A2(new_n33281_), .B(new_n30597_), .ZN(new_n33282_));
  NOR2_X1    g30004(.A1(new_n33279_), .A2(new_n32259_), .ZN(new_n33283_));
  NOR2_X1    g30005(.A1(new_n33283_), .A2(pi1147), .ZN(new_n33284_));
  NOR2_X1    g30006(.A1(new_n33284_), .A2(new_n32257_), .ZN(new_n33285_));
  AOI21_X1   g30007(.A1(new_n33285_), .A2(new_n33282_), .B(pi1150), .ZN(new_n33286_));
  INV_X1     g30008(.I(new_n32105_), .ZN(new_n33287_));
  NOR2_X1    g30009(.A1(new_n32342_), .A2(pi0219), .ZN(new_n33288_));
  AOI21_X1   g30010(.A1(new_n32108_), .A2(new_n33288_), .B(new_n32304_), .ZN(new_n33289_));
  AOI21_X1   g30011(.A1(new_n33287_), .A2(new_n33289_), .B(new_n32259_), .ZN(new_n33290_));
  INV_X1     g30012(.I(new_n33290_), .ZN(new_n33291_));
  NOR4_X1    g30013(.A1(new_n33291_), .A2(new_n31940_), .A3(new_n32258_), .A4(new_n33286_), .ZN(new_n33292_));
  NOR2_X1    g30014(.A1(new_n32349_), .A2(new_n31993_), .ZN(new_n33293_));
  INV_X1     g30015(.I(new_n33293_), .ZN(new_n33294_));
  NOR2_X1    g30016(.A1(new_n33294_), .A2(pi1151), .ZN(new_n33295_));
  NAND2_X1   g30017(.A1(new_n31606_), .A2(new_n31810_), .ZN(new_n33296_));
  AOI21_X1   g30018(.A1(new_n32348_), .A2(new_n32250_), .B(new_n33296_), .ZN(new_n33297_));
  OR2_X2     g30019(.A1(new_n33297_), .A2(pi1147), .Z(new_n33298_));
  OAI21_X1   g30020(.A1(new_n33295_), .A2(new_n33298_), .B(new_n32242_), .ZN(new_n33299_));
  OAI21_X1   g30021(.A1(new_n32108_), .A2(new_n33075_), .B(new_n8739_), .ZN(new_n33300_));
  NAND2_X1   g30022(.A1(new_n33300_), .A2(new_n31691_), .ZN(new_n33301_));
  NAND2_X1   g30023(.A1(new_n33301_), .A2(new_n32249_), .ZN(new_n33302_));
  NAND2_X1   g30024(.A1(new_n33302_), .A2(pi1147), .ZN(new_n33303_));
  NOR2_X1    g30025(.A1(new_n33289_), .A2(new_n31993_), .ZN(new_n33304_));
  AOI21_X1   g30026(.A1(new_n31670_), .A2(new_n33304_), .B(new_n33303_), .ZN(new_n33305_));
  OAI21_X1   g30027(.A1(new_n33292_), .A2(new_n33299_), .B(new_n33305_), .ZN(new_n33306_));
  AOI21_X1   g30028(.A1(new_n33278_), .A2(new_n31941_), .B(new_n33306_), .ZN(new_n33307_));
  NOR2_X1    g30029(.A1(new_n33307_), .A2(new_n28529_), .ZN(new_n33308_));
  XOR2_X1    g30030(.A1(new_n33308_), .A2(new_n31079_), .Z(new_n33309_));
  AOI21_X1   g30031(.A1(new_n33309_), .A2(new_n32159_), .B(new_n30557_), .ZN(new_n33310_));
  NOR2_X1    g30032(.A1(pi1147), .A2(pi1150), .ZN(new_n33311_));
  NAND2_X1   g30033(.A1(new_n33220_), .A2(new_n31670_), .ZN(new_n33312_));
  NAND2_X1   g30034(.A1(new_n33312_), .A2(new_n33311_), .ZN(new_n33313_));
  NAND2_X1   g30035(.A1(new_n33231_), .A2(pi1151), .ZN(new_n33314_));
  NOR4_X1    g30036(.A1(new_n33249_), .A2(new_n31940_), .A3(new_n32224_), .A4(new_n33314_), .ZN(new_n33315_));
  AOI22_X1   g30037(.A1(new_n33313_), .A2(new_n33315_), .B1(new_n33203_), .B2(new_n32144_), .ZN(new_n33316_));
  NOR2_X1    g30038(.A1(new_n32028_), .A2(pi1151), .ZN(new_n33317_));
  INV_X1     g30039(.I(new_n33317_), .ZN(new_n33318_));
  OAI21_X1   g30040(.A1(new_n32358_), .A2(new_n33318_), .B(new_n31940_), .ZN(new_n33319_));
  AOI21_X1   g30041(.A1(new_n32103_), .A2(new_n32165_), .B(new_n33314_), .ZN(new_n33320_));
  AOI21_X1   g30042(.A1(new_n33320_), .A2(new_n33319_), .B(pi1150), .ZN(new_n33321_));
  NOR2_X1    g30043(.A1(new_n32258_), .A2(new_n31940_), .ZN(new_n33322_));
  NOR2_X1    g30044(.A1(new_n31973_), .A2(pi1151), .ZN(new_n33323_));
  INV_X1     g30045(.I(new_n33323_), .ZN(new_n33324_));
  NOR2_X1    g30046(.A1(new_n32145_), .A2(new_n33324_), .ZN(new_n33325_));
  NAND2_X1   g30047(.A1(new_n33322_), .A2(new_n33325_), .ZN(new_n33326_));
  OAI22_X1   g30048(.A1(new_n33326_), .A2(new_n33321_), .B1(new_n31670_), .B2(new_n33316_), .ZN(new_n33327_));
  AOI21_X1   g30049(.A1(new_n33327_), .A2(pi1149), .B(new_n31953_), .ZN(new_n33328_));
  NAND2_X1   g30050(.A1(new_n33242_), .A2(pi1151), .ZN(new_n33329_));
  NAND2_X1   g30051(.A1(new_n33329_), .A2(new_n31940_), .ZN(new_n33330_));
  AOI21_X1   g30052(.A1(new_n33036_), .A2(new_n31993_), .B(new_n32067_), .ZN(new_n33331_));
  NAND2_X1   g30053(.A1(new_n32070_), .A2(pi1151), .ZN(new_n33332_));
  NOR2_X1    g30054(.A1(new_n33331_), .A2(new_n33332_), .ZN(new_n33333_));
  AOI21_X1   g30055(.A1(new_n33333_), .A2(new_n33330_), .B(pi1149), .ZN(new_n33334_));
  NOR2_X1    g30056(.A1(new_n31996_), .A2(new_n31670_), .ZN(new_n33335_));
  OAI21_X1   g30057(.A1(new_n33047_), .A2(new_n32125_), .B(new_n33335_), .ZN(new_n33336_));
  NOR3_X1    g30058(.A1(new_n33217_), .A2(new_n33334_), .A3(new_n33336_), .ZN(new_n33337_));
  NOR2_X1    g30059(.A1(new_n31756_), .A2(pi1151), .ZN(new_n33338_));
  NAND2_X1   g30060(.A1(new_n33255_), .A2(new_n31941_), .ZN(new_n33339_));
  NAND2_X1   g30061(.A1(new_n33107_), .A2(new_n32239_), .ZN(new_n33340_));
  NOR4_X1    g30062(.A1(new_n32135_), .A2(new_n32051_), .A3(new_n31670_), .A4(new_n31939_), .ZN(new_n33341_));
  NAND4_X1   g30063(.A1(new_n33340_), .A2(new_n31940_), .A3(new_n33339_), .A4(new_n33341_), .ZN(new_n33342_));
  AOI21_X1   g30064(.A1(new_n33226_), .A2(new_n33338_), .B(new_n33342_), .ZN(new_n33343_));
  OAI21_X1   g30065(.A1(new_n33337_), .A2(pi1150), .B(new_n33343_), .ZN(new_n33344_));
  NAND2_X1   g30066(.A1(new_n32395_), .A2(new_n31810_), .ZN(new_n33345_));
  INV_X1     g30067(.I(new_n33345_), .ZN(new_n33346_));
  INV_X1     g30068(.I(new_n33335_), .ZN(new_n33347_));
  NOR2_X1    g30069(.A1(new_n33294_), .A2(new_n31670_), .ZN(new_n33348_));
  NOR2_X1    g30070(.A1(new_n33348_), .A2(new_n31942_), .ZN(new_n33349_));
  AOI21_X1   g30071(.A1(new_n33270_), .A2(new_n31670_), .B(pi1147), .ZN(new_n33350_));
  NAND2_X1   g30072(.A1(new_n31992_), .A2(pi1151), .ZN(new_n33351_));
  AOI21_X1   g30073(.A1(new_n32051_), .A2(new_n33351_), .B(new_n30918_), .ZN(new_n33352_));
  NAND2_X1   g30074(.A1(new_n33352_), .A2(new_n33350_), .ZN(new_n33353_));
  OAI21_X1   g30075(.A1(new_n33349_), .A2(new_n33353_), .B(new_n33347_), .ZN(new_n33354_));
  AOI21_X1   g30076(.A1(new_n33354_), .A2(new_n33346_), .B(pi1150), .ZN(new_n33355_));
  NAND2_X1   g30077(.A1(new_n33344_), .A2(new_n33355_), .ZN(new_n33356_));
  NOR3_X1    g30078(.A1(new_n33252_), .A2(new_n31670_), .A3(new_n31758_), .ZN(new_n33357_));
  NOR2_X1    g30079(.A1(new_n33357_), .A2(pi1147), .ZN(new_n33358_));
  OR2_X2     g30080(.A1(new_n33235_), .A2(pi1151), .Z(new_n33359_));
  NAND3_X1   g30081(.A1(new_n33280_), .A2(pi1151), .A3(new_n31955_), .ZN(new_n33360_));
  NAND3_X1   g30082(.A1(new_n32088_), .A2(new_n31940_), .A3(pi1151), .ZN(new_n33361_));
  AOI21_X1   g30083(.A1(new_n33361_), .A2(new_n32242_), .B(pi1147), .ZN(new_n33362_));
  NAND2_X1   g30084(.A1(new_n33360_), .A2(new_n33362_), .ZN(new_n33363_));
  NOR2_X1    g30085(.A1(new_n33247_), .A2(new_n31941_), .ZN(new_n33364_));
  AOI22_X1   g30086(.A1(new_n33359_), .A2(new_n32124_), .B1(new_n33363_), .B2(new_n33364_), .ZN(new_n33365_));
  OAI21_X1   g30087(.A1(new_n33037_), .A2(new_n32066_), .B(new_n31955_), .ZN(new_n33366_));
  INV_X1     g30088(.I(new_n33366_), .ZN(new_n33367_));
  NOR3_X1    g30089(.A1(new_n33263_), .A2(pi1151), .A3(new_n31756_), .ZN(new_n33368_));
  AOI21_X1   g30090(.A1(new_n31756_), .A2(new_n32165_), .B(new_n33074_), .ZN(new_n33369_));
  NOR3_X1    g30091(.A1(new_n32412_), .A2(new_n31670_), .A3(new_n33369_), .ZN(new_n33370_));
  OAI21_X1   g30092(.A1(new_n33368_), .A2(pi1147), .B(new_n33370_), .ZN(new_n33371_));
  NAND2_X1   g30093(.A1(new_n33371_), .A2(new_n31941_), .ZN(new_n33372_));
  NOR4_X1    g30094(.A1(new_n32146_), .A2(new_n31670_), .A3(new_n31939_), .A4(new_n33262_), .ZN(new_n33373_));
  NOR2_X1    g30095(.A1(new_n31953_), .A2(new_n31670_), .ZN(new_n33374_));
  NAND4_X1   g30096(.A1(new_n33367_), .A2(new_n33373_), .A3(new_n33372_), .A4(new_n33374_), .ZN(new_n33375_));
  NOR4_X1    g30097(.A1(new_n33375_), .A2(new_n33303_), .A3(new_n33358_), .A4(new_n33365_), .ZN(new_n33376_));
  NAND2_X1   g30098(.A1(new_n33356_), .A2(new_n33376_), .ZN(new_n33377_));
  OAI21_X1   g30099(.A1(new_n33377_), .A2(new_n33328_), .B(pi0209), .ZN(new_n33378_));
  AOI21_X1   g30100(.A1(new_n33328_), .A2(new_n33377_), .B(new_n33378_), .ZN(new_n33379_));
  XOR2_X1    g30101(.A1(new_n33379_), .A2(new_n31080_), .Z(new_n33380_));
  NOR4_X1    g30102(.A1(new_n33380_), .A2(new_n30557_), .A3(new_n4459_), .A4(new_n32262_), .ZN(new_n33381_));
  XOR2_X1    g30103(.A1(new_n33310_), .A2(new_n33381_), .Z(po0404));
  NOR2_X1    g30104(.A1(new_n33290_), .A2(pi1152), .ZN(new_n33383_));
  NAND2_X1   g30105(.A1(new_n33304_), .A2(pi1151), .ZN(new_n33384_));
  OAI21_X1   g30106(.A1(new_n33383_), .A2(new_n33384_), .B(new_n32242_), .ZN(new_n33385_));
  OAI21_X1   g30107(.A1(new_n32109_), .A2(new_n33324_), .B(pi1152), .ZN(new_n33386_));
  NOR2_X1    g30108(.A1(new_n33386_), .A2(new_n33302_), .ZN(new_n33387_));
  AOI21_X1   g30109(.A1(new_n33385_), .A2(new_n33387_), .B(pi1149), .ZN(new_n33388_));
  AOI21_X1   g30110(.A1(new_n33251_), .A2(new_n31759_), .B(pi1152), .ZN(new_n33389_));
  AOI21_X1   g30111(.A1(new_n33389_), .A2(new_n33329_), .B(new_n32245_), .ZN(new_n33390_));
  OAI21_X1   g30112(.A1(new_n32081_), .A2(new_n33347_), .B(new_n31002_), .ZN(new_n33391_));
  NOR2_X1    g30113(.A1(new_n33391_), .A2(new_n33234_), .ZN(new_n33392_));
  NAND2_X1   g30114(.A1(new_n33233_), .A2(pi1151), .ZN(new_n33393_));
  AOI21_X1   g30115(.A1(new_n31002_), .A2(new_n33216_), .B(new_n33393_), .ZN(new_n33394_));
  INV_X1     g30116(.I(new_n33270_), .ZN(new_n33395_));
  NOR3_X1    g30117(.A1(new_n32091_), .A2(pi1151), .A3(new_n31002_), .ZN(new_n33397_));
  NOR2_X1    g30118(.A1(new_n33397_), .A2(pi1149), .ZN(new_n33398_));
  NOR2_X1    g30119(.A1(new_n33297_), .A2(pi1152), .ZN(new_n33399_));
  NOR2_X1    g30120(.A1(pi1150), .A2(pi1152), .ZN(new_n33400_));
  INV_X1     g30121(.I(new_n33400_), .ZN(new_n33401_));
  NOR2_X1    g30122(.A1(new_n33348_), .A2(new_n33401_), .ZN(new_n33402_));
  NAND3_X1   g30123(.A1(new_n33282_), .A2(new_n33283_), .A3(new_n33323_), .ZN(new_n33403_));
  NOR4_X1    g30124(.A1(new_n33402_), .A2(new_n33398_), .A3(new_n33399_), .A4(new_n33403_), .ZN(new_n33404_));
  NOR2_X1    g30125(.A1(new_n33245_), .A2(pi1152), .ZN(new_n33405_));
  NOR3_X1    g30126(.A1(new_n33254_), .A2(pi1150), .A3(new_n33405_), .ZN(new_n33406_));
  OAI21_X1   g30127(.A1(new_n33404_), .A2(pi1148), .B(new_n33406_), .ZN(new_n33407_));
  NOR4_X1    g30128(.A1(new_n33392_), .A2(new_n33390_), .A3(new_n33394_), .A4(new_n33407_), .ZN(new_n33408_));
  OAI21_X1   g30129(.A1(new_n32242_), .A2(new_n32313_), .B(new_n33347_), .ZN(new_n33409_));
  NAND2_X1   g30130(.A1(new_n33227_), .A2(new_n31002_), .ZN(new_n33410_));
  AOI21_X1   g30131(.A1(new_n33225_), .A2(new_n33409_), .B(new_n33410_), .ZN(new_n33411_));
  NOR2_X1    g30132(.A1(new_n33248_), .A2(new_n33401_), .ZN(new_n33412_));
  NOR2_X1    g30133(.A1(new_n32251_), .A2(new_n31002_), .ZN(new_n33413_));
  NAND2_X1   g30134(.A1(new_n33256_), .A2(new_n33413_), .ZN(new_n33414_));
  OAI21_X1   g30135(.A1(new_n33412_), .A2(new_n33414_), .B(new_n33324_), .ZN(new_n33415_));
  NAND2_X1   g30136(.A1(new_n31953_), .A2(new_n31941_), .ZN(new_n33416_));
  AOI21_X1   g30137(.A1(new_n33415_), .A2(new_n32309_), .B(new_n33416_), .ZN(new_n33417_));
  NOR2_X1    g30138(.A1(new_n32358_), .A2(new_n33318_), .ZN(new_n33418_));
  NAND2_X1   g30139(.A1(new_n33266_), .A2(pi1151), .ZN(new_n33419_));
  NAND2_X1   g30140(.A1(pi1151), .A2(pi1152), .ZN(new_n33420_));
  XOR2_X1    g30141(.A1(new_n33419_), .A2(new_n33420_), .Z(new_n33421_));
  OAI21_X1   g30142(.A1(new_n33263_), .A2(new_n32240_), .B(new_n33400_), .ZN(new_n33422_));
  NAND4_X1   g30143(.A1(new_n33421_), .A2(new_n33087_), .A3(new_n33418_), .A4(new_n33422_), .ZN(new_n33423_));
  NOR4_X1    g30144(.A1(new_n33423_), .A2(new_n33312_), .A3(new_n33411_), .A4(new_n33417_), .ZN(new_n33424_));
  OAI21_X1   g30145(.A1(new_n33408_), .A2(pi0213), .B(new_n33424_), .ZN(new_n33425_));
  OAI21_X1   g30146(.A1(new_n33425_), .A2(new_n33388_), .B(new_n28364_), .ZN(new_n33426_));
  NOR2_X1    g30147(.A1(new_n33125_), .A2(new_n28529_), .ZN(new_n33427_));
  AOI21_X1   g30148(.A1(new_n33427_), .A2(new_n33426_), .B(new_n30557_), .ZN(new_n33428_));
  OAI21_X1   g30149(.A1(pi1152), .A2(new_n33352_), .B(new_n33333_), .ZN(new_n33429_));
  NAND3_X1   g30150(.A1(new_n33242_), .A2(pi1151), .A3(pi1152), .ZN(new_n33430_));
  AOI21_X1   g30151(.A1(new_n33429_), .A2(new_n32242_), .B(new_n33430_), .ZN(new_n33431_));
  NOR4_X1    g30152(.A1(new_n32135_), .A2(new_n32051_), .A3(new_n31670_), .A4(new_n31939_), .ZN(new_n33432_));
  OAI21_X1   g30153(.A1(new_n33373_), .A2(new_n33401_), .B(new_n33432_), .ZN(new_n33433_));
  NOR2_X1    g30154(.A1(new_n33433_), .A2(new_n33301_), .ZN(new_n33434_));
  OAI21_X1   g30155(.A1(new_n33431_), .A2(pi1148), .B(new_n33434_), .ZN(new_n33435_));
  OAI21_X1   g30156(.A1(new_n33357_), .A2(new_n33283_), .B(pi1152), .ZN(new_n33436_));
  NAND3_X1   g30157(.A1(new_n33436_), .A2(new_n31953_), .A3(new_n32242_), .ZN(new_n33437_));
  NAND2_X1   g30158(.A1(new_n33220_), .A2(pi1151), .ZN(new_n33438_));
  NAND2_X1   g30159(.A1(new_n33438_), .A2(new_n33400_), .ZN(new_n33439_));
  AOI21_X1   g30160(.A1(pi1150), .A2(pi1152), .B(pi1151), .ZN(new_n33440_));
  OAI21_X1   g30161(.A1(new_n32087_), .A2(new_n33440_), .B(new_n33234_), .ZN(new_n33441_));
  NOR2_X1    g30162(.A1(new_n31953_), .A2(new_n31002_), .ZN(new_n33442_));
  AOI22_X1   g30163(.A1(new_n33439_), .A2(new_n33418_), .B1(new_n33441_), .B2(new_n33442_), .ZN(new_n33443_));
  OAI21_X1   g30164(.A1(new_n32224_), .A2(new_n33314_), .B(new_n31002_), .ZN(new_n33444_));
  NAND2_X1   g30165(.A1(new_n33320_), .A2(new_n33444_), .ZN(new_n33445_));
  OAI21_X1   g30166(.A1(new_n33445_), .A2(new_n33443_), .B(new_n31941_), .ZN(new_n33446_));
  NAND2_X1   g30167(.A1(pi1150), .A2(pi1151), .ZN(new_n33447_));
  NOR3_X1    g30168(.A1(new_n32143_), .A2(new_n31973_), .A3(new_n33447_), .ZN(new_n33448_));
  OAI21_X1   g30169(.A1(new_n33325_), .A2(pi1152), .B(new_n33448_), .ZN(new_n33449_));
  NAND2_X1   g30170(.A1(new_n33386_), .A2(new_n33449_), .ZN(new_n33450_));
  NAND4_X1   g30171(.A1(new_n32309_), .A2(pi1149), .A3(pi1151), .A4(new_n33203_), .ZN(new_n33452_));
  NOR2_X1    g30172(.A1(new_n33366_), .A2(new_n33452_), .ZN(new_n33453_));
  NAND4_X1   g30173(.A1(new_n33437_), .A2(new_n33450_), .A3(new_n33446_), .A4(new_n33453_), .ZN(new_n33454_));
  NAND2_X1   g30174(.A1(new_n33454_), .A2(new_n33435_), .ZN(new_n33455_));
  NAND3_X1   g30175(.A1(new_n33345_), .A2(new_n31670_), .A3(new_n31002_), .ZN(new_n33456_));
  NAND3_X1   g30176(.A1(new_n33456_), .A2(new_n31996_), .A3(new_n33336_), .ZN(new_n33457_));
  NOR2_X1    g30177(.A1(new_n33391_), .A2(pi1150), .ZN(new_n33458_));
  NAND2_X1   g30178(.A1(new_n33458_), .A2(new_n33457_), .ZN(new_n33459_));
  NAND2_X1   g30179(.A1(new_n33459_), .A2(new_n31670_), .ZN(new_n33460_));
  AOI21_X1   g30180(.A1(new_n33460_), .A2(new_n33395_), .B(pi1148), .ZN(new_n33461_));
  NOR2_X1    g30181(.A1(new_n33410_), .A2(pi1150), .ZN(new_n33462_));
  NAND2_X1   g30182(.A1(new_n33340_), .A2(new_n31002_), .ZN(new_n33463_));
  NAND3_X1   g30183(.A1(new_n33368_), .A2(new_n33463_), .A3(new_n33370_), .ZN(new_n33464_));
  NOR3_X1    g30184(.A1(new_n33461_), .A2(new_n33462_), .A3(new_n33464_), .ZN(new_n33465_));
  AOI21_X1   g30185(.A1(new_n33465_), .A2(new_n33455_), .B(new_n28364_), .ZN(new_n33466_));
  XOR2_X1    g30186(.A1(new_n33466_), .A2(new_n31079_), .Z(new_n33467_));
  OAI21_X1   g30187(.A1(new_n32260_), .A2(pi1152), .B(new_n32253_), .ZN(new_n33468_));
  NAND2_X1   g30188(.A1(new_n33468_), .A2(new_n32242_), .ZN(new_n33469_));
  NOR4_X1    g30189(.A1(new_n32109_), .A2(new_n31002_), .A3(new_n32251_), .A4(new_n33324_), .ZN(new_n33470_));
  NOR3_X1    g30190(.A1(new_n32091_), .A2(pi1151), .A3(new_n32087_), .ZN(new_n33471_));
  OAI21_X1   g30191(.A1(new_n32241_), .A2(pi1152), .B(new_n33471_), .ZN(new_n33472_));
  NAND2_X1   g30192(.A1(new_n33472_), .A2(new_n32242_), .ZN(new_n33473_));
  AOI21_X1   g30193(.A1(new_n33469_), .A2(new_n33470_), .B(new_n33473_), .ZN(new_n33474_));
  NOR4_X1    g30194(.A1(new_n33474_), .A2(new_n31670_), .A3(pi1152), .A4(new_n32082_), .ZN(new_n33475_));
  NAND4_X1   g30195(.A1(new_n33467_), .A2(pi0230), .A3(pi0248), .A4(new_n33475_), .ZN(new_n33476_));
  XNOR2_X1   g30196(.A1(new_n33476_), .A2(new_n33428_), .ZN(po0405));
  NOR2_X1    g30197(.A1(new_n30976_), .A2(new_n8684_), .ZN(new_n33478_));
  NOR2_X1    g30198(.A1(new_n30969_), .A2(new_n31569_), .ZN(new_n33479_));
  NOR2_X1    g30199(.A1(new_n33479_), .A2(new_n30829_), .ZN(new_n33480_));
  AOI22_X1   g30200(.A1(new_n33480_), .A2(new_n30693_), .B1(new_n8545_), .B2(new_n31315_), .ZN(new_n33481_));
  AOI21_X1   g30201(.A1(new_n8684_), .A2(new_n33481_), .B(new_n33478_), .ZN(new_n33482_));
  NAND2_X1   g30202(.A1(new_n33482_), .A2(pi0219), .ZN(new_n33483_));
  XOR2_X1    g30203(.A1(new_n33483_), .A2(new_n31042_), .Z(new_n33484_));
  AOI21_X1   g30204(.A1(new_n33484_), .A2(new_n30976_), .B(po1038), .ZN(new_n33485_));
  NAND2_X1   g30205(.A1(new_n33481_), .A2(new_n8686_), .ZN(new_n33486_));
  NAND2_X1   g30206(.A1(new_n30976_), .A2(new_n8686_), .ZN(new_n33487_));
  XNOR2_X1   g30207(.A1(new_n33487_), .A2(new_n33486_), .ZN(new_n33488_));
  NAND2_X1   g30208(.A1(new_n33488_), .A2(pi0212), .ZN(new_n33489_));
  XOR2_X1    g30209(.A1(new_n33489_), .A2(new_n30916_), .Z(new_n33490_));
  NAND2_X1   g30210(.A1(new_n33490_), .A2(new_n30976_), .ZN(new_n33491_));
  AOI21_X1   g30211(.A1(new_n33491_), .A2(new_n33485_), .B(new_n32259_), .ZN(new_n33492_));
  INV_X1     g30212(.I(new_n33485_), .ZN(new_n33493_));
  NAND2_X1   g30213(.A1(new_n33488_), .A2(new_n8739_), .ZN(new_n33494_));
  NAND2_X1   g30214(.A1(new_n33481_), .A2(pi0211), .ZN(new_n33495_));
  XOR2_X1    g30215(.A1(new_n33495_), .A2(new_n30718_), .Z(new_n33496_));
  NAND2_X1   g30216(.A1(new_n8683_), .A2(pi0212), .ZN(new_n33497_));
  AOI21_X1   g30217(.A1(new_n33496_), .A2(new_n30976_), .B(new_n33497_), .ZN(new_n33498_));
  AOI21_X1   g30218(.A1(new_n33494_), .A2(new_n33498_), .B(pi0214), .ZN(new_n33499_));
  NOR2_X1    g30219(.A1(new_n31993_), .A2(pi1151), .ZN(new_n33500_));
  OR3_X2     g30220(.A1(new_n33499_), .A2(new_n33481_), .A3(new_n33500_), .Z(new_n33501_));
  OAI21_X1   g30221(.A1(new_n33493_), .A2(new_n33501_), .B(new_n31002_), .ZN(new_n33502_));
  OAI21_X1   g30222(.A1(new_n33492_), .A2(new_n33502_), .B(pi1150), .ZN(new_n33503_));
  OAI21_X1   g30223(.A1(new_n33499_), .A2(new_n33482_), .B(new_n7240_), .ZN(new_n33504_));
  NAND2_X1   g30224(.A1(new_n31023_), .A2(new_n8685_), .ZN(new_n33505_));
  OAI21_X1   g30225(.A1(new_n31039_), .A2(new_n31024_), .B(pi0214), .ZN(new_n33506_));
  NAND2_X1   g30226(.A1(new_n31040_), .A2(pi0212), .ZN(new_n33507_));
  XOR2_X1    g30227(.A1(new_n33507_), .A2(new_n30597_), .Z(new_n33508_));
  NAND2_X1   g30228(.A1(new_n31038_), .A2(pi0211), .ZN(new_n33509_));
  NAND2_X1   g30229(.A1(new_n31022_), .A2(new_n8684_), .ZN(new_n33510_));
  AOI21_X1   g30230(.A1(new_n33509_), .A2(new_n33510_), .B(new_n8683_), .ZN(new_n33511_));
  NAND2_X1   g30231(.A1(new_n33508_), .A2(new_n33511_), .ZN(new_n33512_));
  AOI22_X1   g30232(.A1(new_n33512_), .A2(new_n8739_), .B1(new_n33505_), .B2(new_n33506_), .ZN(new_n33513_));
  OAI21_X1   g30233(.A1(new_n33513_), .A2(new_n31044_), .B(new_n33323_), .ZN(new_n33514_));
  NAND2_X1   g30234(.A1(new_n33514_), .A2(new_n31002_), .ZN(new_n33515_));
  INV_X1     g30235(.I(new_n31038_), .ZN(new_n33516_));
  NAND2_X1   g30236(.A1(new_n31040_), .A2(new_n31765_), .ZN(new_n33517_));
  XNOR2_X1   g30237(.A1(new_n33517_), .A2(new_n31768_), .ZN(new_n33518_));
  OAI21_X1   g30238(.A1(new_n33518_), .A2(new_n31022_), .B(new_n33317_), .ZN(new_n33519_));
  NAND2_X1   g30239(.A1(new_n33519_), .A2(new_n31002_), .ZN(new_n33520_));
  NOR2_X1    g30240(.A1(new_n31038_), .A2(new_n8685_), .ZN(new_n33521_));
  XOR2_X1    g30241(.A1(new_n33521_), .A2(new_n8740_), .Z(new_n33522_));
  AOI21_X1   g30242(.A1(new_n33522_), .A2(new_n31023_), .B(pi0219), .ZN(new_n33523_));
  NAND2_X1   g30243(.A1(new_n33508_), .A2(new_n31038_), .ZN(new_n33524_));
  NOR4_X1    g30244(.A1(new_n30977_), .A2(new_n31670_), .A3(new_n31002_), .A4(po1038), .ZN(new_n33525_));
  OAI21_X1   g30245(.A1(new_n31023_), .A2(new_n8683_), .B(new_n33525_), .ZN(new_n33526_));
  AOI21_X1   g30246(.A1(new_n33524_), .A2(new_n33523_), .B(new_n33526_), .ZN(new_n33527_));
  AOI21_X1   g30247(.A1(new_n33520_), .A2(new_n33527_), .B(new_n33335_), .ZN(new_n33528_));
  INV_X1     g30248(.I(new_n33523_), .ZN(new_n33529_));
  NOR2_X1    g30249(.A1(new_n31044_), .A2(new_n33529_), .ZN(new_n33530_));
  NOR2_X1    g30250(.A1(new_n33530_), .A2(pi0212), .ZN(new_n33531_));
  NAND4_X1   g30251(.A1(new_n30976_), .A2(pi0219), .A3(pi1150), .A4(new_n32249_), .ZN(new_n33532_));
  NOR4_X1    g30252(.A1(new_n33528_), .A2(new_n33531_), .A3(new_n33516_), .A4(new_n33532_), .ZN(new_n33533_));
  NAND3_X1   g30253(.A1(new_n33533_), .A2(new_n33504_), .A3(new_n33515_), .ZN(new_n33534_));
  XOR2_X1    g30254(.A1(new_n33534_), .A2(new_n33503_), .Z(new_n33535_));
  NAND2_X1   g30255(.A1(new_n31077_), .A2(pi0209), .ZN(new_n33536_));
  XOR2_X1    g30256(.A1(new_n33536_), .A2(new_n31080_), .Z(new_n33537_));
  AOI21_X1   g30257(.A1(new_n33537_), .A2(new_n33535_), .B(new_n30557_), .ZN(new_n33538_));
  NOR2_X1    g30258(.A1(new_n33475_), .A2(new_n28529_), .ZN(new_n33539_));
  XOR2_X1    g30259(.A1(new_n33539_), .A2(new_n31080_), .Z(new_n33540_));
  OAI22_X1   g30260(.A1(new_n32068_), .A2(new_n30597_), .B1(new_n30989_), .B2(new_n32282_), .ZN(new_n33541_));
  AOI21_X1   g30261(.A1(new_n32071_), .A2(new_n30876_), .B(new_n30829_), .ZN(new_n33542_));
  AOI21_X1   g30262(.A1(new_n33541_), .A2(new_n33542_), .B(new_n32071_), .ZN(new_n33543_));
  NOR2_X1    g30263(.A1(new_n32079_), .A2(pi1151), .ZN(new_n33544_));
  NOR4_X1    g30264(.A1(new_n33543_), .A2(new_n8683_), .A3(new_n30706_), .A4(new_n33544_), .ZN(new_n33545_));
  NAND3_X1   g30265(.A1(new_n30982_), .A2(new_n30597_), .A3(pi0299), .ZN(new_n33546_));
  NOR2_X1    g30266(.A1(new_n31806_), .A2(new_n33546_), .ZN(new_n33547_));
  OAI21_X1   g30267(.A1(new_n31610_), .A2(new_n30984_), .B(new_n33547_), .ZN(new_n33548_));
  NAND2_X1   g30268(.A1(new_n30987_), .A2(new_n33548_), .ZN(new_n33549_));
  OAI21_X1   g30269(.A1(new_n33545_), .A2(new_n33549_), .B(new_n32242_), .ZN(new_n33550_));
  NAND2_X1   g30270(.A1(new_n31691_), .A2(pi0214), .ZN(new_n33551_));
  AOI21_X1   g30271(.A1(new_n33551_), .A2(new_n3098_), .B(new_n30982_), .ZN(new_n33552_));
  AOI21_X1   g30272(.A1(pi0299), .A2(new_n30983_), .B(new_n32344_), .ZN(new_n33553_));
  NOR2_X1    g30273(.A1(new_n33553_), .A2(pi0219), .ZN(new_n33554_));
  OAI21_X1   g30274(.A1(new_n33554_), .A2(new_n33073_), .B(new_n8739_), .ZN(new_n33555_));
  AOI21_X1   g30275(.A1(new_n33551_), .A2(new_n30829_), .B(new_n8684_), .ZN(new_n33556_));
  OAI21_X1   g30276(.A1(new_n33555_), .A2(new_n33552_), .B(new_n33556_), .ZN(new_n33557_));
  NAND3_X1   g30277(.A1(new_n33557_), .A2(new_n31670_), .A3(new_n32107_), .ZN(new_n33558_));
  NOR2_X1    g30278(.A1(new_n31186_), .A2(pi1150), .ZN(new_n33559_));
  AOI21_X1   g30279(.A1(new_n32119_), .A2(pi0212), .B(pi0299), .ZN(new_n33560_));
  NOR3_X1    g30280(.A1(new_n32373_), .A2(new_n30982_), .A3(new_n33560_), .ZN(new_n33561_));
  OR4_X2     g30281(.A1(new_n8739_), .A2(new_n33561_), .A3(new_n32123_), .A4(new_n33554_), .Z(new_n33562_));
  NAND4_X1   g30282(.A1(new_n32141_), .A2(pi1151), .A3(new_n7240_), .A4(new_n33104_), .ZN(new_n33563_));
  NOR2_X1    g30283(.A1(new_n33563_), .A2(new_n32227_), .ZN(new_n33564_));
  NAND2_X1   g30284(.A1(new_n31006_), .A2(new_n33548_), .ZN(new_n33565_));
  OAI21_X1   g30285(.A1(new_n32310_), .A2(new_n31948_), .B(new_n33546_), .ZN(new_n33566_));
  AOI21_X1   g30286(.A1(new_n31001_), .A2(new_n33566_), .B(pi1151), .ZN(new_n33567_));
  NOR2_X1    g30287(.A1(new_n33280_), .A2(new_n33567_), .ZN(new_n33568_));
  NAND4_X1   g30288(.A1(new_n33568_), .A2(new_n33562_), .A3(new_n33564_), .A4(new_n33565_), .ZN(new_n33569_));
  AOI21_X1   g30289(.A1(new_n33558_), .A2(new_n33559_), .B(new_n33569_), .ZN(new_n33570_));
  AOI21_X1   g30290(.A1(new_n33570_), .A2(new_n33550_), .B(pi1152), .ZN(new_n33571_));
  NAND3_X1   g30291(.A1(new_n32133_), .A2(pi0214), .A3(pi0299), .ZN(new_n33572_));
  NAND3_X1   g30292(.A1(new_n32192_), .A2(pi0299), .A3(new_n32220_), .ZN(new_n33573_));
  AOI21_X1   g30293(.A1(new_n33573_), .A2(new_n33572_), .B(new_n30982_), .ZN(new_n33574_));
  NAND4_X1   g30294(.A1(new_n30983_), .A2(pi0212), .A3(new_n10253_), .A4(new_n32364_), .ZN(new_n33575_));
  NOR4_X1    g30295(.A1(new_n31826_), .A2(new_n3098_), .A3(new_n32192_), .A4(new_n33575_), .ZN(new_n33576_));
  OR3_X2     g30296(.A1(new_n33574_), .A2(new_n8739_), .A3(new_n33576_), .Z(new_n33577_));
  OAI21_X1   g30297(.A1(new_n33574_), .A2(new_n8739_), .B(new_n33576_), .ZN(new_n33578_));
  NAND3_X1   g30298(.A1(new_n33577_), .A2(new_n5787_), .A3(new_n33578_), .ZN(new_n33579_));
  NOR2_X1    g30299(.A1(new_n5788_), .A2(new_n8683_), .ZN(new_n33580_));
  XOR2_X1    g30300(.A1(new_n33579_), .A2(new_n33580_), .Z(new_n33581_));
  NOR2_X1    g30301(.A1(new_n30985_), .A2(new_n5787_), .ZN(new_n33582_));
  NAND4_X1   g30302(.A1(new_n32133_), .A2(new_n33582_), .A3(pi0057), .A4(pi1151), .ZN(new_n33583_));
  NOR2_X1    g30303(.A1(new_n33581_), .A2(new_n33583_), .ZN(new_n33584_));
  NOR2_X1    g30304(.A1(new_n30983_), .A2(new_n3098_), .ZN(new_n33585_));
  AOI21_X1   g30305(.A1(new_n31664_), .A2(new_n3098_), .B(new_n33585_), .ZN(new_n33586_));
  NAND2_X1   g30306(.A1(new_n33586_), .A2(pi0214), .ZN(new_n33587_));
  XOR2_X1    g30307(.A1(new_n33587_), .A2(new_n8740_), .Z(new_n33588_));
  OAI21_X1   g30308(.A1(new_n33588_), .A2(new_n31664_), .B(new_n8683_), .ZN(new_n33589_));
  NOR3_X1    g30309(.A1(new_n32136_), .A2(pi0214), .A3(new_n31806_), .ZN(new_n33590_));
  NAND3_X1   g30310(.A1(new_n33589_), .A2(new_n33586_), .A3(new_n33590_), .ZN(new_n33591_));
  NAND4_X1   g30311(.A1(new_n32326_), .A2(pi0057), .A3(pi1151), .A4(new_n33582_), .ZN(new_n33592_));
  AOI21_X1   g30312(.A1(new_n33591_), .A2(new_n5788_), .B(new_n33592_), .ZN(new_n33593_));
  NOR2_X1    g30313(.A1(new_n33584_), .A2(new_n33593_), .ZN(new_n33594_));
  NAND4_X1   g30314(.A1(new_n30986_), .A2(pi0057), .A3(pi0230), .A4(pi0249), .ZN(new_n33595_));
  NOR4_X1    g30315(.A1(new_n33540_), .A2(new_n33571_), .A3(new_n33594_), .A4(new_n33595_), .ZN(new_n33596_));
  XOR2_X1    g30316(.A1(new_n33538_), .A2(new_n33596_), .Z(po0406));
  NAND3_X1   g30317(.A1(new_n12134_), .A2(pi0075), .A3(new_n6285_), .ZN(new_n33598_));
  AOI21_X1   g30318(.A1(new_n9321_), .A2(new_n3213_), .B(new_n33598_), .ZN(new_n33599_));
  XOR2_X1    g30319(.A1(new_n33599_), .A2(new_n7336_), .Z(new_n33600_));
  NOR4_X1    g30320(.A1(new_n33600_), .A2(new_n3455_), .A3(new_n5530_), .A4(new_n7331_), .ZN(po0407));
  NOR2_X1    g30321(.A1(new_n8555_), .A2(pi0476), .ZN(new_n33602_));
  XOR2_X1    g30322(.A1(new_n30722_), .A2(new_n33602_), .Z(new_n33603_));
  NAND2_X1   g30323(.A1(new_n33603_), .A2(pi0897), .ZN(new_n33604_));
  INV_X1     g30324(.I(new_n33604_), .ZN(new_n33605_));
  NAND2_X1   g30325(.A1(new_n33605_), .A2(pi0251), .ZN(new_n33606_));
  INV_X1     g30326(.I(pi1053), .ZN(new_n33607_));
  NAND3_X1   g30327(.A1(pi0199), .A2(pi0200), .A3(pi1039), .ZN(new_n33608_));
  INV_X1     g30328(.I(pi1039), .ZN(new_n33609_));
  NAND3_X1   g30329(.A1(new_n8549_), .A2(new_n33609_), .A3(pi0200), .ZN(new_n33610_));
  AOI21_X1   g30330(.A1(new_n33610_), .A2(new_n33608_), .B(new_n33607_), .ZN(new_n33611_));
  OAI21_X1   g30331(.A1(new_n33605_), .A2(new_n33611_), .B(new_n33606_), .ZN(po0408));
  NOR2_X1    g30332(.A1(new_n7611_), .A2(new_n9380_), .ZN(new_n33613_));
  AND3_X2    g30333(.A1(new_n5405_), .A2(new_n5403_), .A3(pi1001), .Z(new_n33614_));
  NAND3_X1   g30334(.A1(new_n33614_), .A2(pi0835), .A3(pi0950), .ZN(new_n33615_));
  NAND2_X1   g30335(.A1(new_n8930_), .A2(new_n33615_), .ZN(new_n33616_));
  NAND2_X1   g30336(.A1(new_n2979_), .A2(new_n2984_), .ZN(new_n33617_));
  NAND4_X1   g30337(.A1(new_n33616_), .A2(pi0824), .A3(new_n11122_), .A4(new_n33617_), .ZN(new_n33618_));
  NOR2_X1    g30338(.A1(new_n30448_), .A2(new_n33618_), .ZN(new_n33619_));
  AOI21_X1   g30339(.A1(new_n5698_), .A2(new_n33618_), .B(new_n33619_), .ZN(new_n33620_));
  AOI21_X1   g30340(.A1(new_n33620_), .A2(new_n7611_), .B(new_n33613_), .ZN(new_n33621_));
  NAND2_X1   g30341(.A1(new_n33620_), .A2(new_n5385_), .ZN(new_n33622_));
  OAI21_X1   g30342(.A1(new_n5385_), .A2(new_n9380_), .B(new_n33622_), .ZN(new_n33623_));
  NOR2_X1    g30343(.A1(new_n33623_), .A2(new_n5397_), .ZN(new_n33624_));
  XOR2_X1    g30344(.A1(new_n33624_), .A2(new_n8331_), .Z(new_n33625_));
  NOR2_X1    g30345(.A1(new_n33625_), .A2(new_n33621_), .ZN(new_n33626_));
  NOR2_X1    g30346(.A1(new_n33623_), .A2(new_n3098_), .ZN(new_n33627_));
  XOR2_X1    g30347(.A1(new_n33627_), .A2(new_n8338_), .Z(new_n33628_));
  NOR2_X1    g30348(.A1(new_n33628_), .A2(new_n33621_), .ZN(new_n33629_));
  NOR4_X1    g30349(.A1(new_n17124_), .A2(new_n5436_), .A3(new_n8932_), .A4(new_n33615_), .ZN(new_n33630_));
  NOR3_X1    g30350(.A1(new_n33630_), .A2(pi0252), .A3(new_n5679_), .ZN(new_n33631_));
  NOR2_X1    g30351(.A1(pi0057), .A2(pi1092), .ZN(new_n33633_));
  NOR3_X1    g30352(.A1(new_n33631_), .A2(new_n30540_), .A3(new_n33633_), .ZN(new_n33634_));
  NAND2_X1   g30353(.A1(new_n8934_), .A2(new_n9380_), .ZN(new_n33635_));
  NAND2_X1   g30354(.A1(new_n33635_), .A2(new_n10169_), .ZN(new_n33636_));
  NOR2_X1    g30355(.A1(new_n33634_), .A2(new_n33636_), .ZN(new_n33637_));
  NOR4_X1    g30356(.A1(new_n33626_), .A2(new_n33629_), .A3(new_n8934_), .A4(new_n33637_), .ZN(po0409));
  INV_X1     g30357(.I(new_n32773_), .ZN(new_n33639_));
  NOR2_X1    g30358(.A1(new_n31303_), .A2(new_n2726_), .ZN(new_n33640_));
  INV_X1     g30359(.I(new_n33640_), .ZN(new_n33641_));
  NOR2_X1    g30360(.A1(new_n32626_), .A2(new_n2726_), .ZN(new_n33642_));
  INV_X1     g30361(.I(new_n33642_), .ZN(new_n33643_));
  AOI21_X1   g30362(.A1(new_n7240_), .A2(new_n33641_), .B(new_n33643_), .ZN(new_n33644_));
  NOR2_X1    g30363(.A1(new_n10253_), .A2(new_n30659_), .ZN(new_n33645_));
  INV_X1     g30364(.I(new_n33645_), .ZN(new_n33646_));
  NOR2_X1    g30365(.A1(new_n7240_), .A2(new_n33643_), .ZN(new_n33649_));
  NOR2_X1    g30366(.A1(new_n2726_), .A2(pi0211), .ZN(new_n33650_));
  INV_X1     g30367(.I(new_n33650_), .ZN(new_n33651_));
  NAND2_X1   g30368(.A1(new_n33644_), .A2(pi1152), .ZN(new_n33652_));
  NAND2_X1   g30369(.A1(pi0219), .A2(pi1151), .ZN(new_n33653_));
  AOI21_X1   g30370(.A1(new_n33652_), .A2(new_n33651_), .B(new_n33653_), .ZN(new_n33654_));
  OAI21_X1   g30371(.A1(new_n33654_), .A2(new_n33649_), .B(new_n33644_), .ZN(new_n33655_));
  NOR2_X1    g30372(.A1(new_n31936_), .A2(new_n8742_), .ZN(new_n33656_));
  INV_X1     g30373(.I(new_n33656_), .ZN(new_n33657_));
  NAND3_X1   g30374(.A1(new_n30656_), .A2(pi1091), .A3(new_n33657_), .ZN(new_n33658_));
  INV_X1     g30375(.I(new_n30656_), .ZN(new_n33659_));
  NAND3_X1   g30376(.A1(new_n33659_), .A2(new_n2726_), .A3(new_n33657_), .ZN(new_n33660_));
  NAND2_X1   g30377(.A1(new_n33660_), .A2(new_n33658_), .ZN(new_n33661_));
  NAND2_X1   g30378(.A1(new_n33661_), .A2(pi0253), .ZN(new_n33662_));
  NAND3_X1   g30379(.A1(new_n33662_), .A2(new_n33655_), .A3(new_n31651_), .ZN(new_n33663_));
  AOI21_X1   g30380(.A1(pi1153), .A2(new_n30615_), .B(new_n32719_), .ZN(new_n33664_));
  NOR3_X1    g30381(.A1(new_n9259_), .A2(new_n32719_), .A3(pi0253), .ZN(new_n33665_));
  NOR4_X1    g30382(.A1(new_n33659_), .A2(new_n30652_), .A3(new_n33664_), .A4(new_n33665_), .ZN(new_n33666_));
  OAI21_X1   g30383(.A1(new_n33666_), .A2(pi1153), .B(new_n32743_), .ZN(new_n33667_));
  NOR3_X1    g30384(.A1(new_n8684_), .A2(new_n3098_), .A3(new_n2726_), .ZN(new_n33668_));
  NOR2_X1    g30385(.A1(new_n33668_), .A2(pi0253), .ZN(new_n33669_));
  AOI21_X1   g30386(.A1(new_n32754_), .A2(new_n31016_), .B(new_n30616_), .ZN(new_n33670_));
  OAI21_X1   g30387(.A1(new_n31579_), .A2(new_n2726_), .B(new_n33670_), .ZN(new_n33671_));
  AOI21_X1   g30388(.A1(new_n33667_), .A2(new_n33669_), .B(new_n33671_), .ZN(new_n33672_));
  AOI21_X1   g30389(.A1(new_n33663_), .A2(new_n33672_), .B(new_n33639_), .ZN(new_n33673_));
  INV_X1     g30390(.I(new_n33652_), .ZN(new_n33674_));
  NOR2_X1    g30391(.A1(new_n32731_), .A2(pi1153), .ZN(new_n33675_));
  INV_X1     g30392(.I(new_n33675_), .ZN(new_n33676_));
  NAND2_X1   g30393(.A1(new_n32760_), .A2(pi1153), .ZN(new_n33677_));
  NAND4_X1   g30394(.A1(new_n33676_), .A2(pi0253), .A3(new_n33677_), .A4(new_n30615_), .ZN(new_n33678_));
  NAND2_X1   g30395(.A1(new_n33678_), .A2(new_n2726_), .ZN(new_n33679_));
  NOR2_X1    g30396(.A1(new_n7240_), .A2(new_n32626_), .ZN(new_n33680_));
  INV_X1     g30397(.I(new_n33680_), .ZN(new_n33681_));
  NAND2_X1   g30398(.A1(new_n33681_), .A2(new_n2726_), .ZN(new_n33682_));
  AOI21_X1   g30399(.A1(new_n33646_), .A2(pi1153), .B(new_n33643_), .ZN(new_n33683_));
  NAND4_X1   g30400(.A1(new_n33679_), .A2(new_n10256_), .A3(new_n33682_), .A4(new_n33683_), .ZN(new_n33684_));
  NOR3_X1    g30401(.A1(new_n30765_), .A2(new_n8684_), .A3(new_n30660_), .ZN(new_n33685_));
  XOR2_X1    g30402(.A1(new_n33685_), .A2(new_n9260_), .Z(new_n33686_));
  NAND2_X1   g30403(.A1(po1038), .A2(pi1091), .ZN(new_n33687_));
  NOR3_X1    g30404(.A1(new_n30666_), .A2(new_n30588_), .A3(new_n30619_), .ZN(new_n33688_));
  INV_X1     g30405(.I(new_n33688_), .ZN(new_n33689_));
  NOR3_X1    g30406(.A1(new_n33687_), .A2(new_n13614_), .A3(new_n33689_), .ZN(new_n33690_));
  NOR2_X1    g30407(.A1(new_n8684_), .A2(new_n2726_), .ZN(new_n33691_));
  OAI21_X1   g30408(.A1(new_n33691_), .A2(pi0219), .B(pi1153), .ZN(new_n33692_));
  AOI21_X1   g30409(.A1(new_n7240_), .A2(new_n33692_), .B(new_n33643_), .ZN(new_n33693_));
  AOI21_X1   g30410(.A1(new_n33690_), .A2(new_n33693_), .B(pi1151), .ZN(new_n33694_));
  NOR3_X1    g30411(.A1(new_n33684_), .A2(new_n33686_), .A3(new_n33694_), .ZN(new_n33695_));
  OAI21_X1   g30412(.A1(new_n33695_), .A2(pi0219), .B(new_n33674_), .ZN(new_n33696_));
  OAI21_X1   g30413(.A1(new_n33673_), .A2(new_n33696_), .B(pi0230), .ZN(new_n33697_));
  INV_X1     g30414(.I(new_n32576_), .ZN(new_n33698_));
  NOR2_X1    g30415(.A1(new_n33698_), .A2(new_n32559_), .ZN(new_n33699_));
  NAND2_X1   g30416(.A1(new_n33699_), .A2(new_n8684_), .ZN(new_n33700_));
  INV_X1     g30417(.I(new_n33700_), .ZN(new_n33701_));
  NOR2_X1    g30418(.A1(new_n33701_), .A2(new_n32583_), .ZN(new_n33702_));
  INV_X1     g30419(.I(new_n33702_), .ZN(new_n33703_));
  AOI21_X1   g30420(.A1(new_n33703_), .A2(pi1153), .B(new_n32568_), .ZN(new_n33704_));
  INV_X1     g30421(.I(new_n32659_), .ZN(new_n33705_));
  NOR3_X1    g30422(.A1(new_n33705_), .A2(new_n8683_), .A3(new_n13614_), .ZN(new_n33706_));
  NOR3_X1    g30423(.A1(new_n32659_), .A2(pi0219), .A3(new_n13614_), .ZN(new_n33707_));
  OAI21_X1   g30424(.A1(new_n33706_), .A2(new_n33707_), .B(new_n32686_), .ZN(new_n33708_));
  INV_X1     g30425(.I(new_n33708_), .ZN(new_n33709_));
  NOR2_X1    g30426(.A1(new_n32552_), .A2(pi0219), .ZN(new_n33710_));
  NAND2_X1   g30427(.A1(new_n33700_), .A2(new_n32653_), .ZN(new_n33711_));
  NAND2_X1   g30428(.A1(new_n33711_), .A2(new_n33710_), .ZN(new_n33712_));
  INV_X1     g30429(.I(new_n33712_), .ZN(new_n33713_));
  NAND2_X1   g30430(.A1(new_n33713_), .A2(new_n32559_), .ZN(new_n33714_));
  OAI21_X1   g30431(.A1(new_n33714_), .A2(new_n33709_), .B(new_n8683_), .ZN(new_n33715_));
  AOI21_X1   g30432(.A1(new_n33715_), .A2(new_n33704_), .B(new_n32626_), .ZN(new_n33716_));
  XOR2_X1    g30433(.A1(new_n33716_), .A2(new_n33680_), .Z(new_n33717_));
  NOR2_X1    g30434(.A1(new_n8683_), .A2(new_n13614_), .ZN(new_n33718_));
  NOR2_X1    g30435(.A1(new_n32580_), .A2(new_n32598_), .ZN(new_n33719_));
  INV_X1     g30436(.I(new_n33719_), .ZN(new_n33720_));
  AOI21_X1   g30437(.A1(new_n8684_), .A2(new_n32539_), .B(new_n33720_), .ZN(new_n33721_));
  INV_X1     g30438(.I(new_n33721_), .ZN(new_n33722_));
  NOR3_X1    g30439(.A1(new_n33722_), .A2(new_n32588_), .A3(new_n32605_), .ZN(new_n33723_));
  NOR2_X1    g30440(.A1(new_n33723_), .A2(new_n32639_), .ZN(new_n33724_));
  NOR2_X1    g30441(.A1(new_n33724_), .A2(new_n8683_), .ZN(new_n33725_));
  XOR2_X1    g30442(.A1(new_n33725_), .A2(new_n33718_), .Z(new_n33726_));
  INV_X1     g30443(.I(new_n33710_), .ZN(new_n33727_));
  NOR2_X1    g30444(.A1(new_n33722_), .A2(new_n33727_), .ZN(new_n33728_));
  NAND3_X1   g30445(.A1(new_n33726_), .A2(new_n32616_), .A3(new_n33728_), .ZN(new_n33729_));
  INV_X1     g30446(.I(new_n33704_), .ZN(new_n33730_));
  NOR2_X1    g30447(.A1(new_n33723_), .A2(new_n32634_), .ZN(new_n33731_));
  NOR2_X1    g30448(.A1(new_n33731_), .A2(new_n33680_), .ZN(new_n33732_));
  NOR2_X1    g30449(.A1(new_n32678_), .A2(pi1153), .ZN(new_n33733_));
  NAND2_X1   g30450(.A1(new_n32587_), .A2(new_n8683_), .ZN(new_n33736_));
  NOR2_X1    g30451(.A1(new_n32603_), .A2(new_n32598_), .ZN(new_n33737_));
  NAND2_X1   g30452(.A1(new_n33737_), .A2(new_n8683_), .ZN(new_n33738_));
  NOR2_X1    g30453(.A1(new_n32565_), .A2(new_n33640_), .ZN(new_n33739_));
  AOI21_X1   g30454(.A1(new_n33727_), .A2(new_n33739_), .B(new_n7240_), .ZN(new_n33740_));
  XOR2_X1    g30455(.A1(new_n33740_), .A2(new_n33680_), .Z(new_n33741_));
  NOR2_X1    g30456(.A1(new_n32548_), .A2(new_n8683_), .ZN(new_n33742_));
  XOR2_X1    g30457(.A1(new_n33742_), .A2(new_n31936_), .Z(new_n33743_));
  NAND2_X1   g30458(.A1(new_n33743_), .A2(new_n32565_), .ZN(new_n33744_));
  NOR2_X1    g30459(.A1(new_n32538_), .A2(pi0219), .ZN(new_n33745_));
  INV_X1     g30460(.I(new_n33745_), .ZN(new_n33746_));
  NAND4_X1   g30461(.A1(new_n33741_), .A2(new_n33641_), .A3(new_n33744_), .A4(new_n33746_), .ZN(new_n33747_));
  NAND2_X1   g30462(.A1(new_n33747_), .A2(new_n31670_), .ZN(new_n33748_));
  OAI21_X1   g30463(.A1(new_n32568_), .A2(pi1091), .B(new_n13614_), .ZN(new_n33749_));
  NAND4_X1   g30464(.A1(new_n33749_), .A2(new_n33738_), .A3(new_n33748_), .A4(new_n33736_), .ZN(new_n33750_));
  NOR3_X1    g30465(.A1(new_n33730_), .A2(new_n33732_), .A3(new_n33750_), .ZN(new_n33751_));
  INV_X1     g30466(.I(new_n32538_), .ZN(new_n33752_));
  AOI21_X1   g30467(.A1(new_n8684_), .A2(new_n33752_), .B(new_n33727_), .ZN(new_n33753_));
  NOR2_X1    g30468(.A1(new_n33753_), .A2(pi0219), .ZN(new_n33754_));
  NOR2_X1    g30469(.A1(new_n32548_), .A2(new_n7240_), .ZN(new_n33755_));
  AOI21_X1   g30470(.A1(new_n33754_), .A2(new_n33755_), .B(new_n31670_), .ZN(new_n33756_));
  NAND2_X1   g30471(.A1(new_n33747_), .A2(new_n33756_), .ZN(new_n33757_));
  NOR3_X1    g30472(.A1(new_n33757_), .A2(new_n32600_), .A3(new_n32773_), .ZN(new_n33758_));
  OAI21_X1   g30473(.A1(new_n33751_), .A2(pi1152), .B(new_n33758_), .ZN(new_n33759_));
  AOI21_X1   g30474(.A1(new_n33729_), .A2(new_n13614_), .B(new_n33759_), .ZN(new_n33760_));
  AOI21_X1   g30475(.A1(new_n33717_), .A2(new_n33760_), .B(pi1152), .ZN(new_n33761_));
  NOR2_X1    g30476(.A1(new_n33704_), .A2(new_n8683_), .ZN(new_n33762_));
  INV_X1     g30477(.I(new_n32580_), .ZN(new_n33763_));
  NOR2_X1    g30478(.A1(new_n33737_), .A2(pi1153), .ZN(new_n33764_));
  NOR3_X1    g30479(.A1(new_n33722_), .A2(new_n32582_), .A3(new_n33764_), .ZN(new_n33765_));
  INV_X1     g30480(.I(new_n33765_), .ZN(new_n33766_));
  NOR3_X1    g30481(.A1(new_n33766_), .A2(new_n8683_), .A3(new_n33763_), .ZN(new_n33767_));
  INV_X1     g30482(.I(new_n33767_), .ZN(new_n33768_));
  NAND2_X1   g30483(.A1(new_n33762_), .A2(new_n33768_), .ZN(new_n33769_));
  OAI21_X1   g30484(.A1(new_n8683_), .A2(new_n33704_), .B(new_n33767_), .ZN(new_n33770_));
  NAND3_X1   g30485(.A1(new_n33769_), .A2(pi0253), .A3(new_n33770_), .ZN(new_n33771_));
  XOR2_X1    g30486(.A1(new_n33771_), .A2(new_n33680_), .Z(new_n33772_));
  INV_X1     g30487(.I(new_n33723_), .ZN(new_n33773_));
  NOR2_X1    g30488(.A1(new_n32590_), .A2(new_n8683_), .ZN(new_n33774_));
  NOR3_X1    g30489(.A1(new_n33774_), .A2(pi1153), .A3(new_n32634_), .ZN(new_n33775_));
  NOR2_X1    g30490(.A1(new_n33773_), .A2(new_n33775_), .ZN(new_n33776_));
  AOI21_X1   g30491(.A1(new_n33776_), .A2(new_n33713_), .B(new_n33764_), .ZN(new_n33777_));
  NOR4_X1    g30492(.A1(new_n33772_), .A2(new_n32668_), .A3(new_n33757_), .A4(new_n33777_), .ZN(new_n33778_));
  NOR3_X1    g30493(.A1(new_n33773_), .A2(new_n8683_), .A3(new_n13614_), .ZN(new_n33779_));
  NOR3_X1    g30494(.A1(new_n33723_), .A2(new_n8683_), .A3(pi1153), .ZN(new_n33780_));
  OAI21_X1   g30495(.A1(new_n33779_), .A2(new_n33780_), .B(new_n32576_), .ZN(new_n33781_));
  NAND2_X1   g30496(.A1(new_n33708_), .A2(new_n32626_), .ZN(new_n33782_));
  NOR2_X1    g30497(.A1(new_n33730_), .A2(new_n31349_), .ZN(new_n33783_));
  AOI22_X1   g30498(.A1(new_n33783_), .A2(new_n33782_), .B1(new_n33781_), .B2(pi0253), .ZN(new_n33784_));
  AOI21_X1   g30499(.A1(new_n32652_), .A2(new_n32599_), .B(new_n13614_), .ZN(new_n33785_));
  INV_X1     g30500(.I(new_n33785_), .ZN(new_n33786_));
  NAND2_X1   g30501(.A1(new_n33786_), .A2(new_n8683_), .ZN(new_n33787_));
  NAND4_X1   g30502(.A1(new_n33787_), .A2(pi1151), .A3(pi1153), .A4(new_n32687_), .ZN(new_n33788_));
  OAI21_X1   g30503(.A1(new_n33784_), .A2(new_n33788_), .B(new_n33747_), .ZN(new_n33789_));
  INV_X1     g30504(.I(new_n9261_), .ZN(new_n33790_));
  NOR3_X1    g30505(.A1(new_n30619_), .A2(new_n31670_), .A3(new_n9208_), .ZN(new_n33791_));
  AOI21_X1   g30506(.A1(po1038), .A2(new_n33791_), .B(pi1153), .ZN(new_n33792_));
  NOR2_X1    g30507(.A1(new_n30656_), .A2(pi1151), .ZN(new_n33793_));
  NOR4_X1    g30508(.A1(new_n33793_), .A2(new_n33790_), .A3(new_n33646_), .A4(new_n33792_), .ZN(new_n33794_));
  OAI21_X1   g30509(.A1(new_n33794_), .A2(new_n30615_), .B(new_n31578_), .ZN(new_n33795_));
  NAND2_X1   g30510(.A1(new_n33795_), .A2(pi1152), .ZN(new_n33796_));
  NAND4_X1   g30511(.A1(po1038), .A2(pi1151), .A3(new_n9259_), .A4(new_n31303_), .ZN(new_n33800_));
  NAND2_X1   g30512(.A1(new_n33800_), .A2(new_n13614_), .ZN(new_n33801_));
  NOR4_X1    g30513(.A1(new_n7240_), .A2(new_n33689_), .A3(new_n8684_), .A4(new_n8683_), .ZN(new_n33802_));
  NOR2_X1    g30514(.A1(new_n33689_), .A2(new_n8683_), .ZN(new_n33803_));
  NOR3_X1    g30515(.A1(new_n33803_), .A2(pi0211), .A3(new_n7240_), .ZN(new_n33804_));
  NOR2_X1    g30516(.A1(new_n33804_), .A2(new_n33802_), .ZN(new_n33805_));
  INV_X1     g30517(.I(new_n33805_), .ZN(new_n33806_));
  NAND2_X1   g30518(.A1(new_n30980_), .A2(pi1151), .ZN(new_n33807_));
  NAND2_X1   g30519(.A1(new_n30615_), .A2(new_n13614_), .ZN(new_n33808_));
  XOR2_X1    g30520(.A1(new_n33807_), .A2(new_n33808_), .Z(new_n33809_));
  NAND4_X1   g30521(.A1(new_n33806_), .A2(new_n31108_), .A3(new_n33801_), .A4(new_n33809_), .ZN(new_n33810_));
  XNOR2_X1   g30522(.A1(new_n33796_), .A2(new_n33810_), .ZN(new_n33811_));
  AOI21_X1   g30523(.A1(new_n8684_), .A2(new_n32574_), .B(new_n33746_), .ZN(new_n33812_));
  NOR3_X1    g30524(.A1(new_n32574_), .A2(new_n8683_), .A3(new_n7240_), .ZN(new_n33813_));
  INV_X1     g30525(.I(new_n33813_), .ZN(new_n33814_));
  NOR4_X1    g30526(.A1(new_n33811_), .A2(new_n30557_), .A3(new_n32574_), .A4(new_n33814_), .ZN(new_n33815_));
  OAI21_X1   g30527(.A1(new_n33778_), .A2(new_n33789_), .B(new_n33815_), .ZN(new_n33816_));
  NOR2_X1    g30528(.A1(new_n33816_), .A2(new_n33761_), .ZN(new_n33817_));
  XNOR2_X1   g30529(.A1(new_n33817_), .A2(new_n33697_), .ZN(po0410));
  NOR2_X1    g30530(.A1(new_n13817_), .A2(pi0200), .ZN(new_n33819_));
  NOR3_X1    g30531(.A1(new_n30698_), .A2(new_n8683_), .A3(new_n33819_), .ZN(new_n33820_));
  OAI21_X1   g30532(.A1(new_n33820_), .A2(new_n30947_), .B(new_n10253_), .ZN(new_n33821_));
  INV_X1     g30533(.I(new_n33821_), .ZN(new_n33822_));
  NOR3_X1    g30534(.A1(new_n33822_), .A2(pi0219), .A3(new_n30970_), .ZN(new_n33823_));
  NAND2_X1   g30535(.A1(new_n33646_), .A2(pi1154), .ZN(new_n33824_));
  OAI21_X1   g30536(.A1(new_n33823_), .A2(new_n33824_), .B(pi0254), .ZN(new_n33825_));
  OAI21_X1   g30537(.A1(new_n32737_), .A2(new_n13614_), .B(new_n13817_), .ZN(new_n33826_));
  NAND2_X1   g30538(.A1(new_n33676_), .A2(new_n33826_), .ZN(new_n33827_));
  NOR2_X1    g30539(.A1(new_n31683_), .A2(new_n8684_), .ZN(new_n33828_));
  NAND2_X1   g30540(.A1(new_n33650_), .A2(pi1154), .ZN(new_n33829_));
  OAI21_X1   g30541(.A1(new_n30724_), .A2(new_n30947_), .B(new_n30994_), .ZN(new_n33830_));
  AOI21_X1   g30542(.A1(new_n33830_), .A2(new_n31026_), .B(new_n30971_), .ZN(new_n33831_));
  INV_X1     g30543(.I(new_n33831_), .ZN(new_n33832_));
  OAI21_X1   g30544(.A1(new_n33832_), .A2(new_n33829_), .B(new_n2726_), .ZN(new_n33833_));
  AOI22_X1   g30545(.A1(new_n33833_), .A2(pi0219), .B1(new_n33827_), .B2(new_n33828_), .ZN(new_n33834_));
  NAND4_X1   g30546(.A1(new_n30994_), .A2(new_n30735_), .A3(pi0254), .A4(pi1091), .ZN(new_n33835_));
  NOR3_X1    g30547(.A1(new_n33834_), .A2(new_n31644_), .A3(new_n33835_), .ZN(new_n33836_));
  XNOR2_X1   g30548(.A1(new_n33836_), .A2(new_n33825_), .ZN(new_n33837_));
  NOR2_X1    g30549(.A1(new_n31937_), .A2(new_n13614_), .ZN(new_n33838_));
  NAND2_X1   g30550(.A1(new_n30615_), .A2(new_n13817_), .ZN(new_n33839_));
  XOR2_X1    g30551(.A1(new_n33838_), .A2(new_n33839_), .Z(new_n33840_));
  NAND2_X1   g30552(.A1(new_n33840_), .A2(po1038), .ZN(new_n33841_));
  XOR2_X1    g30553(.A1(new_n33841_), .A2(new_n33687_), .Z(new_n33842_));
  NAND2_X1   g30554(.A1(new_n33842_), .A2(pi0254), .ZN(new_n33843_));
  INV_X1     g30555(.I(new_n33843_), .ZN(new_n33844_));
  AOI21_X1   g30556(.A1(new_n8683_), .A2(new_n31002_), .B(new_n7240_), .ZN(new_n33845_));
  NAND2_X1   g30557(.A1(new_n33837_), .A2(new_n33845_), .ZN(new_n33846_));
  NAND2_X1   g30558(.A1(new_n30652_), .A2(pi1153), .ZN(new_n33847_));
  NAND3_X1   g30559(.A1(new_n32724_), .A2(pi1153), .A3(new_n32719_), .ZN(new_n33848_));
  XOR2_X1    g30560(.A1(new_n33848_), .A2(new_n33847_), .Z(new_n33849_));
  NOR3_X1    g30561(.A1(new_n32762_), .A2(new_n30652_), .A3(new_n33664_), .ZN(new_n33850_));
  NOR3_X1    g30562(.A1(new_n33850_), .A2(new_n13817_), .A3(new_n33656_), .ZN(new_n33851_));
  NOR2_X1    g30563(.A1(new_n33849_), .A2(new_n33851_), .ZN(new_n33852_));
  NOR2_X1    g30564(.A1(new_n30653_), .A2(new_n2726_), .ZN(new_n33853_));
  NAND2_X1   g30565(.A1(new_n33853_), .A2(pi1154), .ZN(new_n33854_));
  OAI22_X1   g30566(.A1(new_n33852_), .A2(new_n33854_), .B1(new_n2726_), .B2(new_n9259_), .ZN(new_n33855_));
  AOI21_X1   g30567(.A1(new_n33855_), .A2(new_n30934_), .B(new_n32627_), .ZN(new_n33856_));
  AOI21_X1   g30568(.A1(new_n31017_), .A2(pi1091), .B(new_n13817_), .ZN(new_n33857_));
  INV_X1     g30569(.I(new_n33857_), .ZN(new_n33858_));
  NAND2_X1   g30570(.A1(pi1091), .A2(pi1153), .ZN(new_n33859_));
  AOI21_X1   g30571(.A1(new_n30670_), .A2(pi1091), .B(new_n33859_), .ZN(new_n33860_));
  NOR3_X1    g30572(.A1(new_n30669_), .A2(new_n2726_), .A3(pi1153), .ZN(new_n33861_));
  OAI21_X1   g30573(.A1(new_n33860_), .A2(new_n33861_), .B(new_n32723_), .ZN(new_n33862_));
  AND2_X2    g30574(.A1(new_n33826_), .A2(pi0211), .Z(new_n33863_));
  NAND2_X1   g30575(.A1(new_n13614_), .A2(new_n13817_), .ZN(new_n33864_));
  OAI21_X1   g30576(.A1(new_n9258_), .A2(new_n33864_), .B(pi1091), .ZN(new_n33865_));
  NAND2_X1   g30577(.A1(new_n33865_), .A2(new_n8684_), .ZN(new_n33866_));
  AOI21_X1   g30578(.A1(new_n33862_), .A2(new_n33863_), .B(new_n33866_), .ZN(new_n33867_));
  NAND2_X1   g30579(.A1(new_n33865_), .A2(new_n8683_), .ZN(new_n33868_));
  NOR3_X1    g30580(.A1(new_n30637_), .A2(pi1091), .A3(pi1153), .ZN(new_n33869_));
  NOR4_X1    g30581(.A1(new_n31579_), .A2(new_n2726_), .A3(new_n30813_), .A4(new_n33869_), .ZN(new_n33870_));
  NAND3_X1   g30582(.A1(new_n33870_), .A2(new_n33857_), .A3(new_n33868_), .ZN(new_n33871_));
  OAI22_X1   g30583(.A1(new_n33867_), .A2(new_n33871_), .B1(new_n31937_), .B2(new_n33858_), .ZN(new_n33872_));
  NOR2_X1    g30584(.A1(new_n2726_), .A2(pi1154), .ZN(new_n33873_));
  INV_X1     g30585(.I(new_n33873_), .ZN(new_n33874_));
  NAND2_X1   g30586(.A1(new_n33849_), .A2(new_n9259_), .ZN(new_n33875_));
  NAND2_X1   g30587(.A1(new_n33875_), .A2(new_n33874_), .ZN(new_n33876_));
  NAND4_X1   g30588(.A1(new_n33872_), .A2(pi0254), .A3(new_n30750_), .A4(new_n33876_), .ZN(new_n33877_));
  XNOR2_X1   g30589(.A1(new_n33877_), .A2(new_n33856_), .ZN(new_n33878_));
  AOI21_X1   g30590(.A1(new_n33843_), .A2(new_n31002_), .B(new_n7240_), .ZN(new_n33879_));
  AOI21_X1   g30591(.A1(new_n33878_), .A2(new_n33879_), .B(new_n33639_), .ZN(new_n33880_));
  AOI21_X1   g30592(.A1(new_n33880_), .A2(new_n33846_), .B(new_n30557_), .ZN(new_n33881_));
  INV_X1     g30593(.I(new_n32582_), .ZN(new_n33882_));
  NAND2_X1   g30594(.A1(new_n33882_), .A2(new_n32616_), .ZN(new_n33883_));
  INV_X1     g30595(.I(new_n33883_), .ZN(new_n33884_));
  NAND2_X1   g30596(.A1(new_n33884_), .A2(new_n30637_), .ZN(new_n33885_));
  AOI21_X1   g30597(.A1(new_n33885_), .A2(new_n13614_), .B(new_n33698_), .ZN(new_n33886_));
  INV_X1     g30598(.I(new_n33886_), .ZN(new_n33887_));
  OAI21_X1   g30599(.A1(new_n32586_), .A2(new_n30995_), .B(new_n13614_), .ZN(new_n33888_));
  NOR3_X1    g30600(.A1(new_n32568_), .A2(pi1154), .A3(new_n32570_), .ZN(new_n33889_));
  NOR3_X1    g30601(.A1(new_n33889_), .A2(pi1153), .A3(new_n32619_), .ZN(new_n33890_));
  NAND4_X1   g30602(.A1(new_n33888_), .A2(pi0219), .A3(new_n33890_), .A4(new_n32576_), .ZN(new_n33891_));
  OAI21_X1   g30603(.A1(new_n33891_), .A2(new_n33887_), .B(pi0254), .ZN(new_n33892_));
  NAND3_X1   g30604(.A1(new_n33711_), .A2(pi1153), .A3(new_n32604_), .ZN(new_n33893_));
  NAND2_X1   g30605(.A1(new_n32603_), .A2(pi1154), .ZN(new_n33894_));
  AOI21_X1   g30606(.A1(new_n33893_), .A2(new_n8683_), .B(new_n33894_), .ZN(new_n33895_));
  INV_X1     g30607(.I(new_n32595_), .ZN(new_n33896_));
  INV_X1     g30608(.I(new_n32588_), .ZN(new_n33897_));
  NOR2_X1    g30609(.A1(new_n33897_), .A2(new_n13614_), .ZN(new_n33898_));
  OAI22_X1   g30610(.A1(pi1154), .A2(new_n33896_), .B1(new_n33898_), .B2(new_n32605_), .ZN(new_n33899_));
  AOI21_X1   g30611(.A1(new_n32636_), .A2(new_n30637_), .B(new_n8683_), .ZN(new_n33900_));
  NAND2_X1   g30612(.A1(new_n33899_), .A2(new_n33900_), .ZN(new_n33901_));
  AOI21_X1   g30613(.A1(new_n32539_), .A2(pi0211), .B(pi1154), .ZN(new_n33902_));
  INV_X1     g30614(.I(new_n32686_), .ZN(new_n33903_));
  NOR2_X1    g30615(.A1(new_n33903_), .A2(new_n32570_), .ZN(new_n33904_));
  INV_X1     g30616(.I(new_n33904_), .ZN(new_n33905_));
  NOR3_X1    g30617(.A1(new_n33905_), .A2(pi0219), .A3(new_n33733_), .ZN(new_n33906_));
  OAI21_X1   g30618(.A1(new_n33763_), .A2(new_n33902_), .B(new_n33906_), .ZN(new_n33907_));
  NAND2_X1   g30619(.A1(new_n33907_), .A2(new_n13817_), .ZN(new_n33908_));
  INV_X1     g30620(.I(new_n32687_), .ZN(new_n33909_));
  NOR2_X1    g30621(.A1(new_n33909_), .A2(new_n32559_), .ZN(new_n33910_));
  NAND4_X1   g30622(.A1(new_n33908_), .A2(pi0254), .A3(new_n33901_), .A4(new_n33910_), .ZN(new_n33911_));
  NOR2_X1    g30623(.A1(new_n33911_), .A2(new_n33895_), .ZN(new_n33912_));
  AOI21_X1   g30624(.A1(new_n33912_), .A2(new_n33892_), .B(new_n32626_), .ZN(new_n33913_));
  OAI21_X1   g30625(.A1(new_n33892_), .A2(new_n33912_), .B(new_n33913_), .ZN(new_n33914_));
  XOR2_X1    g30626(.A1(new_n33914_), .A2(new_n33681_), .Z(new_n33915_));
  NAND2_X1   g30627(.A1(new_n33915_), .A2(new_n33878_), .ZN(new_n33916_));
  NAND3_X1   g30628(.A1(new_n33916_), .A2(new_n31002_), .A3(new_n32773_), .ZN(new_n33917_));
  NOR2_X1    g30629(.A1(new_n33727_), .A2(new_n33812_), .ZN(new_n33918_));
  INV_X1     g30630(.I(new_n33918_), .ZN(new_n33919_));
  NOR2_X1    g30631(.A1(pi0254), .A2(pi1091), .ZN(new_n33920_));
  AOI21_X1   g30632(.A1(new_n9260_), .A2(new_n33920_), .B(new_n13614_), .ZN(new_n33921_));
  NOR2_X1    g30633(.A1(new_n32564_), .A2(new_n8684_), .ZN(new_n33922_));
  OAI21_X1   g30634(.A1(new_n32548_), .A2(pi0219), .B(new_n33922_), .ZN(new_n33923_));
  INV_X1     g30635(.I(new_n33923_), .ZN(new_n33924_));
  AOI21_X1   g30636(.A1(new_n8683_), .A2(new_n32538_), .B(new_n33924_), .ZN(new_n33925_));
  NOR2_X1    g30637(.A1(new_n30924_), .A2(new_n2726_), .ZN(new_n33926_));
  OAI21_X1   g30638(.A1(new_n33925_), .A2(new_n33921_), .B(new_n33926_), .ZN(new_n33927_));
  NAND2_X1   g30639(.A1(new_n33812_), .A2(new_n33926_), .ZN(new_n33928_));
  AOI21_X1   g30640(.A1(new_n33744_), .A2(new_n32627_), .B(new_n33928_), .ZN(new_n33929_));
  OAI21_X1   g30641(.A1(new_n33929_), .A2(pi1153), .B(pi1091), .ZN(new_n33930_));
  NOR3_X1    g30642(.A1(new_n33844_), .A2(new_n32626_), .A3(po1038), .ZN(new_n33931_));
  OAI21_X1   g30643(.A1(new_n33930_), .A2(new_n33754_), .B(new_n33931_), .ZN(new_n33932_));
  AOI21_X1   g30644(.A1(new_n33932_), .A2(new_n33927_), .B(new_n33919_), .ZN(new_n33933_));
  NOR2_X1    g30645(.A1(po1038), .A2(new_n33650_), .ZN(new_n33934_));
  AOI21_X1   g30646(.A1(new_n33843_), .A2(new_n33934_), .B(new_n8683_), .ZN(new_n33935_));
  NAND2_X1   g30647(.A1(new_n33927_), .A2(new_n32626_), .ZN(new_n33936_));
  AOI21_X1   g30648(.A1(new_n33681_), .A2(new_n33935_), .B(new_n33936_), .ZN(new_n33937_));
  OAI21_X1   g30649(.A1(new_n33937_), .A2(new_n33930_), .B(new_n31002_), .ZN(new_n33938_));
  AOI21_X1   g30650(.A1(new_n33917_), .A2(new_n33933_), .B(new_n33938_), .ZN(new_n33939_));
  INV_X1     g30651(.I(new_n32568_), .ZN(new_n33940_));
  NAND2_X1   g30652(.A1(new_n30995_), .A2(new_n32627_), .ZN(new_n33941_));
  AOI21_X1   g30653(.A1(new_n32583_), .A2(pi1153), .B(new_n33941_), .ZN(new_n33942_));
  NAND2_X1   g30654(.A1(new_n33890_), .A2(new_n32593_), .ZN(new_n33943_));
  OAI21_X1   g30655(.A1(new_n33943_), .A2(new_n33942_), .B(new_n33940_), .ZN(new_n33944_));
  NAND3_X1   g30656(.A1(new_n33886_), .A2(new_n32559_), .A3(new_n33944_), .ZN(new_n33945_));
  NAND2_X1   g30657(.A1(new_n33945_), .A2(new_n8555_), .ZN(new_n33946_));
  NOR2_X1    g30658(.A1(new_n32576_), .A2(new_n13614_), .ZN(new_n33947_));
  XOR2_X1    g30659(.A1(new_n33947_), .A2(new_n30928_), .Z(new_n33948_));
  NAND2_X1   g30660(.A1(new_n33948_), .A2(new_n32616_), .ZN(new_n33949_));
  NAND2_X1   g30661(.A1(new_n33949_), .A2(new_n32627_), .ZN(new_n33950_));
  AOI21_X1   g30662(.A1(new_n33946_), .A2(new_n32548_), .B(new_n33950_), .ZN(new_n33951_));
  OAI21_X1   g30663(.A1(new_n33773_), .A2(new_n13817_), .B(new_n32640_), .ZN(new_n33952_));
  NAND2_X1   g30664(.A1(new_n33952_), .A2(pi1153), .ZN(new_n33953_));
  OAI21_X1   g30665(.A1(new_n33951_), .A2(new_n33953_), .B(pi0253), .ZN(new_n33954_));
  NOR2_X1    g30666(.A1(new_n8683_), .A2(new_n32626_), .ZN(new_n33955_));
  XOR2_X1    g30667(.A1(new_n33954_), .A2(new_n33955_), .Z(new_n33956_));
  NAND2_X1   g30668(.A1(new_n32687_), .A2(pi1154), .ZN(new_n33957_));
  AOI21_X1   g30669(.A1(new_n33766_), .A2(new_n33957_), .B(new_n13614_), .ZN(new_n33958_));
  AOI21_X1   g30670(.A1(new_n33884_), .A2(pi1154), .B(new_n32686_), .ZN(new_n33959_));
  NAND2_X1   g30671(.A1(new_n32559_), .A2(pi1153), .ZN(new_n33960_));
  AOI21_X1   g30672(.A1(new_n33960_), .A2(new_n8684_), .B(new_n32597_), .ZN(new_n33961_));
  OAI21_X1   g30673(.A1(new_n33959_), .A2(new_n33961_), .B(new_n32627_), .ZN(new_n33962_));
  NOR4_X1    g30674(.A1(new_n33786_), .A2(new_n13817_), .A3(new_n32571_), .A4(new_n33722_), .ZN(new_n33963_));
  OAI21_X1   g30675(.A1(new_n33958_), .A2(new_n33962_), .B(new_n33963_), .ZN(new_n33964_));
  OAI21_X1   g30676(.A1(new_n33956_), .A2(new_n33964_), .B(new_n7240_), .ZN(new_n33965_));
  INV_X1     g30677(.I(new_n33840_), .ZN(new_n33966_));
  NAND4_X1   g30678(.A1(new_n30668_), .A2(new_n3098_), .A3(new_n31704_), .A4(new_n31936_), .ZN(new_n33967_));
  NAND2_X1   g30679(.A1(new_n33967_), .A2(new_n31523_), .ZN(new_n33968_));
  NAND2_X1   g30680(.A1(new_n30951_), .A2(new_n9259_), .ZN(new_n33969_));
  NAND2_X1   g30681(.A1(new_n33969_), .A2(new_n13817_), .ZN(new_n33970_));
  NAND3_X1   g30682(.A1(new_n33968_), .A2(new_n31045_), .A3(new_n33970_), .ZN(new_n33971_));
  NAND2_X1   g30683(.A1(new_n33971_), .A2(new_n13817_), .ZN(new_n33972_));
  AOI21_X1   g30684(.A1(new_n33972_), .A2(new_n30934_), .B(new_n7240_), .ZN(new_n33973_));
  XOR2_X1    g30685(.A1(new_n33973_), .A2(new_n31108_), .Z(new_n33974_));
  NAND2_X1   g30686(.A1(new_n33974_), .A2(new_n33966_), .ZN(new_n33975_));
  AOI21_X1   g30687(.A1(new_n33821_), .A2(new_n7240_), .B(new_n8683_), .ZN(new_n33976_));
  AOI21_X1   g30688(.A1(new_n33831_), .A2(new_n33976_), .B(pi1152), .ZN(new_n33977_));
  OAI21_X1   g30689(.A1(new_n7240_), .A2(new_n30923_), .B(new_n32330_), .ZN(new_n33978_));
  NAND4_X1   g30690(.A1(new_n33837_), .A2(pi0230), .A3(new_n33955_), .A4(new_n33978_), .ZN(new_n33979_));
  AOI21_X1   g30691(.A1(new_n33975_), .A2(new_n33977_), .B(new_n33979_), .ZN(new_n33980_));
  NAND2_X1   g30692(.A1(new_n33965_), .A2(new_n33980_), .ZN(new_n33981_));
  NOR2_X1    g30693(.A1(new_n33939_), .A2(new_n33981_), .ZN(new_n33982_));
  XOR2_X1    g30694(.A1(new_n33982_), .A2(new_n33881_), .Z(po0411));
  NAND2_X1   g30695(.A1(new_n33605_), .A2(pi0255), .ZN(new_n33984_));
  INV_X1     g30696(.I(pi1036), .ZN(new_n33985_));
  NOR2_X1    g30697(.A1(pi0200), .A2(pi1049), .ZN(new_n33986_));
  AOI21_X1   g30698(.A1(pi0200), .A2(new_n33985_), .B(new_n33986_), .ZN(new_n33987_));
  NAND2_X1   g30699(.A1(new_n33604_), .A2(new_n33987_), .ZN(new_n33988_));
  NAND2_X1   g30700(.A1(new_n33984_), .A2(new_n33988_), .ZN(po0412));
  NAND2_X1   g30701(.A1(new_n33605_), .A2(pi0256), .ZN(new_n33990_));
  INV_X1     g30702(.I(pi1070), .ZN(new_n33991_));
  NOR2_X1    g30703(.A1(pi0200), .A2(pi1048), .ZN(new_n33992_));
  AOI21_X1   g30704(.A1(pi0200), .A2(new_n33991_), .B(new_n33992_), .ZN(new_n33993_));
  NAND2_X1   g30705(.A1(new_n33604_), .A2(new_n33993_), .ZN(new_n33994_));
  NAND2_X1   g30706(.A1(new_n33990_), .A2(new_n33994_), .ZN(po0413));
  NAND2_X1   g30707(.A1(new_n33605_), .A2(pi0257), .ZN(new_n33996_));
  INV_X1     g30708(.I(pi1065), .ZN(new_n33997_));
  NOR2_X1    g30709(.A1(pi0200), .A2(pi1084), .ZN(new_n33998_));
  AOI21_X1   g30710(.A1(pi0200), .A2(new_n33997_), .B(new_n33998_), .ZN(new_n33999_));
  NAND2_X1   g30711(.A1(new_n33604_), .A2(new_n33999_), .ZN(new_n34000_));
  NAND2_X1   g30712(.A1(new_n33996_), .A2(new_n34000_), .ZN(po0414));
  INV_X1     g30713(.I(pi0258), .ZN(new_n34002_));
  INV_X1     g30714(.I(pi1062), .ZN(new_n34003_));
  NOR2_X1    g30715(.A1(pi0200), .A2(pi1072), .ZN(new_n34004_));
  AOI21_X1   g30716(.A1(pi0200), .A2(new_n34003_), .B(new_n34004_), .ZN(new_n34005_));
  NAND2_X1   g30717(.A1(new_n33604_), .A2(new_n34005_), .ZN(new_n34006_));
  OAI21_X1   g30718(.A1(new_n34002_), .A2(new_n33604_), .B(new_n34006_), .ZN(po0415));
  NAND2_X1   g30719(.A1(new_n33605_), .A2(pi0259), .ZN(new_n34008_));
  INV_X1     g30720(.I(pi1069), .ZN(new_n34009_));
  NAND2_X1   g30721(.A1(new_n34009_), .A2(pi0200), .ZN(new_n34010_));
  OAI21_X1   g30722(.A1(pi0200), .A2(pi1059), .B(new_n34010_), .ZN(new_n34011_));
  OAI21_X1   g30723(.A1(new_n33605_), .A2(new_n34011_), .B(new_n34008_), .ZN(po0416));
  NAND2_X1   g30724(.A1(new_n33605_), .A2(pi0260), .ZN(new_n34013_));
  INV_X1     g30725(.I(pi1044), .ZN(new_n34014_));
  NAND3_X1   g30726(.A1(pi0199), .A2(pi0200), .A3(pi1067), .ZN(new_n34015_));
  INV_X1     g30727(.I(pi1067), .ZN(new_n34016_));
  NAND3_X1   g30728(.A1(new_n8549_), .A2(new_n34016_), .A3(pi0200), .ZN(new_n34017_));
  AOI21_X1   g30729(.A1(new_n34017_), .A2(new_n34015_), .B(new_n34014_), .ZN(new_n34018_));
  OAI21_X1   g30730(.A1(new_n33605_), .A2(new_n34018_), .B(new_n34013_), .ZN(po0417));
  NAND2_X1   g30731(.A1(new_n33605_), .A2(pi0261), .ZN(new_n34020_));
  INV_X1     g30732(.I(pi1037), .ZN(new_n34021_));
  NAND3_X1   g30733(.A1(pi0199), .A2(pi0200), .A3(pi1040), .ZN(new_n34022_));
  INV_X1     g30734(.I(pi1040), .ZN(new_n34023_));
  NAND3_X1   g30735(.A1(new_n8549_), .A2(new_n34023_), .A3(pi0200), .ZN(new_n34024_));
  AOI21_X1   g30736(.A1(new_n34024_), .A2(new_n34022_), .B(new_n34021_), .ZN(new_n34025_));
  OAI21_X1   g30737(.A1(new_n33605_), .A2(new_n34025_), .B(new_n34020_), .ZN(po0418));
  INV_X1     g30738(.I(pi0123), .ZN(new_n34027_));
  NOR2_X1    g30739(.A1(new_n2984_), .A2(pi0228), .ZN(new_n34028_));
  AOI21_X1   g30740(.A1(new_n34027_), .A2(pi0228), .B(new_n34028_), .ZN(new_n34029_));
  INV_X1     g30741(.I(new_n34029_), .ZN(new_n34030_));
  NOR2_X1    g30742(.A1(new_n34030_), .A2(pi0262), .ZN(new_n34031_));
  INV_X1     g30743(.I(new_n34031_), .ZN(new_n34032_));
  NAND3_X1   g30744(.A1(new_n34032_), .A2(new_n32350_), .A3(new_n30568_), .ZN(new_n34033_));
  NOR2_X1    g30745(.A1(new_n34029_), .A2(new_n8545_), .ZN(new_n34034_));
  OAI21_X1   g30746(.A1(new_n34032_), .A2(pi0208), .B(new_n34034_), .ZN(new_n34035_));
  AOI21_X1   g30747(.A1(new_n34033_), .A2(new_n8549_), .B(new_n34035_), .ZN(new_n34036_));
  NOR3_X1    g30748(.A1(new_n3005_), .A2(new_n3811_), .A3(new_n2984_), .ZN(new_n34037_));
  NOR3_X1    g30749(.A1(new_n2984_), .A2(pi0228), .A3(pi0262), .ZN(new_n34038_));
  OAI21_X1   g30750(.A1(new_n34037_), .A2(new_n34038_), .B(pi1142), .ZN(new_n34039_));
  NOR3_X1    g30751(.A1(new_n34027_), .A2(new_n3005_), .A3(new_n3811_), .ZN(new_n34040_));
  NOR3_X1    g30752(.A1(new_n3005_), .A2(pi0123), .A3(pi0262), .ZN(new_n34041_));
  OAI21_X1   g30753(.A1(new_n34040_), .A2(new_n34041_), .B(pi1142), .ZN(new_n34042_));
  NAND2_X1   g30754(.A1(new_n34039_), .A2(new_n34042_), .ZN(new_n34043_));
  NAND2_X1   g30755(.A1(new_n31741_), .A2(new_n34030_), .ZN(new_n34044_));
  AOI21_X1   g30756(.A1(new_n7240_), .A2(new_n34043_), .B(new_n34044_), .ZN(new_n34045_));
  NOR2_X1    g30757(.A1(new_n32350_), .A2(new_n34043_), .ZN(new_n34046_));
  NOR4_X1    g30758(.A1(new_n34036_), .A2(po1038), .A3(new_n34045_), .A4(new_n34046_), .ZN(new_n34047_));
  AOI21_X1   g30759(.A1(new_n34039_), .A2(new_n34042_), .B(pi0299), .ZN(new_n34048_));
  NAND3_X1   g30760(.A1(new_n34030_), .A2(new_n8549_), .A3(new_n31640_), .ZN(new_n34049_));
  OAI21_X1   g30761(.A1(new_n34049_), .A2(new_n34048_), .B(new_n8546_), .ZN(new_n34050_));
  NAND4_X1   g30762(.A1(new_n34050_), .A2(pi0299), .A3(new_n31740_), .A4(new_n34032_), .ZN(new_n34051_));
  NOR2_X1    g30763(.A1(new_n34047_), .A2(new_n34051_), .ZN(po0419));
  AOI21_X1   g30764(.A1(new_n33909_), .A2(pi1155), .B(new_n13817_), .ZN(new_n34053_));
  NAND2_X1   g30765(.A1(new_n34053_), .A2(new_n32669_), .ZN(new_n34054_));
  NOR2_X1    g30766(.A1(new_n32605_), .A2(new_n32597_), .ZN(new_n34055_));
  INV_X1     g30767(.I(new_n34055_), .ZN(new_n34056_));
  AOI21_X1   g30768(.A1(new_n32667_), .A2(pi1155), .B(pi1154), .ZN(new_n34057_));
  AOI21_X1   g30769(.A1(new_n34057_), .A2(new_n34056_), .B(new_n13969_), .ZN(new_n34058_));
  NAND2_X1   g30770(.A1(new_n32605_), .A2(new_n13817_), .ZN(new_n34059_));
  NAND3_X1   g30771(.A1(new_n34059_), .A2(new_n32589_), .A3(pi1155), .ZN(new_n34060_));
  OAI21_X1   g30772(.A1(new_n34060_), .A2(new_n34054_), .B(new_n8555_), .ZN(new_n34061_));
  NAND3_X1   g30773(.A1(new_n34061_), .A2(new_n34058_), .A3(new_n32534_), .ZN(new_n34062_));
  NOR2_X1    g30774(.A1(new_n32568_), .A2(pi1091), .ZN(new_n34063_));
  AOI21_X1   g30775(.A1(new_n32590_), .A2(pi1155), .B(new_n30769_), .ZN(new_n34064_));
  NOR3_X1    g30776(.A1(new_n32589_), .A2(pi1154), .A3(new_n13778_), .ZN(new_n34065_));
  OAI21_X1   g30777(.A1(new_n34064_), .A2(new_n34065_), .B(new_n34063_), .ZN(new_n34066_));
  NOR3_X1    g30778(.A1(new_n32653_), .A2(new_n13817_), .A3(new_n13778_), .ZN(new_n34067_));
  OAI21_X1   g30779(.A1(pi1156), .A2(new_n34067_), .B(new_n34066_), .ZN(new_n34068_));
  AOI21_X1   g30780(.A1(new_n34062_), .A2(new_n8684_), .B(new_n34068_), .ZN(new_n34069_));
  OAI21_X1   g30781(.A1(new_n34069_), .A2(new_n34054_), .B(new_n8683_), .ZN(new_n34070_));
  OR3_X2     g30782(.A1(new_n34067_), .A2(new_n8684_), .A3(pi1156), .Z(new_n34071_));
  NAND3_X1   g30783(.A1(new_n34058_), .A2(new_n32600_), .A3(new_n34053_), .ZN(new_n34072_));
  AOI21_X1   g30784(.A1(new_n34071_), .A2(new_n33720_), .B(new_n34072_), .ZN(new_n34073_));
  INV_X1     g30785(.I(pi0263), .ZN(new_n34074_));
  NAND2_X1   g30786(.A1(new_n32631_), .A2(new_n34074_), .ZN(new_n34075_));
  AOI21_X1   g30787(.A1(new_n34070_), .A2(new_n34073_), .B(new_n34075_), .ZN(new_n34076_));
  NOR2_X1    g30788(.A1(new_n33897_), .A2(new_n13778_), .ZN(new_n34077_));
  OAI21_X1   g30789(.A1(pi1154), .A2(new_n32616_), .B(new_n34077_), .ZN(new_n34078_));
  NAND2_X1   g30790(.A1(new_n34066_), .A2(new_n34078_), .ZN(new_n34079_));
  OAI21_X1   g30791(.A1(new_n34060_), .A2(new_n32774_), .B(new_n34078_), .ZN(new_n34080_));
  NAND2_X1   g30792(.A1(new_n32639_), .A2(new_n30625_), .ZN(new_n34081_));
  OAI21_X1   g30793(.A1(new_n34077_), .A2(new_n34081_), .B(new_n33940_), .ZN(new_n34082_));
  NOR2_X1    g30794(.A1(new_n8683_), .A2(pi1156), .ZN(new_n34083_));
  INV_X1     g30795(.I(new_n34083_), .ZN(new_n34084_));
  NOR3_X1    g30796(.A1(new_n32571_), .A2(new_n13817_), .A3(new_n34084_), .ZN(new_n34085_));
  NAND4_X1   g30797(.A1(new_n34079_), .A2(new_n34080_), .A3(new_n34082_), .A4(new_n34085_), .ZN(new_n34086_));
  NOR2_X1    g30798(.A1(new_n32583_), .A2(new_n33763_), .ZN(new_n34087_));
  AOI21_X1   g30799(.A1(pi1155), .A2(new_n32568_), .B(new_n32644_), .ZN(new_n34088_));
  NAND2_X1   g30800(.A1(new_n34088_), .A2(new_n32580_), .ZN(new_n34089_));
  XOR2_X1    g30801(.A1(new_n34087_), .A2(new_n34089_), .Z(new_n34090_));
  NOR3_X1    g30802(.A1(new_n34090_), .A2(new_n13817_), .A3(new_n32567_), .ZN(new_n34091_));
  NOR2_X1    g30803(.A1(new_n34090_), .A2(new_n13817_), .ZN(new_n34092_));
  NOR2_X1    g30804(.A1(new_n34092_), .A2(new_n32774_), .ZN(new_n34093_));
  OAI22_X1   g30805(.A1(new_n34093_), .A2(new_n8683_), .B1(pi1156), .B2(new_n34091_), .ZN(new_n34094_));
  NOR2_X1    g30806(.A1(new_n33699_), .A2(new_n13778_), .ZN(new_n34095_));
  XOR2_X1    g30807(.A1(new_n34095_), .A2(new_n30769_), .Z(new_n34096_));
  NOR2_X1    g30808(.A1(new_n34088_), .A2(new_n13817_), .ZN(new_n34097_));
  NOR4_X1    g30809(.A1(new_n34096_), .A2(new_n31401_), .A3(new_n33883_), .A4(new_n34097_), .ZN(new_n34098_));
  AOI21_X1   g30810(.A1(new_n34094_), .A2(new_n34098_), .B(pi0263), .ZN(new_n34099_));
  OAI21_X1   g30811(.A1(new_n34076_), .A2(new_n34086_), .B(new_n34099_), .ZN(new_n34100_));
  NOR2_X1    g30812(.A1(new_n32659_), .A2(new_n13817_), .ZN(new_n34101_));
  XOR2_X1    g30813(.A1(new_n34101_), .A2(new_n30769_), .Z(new_n34102_));
  NOR2_X1    g30814(.A1(new_n34102_), .A2(new_n32691_), .ZN(new_n34103_));
  NOR2_X1    g30815(.A1(new_n34103_), .A2(pi1156), .ZN(new_n34104_));
  NOR2_X1    g30816(.A1(new_n34104_), .A2(new_n33894_), .ZN(new_n34105_));
  INV_X1     g30817(.I(new_n33910_), .ZN(new_n34106_));
  OAI21_X1   g30818(.A1(new_n32662_), .A2(new_n32567_), .B(pi1155), .ZN(new_n34107_));
  XOR2_X1    g30819(.A1(new_n34107_), .A2(new_n30769_), .Z(new_n34108_));
  NAND3_X1   g30820(.A1(new_n34108_), .A2(new_n32678_), .A3(new_n34106_), .ZN(new_n34109_));
  NOR2_X1    g30821(.A1(new_n34103_), .A2(new_n13969_), .ZN(new_n34110_));
  AOI21_X1   g30822(.A1(new_n34110_), .A2(new_n34109_), .B(new_n30616_), .ZN(new_n34111_));
  AND3_X2    g30823(.A1(new_n34108_), .A2(pi0211), .A3(new_n32678_), .Z(new_n34112_));
  OAI21_X1   g30824(.A1(new_n34111_), .A2(new_n34105_), .B(new_n34112_), .ZN(new_n34113_));
  NOR2_X1    g30825(.A1(new_n33904_), .A2(new_n13778_), .ZN(new_n34114_));
  XOR2_X1    g30826(.A1(new_n34114_), .A2(new_n30768_), .Z(new_n34115_));
  NOR2_X1    g30827(.A1(new_n34106_), .A2(new_n32698_), .ZN(new_n34116_));
  NAND2_X1   g30828(.A1(new_n34106_), .A2(new_n13969_), .ZN(new_n34117_));
  AOI22_X1   g30829(.A1(new_n34105_), .A2(new_n34117_), .B1(new_n34115_), .B2(new_n34116_), .ZN(new_n34118_));
  OR2_X2     g30830(.A1(new_n34102_), .A2(new_n32696_), .Z(new_n34119_));
  AOI21_X1   g30831(.A1(new_n34118_), .A2(new_n34113_), .B(new_n34119_), .ZN(new_n34120_));
  AOI21_X1   g30832(.A1(new_n34100_), .A2(new_n34120_), .B(po1038), .ZN(new_n34121_));
  NAND2_X1   g30833(.A1(new_n31480_), .A2(new_n30927_), .ZN(new_n34122_));
  AOI21_X1   g30834(.A1(new_n34122_), .A2(new_n8555_), .B(new_n13778_), .ZN(new_n34123_));
  OAI21_X1   g30835(.A1(new_n34123_), .A2(pi0211), .B(new_n8683_), .ZN(new_n34124_));
  OAI21_X1   g30836(.A1(new_n30677_), .A2(new_n34084_), .B(new_n33874_), .ZN(new_n34125_));
  NOR2_X1    g30837(.A1(new_n30674_), .A2(new_n13817_), .ZN(new_n34126_));
  OAI21_X1   g30838(.A1(new_n34126_), .A2(pi1155), .B(pi0199), .ZN(new_n34127_));
  NOR2_X1    g30839(.A1(new_n31401_), .A2(new_n2726_), .ZN(new_n34128_));
  NAND4_X1   g30840(.A1(new_n34125_), .A2(new_n34127_), .A3(new_n32731_), .A4(new_n34128_), .ZN(new_n34129_));
  AOI21_X1   g30841(.A1(new_n13817_), .A2(new_n34129_), .B(new_n31502_), .ZN(new_n34130_));
  INV_X1     g30842(.I(new_n33853_), .ZN(new_n34131_));
  NOR2_X1    g30843(.A1(new_n31052_), .A2(new_n13778_), .ZN(new_n34132_));
  INV_X1     g30844(.I(new_n34132_), .ZN(new_n34133_));
  OAI22_X1   g30845(.A1(new_n34131_), .A2(new_n34133_), .B1(new_n13817_), .B2(new_n32760_), .ZN(new_n34134_));
  NAND2_X1   g30846(.A1(new_n33691_), .A2(new_n30659_), .ZN(new_n34135_));
  AOI21_X1   g30847(.A1(new_n34135_), .A2(new_n13817_), .B(new_n8549_), .ZN(new_n34136_));
  NAND2_X1   g30848(.A1(new_n34134_), .A2(new_n34136_), .ZN(new_n34137_));
  AOI21_X1   g30849(.A1(new_n30805_), .A2(pi0211), .B(new_n13969_), .ZN(new_n34138_));
  NAND2_X1   g30850(.A1(new_n34137_), .A2(new_n34138_), .ZN(new_n34139_));
  NOR2_X1    g30851(.A1(new_n8683_), .A2(new_n13969_), .ZN(new_n34140_));
  XOR2_X1    g30852(.A1(new_n34139_), .A2(new_n34140_), .Z(new_n34141_));
  NOR2_X1    g30853(.A1(new_n30677_), .A2(new_n30927_), .ZN(new_n34142_));
  NOR2_X1    g30854(.A1(new_n34142_), .A2(new_n8684_), .ZN(new_n34143_));
  INV_X1     g30855(.I(new_n33691_), .ZN(new_n34144_));
  OAI21_X1   g30856(.A1(new_n32731_), .A2(new_n33873_), .B(new_n31281_), .ZN(new_n34145_));
  NOR2_X1    g30857(.A1(new_n34145_), .A2(new_n34144_), .ZN(new_n34146_));
  XNOR2_X1   g30858(.A1(new_n34146_), .A2(new_n34143_), .ZN(new_n34147_));
  NOR3_X1    g30859(.A1(new_n34141_), .A2(new_n34074_), .A3(new_n34147_), .ZN(new_n34148_));
  NAND2_X1   g30860(.A1(new_n34134_), .A2(new_n30621_), .ZN(new_n34149_));
  AOI21_X1   g30861(.A1(new_n13817_), .A2(new_n30743_), .B(new_n30855_), .ZN(new_n34150_));
  NAND3_X1   g30862(.A1(new_n30855_), .A2(new_n13817_), .A3(new_n8774_), .ZN(new_n34151_));
  NAND3_X1   g30863(.A1(new_n34151_), .A2(new_n13969_), .A3(new_n31800_), .ZN(new_n34152_));
  INV_X1     g30864(.I(new_n10254_), .ZN(new_n34153_));
  NOR2_X1    g30865(.A1(pi0263), .A2(pi1091), .ZN(new_n34154_));
  NOR2_X1    g30866(.A1(new_n34153_), .A2(new_n34154_), .ZN(new_n34155_));
  NAND4_X1   g30867(.A1(new_n34152_), .A2(new_n34150_), .A3(new_n34142_), .A4(new_n34155_), .ZN(new_n34156_));
  AOI21_X1   g30868(.A1(new_n34149_), .A2(new_n2726_), .B(new_n34156_), .ZN(new_n34157_));
  OAI21_X1   g30869(.A1(new_n34148_), .A2(new_n34130_), .B(new_n34157_), .ZN(new_n34158_));
  NOR2_X1    g30870(.A1(new_n8775_), .A2(new_n13778_), .ZN(new_n34159_));
  OAI21_X1   g30871(.A1(new_n30671_), .A2(pi1154), .B(new_n34159_), .ZN(new_n34160_));
  OR3_X2     g30872(.A1(new_n30657_), .A2(new_n13817_), .A3(new_n30659_), .Z(new_n34161_));
  AOI21_X1   g30873(.A1(new_n34160_), .A2(new_n13969_), .B(new_n34161_), .ZN(new_n34162_));
  NOR2_X1    g30874(.A1(new_n34145_), .A2(new_n13969_), .ZN(new_n34163_));
  OAI21_X1   g30875(.A1(new_n34162_), .A2(pi0211), .B(new_n34163_), .ZN(new_n34164_));
  AOI21_X1   g30876(.A1(new_n34158_), .A2(new_n34124_), .B(new_n34164_), .ZN(new_n34165_));
  NAND2_X1   g30877(.A1(new_n34165_), .A2(new_n32630_), .ZN(new_n34166_));
  INV_X1     g30878(.I(new_n33744_), .ZN(new_n34167_));
  NOR2_X1    g30879(.A1(new_n34167_), .A2(pi0263), .ZN(new_n34168_));
  NAND2_X1   g30880(.A1(new_n33923_), .A2(new_n34074_), .ZN(new_n34169_));
  NOR2_X1    g30881(.A1(new_n8684_), .A2(pi1155), .ZN(new_n34170_));
  AOI21_X1   g30882(.A1(new_n8684_), .A2(new_n33873_), .B(new_n34170_), .ZN(new_n34171_));
  OAI21_X1   g30883(.A1(new_n33752_), .A2(new_n34171_), .B(new_n8684_), .ZN(new_n34172_));
  NAND3_X1   g30884(.A1(new_n31401_), .A2(pi0219), .A3(pi1091), .ZN(new_n34173_));
  NAND2_X1   g30885(.A1(new_n32631_), .A2(new_n34173_), .ZN(new_n34174_));
  NAND4_X1   g30886(.A1(new_n34174_), .A2(new_n13778_), .A3(new_n31936_), .A4(new_n33829_), .ZN(new_n34175_));
  NOR4_X1    g30887(.A1(new_n33746_), .A2(pi0211), .A3(new_n32574_), .A4(new_n34175_), .ZN(new_n34176_));
  NAND3_X1   g30888(.A1(new_n34176_), .A2(new_n34169_), .A3(new_n34172_), .ZN(new_n34177_));
  OAI21_X1   g30889(.A1(new_n34168_), .A2(new_n34177_), .B(new_n7240_), .ZN(new_n34178_));
  NOR2_X1    g30890(.A1(new_n30919_), .A2(new_n8683_), .ZN(new_n34179_));
  NAND3_X1   g30891(.A1(new_n30625_), .A2(new_n30637_), .A3(pi0219), .ZN(new_n34180_));
  XOR2_X1    g30892(.A1(new_n34180_), .A2(new_n34179_), .Z(new_n34181_));
  NOR2_X1    g30893(.A1(new_n34181_), .A2(new_n2726_), .ZN(new_n34182_));
  NOR2_X1    g30894(.A1(new_n34182_), .A2(new_n34154_), .ZN(new_n34183_));
  NOR2_X1    g30895(.A1(new_n34183_), .A2(new_n32631_), .ZN(new_n34184_));
  AOI21_X1   g30896(.A1(new_n34178_), .A2(new_n34184_), .B(new_n32773_), .ZN(new_n34185_));
  OAI21_X1   g30897(.A1(new_n34121_), .A2(new_n34166_), .B(new_n34185_), .ZN(new_n34186_));
  NOR4_X1    g30898(.A1(new_n31084_), .A2(new_n30685_), .A3(pi0299), .A4(new_n13969_), .ZN(new_n34187_));
  OAI21_X1   g30899(.A1(new_n34187_), .A2(new_n30681_), .B(new_n30678_), .ZN(new_n34188_));
  NAND2_X1   g30900(.A1(new_n34188_), .A2(new_n8683_), .ZN(new_n34189_));
  NOR2_X1    g30901(.A1(new_n31800_), .A2(new_n13969_), .ZN(new_n34190_));
  AOI21_X1   g30902(.A1(new_n34189_), .A2(new_n34190_), .B(po1038), .ZN(new_n34191_));
  AND2_X2    g30903(.A1(new_n34188_), .A2(new_n30611_), .Z(new_n34192_));
  NOR4_X1    g30904(.A1(new_n34124_), .A2(new_n8684_), .A3(new_n34191_), .A4(new_n34192_), .ZN(new_n34193_));
  NOR2_X1    g30905(.A1(new_n34181_), .A2(new_n7240_), .ZN(new_n34194_));
  AOI21_X1   g30906(.A1(new_n34193_), .A2(new_n34194_), .B(pi0230), .ZN(new_n34195_));
  NOR2_X1    g30907(.A1(new_n34165_), .A2(new_n7240_), .ZN(new_n34196_));
  XOR2_X1    g30908(.A1(new_n34196_), .A2(new_n32805_), .Z(new_n34197_));
  OAI21_X1   g30909(.A1(new_n34154_), .A2(new_n34182_), .B(new_n34197_), .ZN(new_n34198_));
  AOI21_X1   g30910(.A1(new_n34186_), .A2(new_n34195_), .B(new_n34198_), .ZN(po0420));
  INV_X1     g30911(.I(pi0796), .ZN(new_n34200_));
  NOR3_X1    g30912(.A1(new_n32530_), .A2(new_n34200_), .A3(new_n2726_), .ZN(new_n34201_));
  NOR3_X1    g30913(.A1(new_n32530_), .A2(pi0796), .A3(pi1091), .ZN(new_n34202_));
  OAI21_X1   g30914(.A1(new_n34201_), .A2(new_n34202_), .B(pi0264), .ZN(new_n34203_));
  NAND2_X1   g30915(.A1(pi1091), .A2(pi1142), .ZN(new_n34204_));
  NAND2_X1   g30916(.A1(new_n34203_), .A2(new_n34204_), .ZN(new_n34205_));
  NAND2_X1   g30917(.A1(pi1091), .A2(pi1141), .ZN(new_n34206_));
  NAND2_X1   g30918(.A1(new_n34203_), .A2(new_n34206_), .ZN(new_n34207_));
  NAND2_X1   g30919(.A1(new_n34207_), .A2(pi0200), .ZN(new_n34208_));
  XOR2_X1    g30920(.A1(new_n34208_), .A2(new_n30722_), .Z(new_n34209_));
  OAI21_X1   g30921(.A1(new_n34209_), .A2(new_n34205_), .B(new_n12655_), .ZN(new_n34210_));
  NOR3_X1    g30922(.A1(new_n32541_), .A2(new_n34200_), .A3(new_n2726_), .ZN(new_n34211_));
  NOR3_X1    g30923(.A1(new_n32541_), .A2(pi0796), .A3(pi1091), .ZN(new_n34212_));
  OAI21_X1   g30924(.A1(new_n34211_), .A2(new_n34212_), .B(pi0264), .ZN(new_n34213_));
  NOR2_X1    g30925(.A1(pi0199), .A2(pi1091), .ZN(new_n34214_));
  INV_X1     g30926(.I(new_n34214_), .ZN(new_n34215_));
  OAI21_X1   g30927(.A1(new_n34215_), .A2(pi1143), .B(pi0200), .ZN(new_n34216_));
  NOR2_X1    g30928(.A1(new_n34213_), .A2(new_n34216_), .ZN(new_n34217_));
  NAND2_X1   g30929(.A1(pi0200), .A2(pi1141), .ZN(new_n34218_));
  OAI21_X1   g30930(.A1(new_n31371_), .A2(new_n34218_), .B(new_n3814_), .ZN(new_n34219_));
  AOI21_X1   g30931(.A1(new_n34219_), .A2(pi0199), .B(new_n30557_), .ZN(new_n34220_));
  XOR2_X1    g30932(.A1(new_n34220_), .A2(new_n32800_), .Z(new_n34221_));
  NAND3_X1   g30933(.A1(pi0211), .A2(pi0219), .A3(pi1142), .ZN(new_n34222_));
  NAND3_X1   g30934(.A1(new_n8683_), .A2(new_n3814_), .A3(pi0211), .ZN(new_n34223_));
  AOI21_X1   g30935(.A1(new_n34223_), .A2(new_n34222_), .B(new_n3980_), .ZN(new_n34224_));
  NOR3_X1    g30936(.A1(new_n34224_), .A2(new_n30557_), .A3(new_n32828_), .ZN(new_n34225_));
  AOI22_X1   g30937(.A1(new_n34210_), .A2(new_n34217_), .B1(new_n34221_), .B2(new_n34225_), .ZN(new_n34226_));
  NAND2_X1   g30938(.A1(new_n34207_), .A2(pi0211), .ZN(new_n34227_));
  XOR2_X1    g30939(.A1(new_n34227_), .A2(new_n31936_), .Z(new_n34228_));
  OAI21_X1   g30940(.A1(new_n34228_), .A2(new_n34205_), .B(new_n12655_), .ZN(new_n34229_));
  NOR2_X1    g30941(.A1(new_n33650_), .A2(new_n8683_), .ZN(new_n34230_));
  NOR3_X1    g30942(.A1(new_n34213_), .A2(new_n32828_), .A3(new_n34230_), .ZN(new_n34231_));
  NAND2_X1   g30943(.A1(new_n34229_), .A2(new_n34231_), .ZN(new_n34232_));
  NOR2_X1    g30944(.A1(new_n34226_), .A2(new_n34232_), .ZN(po0421));
  XNOR2_X1   g30945(.A1(new_n31936_), .A2(new_n30558_), .ZN(new_n34234_));
  OAI21_X1   g30946(.A1(new_n34234_), .A2(new_n3814_), .B(new_n32520_), .ZN(new_n34235_));
  AOI21_X1   g30947(.A1(new_n12655_), .A2(new_n34235_), .B(new_n30557_), .ZN(new_n34236_));
  NAND2_X1   g30948(.A1(new_n32529_), .A2(pi1091), .ZN(new_n34237_));
  INV_X1     g30949(.I(pi0819), .ZN(new_n34238_));
  NAND2_X1   g30950(.A1(new_n32529_), .A2(new_n34238_), .ZN(new_n34239_));
  XOR2_X1    g30951(.A1(new_n34237_), .A2(new_n34239_), .Z(new_n34240_));
  NAND2_X1   g30952(.A1(new_n34240_), .A2(pi0265), .ZN(new_n34241_));
  NAND2_X1   g30953(.A1(new_n34241_), .A2(new_n34204_), .ZN(new_n34242_));
  NAND2_X1   g30954(.A1(new_n34242_), .A2(pi0211), .ZN(new_n34243_));
  XOR2_X1    g30955(.A1(new_n34243_), .A2(new_n31936_), .Z(new_n34244_));
  NAND2_X1   g30956(.A1(pi1091), .A2(pi1143), .ZN(new_n34245_));
  NAND2_X1   g30957(.A1(new_n34241_), .A2(new_n34245_), .ZN(new_n34246_));
  INV_X1     g30958(.I(pi0265), .ZN(new_n34247_));
  NAND3_X1   g30959(.A1(new_n32540_), .A2(pi0819), .A3(pi1091), .ZN(new_n34248_));
  NAND3_X1   g30960(.A1(new_n32540_), .A2(new_n34238_), .A3(new_n2726_), .ZN(new_n34249_));
  AOI21_X1   g30961(.A1(new_n34248_), .A2(new_n34249_), .B(new_n34247_), .ZN(new_n34250_));
  OAI21_X1   g30962(.A1(new_n34215_), .A2(pi1144), .B(pi0200), .ZN(new_n34251_));
  NOR2_X1    g30963(.A1(new_n34250_), .A2(new_n34251_), .ZN(new_n34252_));
  NOR4_X1    g30964(.A1(new_n34244_), .A2(new_n12655_), .A3(new_n34246_), .A4(new_n34252_), .ZN(new_n34253_));
  INV_X1     g30965(.I(new_n34230_), .ZN(new_n34254_));
  NAND2_X1   g30966(.A1(new_n34242_), .A2(pi0200), .ZN(new_n34255_));
  XOR2_X1    g30967(.A1(new_n34255_), .A2(new_n30722_), .Z(new_n34256_));
  AOI21_X1   g30968(.A1(new_n12654_), .A2(new_n34250_), .B(new_n32490_), .ZN(new_n34257_));
  NOR4_X1    g30969(.A1(new_n34256_), .A2(new_n34254_), .A3(new_n34246_), .A4(new_n34257_), .ZN(new_n34258_));
  NOR2_X1    g30970(.A1(new_n34253_), .A2(new_n34258_), .ZN(new_n34259_));
  NAND2_X1   g30971(.A1(new_n8549_), .A2(pi1142), .ZN(new_n34260_));
  AOI21_X1   g30972(.A1(new_n32459_), .A2(new_n34260_), .B(new_n30564_), .ZN(new_n34261_));
  NOR4_X1    g30973(.A1(new_n34259_), .A2(new_n30557_), .A3(new_n12655_), .A4(new_n34261_), .ZN(new_n34262_));
  XOR2_X1    g30974(.A1(new_n34262_), .A2(new_n34236_), .Z(po0422));
  NAND2_X1   g30975(.A1(new_n32540_), .A2(pi1091), .ZN(new_n34264_));
  INV_X1     g30976(.I(pi0948), .ZN(new_n34265_));
  NAND2_X1   g30977(.A1(new_n32540_), .A2(new_n34265_), .ZN(new_n34266_));
  XOR2_X1    g30978(.A1(new_n34264_), .A2(new_n34266_), .Z(new_n34267_));
  NAND2_X1   g30979(.A1(new_n34267_), .A2(pi0266), .ZN(new_n34268_));
  NAND2_X1   g30980(.A1(new_n34268_), .A2(pi0199), .ZN(new_n34269_));
  NAND3_X1   g30981(.A1(new_n32529_), .A2(pi0948), .A3(pi1091), .ZN(new_n34270_));
  NAND3_X1   g30982(.A1(new_n32529_), .A2(new_n34265_), .A3(new_n2726_), .ZN(new_n34271_));
  AOI21_X1   g30983(.A1(new_n34270_), .A2(new_n34271_), .B(new_n4786_), .ZN(new_n34272_));
  NAND4_X1   g30984(.A1(new_n34272_), .A2(pi0199), .A3(pi1091), .A4(pi1136), .ZN(new_n34273_));
  XNOR2_X1   g30985(.A1(new_n34269_), .A2(new_n34273_), .ZN(new_n34274_));
  OR2_X2     g30986(.A1(new_n34274_), .A2(new_n8555_), .Z(new_n34275_));
  AOI21_X1   g30987(.A1(new_n34275_), .A2(new_n2726_), .B(new_n8549_), .ZN(new_n34276_));
  NOR2_X1    g30988(.A1(new_n2726_), .A2(new_n4959_), .ZN(new_n34277_));
  OAI21_X1   g30989(.A1(new_n34272_), .A2(pi0199), .B(new_n34277_), .ZN(new_n34278_));
  AND2_X2    g30990(.A1(new_n34278_), .A2(new_n8555_), .Z(new_n34279_));
  NOR3_X1    g30991(.A1(new_n34279_), .A2(new_n8549_), .A3(new_n34268_), .ZN(new_n34280_));
  OAI21_X1   g30992(.A1(new_n34276_), .A2(new_n34280_), .B(new_n12654_), .ZN(new_n34281_));
  NOR2_X1    g30993(.A1(new_n34272_), .A2(pi0219), .ZN(new_n34282_));
  NAND2_X1   g30994(.A1(new_n34282_), .A2(pi1091), .ZN(new_n34283_));
  NAND2_X1   g30995(.A1(new_n34283_), .A2(new_n8684_), .ZN(new_n34284_));
  NAND2_X1   g30996(.A1(new_n8683_), .A2(new_n2726_), .ZN(new_n34285_));
  OAI21_X1   g30997(.A1(new_n34285_), .A2(pi1136), .B(pi0211), .ZN(new_n34286_));
  AOI21_X1   g30998(.A1(new_n34268_), .A2(new_n34286_), .B(new_n12654_), .ZN(new_n34287_));
  NAND3_X1   g30999(.A1(new_n34287_), .A2(new_n34284_), .A3(pi1135), .ZN(new_n34288_));
  AOI21_X1   g31000(.A1(new_n34281_), .A2(new_n30557_), .B(new_n34288_), .ZN(new_n34289_));
  NOR2_X1    g31001(.A1(new_n34289_), .A2(new_n5132_), .ZN(new_n34290_));
  NAND2_X1   g31002(.A1(new_n34280_), .A2(new_n12654_), .ZN(new_n34291_));
  NAND2_X1   g31003(.A1(new_n34274_), .A2(new_n34291_), .ZN(new_n34292_));
  AOI21_X1   g31004(.A1(new_n34287_), .A2(new_n34282_), .B(pi1135), .ZN(new_n34293_));
  NAND2_X1   g31005(.A1(new_n8549_), .A2(pi1135), .ZN(new_n34294_));
  AOI21_X1   g31006(.A1(new_n34294_), .A2(pi0200), .B(new_n3098_), .ZN(new_n34295_));
  AOI22_X1   g31007(.A1(pi0211), .A2(pi1136), .B1(pi0219), .B2(pi1135), .ZN(new_n34296_));
  NOR2_X1    g31008(.A1(new_n8549_), .A2(new_n4785_), .ZN(new_n34297_));
  NOR4_X1    g31009(.A1(new_n34297_), .A2(new_n34296_), .A3(pi0200), .A4(new_n3098_), .ZN(new_n34298_));
  XOR2_X1    g31010(.A1(new_n34298_), .A2(new_n34295_), .Z(new_n34299_));
  NAND2_X1   g31011(.A1(new_n34296_), .A2(pi0230), .ZN(new_n34300_));
  NOR2_X1    g31012(.A1(new_n7240_), .A2(new_n30557_), .ZN(new_n34301_));
  XNOR2_X1   g31013(.A1(new_n34301_), .A2(new_n34300_), .ZN(new_n34302_));
  AOI21_X1   g31014(.A1(new_n34302_), .A2(new_n34299_), .B(pi0230), .ZN(new_n34303_));
  OAI21_X1   g31015(.A1(new_n34293_), .A2(new_n34144_), .B(new_n34303_), .ZN(new_n34304_));
  NOR2_X1    g31016(.A1(pi0211), .A2(pi1135), .ZN(new_n34305_));
  INV_X1     g31017(.I(new_n34305_), .ZN(new_n34306_));
  AOI22_X1   g31018(.A1(new_n34306_), .A2(pi1136), .B1(pi0219), .B2(pi1135), .ZN(new_n34307_));
  OAI21_X1   g31019(.A1(pi0199), .A2(pi1136), .B(pi1135), .ZN(new_n34308_));
  NAND2_X1   g31020(.A1(pi0200), .A2(pi1136), .ZN(new_n34309_));
  NAND3_X1   g31021(.A1(new_n34308_), .A2(new_n34309_), .A3(pi0230), .ZN(new_n34310_));
  XOR2_X1    g31022(.A1(new_n32800_), .A2(new_n34310_), .Z(new_n34311_));
  NOR4_X1    g31023(.A1(new_n34311_), .A2(new_n8555_), .A3(new_n5132_), .A4(new_n34307_), .ZN(new_n34312_));
  NAND3_X1   g31024(.A1(new_n34292_), .A2(new_n34304_), .A3(new_n34312_), .ZN(new_n34313_));
  XNOR2_X1   g31025(.A1(new_n34290_), .A2(new_n34313_), .ZN(po0423));
  NOR2_X1    g31026(.A1(new_n34132_), .A2(pi1091), .ZN(new_n34315_));
  AOI21_X1   g31027(.A1(new_n34315_), .A2(new_n13817_), .B(new_n33676_), .ZN(new_n34316_));
  NOR2_X1    g31028(.A1(new_n9208_), .A2(new_n30767_), .ZN(new_n34317_));
  NOR3_X1    g31029(.A1(new_n34316_), .A2(pi1091), .A3(new_n34317_), .ZN(new_n34318_));
  NOR2_X1    g31030(.A1(new_n34318_), .A2(new_n13778_), .ZN(new_n34319_));
  NAND2_X1   g31031(.A1(new_n34319_), .A2(pi0211), .ZN(new_n34320_));
  AOI21_X1   g31032(.A1(new_n31008_), .A2(pi1155), .B(new_n13817_), .ZN(new_n34321_));
  INV_X1     g31033(.I(new_n34126_), .ZN(new_n34322_));
  AOI21_X1   g31034(.A1(new_n31683_), .A2(new_n30701_), .B(new_n34322_), .ZN(new_n34323_));
  NAND2_X1   g31035(.A1(new_n31937_), .A2(new_n2726_), .ZN(new_n34324_));
  NAND3_X1   g31036(.A1(new_n34321_), .A2(new_n34323_), .A3(new_n34324_), .ZN(new_n34325_));
  AOI21_X1   g31037(.A1(new_n34320_), .A2(new_n34133_), .B(new_n34325_), .ZN(new_n34326_));
  INV_X1     g31038(.I(new_n34319_), .ZN(new_n34327_));
  NOR3_X1    g31039(.A1(new_n30667_), .A2(pi0211), .A3(new_n33873_), .ZN(new_n34328_));
  NOR3_X1    g31040(.A1(new_n31706_), .A2(new_n34328_), .A3(new_n8683_), .ZN(new_n34329_));
  NAND3_X1   g31041(.A1(new_n30995_), .A2(new_n2726_), .A3(new_n13778_), .ZN(new_n34330_));
  NAND2_X1   g31042(.A1(new_n31031_), .A2(new_n34330_), .ZN(new_n34331_));
  AOI21_X1   g31043(.A1(new_n34331_), .A2(new_n34315_), .B(new_n33676_), .ZN(new_n34332_));
  OAI21_X1   g31044(.A1(pi1154), .A2(new_n34329_), .B(new_n34332_), .ZN(new_n34333_));
  OAI21_X1   g31045(.A1(new_n34327_), .A2(new_n34333_), .B(pi0267), .ZN(new_n34334_));
  NOR2_X1    g31046(.A1(new_n34326_), .A2(new_n34334_), .ZN(new_n34335_));
  NOR2_X1    g31047(.A1(new_n13614_), .A2(new_n13778_), .ZN(new_n34336_));
  NOR2_X1    g31048(.A1(new_n32724_), .A2(new_n13778_), .ZN(new_n34337_));
  XOR2_X1    g31049(.A1(new_n34337_), .A2(new_n34336_), .Z(new_n34338_));
  NOR2_X1    g31050(.A1(new_n30969_), .A2(pi1155), .ZN(new_n34339_));
  AOI22_X1   g31051(.A1(new_n34338_), .A2(new_n32754_), .B1(pi1091), .B2(new_n34339_), .ZN(new_n34340_));
  NOR2_X1    g31052(.A1(new_n34340_), .A2(new_n13817_), .ZN(new_n34341_));
  NOR2_X1    g31053(.A1(new_n8683_), .A2(new_n13817_), .ZN(new_n34342_));
  XOR2_X1    g31054(.A1(new_n34341_), .A2(new_n34342_), .Z(new_n34343_));
  NOR3_X1    g31055(.A1(new_n32744_), .A2(new_n13614_), .A3(new_n13778_), .ZN(new_n34344_));
  NOR3_X1    g31056(.A1(new_n32743_), .A2(new_n13614_), .A3(pi1155), .ZN(new_n34345_));
  OAI21_X1   g31057(.A1(new_n34344_), .A2(new_n34345_), .B(new_n32737_), .ZN(new_n34346_));
  NOR2_X1    g31058(.A1(new_n33853_), .A2(pi1155), .ZN(new_n34347_));
  AOI21_X1   g31059(.A1(new_n34346_), .A2(new_n34347_), .B(new_n33677_), .ZN(new_n34348_));
  NAND2_X1   g31060(.A1(new_n34343_), .A2(new_n34348_), .ZN(new_n34349_));
  NOR2_X1    g31061(.A1(new_n31013_), .A2(new_n13614_), .ZN(new_n34350_));
  NOR2_X1    g31062(.A1(new_n34350_), .A2(new_n33874_), .ZN(new_n34351_));
  AOI21_X1   g31063(.A1(new_n34351_), .A2(pi0211), .B(new_n32724_), .ZN(new_n34352_));
  NOR3_X1    g31064(.A1(new_n34352_), .A2(pi1155), .A3(new_n30666_), .ZN(new_n34353_));
  OR2_X2     g31065(.A1(new_n34321_), .A2(pi1091), .Z(new_n34354_));
  NOR2_X1    g31066(.A1(new_n30670_), .A2(new_n13778_), .ZN(new_n34355_));
  NOR2_X1    g31067(.A1(new_n31032_), .A2(pi1155), .ZN(new_n34356_));
  NOR4_X1    g31068(.A1(new_n34355_), .A2(new_n8684_), .A3(new_n10254_), .A4(new_n34356_), .ZN(new_n34357_));
  OAI21_X1   g31069(.A1(new_n34353_), .A2(new_n34354_), .B(new_n34357_), .ZN(new_n34358_));
  NAND2_X1   g31070(.A1(new_n34349_), .A2(new_n34358_), .ZN(new_n34359_));
  INV_X1     g31071(.I(new_n31706_), .ZN(new_n34360_));
  NOR3_X1    g31072(.A1(new_n34350_), .A2(new_n8683_), .A3(new_n33874_), .ZN(new_n34361_));
  OAI21_X1   g31073(.A1(new_n34361_), .A2(pi1155), .B(new_n34360_), .ZN(new_n34362_));
  NOR2_X1    g31074(.A1(new_n34316_), .A2(pi1091), .ZN(new_n34363_));
  XNOR2_X1   g31075(.A1(new_n32724_), .A2(new_n33859_), .ZN(new_n34364_));
  NOR3_X1    g31076(.A1(new_n30735_), .A2(new_n32625_), .A3(new_n30981_), .ZN(new_n34365_));
  NAND4_X1   g31077(.A1(new_n34364_), .A2(new_n34317_), .A3(new_n34339_), .A4(new_n34365_), .ZN(new_n34366_));
  AOI21_X1   g31078(.A1(new_n34362_), .A2(new_n34363_), .B(new_n34366_), .ZN(new_n34367_));
  NAND2_X1   g31079(.A1(new_n34359_), .A2(new_n34367_), .ZN(new_n34368_));
  XOR2_X1    g31080(.A1(new_n34368_), .A2(new_n34335_), .Z(new_n34369_));
  AOI21_X1   g31081(.A1(new_n32589_), .A2(new_n33719_), .B(new_n32686_), .ZN(new_n34370_));
  NOR2_X1    g31082(.A1(new_n33884_), .A2(pi1155), .ZN(new_n34371_));
  NOR4_X1    g31083(.A1(new_n34371_), .A2(new_n13614_), .A3(new_n32653_), .A4(new_n34370_), .ZN(new_n34372_));
  OAI21_X1   g31084(.A1(new_n34106_), .A2(new_n13778_), .B(new_n13614_), .ZN(new_n34373_));
  NAND2_X1   g31085(.A1(new_n34373_), .A2(new_n32644_), .ZN(new_n34374_));
  OAI21_X1   g31086(.A1(new_n33733_), .A2(new_n32559_), .B(new_n13778_), .ZN(new_n34375_));
  NOR2_X1    g31087(.A1(new_n33903_), .A2(new_n13614_), .ZN(new_n34376_));
  AOI21_X1   g31088(.A1(new_n34376_), .A2(new_n34375_), .B(pi1154), .ZN(new_n34377_));
  NAND2_X1   g31089(.A1(new_n8684_), .A2(new_n32625_), .ZN(new_n34378_));
  AOI21_X1   g31090(.A1(new_n34374_), .A2(new_n34377_), .B(new_n34378_), .ZN(new_n34379_));
  NOR2_X1    g31091(.A1(new_n32686_), .A2(new_n13614_), .ZN(new_n34380_));
  XNOR2_X1   g31092(.A1(new_n34380_), .A2(new_n34336_), .ZN(new_n34381_));
  NOR3_X1    g31093(.A1(new_n33904_), .A2(pi0211), .A3(pi1155), .ZN(new_n34382_));
  NOR2_X1    g31094(.A1(new_n32619_), .A2(pi1153), .ZN(new_n34383_));
  NOR3_X1    g31095(.A1(new_n33940_), .A2(new_n32559_), .A3(new_n34383_), .ZN(new_n34384_));
  NAND4_X1   g31096(.A1(new_n34384_), .A2(new_n30768_), .A3(new_n32613_), .A4(new_n32661_), .ZN(new_n34385_));
  OR4_X2     g31097(.A1(new_n34374_), .A2(new_n34381_), .A3(new_n34382_), .A4(new_n34385_), .Z(new_n34386_));
  OAI22_X1   g31098(.A1(new_n34386_), .A2(new_n34379_), .B1(new_n13817_), .B2(new_n34372_), .ZN(new_n34387_));
  NAND2_X1   g31099(.A1(new_n33909_), .A2(new_n30769_), .ZN(new_n34388_));
  AOI21_X1   g31100(.A1(new_n34388_), .A2(pi1153), .B(new_n32696_), .ZN(new_n34389_));
  AOI21_X1   g31101(.A1(new_n34387_), .A2(new_n34389_), .B(new_n8683_), .ZN(new_n34390_));
  AOI21_X1   g31102(.A1(new_n32600_), .A2(pi1153), .B(new_n13778_), .ZN(new_n34391_));
  OR3_X2     g31103(.A1(new_n33731_), .A2(pi0267), .A3(new_n34391_), .Z(new_n34392_));
  NAND2_X1   g31104(.A1(new_n32568_), .A2(new_n13817_), .ZN(new_n34393_));
  NAND3_X1   g31105(.A1(new_n34393_), .A2(new_n32588_), .A3(new_n32616_), .ZN(new_n34394_));
  AOI21_X1   g31106(.A1(new_n30852_), .A2(new_n33749_), .B(new_n34394_), .ZN(new_n34395_));
  AOI21_X1   g31107(.A1(new_n34392_), .A2(new_n34395_), .B(pi1154), .ZN(new_n34396_));
  INV_X1     g31108(.I(new_n34370_), .ZN(new_n34397_));
  NOR3_X1    g31109(.A1(new_n34384_), .A2(pi0267), .A3(pi1155), .ZN(new_n34398_));
  INV_X1     g31110(.I(new_n30928_), .ZN(new_n34399_));
  NOR4_X1    g31111(.A1(new_n33940_), .A2(new_n32647_), .A3(new_n34399_), .A4(new_n32570_), .ZN(new_n34400_));
  OAI21_X1   g31112(.A1(new_n31304_), .A2(new_n33699_), .B(new_n34400_), .ZN(new_n34401_));
  OAI21_X1   g31113(.A1(new_n34401_), .A2(new_n34398_), .B(new_n13817_), .ZN(new_n34402_));
  NAND4_X1   g31114(.A1(new_n34402_), .A2(pi1153), .A3(new_n33884_), .A4(new_n34397_), .ZN(new_n34403_));
  OAI21_X1   g31115(.A1(new_n34396_), .A2(new_n34403_), .B(new_n8684_), .ZN(new_n34404_));
  AOI21_X1   g31116(.A1(new_n13614_), .A2(new_n32675_), .B(new_n32687_), .ZN(new_n34405_));
  NAND2_X1   g31117(.A1(new_n32668_), .A2(new_n13817_), .ZN(new_n34406_));
  OAI21_X1   g31118(.A1(new_n34406_), .A2(new_n34391_), .B(new_n32539_), .ZN(new_n34407_));
  NAND3_X1   g31119(.A1(new_n34407_), .A2(new_n13778_), .A3(new_n32653_), .ZN(new_n34408_));
  NAND2_X1   g31120(.A1(new_n34408_), .A2(new_n34405_), .ZN(new_n34409_));
  AOI21_X1   g31121(.A1(new_n32686_), .A2(new_n13614_), .B(pi1154), .ZN(new_n34410_));
  NOR2_X1    g31122(.A1(new_n34410_), .A2(new_n32599_), .ZN(new_n34411_));
  NAND2_X1   g31123(.A1(new_n34409_), .A2(new_n34411_), .ZN(new_n34412_));
  NOR2_X1    g31124(.A1(new_n33897_), .A2(new_n13817_), .ZN(new_n34413_));
  NAND2_X1   g31125(.A1(new_n32661_), .A2(pi1155), .ZN(new_n34414_));
  OAI21_X1   g31126(.A1(new_n34413_), .A2(new_n34414_), .B(new_n32605_), .ZN(new_n34415_));
  AOI21_X1   g31127(.A1(new_n34415_), .A2(pi1153), .B(pi0211), .ZN(new_n34416_));
  AOI21_X1   g31128(.A1(new_n34410_), .A2(new_n32670_), .B(pi1155), .ZN(new_n34417_));
  NAND3_X1   g31129(.A1(new_n34417_), .A2(pi1154), .A3(new_n34405_), .ZN(new_n34418_));
  OAI21_X1   g31130(.A1(new_n34416_), .A2(new_n34418_), .B(new_n32625_), .ZN(new_n34419_));
  INV_X1     g31131(.I(new_n34417_), .ZN(new_n34420_));
  NOR4_X1    g31132(.A1(new_n32584_), .A2(new_n13614_), .A3(new_n30769_), .A4(new_n32580_), .ZN(new_n34421_));
  NOR3_X1    g31133(.A1(new_n34421_), .A2(pi1154), .A3(new_n34384_), .ZN(new_n34422_));
  NOR4_X1    g31134(.A1(new_n34422_), .A2(new_n31937_), .A3(new_n33896_), .A4(new_n34420_), .ZN(new_n34423_));
  NAND4_X1   g31135(.A1(new_n34404_), .A2(new_n34412_), .A3(new_n34419_), .A4(new_n34423_), .ZN(new_n34424_));
  OAI21_X1   g31136(.A1(new_n34424_), .A2(new_n34390_), .B(new_n32628_), .ZN(new_n34425_));
  AOI21_X1   g31137(.A1(new_n34390_), .A2(new_n34424_), .B(new_n34425_), .ZN(new_n34426_));
  NAND2_X1   g31138(.A1(po1038), .A2(new_n32628_), .ZN(new_n34427_));
  XOR2_X1    g31139(.A1(new_n34426_), .A2(new_n34427_), .Z(new_n34428_));
  OAI21_X1   g31140(.A1(new_n34428_), .A2(new_n34369_), .B(new_n32773_), .ZN(new_n34429_));
  NAND3_X1   g31141(.A1(new_n32551_), .A2(new_n32625_), .A3(new_n32629_), .ZN(new_n34430_));
  NOR2_X1    g31142(.A1(new_n32628_), .A2(new_n2726_), .ZN(new_n34431_));
  NOR2_X1    g31143(.A1(new_n30994_), .A2(new_n8683_), .ZN(new_n34432_));
  NAND3_X1   g31144(.A1(new_n31304_), .A2(new_n30635_), .A3(pi0219), .ZN(new_n34433_));
  XOR2_X1    g31145(.A1(new_n34433_), .A2(new_n34432_), .Z(new_n34434_));
  NOR3_X1    g31146(.A1(new_n34434_), .A2(new_n32625_), .A3(new_n2726_), .ZN(new_n34435_));
  XOR2_X1    g31147(.A1(new_n34435_), .A2(new_n34431_), .Z(new_n34436_));
  NAND2_X1   g31148(.A1(new_n34430_), .A2(new_n34436_), .ZN(new_n34437_));
  OAI21_X1   g31149(.A1(new_n33744_), .A2(new_n34437_), .B(new_n32625_), .ZN(new_n34438_));
  NAND4_X1   g31150(.A1(new_n34429_), .A2(po1038), .A3(new_n33925_), .A4(new_n34438_), .ZN(new_n34439_));
  NOR2_X1    g31151(.A1(new_n34323_), .A2(new_n8683_), .ZN(new_n34440_));
  XOR2_X1    g31152(.A1(new_n34440_), .A2(new_n31936_), .Z(new_n34441_));
  NAND4_X1   g31153(.A1(new_n30783_), .A2(new_n8549_), .A3(new_n8555_), .A4(pi1153), .ZN(new_n34443_));
  NAND3_X1   g31154(.A1(new_n34441_), .A2(new_n30611_), .A3(new_n34443_), .ZN(new_n34444_));
  NOR4_X1    g31155(.A1(new_n31009_), .A2(new_n13778_), .A3(new_n30735_), .A4(new_n31016_), .ZN(new_n34445_));
  AOI21_X1   g31156(.A1(pi1154), .A2(new_n31031_), .B(new_n34350_), .ZN(new_n34446_));
  NOR3_X1    g31157(.A1(new_n34446_), .A2(new_n8683_), .A3(new_n13778_), .ZN(new_n34447_));
  OAI21_X1   g31158(.A1(new_n34447_), .A2(new_n34445_), .B(pi0211), .ZN(new_n34448_));
  AOI21_X1   g31159(.A1(new_n34444_), .A2(new_n7240_), .B(new_n34448_), .ZN(new_n34449_));
  NOR2_X1    g31160(.A1(new_n34434_), .A2(new_n7240_), .ZN(new_n34450_));
  AOI21_X1   g31161(.A1(new_n34449_), .A2(new_n34450_), .B(pi0230), .ZN(new_n34451_));
  NAND2_X1   g31162(.A1(new_n2726_), .A2(pi0267), .ZN(new_n34452_));
  OAI21_X1   g31163(.A1(new_n34434_), .A2(new_n2726_), .B(new_n34452_), .ZN(new_n34453_));
  NAND2_X1   g31164(.A1(new_n34369_), .A2(po1038), .ZN(new_n34454_));
  XNOR2_X1   g31165(.A1(new_n34454_), .A2(new_n32805_), .ZN(new_n34455_));
  NAND2_X1   g31166(.A1(new_n34455_), .A2(new_n34453_), .ZN(new_n34456_));
  AOI21_X1   g31167(.A1(new_n34439_), .A2(new_n34451_), .B(new_n34456_), .ZN(po0424));
  NOR2_X1    g31168(.A1(new_n33924_), .A2(new_n7240_), .ZN(new_n34458_));
  NAND3_X1   g31169(.A1(new_n32687_), .A2(pi0219), .A3(po1038), .ZN(new_n34459_));
  NAND3_X1   g31170(.A1(new_n33909_), .A2(pi0219), .A3(new_n7240_), .ZN(new_n34460_));
  AOI21_X1   g31171(.A1(new_n34460_), .A2(new_n34459_), .B(new_n33698_), .ZN(new_n34461_));
  NAND2_X1   g31172(.A1(new_n34461_), .A2(new_n34458_), .ZN(new_n34462_));
  NAND2_X1   g31173(.A1(new_n34462_), .A2(new_n33752_), .ZN(new_n34463_));
  NAND2_X1   g31174(.A1(new_n34463_), .A2(pi0219), .ZN(new_n34464_));
  AOI21_X1   g31175(.A1(new_n32543_), .A2(new_n2726_), .B(po1038), .ZN(new_n34465_));
  AOI21_X1   g31176(.A1(new_n34464_), .A2(new_n34465_), .B(new_n33773_), .ZN(new_n34466_));
  INV_X1     g31177(.I(new_n34458_), .ZN(new_n34467_));
  NOR3_X1    g31178(.A1(new_n33702_), .A2(new_n8683_), .A3(new_n32580_), .ZN(new_n34468_));
  AOI21_X1   g31179(.A1(new_n33882_), .A2(new_n33728_), .B(new_n34468_), .ZN(new_n34469_));
  NAND2_X1   g31180(.A1(new_n34469_), .A2(po1038), .ZN(new_n34470_));
  AOI21_X1   g31181(.A1(new_n34470_), .A2(new_n32640_), .B(new_n33738_), .ZN(new_n34471_));
  OAI21_X1   g31182(.A1(new_n32565_), .A2(new_n33724_), .B(new_n34471_), .ZN(new_n34472_));
  OAI21_X1   g31183(.A1(new_n33753_), .A2(new_n34467_), .B(new_n34472_), .ZN(new_n34473_));
  NAND2_X1   g31184(.A1(new_n34473_), .A2(pi0268), .ZN(new_n34474_));
  NAND2_X1   g31185(.A1(pi0268), .A2(pi1151), .ZN(new_n34475_));
  XOR2_X1    g31186(.A1(new_n34474_), .A2(new_n34475_), .Z(new_n34476_));
  AOI21_X1   g31187(.A1(new_n34476_), .A2(new_n34466_), .B(new_n31002_), .ZN(new_n34477_));
  NOR2_X1    g31188(.A1(new_n33909_), .A2(new_n8683_), .ZN(new_n34478_));
  OAI21_X1   g31189(.A1(po1038), .A2(new_n32619_), .B(new_n34478_), .ZN(new_n34479_));
  NOR2_X1    g31190(.A1(new_n32565_), .A2(new_n31349_), .ZN(new_n34480_));
  INV_X1     g31191(.I(new_n34480_), .ZN(new_n34481_));
  AND3_X2    g31192(.A1(new_n34479_), .A2(new_n33746_), .A3(new_n34481_), .Z(new_n34482_));
  NOR2_X1    g31193(.A1(new_n33755_), .A2(new_n31349_), .ZN(new_n34483_));
  INV_X1     g31194(.I(new_n34483_), .ZN(new_n34484_));
  NAND2_X1   g31195(.A1(new_n33755_), .A2(new_n31349_), .ZN(new_n34485_));
  AOI21_X1   g31196(.A1(new_n34484_), .A2(new_n34485_), .B(new_n33752_), .ZN(new_n34486_));
  NOR2_X1    g31197(.A1(new_n34461_), .A2(new_n34486_), .ZN(new_n34487_));
  NOR2_X1    g31198(.A1(new_n34487_), .A2(new_n32548_), .ZN(new_n34488_));
  NOR2_X1    g31199(.A1(new_n34482_), .A2(new_n34488_), .ZN(new_n34489_));
  INV_X1     g31200(.I(new_n32566_), .ZN(new_n34490_));
  AOI21_X1   g31201(.A1(new_n33714_), .A2(new_n8683_), .B(new_n34490_), .ZN(new_n34491_));
  INV_X1     g31202(.I(new_n34491_), .ZN(new_n34492_));
  NOR2_X1    g31203(.A1(new_n5788_), .A2(pi0057), .ZN(new_n34494_));
  AOI21_X1   g31204(.A1(new_n34492_), .A2(new_n34494_), .B(new_n32613_), .ZN(new_n34495_));
  NOR2_X1    g31205(.A1(new_n34495_), .A2(new_n31670_), .ZN(new_n34496_));
  XNOR2_X1   g31206(.A1(new_n34496_), .A2(new_n34475_), .ZN(new_n34497_));
  NAND2_X1   g31207(.A1(new_n34497_), .A2(new_n34489_), .ZN(new_n34498_));
  OR3_X2     g31208(.A1(new_n34167_), .A2(new_n7240_), .A3(new_n33812_), .Z(new_n34499_));
  AOI21_X1   g31209(.A1(new_n34492_), .A2(new_n34499_), .B(new_n33700_), .ZN(new_n34500_));
  INV_X1     g31210(.I(new_n34500_), .ZN(new_n34501_));
  NAND2_X1   g31211(.A1(new_n34501_), .A2(pi1151), .ZN(new_n34502_));
  XOR2_X1    g31212(.A1(new_n34502_), .A2(new_n34475_), .Z(new_n34503_));
  INV_X1     g31213(.I(new_n34469_), .ZN(new_n34504_));
  NOR2_X1    g31214(.A1(new_n32574_), .A2(new_n8683_), .ZN(new_n34505_));
  AOI21_X1   g31215(.A1(new_n33753_), .A2(new_n34505_), .B(po1038), .ZN(new_n34506_));
  NAND2_X1   g31216(.A1(new_n34504_), .A2(new_n34506_), .ZN(new_n34507_));
  NAND2_X1   g31217(.A1(new_n34507_), .A2(new_n33723_), .ZN(new_n34508_));
  NAND2_X1   g31218(.A1(new_n34508_), .A2(pi0268), .ZN(new_n34509_));
  XOR2_X1    g31219(.A1(new_n34509_), .A2(new_n34475_), .Z(new_n34510_));
  NAND2_X1   g31220(.A1(new_n34510_), .A2(new_n34487_), .ZN(new_n34511_));
  NAND3_X1   g31221(.A1(new_n33702_), .A2(pi0219), .A3(po1038), .ZN(new_n34512_));
  NAND3_X1   g31222(.A1(new_n33703_), .A2(pi0219), .A3(new_n7240_), .ZN(new_n34513_));
  AOI21_X1   g31223(.A1(new_n34513_), .A2(new_n34512_), .B(new_n33705_), .ZN(new_n34514_));
  OAI21_X1   g31224(.A1(po1038), .A2(new_n34167_), .B(new_n33754_), .ZN(new_n34515_));
  NOR3_X1    g31225(.A1(new_n34514_), .A2(new_n31002_), .A3(new_n34515_), .ZN(new_n34516_));
  NAND4_X1   g31226(.A1(new_n34511_), .A2(new_n34498_), .A3(new_n34503_), .A4(new_n34516_), .ZN(new_n34517_));
  XNOR2_X1   g31227(.A1(new_n34477_), .A2(new_n34517_), .ZN(new_n34518_));
  NOR2_X1    g31228(.A1(new_n34471_), .A2(new_n34480_), .ZN(new_n34519_));
  NOR4_X1    g31229(.A1(new_n34519_), .A2(pi0219), .A3(new_n7240_), .A4(new_n33753_), .ZN(new_n34520_));
  NOR2_X1    g31230(.A1(new_n34520_), .A2(new_n31670_), .ZN(new_n34521_));
  XNOR2_X1   g31231(.A1(new_n34521_), .A2(new_n33420_), .ZN(new_n34522_));
  NAND2_X1   g31232(.A1(new_n34522_), .A2(new_n34482_), .ZN(new_n34523_));
  INV_X1     g31233(.I(new_n33731_), .ZN(new_n34524_));
  NAND2_X1   g31234(.A1(po1038), .A2(pi0219), .ZN(new_n34525_));
  OAI22_X1   g31235(.A1(new_n34524_), .A2(new_n34525_), .B1(new_n33710_), .B2(new_n34467_), .ZN(new_n34526_));
  NAND2_X1   g31236(.A1(new_n33919_), .A2(po1038), .ZN(new_n34527_));
  AOI21_X1   g31237(.A1(new_n33713_), .A2(new_n32667_), .B(pi0219), .ZN(new_n34528_));
  NOR4_X1    g31238(.A1(new_n34528_), .A2(new_n7240_), .A3(new_n34524_), .A4(new_n33923_), .ZN(new_n34529_));
  XOR2_X1    g31239(.A1(new_n34529_), .A2(new_n34527_), .Z(new_n34530_));
  NAND2_X1   g31240(.A1(new_n34530_), .A2(pi1152), .ZN(new_n34531_));
  XNOR2_X1   g31241(.A1(new_n34531_), .A2(new_n33420_), .ZN(new_n34532_));
  NOR2_X1    g31242(.A1(new_n34532_), .A2(new_n34526_), .ZN(new_n34533_));
  INV_X1     g31243(.I(pi0268), .ZN(new_n34534_));
  NAND2_X1   g31244(.A1(new_n34534_), .A2(new_n32242_), .ZN(new_n34535_));
  NAND2_X1   g31245(.A1(new_n33814_), .A2(new_n7240_), .ZN(new_n34536_));
  OAI21_X1   g31246(.A1(new_n33713_), .A2(new_n34536_), .B(new_n33774_), .ZN(new_n34537_));
  NAND2_X1   g31247(.A1(new_n34537_), .A2(pi1151), .ZN(new_n34538_));
  XNOR2_X1   g31248(.A1(new_n34538_), .A2(new_n33420_), .ZN(new_n34539_));
  INV_X1     g31249(.I(new_n34487_), .ZN(new_n34540_));
  NAND2_X1   g31250(.A1(new_n34540_), .A2(new_n32548_), .ZN(new_n34541_));
  NOR3_X1    g31251(.A1(new_n34539_), .A2(new_n34534_), .A3(new_n34541_), .ZN(new_n34542_));
  OAI21_X1   g31252(.A1(new_n34533_), .A2(new_n34535_), .B(new_n34542_), .ZN(new_n34543_));
  NOR2_X1    g31253(.A1(new_n32696_), .A2(new_n8683_), .ZN(new_n34544_));
  OAI21_X1   g31254(.A1(new_n34514_), .A2(new_n32573_), .B(new_n34544_), .ZN(new_n34545_));
  NAND3_X1   g31255(.A1(new_n34545_), .A2(new_n7240_), .A3(new_n33746_), .ZN(new_n34546_));
  NAND2_X1   g31256(.A1(new_n34546_), .A2(new_n34167_), .ZN(new_n34547_));
  NAND2_X1   g31257(.A1(new_n34547_), .A2(pi1152), .ZN(new_n34548_));
  XOR2_X1    g31258(.A1(new_n34548_), .A2(new_n33420_), .Z(new_n34549_));
  NOR2_X1    g31259(.A1(new_n33754_), .A2(new_n7240_), .ZN(new_n34550_));
  NOR3_X1    g31260(.A1(new_n34504_), .A2(new_n7240_), .A3(new_n33744_), .ZN(new_n34551_));
  XNOR2_X1   g31261(.A1(new_n34551_), .A2(new_n34550_), .ZN(new_n34552_));
  INV_X1     g31262(.I(new_n34552_), .ZN(new_n34553_));
  NAND3_X1   g31263(.A1(new_n34549_), .A2(new_n32772_), .A3(new_n34553_), .ZN(new_n34554_));
  AOI21_X1   g31264(.A1(new_n34523_), .A2(new_n34543_), .B(new_n34554_), .ZN(new_n34555_));
  OAI21_X1   g31265(.A1(new_n34555_), .A2(pi1150), .B(new_n34518_), .ZN(new_n34556_));
  NAND3_X1   g31266(.A1(new_n32522_), .A2(new_n30668_), .A3(new_n33657_), .ZN(new_n34557_));
  NAND3_X1   g31267(.A1(new_n32522_), .A2(new_n30652_), .A3(new_n33656_), .ZN(new_n34558_));
  NAND2_X1   g31268(.A1(new_n34557_), .A2(new_n34558_), .ZN(new_n34559_));
  NOR2_X1    g31269(.A1(new_n7240_), .A2(new_n9259_), .ZN(new_n34560_));
  AOI21_X1   g31270(.A1(new_n7240_), .A2(new_n9262_), .B(new_n34560_), .ZN(new_n34561_));
  AOI21_X1   g31271(.A1(pi1150), .A2(pi1152), .B(pi1151), .ZN(new_n34562_));
  OAI22_X1   g31272(.A1(new_n34559_), .A2(new_n33420_), .B1(new_n34561_), .B2(new_n34562_), .ZN(new_n34563_));
  NAND3_X1   g31273(.A1(new_n34563_), .A2(pi1151), .A3(new_n33806_), .ZN(new_n34564_));
  NAND2_X1   g31274(.A1(new_n12655_), .A2(new_n8684_), .ZN(new_n34565_));
  OAI21_X1   g31275(.A1(po1038), .A2(new_n30735_), .B(new_n34565_), .ZN(new_n34566_));
  INV_X1     g31276(.I(new_n34566_), .ZN(new_n34567_));
  NOR2_X1    g31277(.A1(new_n12655_), .A2(pi0199), .ZN(new_n34568_));
  NOR2_X1    g31278(.A1(new_n34568_), .A2(new_n32089_), .ZN(new_n34569_));
  NAND2_X1   g31279(.A1(new_n34569_), .A2(pi1150), .ZN(new_n34570_));
  AOI21_X1   g31280(.A1(new_n34567_), .A2(new_n31670_), .B(new_n34570_), .ZN(new_n34571_));
  OAI21_X1   g31281(.A1(new_n34571_), .A2(pi1152), .B(new_n34567_), .ZN(new_n34572_));
  AND2_X2    g31282(.A1(new_n34572_), .A2(pi0230), .Z(new_n34573_));
  AOI21_X1   g31283(.A1(new_n34573_), .A2(new_n34564_), .B(pi0230), .ZN(new_n34574_));
  OAI21_X1   g31284(.A1(new_n34534_), .A2(new_n2726_), .B(new_n31002_), .ZN(new_n34575_));
  NAND2_X1   g31285(.A1(new_n32772_), .A2(new_n34575_), .ZN(new_n34576_));
  OAI21_X1   g31286(.A1(new_n34572_), .A2(new_n34576_), .B(new_n2726_), .ZN(new_n34577_));
  OAI21_X1   g31287(.A1(new_n34572_), .A2(new_n34564_), .B(new_n31002_), .ZN(new_n34578_));
  NAND3_X1   g31288(.A1(new_n34577_), .A2(new_n34578_), .A3(pi0268), .ZN(new_n34579_));
  AOI21_X1   g31289(.A1(new_n34556_), .A2(new_n34574_), .B(new_n34579_), .ZN(po0425));
  NAND2_X1   g31290(.A1(new_n12655_), .A2(new_n8549_), .ZN(new_n34581_));
  NOR2_X1    g31291(.A1(new_n12654_), .A2(new_n8683_), .ZN(new_n34582_));
  NOR2_X1    g31292(.A1(new_n2726_), .A2(pi0200), .ZN(new_n34583_));
  NAND4_X1   g31293(.A1(new_n34581_), .A2(pi1138), .A3(new_n34582_), .A4(new_n34583_), .ZN(new_n34584_));
  NAND2_X1   g31294(.A1(new_n34584_), .A2(new_n4465_), .ZN(new_n34585_));
  INV_X1     g31295(.I(pi0269), .ZN(new_n34586_));
  INV_X1     g31296(.I(pi0817), .ZN(new_n34587_));
  NAND2_X1   g31297(.A1(new_n32529_), .A2(new_n34587_), .ZN(new_n34588_));
  XNOR2_X1   g31298(.A1(new_n34237_), .A2(new_n34588_), .ZN(new_n34589_));
  NOR3_X1    g31299(.A1(new_n34589_), .A2(new_n34586_), .A3(new_n33651_), .ZN(new_n34590_));
  INV_X1     g31300(.I(new_n34568_), .ZN(new_n34591_));
  NOR2_X1    g31301(.A1(new_n2726_), .A2(pi1137), .ZN(new_n34592_));
  NAND2_X1   g31302(.A1(pi0200), .A2(pi1091), .ZN(new_n34593_));
  XOR2_X1    g31303(.A1(new_n34592_), .A2(new_n34593_), .Z(new_n34594_));
  NOR2_X1    g31304(.A1(pi0211), .A2(pi1136), .ZN(new_n34595_));
  AOI21_X1   g31305(.A1(pi0211), .A2(new_n4626_), .B(new_n34595_), .ZN(new_n34596_));
  NAND3_X1   g31306(.A1(new_n34596_), .A2(pi1091), .A3(pi1136), .ZN(new_n34597_));
  OAI22_X1   g31307(.A1(new_n34591_), .A2(new_n32090_), .B1(new_n34594_), .B2(new_n34597_), .ZN(new_n34598_));
  NAND3_X1   g31308(.A1(new_n32540_), .A2(pi0817), .A3(pi1091), .ZN(new_n34599_));
  NAND3_X1   g31309(.A1(new_n32540_), .A2(new_n34587_), .A3(new_n2726_), .ZN(new_n34600_));
  AOI21_X1   g31310(.A1(new_n34599_), .A2(new_n34600_), .B(new_n34586_), .ZN(new_n34601_));
  AOI22_X1   g31311(.A1(new_n34585_), .A2(new_n34590_), .B1(new_n34598_), .B2(new_n34601_), .ZN(new_n34602_));
  NAND4_X1   g31312(.A1(pi0199), .A2(pi0200), .A3(pi1136), .A4(pi1138), .ZN(new_n34603_));
  NOR2_X1    g31313(.A1(new_n12655_), .A2(new_n8549_), .ZN(new_n34604_));
  INV_X1     g31314(.I(new_n34604_), .ZN(new_n34605_));
  AOI21_X1   g31315(.A1(new_n4626_), .A2(new_n34603_), .B(new_n34605_), .ZN(new_n34606_));
  NOR3_X1    g31316(.A1(new_n34596_), .A2(new_n8683_), .A3(new_n4465_), .ZN(new_n34607_));
  XOR2_X1    g31317(.A1(new_n34607_), .A2(new_n30615_), .Z(new_n34608_));
  NOR2_X1    g31318(.A1(new_n34608_), .A2(new_n12654_), .ZN(new_n34609_));
  OAI21_X1   g31319(.A1(new_n34606_), .A2(new_n34609_), .B(pi0230), .ZN(new_n34610_));
  OAI21_X1   g31320(.A1(new_n34602_), .A2(pi0230), .B(new_n34610_), .ZN(po0426));
  NAND2_X1   g31321(.A1(new_n2726_), .A2(new_n3980_), .ZN(new_n34612_));
  NOR2_X1    g31322(.A1(new_n34612_), .A2(pi0199), .ZN(new_n34613_));
  NOR2_X1    g31323(.A1(new_n34582_), .A2(new_n34612_), .ZN(new_n34614_));
  INV_X1     g31324(.I(pi0805), .ZN(new_n34615_));
  NAND2_X1   g31325(.A1(new_n32540_), .A2(new_n34615_), .ZN(new_n34616_));
  XOR2_X1    g31326(.A1(new_n34264_), .A2(new_n34616_), .Z(new_n34617_));
  NAND3_X1   g31327(.A1(new_n34617_), .A2(pi0211), .A3(pi0270), .ZN(new_n34618_));
  OAI22_X1   g31328(.A1(new_n34614_), .A2(new_n34618_), .B1(new_n8555_), .B2(new_n34613_), .ZN(new_n34619_));
  NAND2_X1   g31329(.A1(new_n4141_), .A2(pi0211), .ZN(new_n34620_));
  OAI21_X1   g31330(.A1(pi0211), .A2(pi1139), .B(new_n34620_), .ZN(new_n34621_));
  AOI21_X1   g31331(.A1(new_n34619_), .A2(new_n12654_), .B(pi0230), .ZN(new_n34626_));
  NAND3_X1   g31332(.A1(pi0200), .A2(pi1091), .A3(pi1140), .ZN(new_n34627_));
  NAND3_X1   g31333(.A1(new_n8555_), .A2(new_n4141_), .A3(pi1091), .ZN(new_n34628_));
  AOI21_X1   g31334(.A1(new_n34628_), .A2(new_n34627_), .B(new_n4300_), .ZN(new_n34629_));
  INV_X1     g31335(.I(pi0270), .ZN(new_n34630_));
  NAND2_X1   g31336(.A1(new_n32529_), .A2(new_n34615_), .ZN(new_n34631_));
  XNOR2_X1   g31337(.A1(new_n34237_), .A2(new_n34631_), .ZN(new_n34632_));
  NOR2_X1    g31338(.A1(new_n34621_), .A2(new_n2726_), .ZN(new_n34633_));
  NOR4_X1    g31339(.A1(new_n32090_), .A2(new_n34630_), .A3(new_n34632_), .A4(new_n34633_), .ZN(new_n34634_));
  OAI21_X1   g31340(.A1(new_n34634_), .A2(new_n34629_), .B(new_n34568_), .ZN(new_n34635_));
  NOR2_X1    g31341(.A1(new_n34626_), .A2(new_n34635_), .ZN(po0427));
  NAND4_X1   g31342(.A1(pi0211), .A2(pi0219), .A3(pi1145), .A4(pi1146), .ZN(new_n34637_));
  NAND2_X1   g31343(.A1(new_n34637_), .A2(new_n31940_), .ZN(new_n34638_));
  AOI21_X1   g31344(.A1(new_n34638_), .A2(pi0211), .B(new_n30557_), .ZN(new_n34639_));
  XNOR2_X1   g31345(.A1(new_n34301_), .A2(new_n34639_), .ZN(new_n34640_));
  NAND3_X1   g31346(.A1(new_n31503_), .A2(pi0211), .A3(pi0219), .ZN(new_n34641_));
  NAND3_X1   g31347(.A1(new_n31511_), .A2(pi0211), .A3(new_n8683_), .ZN(new_n34642_));
  NAND2_X1   g31348(.A1(new_n34642_), .A2(new_n34641_), .ZN(new_n34643_));
  NAND2_X1   g31349(.A1(new_n31902_), .A2(pi0200), .ZN(new_n34644_));
  NAND2_X1   g31350(.A1(new_n34644_), .A2(new_n3518_), .ZN(new_n34645_));
  AOI22_X1   g31351(.A1(new_n34645_), .A2(pi0199), .B1(new_n34643_), .B2(new_n31912_), .ZN(new_n34646_));
  NOR4_X1    g31352(.A1(new_n34640_), .A2(new_n31940_), .A3(new_n33689_), .A4(new_n34646_), .ZN(new_n34647_));
  NOR2_X1    g31353(.A1(new_n32533_), .A2(pi0271), .ZN(new_n34648_));
  INV_X1     g31354(.I(pi0271), .ZN(new_n34649_));
  NOR2_X1    g31355(.A1(new_n32532_), .A2(new_n34649_), .ZN(new_n34650_));
  OAI21_X1   g31356(.A1(new_n34648_), .A2(new_n34650_), .B(new_n2726_), .ZN(new_n34651_));
  OAI21_X1   g31357(.A1(new_n2726_), .A2(new_n3350_), .B(new_n34651_), .ZN(new_n34652_));
  NOR2_X1    g31358(.A1(new_n33651_), .A2(new_n3350_), .ZN(new_n34653_));
  INV_X1     g31359(.I(new_n34653_), .ZN(new_n34654_));
  AOI21_X1   g31360(.A1(new_n34652_), .A2(new_n34654_), .B(new_n8683_), .ZN(new_n34655_));
  NAND2_X1   g31361(.A1(new_n32542_), .A2(new_n34649_), .ZN(new_n34656_));
  NAND2_X1   g31362(.A1(new_n32543_), .A2(pi0271), .ZN(new_n34657_));
  AOI21_X1   g31363(.A1(new_n34657_), .A2(new_n34656_), .B(pi1091), .ZN(new_n34658_));
  NOR2_X1    g31364(.A1(new_n33651_), .A2(new_n3518_), .ZN(new_n34659_));
  NAND3_X1   g31365(.A1(new_n34658_), .A2(pi0219), .A3(new_n34659_), .ZN(new_n34660_));
  NAND2_X1   g31366(.A1(new_n34655_), .A2(new_n34660_), .ZN(new_n34661_));
  OR2_X2     g31367(.A1(new_n34655_), .A2(new_n34660_), .Z(new_n34662_));
  NAND3_X1   g31368(.A1(new_n34662_), .A2(new_n12654_), .A3(new_n34661_), .ZN(new_n34663_));
  NAND3_X1   g31369(.A1(pi0199), .A2(pi1091), .A3(pi1145), .ZN(new_n34664_));
  INV_X1     g31370(.I(new_n34658_), .ZN(new_n34665_));
  NAND2_X1   g31371(.A1(new_n34652_), .A2(pi0200), .ZN(new_n34666_));
  XOR2_X1    g31372(.A1(new_n34666_), .A2(new_n30722_), .Z(new_n34667_));
  NOR2_X1    g31373(.A1(new_n34667_), .A2(new_n34665_), .ZN(new_n34668_));
  NOR2_X1    g31374(.A1(pi0200), .A2(pi1091), .ZN(new_n34669_));
  AOI21_X1   g31375(.A1(new_n34669_), .A2(new_n31940_), .B(new_n8549_), .ZN(new_n34670_));
  NAND2_X1   g31376(.A1(new_n34668_), .A2(new_n34670_), .ZN(new_n34671_));
  NOR3_X1    g31377(.A1(new_n8549_), .A2(new_n8683_), .A3(new_n31940_), .ZN(new_n34672_));
  NAND4_X1   g31378(.A1(new_n34665_), .A2(new_n12654_), .A3(new_n33691_), .A4(new_n34672_), .ZN(new_n34673_));
  AOI21_X1   g31379(.A1(new_n34671_), .A2(new_n34664_), .B(new_n34673_), .ZN(new_n34674_));
  OR2_X2     g31380(.A1(new_n34674_), .A2(new_n34663_), .Z(new_n34675_));
  AOI21_X1   g31381(.A1(new_n34674_), .A2(new_n34663_), .B(pi0230), .ZN(new_n34676_));
  AOI21_X1   g31382(.A1(new_n34675_), .A2(new_n34676_), .B(new_n34647_), .ZN(po0428));
  NOR2_X1    g31383(.A1(new_n7240_), .A2(pi0211), .ZN(new_n34678_));
  INV_X1     g31384(.I(new_n10256_), .ZN(new_n34679_));
  NAND2_X1   g31385(.A1(new_n34679_), .A2(new_n9213_), .ZN(new_n34680_));
  XOR2_X1    g31386(.A1(new_n34680_), .A2(new_n34678_), .Z(new_n34681_));
  OAI21_X1   g31387(.A1(new_n31941_), .A2(new_n34566_), .B(new_n34681_), .ZN(new_n34682_));
  AOI22_X1   g31388(.A1(new_n34682_), .A2(pi1150), .B1(pi1091), .B2(pi1148), .ZN(new_n34683_));
  INV_X1     g31389(.I(new_n34569_), .ZN(new_n34684_));
  OAI21_X1   g31390(.A1(new_n34684_), .A2(new_n34566_), .B(new_n31941_), .ZN(new_n34685_));
  NAND2_X1   g31391(.A1(new_n34685_), .A2(pi1150), .ZN(new_n34686_));
  NOR2_X1    g31392(.A1(pi0272), .A2(pi0283), .ZN(new_n34687_));
  OAI21_X1   g31393(.A1(new_n34683_), .A2(new_n34686_), .B(new_n34687_), .ZN(new_n34688_));
  NOR2_X1    g31394(.A1(new_n9259_), .A2(new_n2726_), .ZN(new_n34689_));
  NOR4_X1    g31395(.A1(po1038), .A2(pi0299), .A3(new_n32734_), .A4(new_n34689_), .ZN(new_n34690_));
  OAI21_X1   g31396(.A1(new_n34559_), .A2(new_n2726_), .B(pi1149), .ZN(new_n34691_));
  XOR2_X1    g31397(.A1(new_n34691_), .A2(new_n33113_), .Z(new_n34692_));
  NAND2_X1   g31398(.A1(new_n34692_), .A2(new_n34690_), .ZN(new_n34693_));
  AOI21_X1   g31399(.A1(new_n2726_), .A2(new_n31941_), .B(new_n32242_), .ZN(new_n34694_));
  NAND2_X1   g31400(.A1(new_n33806_), .A2(new_n34694_), .ZN(new_n34695_));
  NAND4_X1   g31401(.A1(new_n34688_), .A2(new_n31953_), .A3(new_n34693_), .A4(new_n34695_), .ZN(new_n34696_));
  NOR2_X1    g31402(.A1(new_n34520_), .A2(new_n31941_), .ZN(new_n34697_));
  XNOR2_X1   g31403(.A1(new_n34697_), .A2(new_n33113_), .ZN(new_n34698_));
  AOI21_X1   g31404(.A1(new_n34698_), .A2(new_n34553_), .B(new_n31953_), .ZN(new_n34699_));
  NAND2_X1   g31405(.A1(new_n34547_), .A2(pi1150), .ZN(new_n34700_));
  XOR2_X1    g31406(.A1(new_n34700_), .A2(new_n33113_), .Z(new_n34701_));
  NOR2_X1    g31407(.A1(new_n34495_), .A2(new_n32242_), .ZN(new_n34702_));
  XNOR2_X1   g31408(.A1(new_n34702_), .A2(new_n33113_), .ZN(new_n34703_));
  NAND2_X1   g31409(.A1(new_n34703_), .A2(new_n34500_), .ZN(new_n34704_));
  INV_X1     g31410(.I(new_n34482_), .ZN(new_n34705_));
  NOR2_X1    g31411(.A1(new_n34514_), .A2(new_n34515_), .ZN(new_n34706_));
  NOR2_X1    g31412(.A1(new_n34705_), .A2(new_n31953_), .ZN(new_n34709_));
  NAND3_X1   g31413(.A1(new_n34701_), .A2(new_n34704_), .A3(new_n34709_), .ZN(new_n34710_));
  XOR2_X1    g31414(.A1(new_n34699_), .A2(new_n34710_), .Z(new_n34711_));
  NOR2_X1    g31415(.A1(new_n34559_), .A2(new_n31941_), .ZN(new_n34712_));
  XOR2_X1    g31416(.A1(new_n34712_), .A2(new_n33113_), .Z(new_n34713_));
  INV_X1     g31417(.I(new_n34561_), .ZN(new_n34714_));
  AOI21_X1   g31418(.A1(new_n32242_), .A2(new_n31976_), .B(new_n33805_), .ZN(new_n34715_));
  INV_X1     g31419(.I(new_n34715_), .ZN(new_n34716_));
  NAND3_X1   g31420(.A1(new_n34716_), .A2(new_n32771_), .A3(new_n2726_), .ZN(new_n34717_));
  NAND3_X1   g31421(.A1(new_n34717_), .A2(pi0272), .A3(new_n34714_), .ZN(new_n34718_));
  OAI21_X1   g31422(.A1(new_n34718_), .A2(new_n34713_), .B(new_n2726_), .ZN(new_n34719_));
  AOI21_X1   g31423(.A1(new_n34682_), .A2(pi1150), .B(pi1148), .ZN(new_n34720_));
  NAND2_X1   g31424(.A1(new_n32090_), .A2(new_n34565_), .ZN(new_n34721_));
  NOR2_X1    g31425(.A1(new_n7240_), .A2(new_n30738_), .ZN(new_n34722_));
  AOI21_X1   g31426(.A1(new_n34721_), .A2(new_n34722_), .B(new_n32242_), .ZN(new_n34723_));
  NOR4_X1    g31427(.A1(new_n34720_), .A2(new_n31941_), .A3(new_n34684_), .A4(new_n34723_), .ZN(new_n34724_));
  AND2_X2    g31428(.A1(new_n34724_), .A2(pi0230), .Z(new_n34725_));
  AOI21_X1   g31429(.A1(new_n34725_), .A2(new_n34719_), .B(pi0283), .ZN(new_n34726_));
  NAND2_X1   g31430(.A1(new_n34712_), .A2(new_n34714_), .ZN(new_n34727_));
  NAND4_X1   g31431(.A1(new_n34721_), .A2(pi1149), .A3(pi1150), .A4(new_n34722_), .ZN(new_n34728_));
  AOI21_X1   g31432(.A1(new_n34727_), .A2(new_n34728_), .B(new_n34716_), .ZN(new_n34729_));
  OAI21_X1   g31433(.A1(new_n34724_), .A2(pi0230), .B(new_n34729_), .ZN(new_n34730_));
  OR3_X2     g31434(.A1(new_n34711_), .A2(new_n34726_), .A3(new_n34730_), .Z(new_n34731_));
  NAND2_X1   g31435(.A1(new_n34473_), .A2(pi1150), .ZN(new_n34732_));
  XNOR2_X1   g31436(.A1(new_n34732_), .A2(new_n33113_), .ZN(new_n34733_));
  NOR2_X1    g31437(.A1(new_n34733_), .A2(new_n34508_), .ZN(new_n34734_));
  NAND2_X1   g31438(.A1(new_n34530_), .A2(pi1149), .ZN(new_n34735_));
  XNOR2_X1   g31439(.A1(new_n34735_), .A2(new_n33113_), .ZN(new_n34736_));
  NAND2_X1   g31440(.A1(new_n34526_), .A2(pi1150), .ZN(new_n34737_));
  XNOR2_X1   g31441(.A1(new_n34737_), .A2(new_n33113_), .ZN(new_n34738_));
  NOR2_X1    g31442(.A1(new_n34738_), .A2(new_n34541_), .ZN(new_n34739_));
  AOI21_X1   g31443(.A1(pi0283), .A2(pi1148), .B(new_n34739_), .ZN(new_n34740_));
  NOR4_X1    g31444(.A1(new_n34736_), .A2(new_n31953_), .A3(new_n34537_), .A4(new_n34740_), .ZN(new_n34741_));
  NOR2_X1    g31445(.A1(new_n34466_), .A2(new_n31941_), .ZN(new_n34742_));
  XOR2_X1    g31446(.A1(new_n34742_), .A2(new_n33113_), .Z(new_n34743_));
  NOR2_X1    g31447(.A1(new_n34743_), .A2(new_n34540_), .ZN(new_n34744_));
  OAI21_X1   g31448(.A1(new_n34734_), .A2(new_n34741_), .B(new_n34744_), .ZN(new_n34745_));
  AOI21_X1   g31449(.A1(new_n34731_), .A2(new_n34696_), .B(new_n34745_), .ZN(po0429));
  AOI21_X1   g31450(.A1(new_n32545_), .A2(pi0273), .B(new_n34649_), .ZN(new_n34747_));
  NAND2_X1   g31451(.A1(new_n34747_), .A2(new_n32534_), .ZN(new_n34748_));
  AOI21_X1   g31452(.A1(new_n34214_), .A2(new_n3350_), .B(new_n8555_), .ZN(new_n34749_));
  NAND2_X1   g31453(.A1(new_n34748_), .A2(new_n34749_), .ZN(new_n34750_));
  XOR2_X1    g31454(.A1(new_n32544_), .A2(pi0271), .Z(new_n34751_));
  OAI21_X1   g31455(.A1(new_n32543_), .A2(new_n34751_), .B(pi0199), .ZN(new_n34752_));
  NAND3_X1   g31456(.A1(new_n34750_), .A2(new_n3098_), .A3(new_n34752_), .ZN(new_n34753_));
  NAND2_X1   g31457(.A1(new_n34748_), .A2(pi0219), .ZN(new_n34754_));
  NOR4_X1    g31458(.A1(new_n32543_), .A2(new_n8683_), .A3(new_n34654_), .A4(new_n34751_), .ZN(new_n34755_));
  XOR2_X1    g31459(.A1(new_n34754_), .A2(new_n34755_), .Z(new_n34756_));
  OAI21_X1   g31460(.A1(new_n34756_), .A2(new_n3098_), .B(new_n34753_), .ZN(new_n34757_));
  NOR2_X1    g31461(.A1(new_n34757_), .A2(new_n7240_), .ZN(new_n34758_));
  AOI22_X1   g31462(.A1(new_n32568_), .A2(new_n9259_), .B1(pi0299), .B2(new_n32570_), .ZN(new_n34759_));
  NOR2_X1    g31463(.A1(new_n34759_), .A2(new_n31940_), .ZN(new_n34760_));
  AOI21_X1   g31464(.A1(new_n34760_), .A2(new_n34758_), .B(pi1091), .ZN(new_n34761_));
  OAI21_X1   g31465(.A1(new_n34756_), .A2(new_n3098_), .B(new_n2726_), .ZN(new_n34762_));
  NAND2_X1   g31466(.A1(new_n34762_), .A2(new_n30615_), .ZN(new_n34763_));
  NAND3_X1   g31467(.A1(po1038), .A2(pi1091), .A3(new_n31936_), .ZN(new_n34764_));
  NAND2_X1   g31468(.A1(new_n34764_), .A2(new_n31953_), .ZN(new_n34765_));
  NAND4_X1   g31469(.A1(new_n34668_), .A2(po1038), .A3(new_n32737_), .A4(new_n34765_), .ZN(new_n34766_));
  AOI21_X1   g31470(.A1(new_n34753_), .A2(new_n34763_), .B(new_n34766_), .ZN(new_n34767_));
  AND2_X2    g31471(.A1(new_n34757_), .A2(new_n32836_), .Z(new_n34768_));
  OR2_X2     g31472(.A1(new_n34756_), .A2(pi1148), .Z(new_n34769_));
  NAND3_X1   g31473(.A1(new_n34681_), .A2(pi1146), .A3(new_n33146_), .ZN(new_n34770_));
  OAI21_X1   g31474(.A1(pi1146), .A2(new_n8773_), .B(new_n32089_), .ZN(new_n34771_));
  OAI21_X1   g31475(.A1(new_n34591_), .A2(new_n34771_), .B(new_n8684_), .ZN(new_n34772_));
  NAND3_X1   g31476(.A1(new_n34772_), .A2(pi1147), .A3(new_n31912_), .ZN(new_n34773_));
  AOI21_X1   g31477(.A1(new_n34770_), .A2(new_n31953_), .B(new_n34773_), .ZN(new_n34774_));
  NAND4_X1   g31478(.A1(new_n12655_), .A2(new_n8684_), .A3(new_n8683_), .A4(new_n3350_), .ZN(new_n34775_));
  NAND4_X1   g31479(.A1(new_n12655_), .A2(new_n8683_), .A3(pi0230), .A4(pi1148), .ZN(new_n34779_));
  AOI21_X1   g31480(.A1(new_n31940_), .A2(new_n34775_), .B(new_n34779_), .ZN(new_n34780_));
  OAI21_X1   g31481(.A1(new_n34774_), .A2(pi0230), .B(new_n34780_), .ZN(new_n34781_));
  OAI21_X1   g31482(.A1(new_n34768_), .A2(new_n34769_), .B(new_n34781_), .ZN(new_n34782_));
  OAI21_X1   g31483(.A1(new_n34767_), .A2(new_n34782_), .B(new_n33813_), .ZN(new_n34783_));
  NOR2_X1    g31484(.A1(new_n34761_), .A2(new_n34783_), .ZN(po0430));
  INV_X1     g31485(.I(pi0659), .ZN(new_n34785_));
  NOR3_X1    g31486(.A1(new_n32530_), .A2(new_n34785_), .A3(new_n2726_), .ZN(new_n34786_));
  NOR3_X1    g31487(.A1(new_n32530_), .A2(pi0659), .A3(pi1091), .ZN(new_n34787_));
  OAI21_X1   g31488(.A1(new_n34786_), .A2(new_n34787_), .B(pi0274), .ZN(new_n34788_));
  NAND2_X1   g31489(.A1(new_n34788_), .A2(new_n34245_), .ZN(new_n34789_));
  OAI21_X1   g31490(.A1(new_n2726_), .A2(new_n3057_), .B(new_n34788_), .ZN(new_n34790_));
  NAND2_X1   g31491(.A1(new_n34790_), .A2(pi0200), .ZN(new_n34791_));
  XOR2_X1    g31492(.A1(new_n34791_), .A2(new_n30722_), .Z(new_n34792_));
  OAI21_X1   g31493(.A1(new_n34792_), .A2(new_n34789_), .B(new_n12655_), .ZN(new_n34793_));
  NOR3_X1    g31494(.A1(new_n32541_), .A2(new_n34785_), .A3(new_n2726_), .ZN(new_n34794_));
  NOR3_X1    g31495(.A1(new_n32541_), .A2(pi0659), .A3(pi1091), .ZN(new_n34795_));
  OAI21_X1   g31496(.A1(new_n34794_), .A2(new_n34795_), .B(pi0274), .ZN(new_n34796_));
  OAI21_X1   g31497(.A1(new_n34215_), .A2(pi1145), .B(pi0200), .ZN(new_n34797_));
  NOR2_X1    g31498(.A1(new_n34796_), .A2(new_n34797_), .ZN(new_n34798_));
  NAND2_X1   g31499(.A1(new_n34793_), .A2(new_n34798_), .ZN(new_n34799_));
  NOR2_X1    g31500(.A1(new_n31937_), .A2(new_n31383_), .ZN(new_n34800_));
  NOR2_X1    g31501(.A1(new_n31384_), .A2(new_n31936_), .ZN(new_n34801_));
  OAI21_X1   g31502(.A1(new_n34800_), .A2(new_n34801_), .B(pi1143), .ZN(new_n34802_));
  OAI21_X1   g31503(.A1(new_n27298_), .A2(pi1144), .B(pi0199), .ZN(new_n34803_));
  OAI21_X1   g31504(.A1(new_n31899_), .A2(new_n34803_), .B(new_n3650_), .ZN(new_n34804_));
  NAND2_X1   g31505(.A1(new_n26962_), .A2(new_n34804_), .ZN(new_n34805_));
  OAI21_X1   g31506(.A1(new_n31511_), .A2(pi0211), .B(new_n30620_), .ZN(new_n34806_));
  AOI21_X1   g31507(.A1(new_n34805_), .A2(new_n34802_), .B(new_n34806_), .ZN(new_n34807_));
  INV_X1     g31508(.I(new_n32020_), .ZN(new_n34808_));
  NOR2_X1    g31509(.A1(new_n34808_), .A2(new_n34802_), .ZN(new_n34809_));
  AOI21_X1   g31510(.A1(new_n34809_), .A2(new_n34807_), .B(pi0230), .ZN(new_n34810_));
  NAND2_X1   g31511(.A1(new_n34790_), .A2(pi0211), .ZN(new_n34811_));
  XOR2_X1    g31512(.A1(new_n34811_), .A2(new_n31936_), .Z(new_n34812_));
  OAI21_X1   g31513(.A1(new_n34812_), .A2(new_n34789_), .B(new_n12655_), .ZN(new_n34813_));
  NOR3_X1    g31514(.A1(new_n34796_), .A2(new_n8683_), .A3(new_n34659_), .ZN(new_n34814_));
  NAND2_X1   g31515(.A1(new_n34813_), .A2(new_n34814_), .ZN(new_n34815_));
  AOI21_X1   g31516(.A1(new_n34799_), .A2(new_n34810_), .B(new_n34815_), .ZN(po0431));
  INV_X1     g31517(.I(new_n34681_), .ZN(new_n34817_));
  NAND2_X1   g31518(.A1(new_n34566_), .A2(new_n31941_), .ZN(new_n34818_));
  NAND3_X1   g31519(.A1(new_n34817_), .A2(pi1151), .A3(new_n34818_), .ZN(new_n34819_));
  NAND2_X1   g31520(.A1(new_n34819_), .A2(pi1150), .ZN(new_n34820_));
  NAND2_X1   g31521(.A1(new_n31941_), .A2(new_n31670_), .ZN(new_n34821_));
  NOR3_X1    g31522(.A1(new_n32242_), .A2(new_n31670_), .A3(pi1149), .ZN(new_n34822_));
  NAND4_X1   g31523(.A1(new_n34559_), .A2(new_n33805_), .A3(new_n34821_), .A4(new_n34822_), .ZN(new_n34823_));
  XNOR2_X1   g31524(.A1(new_n34820_), .A2(new_n34823_), .ZN(new_n34824_));
  NOR3_X1    g31525(.A1(new_n33447_), .A2(new_n32770_), .A3(new_n31941_), .ZN(new_n34825_));
  AOI21_X1   g31526(.A1(new_n34690_), .A2(new_n34825_), .B(pi1091), .ZN(new_n34826_));
  NOR2_X1    g31527(.A1(new_n34559_), .A2(new_n32242_), .ZN(new_n34827_));
  XNOR2_X1   g31528(.A1(new_n34827_), .A2(new_n33447_), .ZN(new_n34828_));
  NAND2_X1   g31529(.A1(new_n34828_), .A2(new_n34714_), .ZN(new_n34829_));
  NOR2_X1    g31530(.A1(new_n33805_), .A2(new_n32246_), .ZN(new_n34830_));
  NOR2_X1    g31531(.A1(new_n34569_), .A2(pi1149), .ZN(new_n34831_));
  NOR3_X1    g31532(.A1(new_n34831_), .A2(new_n31670_), .A3(new_n34566_), .ZN(new_n34832_));
  OAI21_X1   g31533(.A1(new_n34832_), .A2(new_n34818_), .B(pi1150), .ZN(new_n34833_));
  AOI21_X1   g31534(.A1(new_n34829_), .A2(new_n34830_), .B(new_n34833_), .ZN(new_n34834_));
  AND2_X2    g31535(.A1(new_n34834_), .A2(pi1091), .Z(new_n34835_));
  OAI22_X1   g31536(.A1(new_n34835_), .A2(pi0275), .B1(new_n34824_), .B2(new_n34826_), .ZN(new_n34836_));
  NOR2_X1    g31537(.A1(new_n32769_), .A2(new_n32771_), .ZN(new_n34837_));
  AOI21_X1   g31538(.A1(new_n34836_), .A2(new_n34837_), .B(new_n30557_), .ZN(new_n34838_));
  NAND2_X1   g31539(.A1(new_n32770_), .A2(new_n31941_), .ZN(new_n34839_));
  XOR2_X1    g31540(.A1(new_n34502_), .A2(new_n33447_), .Z(new_n34840_));
  AOI21_X1   g31541(.A1(new_n34840_), .A2(new_n34706_), .B(new_n34839_), .ZN(new_n34841_));
  XOR2_X1    g31542(.A1(new_n34702_), .A2(new_n33447_), .Z(new_n34842_));
  NOR4_X1    g31543(.A1(new_n34841_), .A2(new_n34482_), .A3(new_n34488_), .A4(new_n34842_), .ZN(new_n34843_));
  NOR2_X1    g31544(.A1(new_n34466_), .A2(new_n32242_), .ZN(new_n34844_));
  XOR2_X1    g31545(.A1(new_n34844_), .A2(new_n33447_), .Z(new_n34845_));
  OAI21_X1   g31546(.A1(new_n34845_), .A2(new_n34540_), .B(new_n32770_), .ZN(new_n34846_));
  NOR2_X1    g31547(.A1(new_n34843_), .A2(new_n34846_), .ZN(new_n34847_));
  NOR2_X1    g31548(.A1(new_n34520_), .A2(new_n32242_), .ZN(new_n34848_));
  XOR2_X1    g31549(.A1(new_n34848_), .A2(new_n33447_), .Z(new_n34849_));
  NOR2_X1    g31550(.A1(new_n34849_), .A2(new_n34705_), .ZN(new_n34850_));
  NAND2_X1   g31551(.A1(new_n34530_), .A2(pi1151), .ZN(new_n34851_));
  XNOR2_X1   g31552(.A1(new_n34851_), .A2(new_n33447_), .ZN(new_n34852_));
  NOR2_X1    g31553(.A1(new_n34852_), .A2(new_n34526_), .ZN(new_n34853_));
  NOR2_X1    g31554(.A1(new_n34853_), .A2(new_n34839_), .ZN(new_n34854_));
  NAND2_X1   g31555(.A1(new_n34537_), .A2(pi1150), .ZN(new_n34855_));
  XNOR2_X1   g31556(.A1(new_n34855_), .A2(new_n33447_), .ZN(new_n34856_));
  NOR4_X1    g31557(.A1(new_n34854_), .A2(new_n32770_), .A3(new_n34541_), .A4(new_n34856_), .ZN(new_n34857_));
  NAND2_X1   g31558(.A1(new_n34547_), .A2(pi1151), .ZN(new_n34858_));
  XNOR2_X1   g31559(.A1(new_n34858_), .A2(new_n33447_), .ZN(new_n34859_));
  NAND2_X1   g31560(.A1(new_n34473_), .A2(pi1151), .ZN(new_n34860_));
  XNOR2_X1   g31561(.A1(new_n34860_), .A2(new_n33447_), .ZN(new_n34861_));
  NOR3_X1    g31562(.A1(new_n30557_), .A2(new_n32769_), .A3(new_n32771_), .ZN(new_n34862_));
  NAND4_X1   g31563(.A1(new_n34507_), .A2(new_n33723_), .A3(new_n34834_), .A4(new_n34862_), .ZN(new_n34863_));
  NOR4_X1    g31564(.A1(new_n34861_), .A2(new_n34552_), .A3(new_n34859_), .A4(new_n34863_), .ZN(new_n34864_));
  OAI21_X1   g31565(.A1(new_n34857_), .A2(new_n34850_), .B(new_n34864_), .ZN(new_n34865_));
  NOR2_X1    g31566(.A1(new_n34865_), .A2(new_n34847_), .ZN(new_n34866_));
  XOR2_X1    g31567(.A1(new_n34866_), .A2(new_n34838_), .Z(po0432));
  NAND3_X1   g31568(.A1(pi0200), .A2(pi1091), .A3(pi1145), .ZN(new_n34868_));
  NAND3_X1   g31569(.A1(new_n8555_), .A2(new_n3518_), .A3(pi1091), .ZN(new_n34869_));
  AOI21_X1   g31570(.A1(new_n34869_), .A2(new_n34868_), .B(new_n3057_), .ZN(new_n34870_));
  NOR3_X1    g31571(.A1(new_n32002_), .A2(new_n2726_), .A3(new_n30559_), .ZN(new_n34871_));
  NAND2_X1   g31572(.A1(pi0276), .A2(pi1091), .ZN(new_n34872_));
  XOR2_X1    g31573(.A1(new_n34872_), .A2(pi0802), .Z(new_n34873_));
  NOR4_X1    g31574(.A1(new_n32090_), .A2(new_n32530_), .A3(new_n34871_), .A4(new_n34873_), .ZN(new_n34874_));
  OAI21_X1   g31575(.A1(new_n34874_), .A2(new_n34870_), .B(new_n34568_), .ZN(new_n34875_));
  NOR2_X1    g31576(.A1(new_n32002_), .A2(new_n30559_), .ZN(new_n34876_));
  NOR3_X1    g31577(.A1(new_n34876_), .A2(new_n8683_), .A3(new_n3350_), .ZN(new_n34877_));
  XOR2_X1    g31578(.A1(new_n34877_), .A2(new_n30615_), .Z(new_n34878_));
  AOI21_X1   g31579(.A1(new_n32800_), .A2(new_n34878_), .B(pi0230), .ZN(new_n34882_));
  INV_X1     g31580(.I(new_n34749_), .ZN(new_n34883_));
  NOR4_X1    g31581(.A1(new_n12655_), .A2(new_n32541_), .A3(new_n34883_), .A4(new_n34873_), .ZN(new_n34884_));
  OAI21_X1   g31582(.A1(new_n34884_), .A2(new_n34582_), .B(new_n34653_), .ZN(new_n34885_));
  AOI21_X1   g31583(.A1(new_n34875_), .A2(new_n34882_), .B(new_n34885_), .ZN(po0433));
  INV_X1     g31584(.I(pi0820), .ZN(new_n34887_));
  NOR3_X1    g31585(.A1(new_n32530_), .A2(new_n34887_), .A3(new_n2726_), .ZN(new_n34888_));
  NOR3_X1    g31586(.A1(new_n32530_), .A2(pi0820), .A3(pi1091), .ZN(new_n34889_));
  OAI21_X1   g31587(.A1(new_n34888_), .A2(new_n34889_), .B(pi0277), .ZN(new_n34890_));
  NAND2_X1   g31588(.A1(new_n34890_), .A2(new_n34206_), .ZN(new_n34891_));
  OAI21_X1   g31589(.A1(new_n2726_), .A2(new_n4141_), .B(new_n34890_), .ZN(new_n34892_));
  NAND2_X1   g31590(.A1(new_n34892_), .A2(pi0200), .ZN(new_n34893_));
  XOR2_X1    g31591(.A1(new_n34893_), .A2(new_n30722_), .Z(new_n34894_));
  OAI21_X1   g31592(.A1(new_n34894_), .A2(new_n34891_), .B(new_n12655_), .ZN(new_n34895_));
  NOR3_X1    g31593(.A1(new_n32541_), .A2(new_n34887_), .A3(new_n2726_), .ZN(new_n34896_));
  NOR3_X1    g31594(.A1(new_n32541_), .A2(pi0820), .A3(pi1091), .ZN(new_n34897_));
  OAI21_X1   g31595(.A1(new_n34896_), .A2(new_n34897_), .B(pi0277), .ZN(new_n34898_));
  NAND2_X1   g31596(.A1(new_n2726_), .A2(new_n3814_), .ZN(new_n34899_));
  OAI21_X1   g31597(.A1(new_n34899_), .A2(pi0199), .B(pi0200), .ZN(new_n34900_));
  NOR2_X1    g31598(.A1(new_n34898_), .A2(new_n34900_), .ZN(new_n34901_));
  NAND2_X1   g31599(.A1(new_n34895_), .A2(new_n34901_), .ZN(new_n34902_));
  OAI21_X1   g31600(.A1(new_n3980_), .A2(pi0199), .B(pi0200), .ZN(new_n34903_));
  OAI21_X1   g31601(.A1(new_n30571_), .A2(new_n34903_), .B(new_n4141_), .ZN(new_n34904_));
  AOI21_X1   g31602(.A1(new_n34904_), .A2(pi0199), .B(new_n30557_), .ZN(new_n34905_));
  XOR2_X1    g31603(.A1(new_n32800_), .A2(new_n34905_), .Z(new_n34906_));
  NAND4_X1   g31604(.A1(pi0211), .A2(pi0219), .A3(pi1140), .A4(pi1141), .ZN(new_n34907_));
  NAND2_X1   g31605(.A1(new_n34907_), .A2(new_n3814_), .ZN(new_n34908_));
  NAND4_X1   g31606(.A1(new_n34906_), .A2(pi0211), .A3(pi0230), .A4(new_n34908_), .ZN(new_n34909_));
  NAND2_X1   g31607(.A1(new_n34892_), .A2(pi0211), .ZN(new_n34910_));
  XOR2_X1    g31608(.A1(new_n34910_), .A2(new_n31936_), .Z(new_n34911_));
  OAI21_X1   g31609(.A1(new_n34911_), .A2(new_n34891_), .B(new_n12655_), .ZN(new_n34912_));
  OAI21_X1   g31610(.A1(new_n34899_), .A2(pi0219), .B(pi0211), .ZN(new_n34913_));
  NOR2_X1    g31611(.A1(new_n34898_), .A2(new_n34913_), .ZN(new_n34914_));
  NAND2_X1   g31612(.A1(new_n34912_), .A2(new_n34914_), .ZN(new_n34915_));
  AOI21_X1   g31613(.A1(new_n34902_), .A2(new_n34909_), .B(new_n34915_), .ZN(po0434));
  INV_X1     g31614(.I(pi0278), .ZN(po1130));
  NAND3_X1   g31615(.A1(new_n32540_), .A2(pi0976), .A3(pi1091), .ZN(new_n34918_));
  NOR2_X1    g31616(.A1(new_n32541_), .A2(pi0976), .ZN(new_n34919_));
  NAND2_X1   g31617(.A1(new_n34919_), .A2(new_n34264_), .ZN(new_n34920_));
  AOI21_X1   g31618(.A1(new_n34920_), .A2(new_n34918_), .B(po1130), .ZN(new_n34921_));
  INV_X1     g31619(.I(new_n34921_), .ZN(new_n34922_));
  NOR2_X1    g31620(.A1(new_n32530_), .A2(pi0976), .ZN(new_n34923_));
  XNOR2_X1   g31621(.A1(new_n34923_), .A2(new_n34237_), .ZN(new_n34924_));
  NAND2_X1   g31622(.A1(new_n34924_), .A2(pi0278), .ZN(new_n34925_));
  INV_X1     g31623(.I(pi1132), .ZN(new_n34926_));
  NAND2_X1   g31624(.A1(new_n34926_), .A2(pi1091), .ZN(new_n34927_));
  AOI21_X1   g31625(.A1(new_n34925_), .A2(new_n34927_), .B(new_n8549_), .ZN(new_n34928_));
  XOR2_X1    g31626(.A1(new_n34928_), .A2(new_n32795_), .Z(new_n34929_));
  NOR2_X1    g31627(.A1(new_n34929_), .A2(new_n34922_), .ZN(new_n34930_));
  NAND2_X1   g31628(.A1(new_n34925_), .A2(pi0199), .ZN(new_n34931_));
  NOR4_X1    g31629(.A1(new_n34922_), .A2(new_n8549_), .A3(new_n2726_), .A4(pi1133), .ZN(new_n34932_));
  OR2_X2     g31630(.A1(new_n34931_), .A2(new_n34932_), .Z(new_n34933_));
  AOI21_X1   g31631(.A1(new_n34931_), .A2(new_n34932_), .B(new_n8555_), .ZN(new_n34934_));
  AOI21_X1   g31632(.A1(new_n34933_), .A2(new_n34934_), .B(pi0299), .ZN(new_n34935_));
  AOI21_X1   g31633(.A1(new_n34930_), .A2(new_n34935_), .B(pi1091), .ZN(new_n34936_));
  OAI22_X1   g31634(.A1(new_n34936_), .A2(new_n8549_), .B1(new_n34153_), .B2(new_n33651_), .ZN(new_n34937_));
  NAND2_X1   g31635(.A1(new_n34925_), .A2(pi0219), .ZN(new_n34938_));
  INV_X1     g31636(.I(pi1133), .ZN(new_n34939_));
  NOR2_X1    g31637(.A1(new_n8684_), .A2(new_n34939_), .ZN(new_n34940_));
  AOI21_X1   g31638(.A1(new_n8684_), .A2(pi1132), .B(new_n34940_), .ZN(new_n34941_));
  NAND4_X1   g31639(.A1(new_n34921_), .A2(pi0219), .A3(pi1091), .A4(new_n34941_), .ZN(new_n34942_));
  XOR2_X1    g31640(.A1(new_n34938_), .A2(new_n34942_), .Z(new_n34943_));
  AOI21_X1   g31641(.A1(new_n34943_), .A2(po1038), .B(pi0230), .ZN(new_n34944_));
  INV_X1     g31642(.I(new_n34944_), .ZN(new_n34945_));
  NAND2_X1   g31643(.A1(new_n34943_), .A2(new_n32522_), .ZN(new_n34946_));
  AOI21_X1   g31644(.A1(new_n34945_), .A2(new_n34764_), .B(new_n34946_), .ZN(new_n34947_));
  AOI21_X1   g31645(.A1(new_n34937_), .A2(new_n34947_), .B(new_n5132_), .ZN(new_n34948_));
  NOR3_X1    g31646(.A1(new_n7240_), .A2(pi0219), .A3(new_n34941_), .ZN(new_n34949_));
  NOR2_X1    g31647(.A1(new_n34941_), .A2(new_n30620_), .ZN(new_n34950_));
  NOR2_X1    g31648(.A1(new_n34301_), .A2(new_n34950_), .ZN(new_n34951_));
  AOI21_X1   g31649(.A1(new_n27299_), .A2(new_n34939_), .B(new_n8549_), .ZN(new_n34952_));
  AOI21_X1   g31650(.A1(new_n34952_), .A2(pi0200), .B(pi1132), .ZN(new_n34953_));
  NOR4_X1    g31651(.A1(new_n34951_), .A2(new_n8549_), .A3(new_n34949_), .A4(new_n34953_), .ZN(new_n34954_));
  AOI21_X1   g31652(.A1(new_n34944_), .A2(new_n34954_), .B(po1038), .ZN(new_n34955_));
  AOI22_X1   g31653(.A1(new_n34930_), .A2(pi0299), .B1(new_n34935_), .B2(new_n34943_), .ZN(new_n34956_));
  NAND2_X1   g31654(.A1(po1038), .A2(new_n34941_), .ZN(new_n34957_));
  XOR2_X1    g31655(.A1(new_n9213_), .A2(new_n34957_), .Z(new_n34958_));
  OAI21_X1   g31656(.A1(new_n34958_), .A2(new_n8684_), .B(new_n30557_), .ZN(new_n34959_));
  INV_X1     g31657(.I(new_n34950_), .ZN(new_n34960_));
  NAND2_X1   g31658(.A1(new_n8555_), .A2(new_n34926_), .ZN(new_n34961_));
  OAI21_X1   g31659(.A1(new_n34952_), .A2(new_n34961_), .B(pi0199), .ZN(new_n34962_));
  NAND4_X1   g31660(.A1(po1038), .A2(pi0299), .A3(pi1134), .A4(new_n30615_), .ZN(new_n34963_));
  AOI21_X1   g31661(.A1(new_n34960_), .A2(new_n34962_), .B(new_n34963_), .ZN(new_n34964_));
  NAND2_X1   g31662(.A1(new_n34959_), .A2(new_n34964_), .ZN(new_n34965_));
  NOR3_X1    g31663(.A1(new_n34956_), .A2(new_n34955_), .A3(new_n34965_), .ZN(new_n34966_));
  XOR2_X1    g31664(.A1(new_n34948_), .A2(new_n34966_), .Z(po0435));
  NAND3_X1   g31665(.A1(new_n32529_), .A2(pi0958), .A3(pi1091), .ZN(new_n34968_));
  OR3_X2     g31666(.A1(new_n32530_), .A2(pi0958), .A3(pi1091), .Z(new_n34969_));
  AOI21_X1   g31667(.A1(new_n34969_), .A2(new_n34968_), .B(new_n4964_), .ZN(new_n34970_));
  INV_X1     g31668(.I(new_n34583_), .ZN(new_n34971_));
  NOR3_X1    g31669(.A1(new_n12655_), .A2(new_n34939_), .A3(new_n34971_), .ZN(new_n34972_));
  AOI21_X1   g31670(.A1(new_n34972_), .A2(new_n34970_), .B(pi0199), .ZN(new_n34973_));
  NOR2_X1    g31671(.A1(new_n32541_), .A2(pi0958), .ZN(new_n34974_));
  XNOR2_X1   g31672(.A1(new_n34974_), .A2(new_n34264_), .ZN(new_n34975_));
  NAND2_X1   g31673(.A1(new_n34975_), .A2(pi0279), .ZN(new_n34976_));
  OAI21_X1   g31674(.A1(new_n4959_), .A2(new_n34971_), .B(new_n34976_), .ZN(new_n34977_));
  NOR2_X1    g31675(.A1(new_n34977_), .A2(new_n34973_), .ZN(new_n34978_));
  NAND2_X1   g31676(.A1(new_n33650_), .A2(pi1135), .ZN(new_n34979_));
  AOI21_X1   g31677(.A1(new_n34976_), .A2(new_n8683_), .B(new_n34979_), .ZN(new_n34980_));
  NOR3_X1    g31678(.A1(new_n34980_), .A2(pi0230), .A3(new_n12654_), .ZN(new_n34981_));
  OAI21_X1   g31679(.A1(new_n2726_), .A2(pi1133), .B(new_n8683_), .ZN(new_n34982_));
  OAI21_X1   g31680(.A1(new_n34970_), .A2(new_n34982_), .B(new_n33691_), .ZN(new_n34983_));
  NOR2_X1    g31681(.A1(new_n34981_), .A2(new_n34983_), .ZN(new_n34984_));
  NAND2_X1   g31682(.A1(new_n34984_), .A2(new_n34978_), .ZN(new_n34985_));
  NAND2_X1   g31683(.A1(new_n34985_), .A2(new_n2726_), .ZN(new_n34986_));
  AOI21_X1   g31684(.A1(new_n34986_), .A2(pi0200), .B(new_n5132_), .ZN(new_n34987_));
  INV_X1     g31685(.I(new_n34984_), .ZN(new_n34988_));
  NAND3_X1   g31686(.A1(new_n8684_), .A2(new_n34939_), .A3(pi0219), .ZN(new_n34989_));
  NAND4_X1   g31687(.A1(new_n30616_), .A2(pi0211), .A3(new_n34939_), .A4(pi1135), .ZN(new_n34990_));
  NAND2_X1   g31688(.A1(new_n34990_), .A2(new_n34989_), .ZN(new_n34991_));
  NAND4_X1   g31689(.A1(new_n31420_), .A2(pi0200), .A3(pi1133), .A4(new_n4959_), .ZN(new_n34992_));
  NAND2_X1   g31690(.A1(pi0200), .A2(pi1133), .ZN(new_n34993_));
  NAND3_X1   g31691(.A1(new_n30651_), .A2(new_n4959_), .A3(new_n34993_), .ZN(new_n34994_));
  NAND3_X1   g31692(.A1(new_n34992_), .A2(new_n34994_), .A3(pi0230), .ZN(new_n34995_));
  XNOR2_X1   g31693(.A1(new_n32800_), .A2(new_n34995_), .ZN(new_n34996_));
  NAND2_X1   g31694(.A1(new_n32090_), .A2(new_n2726_), .ZN(new_n34997_));
  AOI22_X1   g31695(.A1(new_n34996_), .A2(new_n34991_), .B1(new_n34940_), .B2(new_n34997_), .ZN(new_n34998_));
  NOR2_X1    g31696(.A1(new_n8683_), .A2(pi1135), .ZN(new_n34999_));
  XOR2_X1    g31697(.A1(new_n31936_), .A2(new_n34999_), .Z(new_n35000_));
  NAND2_X1   g31698(.A1(new_n35000_), .A2(pi1133), .ZN(new_n35001_));
  NAND2_X1   g31699(.A1(new_n35001_), .A2(pi0230), .ZN(new_n35002_));
  XNOR2_X1   g31700(.A1(new_n35002_), .A2(new_n34301_), .ZN(new_n35003_));
  OAI21_X1   g31701(.A1(new_n8549_), .A2(pi1135), .B(pi0299), .ZN(new_n35004_));
  AOI21_X1   g31702(.A1(new_n8549_), .A2(new_n34939_), .B(new_n35004_), .ZN(new_n35005_));
  NOR2_X1    g31703(.A1(new_n35001_), .A2(new_n27299_), .ZN(new_n35006_));
  XOR2_X1    g31704(.A1(new_n35006_), .A2(new_n35005_), .Z(new_n35007_));
  NAND4_X1   g31705(.A1(new_n34978_), .A2(pi1134), .A3(new_n35003_), .A4(new_n35007_), .ZN(new_n35008_));
  AOI21_X1   g31706(.A1(new_n34988_), .A2(new_n34998_), .B(new_n35008_), .ZN(new_n35009_));
  XOR2_X1    g31707(.A1(new_n34987_), .A2(new_n35009_), .Z(po0436));
  AOI21_X1   g31708(.A1(pi0211), .A2(new_n4785_), .B(new_n34305_), .ZN(new_n35011_));
  NOR3_X1    g31709(.A1(new_n35011_), .A2(new_n8683_), .A3(new_n4626_), .ZN(new_n35012_));
  XOR2_X1    g31710(.A1(new_n35012_), .A2(new_n30615_), .Z(new_n35013_));
  NAND4_X1   g31711(.A1(pi0199), .A2(pi0200), .A3(pi1135), .A4(pi1137), .ZN(new_n35014_));
  NAND2_X1   g31712(.A1(new_n35014_), .A2(new_n4785_), .ZN(new_n35015_));
  AOI21_X1   g31713(.A1(new_n35015_), .A2(pi0199), .B(new_n30557_), .ZN(new_n35016_));
  XOR2_X1    g31714(.A1(new_n32800_), .A2(new_n35016_), .Z(new_n35017_));
  INV_X1     g31715(.I(pi0914), .ZN(new_n35018_));
  NOR3_X1    g31716(.A1(new_n32541_), .A2(new_n35018_), .A3(new_n2726_), .ZN(new_n35019_));
  NOR3_X1    g31717(.A1(new_n32541_), .A2(pi0914), .A3(pi1091), .ZN(new_n35020_));
  OAI21_X1   g31718(.A1(new_n35019_), .A2(new_n35020_), .B(pi0280), .ZN(new_n35021_));
  NOR2_X1    g31719(.A1(new_n35021_), .A2(new_n8549_), .ZN(new_n35022_));
  OAI21_X1   g31720(.A1(new_n35022_), .A2(pi1137), .B(new_n34583_), .ZN(new_n35023_));
  NAND2_X1   g31721(.A1(new_n35023_), .A2(new_n12654_), .ZN(new_n35024_));
  INV_X1     g31722(.I(new_n35011_), .ZN(new_n35025_));
  NAND2_X1   g31723(.A1(new_n32529_), .A2(new_n35018_), .ZN(new_n35026_));
  XOR2_X1    g31724(.A1(new_n34237_), .A2(new_n35026_), .Z(new_n35027_));
  NAND2_X1   g31725(.A1(new_n35027_), .A2(pi0280), .ZN(new_n35028_));
  OAI21_X1   g31726(.A1(new_n35028_), .A2(new_n8683_), .B(new_n2726_), .ZN(new_n35029_));
  OAI21_X1   g31727(.A1(new_n34285_), .A2(pi1137), .B(pi0211), .ZN(new_n35030_));
  NAND2_X1   g31728(.A1(new_n35021_), .A2(new_n35030_), .ZN(new_n35031_));
  NAND3_X1   g31729(.A1(pi0200), .A2(pi1091), .A3(pi1136), .ZN(new_n35032_));
  NAND3_X1   g31730(.A1(new_n8555_), .A2(new_n4785_), .A3(pi1091), .ZN(new_n35033_));
  NAND2_X1   g31731(.A1(new_n35033_), .A2(new_n35032_), .ZN(new_n35034_));
  AOI21_X1   g31732(.A1(new_n35034_), .A2(pi1135), .B(pi0199), .ZN(new_n35035_));
  NAND4_X1   g31733(.A1(new_n35028_), .A2(new_n12654_), .A3(new_n35031_), .A4(new_n35035_), .ZN(new_n35036_));
  AOI21_X1   g31734(.A1(new_n35025_), .A2(new_n35029_), .B(new_n35036_), .ZN(new_n35037_));
  OR2_X2     g31735(.A1(new_n35037_), .A2(new_n35024_), .Z(new_n35038_));
  AOI21_X1   g31736(.A1(new_n35037_), .A2(new_n35024_), .B(pi0230), .ZN(new_n35039_));
  AOI22_X1   g31737(.A1(new_n35038_), .A2(new_n35039_), .B1(new_n35013_), .B2(new_n35017_), .ZN(po0437));
  NAND4_X1   g31738(.A1(new_n34581_), .A2(pi1139), .A3(new_n34582_), .A4(new_n34583_), .ZN(new_n35041_));
  NAND2_X1   g31739(.A1(new_n35041_), .A2(new_n4300_), .ZN(new_n35042_));
  INV_X1     g31740(.I(pi0281), .ZN(new_n35043_));
  INV_X1     g31741(.I(pi0830), .ZN(new_n35044_));
  NAND2_X1   g31742(.A1(new_n32529_), .A2(new_n35044_), .ZN(new_n35045_));
  XNOR2_X1   g31743(.A1(new_n34237_), .A2(new_n35045_), .ZN(new_n35046_));
  NOR3_X1    g31744(.A1(new_n35046_), .A2(new_n35043_), .A3(new_n33651_), .ZN(new_n35047_));
  NOR2_X1    g31745(.A1(new_n2726_), .A2(pi1138), .ZN(new_n35048_));
  XOR2_X1    g31746(.A1(new_n35048_), .A2(new_n34593_), .Z(new_n35049_));
  NOR2_X1    g31747(.A1(pi0211), .A2(pi1137), .ZN(new_n35050_));
  AOI21_X1   g31748(.A1(pi0211), .A2(new_n4465_), .B(new_n35050_), .ZN(new_n35051_));
  NAND3_X1   g31749(.A1(new_n35051_), .A2(pi1091), .A3(pi1137), .ZN(new_n35052_));
  OAI22_X1   g31750(.A1(new_n34591_), .A2(new_n32090_), .B1(new_n35049_), .B2(new_n35052_), .ZN(new_n35053_));
  NAND3_X1   g31751(.A1(new_n32540_), .A2(pi0830), .A3(pi1091), .ZN(new_n35054_));
  NAND3_X1   g31752(.A1(new_n32540_), .A2(new_n35044_), .A3(new_n2726_), .ZN(new_n35055_));
  AOI21_X1   g31753(.A1(new_n35054_), .A2(new_n35055_), .B(new_n35043_), .ZN(new_n35056_));
  AOI22_X1   g31754(.A1(new_n35042_), .A2(new_n35047_), .B1(new_n35053_), .B2(new_n35056_), .ZN(new_n35057_));
  NAND4_X1   g31755(.A1(pi0199), .A2(pi0200), .A3(pi1137), .A4(pi1139), .ZN(new_n35058_));
  AOI21_X1   g31756(.A1(new_n4465_), .A2(new_n35058_), .B(new_n34605_), .ZN(new_n35059_));
  NOR3_X1    g31757(.A1(new_n35051_), .A2(new_n8683_), .A3(new_n4300_), .ZN(new_n35060_));
  XOR2_X1    g31758(.A1(new_n35060_), .A2(new_n30615_), .Z(new_n35061_));
  NOR2_X1    g31759(.A1(new_n35061_), .A2(new_n12654_), .ZN(new_n35062_));
  OAI21_X1   g31760(.A1(new_n35059_), .A2(new_n35062_), .B(pi0230), .ZN(new_n35063_));
  OAI21_X1   g31761(.A1(new_n35057_), .A2(pi0230), .B(new_n35063_), .ZN(po0438));
  INV_X1     g31762(.I(new_n34582_), .ZN(new_n35065_));
  NOR2_X1    g31763(.A1(new_n34215_), .A2(pi1140), .ZN(new_n35066_));
  INV_X1     g31764(.I(pi0836), .ZN(new_n35067_));
  NOR3_X1    g31765(.A1(new_n32541_), .A2(new_n35067_), .A3(new_n2726_), .ZN(new_n35068_));
  NOR3_X1    g31766(.A1(new_n32541_), .A2(pi0836), .A3(pi1091), .ZN(new_n35069_));
  INV_X1     g31767(.I(pi0282), .ZN(new_n35070_));
  AOI21_X1   g31768(.A1(new_n33650_), .A2(pi1140), .B(new_n35070_), .ZN(new_n35071_));
  OAI21_X1   g31769(.A1(new_n35068_), .A2(new_n35069_), .B(new_n35071_), .ZN(new_n35072_));
  OAI22_X1   g31770(.A1(new_n35065_), .A2(new_n35072_), .B1(new_n8555_), .B2(new_n35066_), .ZN(new_n35073_));
  AOI21_X1   g31771(.A1(new_n35073_), .A2(new_n12654_), .B(new_n30557_), .ZN(new_n35074_));
  NOR2_X1    g31772(.A1(new_n2726_), .A2(pi1139), .ZN(new_n35075_));
  XOR2_X1    g31773(.A1(new_n35075_), .A2(new_n34593_), .Z(new_n35076_));
  NAND2_X1   g31774(.A1(new_n32529_), .A2(new_n35067_), .ZN(new_n35077_));
  XNOR2_X1   g31775(.A1(new_n34237_), .A2(new_n35077_), .ZN(new_n35078_));
  NOR2_X1    g31776(.A1(pi0211), .A2(pi1138), .ZN(new_n35079_));
  AOI21_X1   g31777(.A1(pi0211), .A2(new_n4300_), .B(new_n35079_), .ZN(new_n35080_));
  AOI21_X1   g31778(.A1(new_n35080_), .A2(pi1091), .B(new_n35070_), .ZN(new_n35081_));
  NAND2_X1   g31779(.A1(new_n32089_), .A2(new_n35081_), .ZN(new_n35082_));
  OAI22_X1   g31780(.A1(new_n35082_), .A2(new_n35078_), .B1(new_n4465_), .B2(new_n35076_), .ZN(new_n35083_));
  NOR4_X1    g31781(.A1(new_n8549_), .A2(new_n8555_), .A3(new_n4465_), .A4(new_n4141_), .ZN(new_n35084_));
  OAI21_X1   g31782(.A1(pi1139), .A2(new_n35084_), .B(new_n34604_), .ZN(new_n35085_));
  NOR4_X1    g31783(.A1(new_n35085_), .A2(pi0199), .A3(new_n30557_), .A4(new_n12655_), .ZN(new_n35088_));
  NAND2_X1   g31784(.A1(new_n35088_), .A2(new_n35083_), .ZN(new_n35089_));
  XNOR2_X1   g31785(.A1(new_n35089_), .A2(new_n35074_), .ZN(po0439));
  NAND2_X1   g31786(.A1(pi1147), .A2(pi1148), .ZN(new_n35091_));
  NAND2_X1   g31787(.A1(new_n34530_), .A2(pi1148), .ZN(new_n35092_));
  XOR2_X1    g31788(.A1(new_n35092_), .A2(new_n35091_), .Z(new_n35093_));
  NAND2_X1   g31789(.A1(new_n35093_), .A2(new_n34466_), .ZN(new_n35094_));
  NAND2_X1   g31790(.A1(new_n34508_), .A2(pi1147), .ZN(new_n35095_));
  XNOR2_X1   g31791(.A1(new_n35095_), .A2(new_n35091_), .ZN(new_n35096_));
  NOR2_X1    g31792(.A1(new_n35096_), .A2(new_n34541_), .ZN(new_n35097_));
  NAND2_X1   g31793(.A1(new_n32771_), .A2(new_n31941_), .ZN(new_n35098_));
  NAND2_X1   g31794(.A1(new_n34537_), .A2(pi1148), .ZN(new_n35099_));
  XNOR2_X1   g31795(.A1(new_n35099_), .A2(new_n35091_), .ZN(new_n35100_));
  NOR2_X1    g31796(.A1(new_n35100_), .A2(new_n34540_), .ZN(new_n35101_));
  OAI21_X1   g31797(.A1(new_n35097_), .A2(new_n35098_), .B(new_n35101_), .ZN(new_n35102_));
  NAND3_X1   g31798(.A1(new_n35102_), .A2(new_n35094_), .A3(new_n31941_), .ZN(new_n35103_));
  NAND2_X1   g31799(.A1(new_n34473_), .A2(pi1147), .ZN(new_n35104_));
  XNOR2_X1   g31800(.A1(new_n35104_), .A2(new_n35091_), .ZN(new_n35105_));
  NOR2_X1    g31801(.A1(new_n35105_), .A2(new_n34526_), .ZN(new_n35106_));
  AOI21_X1   g31802(.A1(new_n33806_), .A2(pi1147), .B(pi1148), .ZN(new_n35107_));
  OAI21_X1   g31803(.A1(new_n31941_), .A2(new_n34681_), .B(new_n35107_), .ZN(new_n35108_));
  NOR2_X1    g31804(.A1(new_n34714_), .A2(pi1149), .ZN(new_n35109_));
  NAND2_X1   g31805(.A1(new_n34569_), .A2(pi1147), .ZN(new_n35110_));
  OAI21_X1   g31806(.A1(new_n35109_), .A2(new_n35110_), .B(new_n31953_), .ZN(new_n35111_));
  AOI21_X1   g31807(.A1(new_n35108_), .A2(pi0230), .B(new_n35111_), .ZN(new_n35112_));
  OAI21_X1   g31808(.A1(new_n34817_), .A2(new_n31940_), .B(new_n34712_), .ZN(new_n35113_));
  OAI21_X1   g31809(.A1(new_n35112_), .A2(new_n35113_), .B(new_n30557_), .ZN(new_n35114_));
  AOI21_X1   g31810(.A1(new_n35103_), .A2(new_n35106_), .B(new_n35114_), .ZN(new_n35115_));
  NOR2_X1    g31811(.A1(new_n34520_), .A2(new_n31940_), .ZN(new_n35116_));
  XNOR2_X1   g31812(.A1(new_n35116_), .A2(new_n32084_), .ZN(new_n35117_));
  NAND2_X1   g31813(.A1(new_n35117_), .A2(new_n34489_), .ZN(new_n35118_));
  NOR2_X1    g31814(.A1(pi0283), .A2(pi1148), .ZN(new_n35119_));
  NAND2_X1   g31815(.A1(new_n34552_), .A2(pi1149), .ZN(new_n35120_));
  XOR2_X1    g31816(.A1(new_n35120_), .A2(new_n32084_), .Z(new_n35121_));
  NAND2_X1   g31817(.A1(new_n35121_), .A2(new_n34706_), .ZN(new_n35122_));
  AOI21_X1   g31818(.A1(new_n35118_), .A2(new_n35119_), .B(new_n35122_), .ZN(new_n35123_));
  NOR2_X1    g31819(.A1(new_n34495_), .A2(new_n31940_), .ZN(new_n35124_));
  XOR2_X1    g31820(.A1(new_n35124_), .A2(new_n32084_), .Z(new_n35125_));
  OAI21_X1   g31821(.A1(new_n35125_), .A2(new_n34705_), .B(new_n31953_), .ZN(new_n35126_));
  NOR2_X1    g31822(.A1(new_n35123_), .A2(new_n35126_), .ZN(new_n35127_));
  NAND2_X1   g31823(.A1(new_n34547_), .A2(pi1149), .ZN(new_n35128_));
  XNOR2_X1   g31824(.A1(new_n35128_), .A2(new_n32084_), .ZN(new_n35129_));
  NOR4_X1    g31825(.A1(new_n35127_), .A2(new_n34501_), .A3(new_n35115_), .A4(new_n35129_), .ZN(po0440));
  NOR2_X1    g31826(.A1(new_n32092_), .A2(new_n34029_), .ZN(new_n35131_));
  NOR3_X1    g31827(.A1(new_n34029_), .A2(new_n3682_), .A3(new_n3650_), .ZN(new_n35132_));
  XOR2_X1    g31828(.A1(new_n35131_), .A2(new_n35132_), .Z(po0441));
  NAND2_X1   g31829(.A1(new_n8532_), .A2(new_n3291_), .ZN(new_n35134_));
  NOR3_X1    g31830(.A1(new_n35134_), .A2(new_n6663_), .A3(new_n9863_), .ZN(new_n35135_));
  NAND2_X1   g31831(.A1(new_n35135_), .A2(new_n6666_), .ZN(new_n35136_));
  NOR3_X1    g31832(.A1(new_n6407_), .A2(pi0286), .A3(pi0288), .ZN(new_n35137_));
  AOI21_X1   g31833(.A1(new_n35137_), .A2(new_n6665_), .B(pi0285), .ZN(new_n35138_));
  OR3_X2     g31834(.A1(new_n35136_), .A2(new_n7240_), .A3(new_n35138_), .Z(new_n35139_));
  INV_X1     g31835(.I(new_n35136_), .ZN(new_n35140_));
  NOR2_X1    g31836(.A1(new_n35140_), .A2(po1038), .ZN(new_n35141_));
  NOR2_X1    g31837(.A1(new_n35140_), .A2(new_n6662_), .ZN(new_n35142_));
  NOR2_X1    g31838(.A1(new_n35136_), .A2(pi0285), .ZN(new_n35143_));
  OAI22_X1   g31839(.A1(new_n35134_), .A2(new_n35141_), .B1(new_n35142_), .B2(new_n35143_), .ZN(new_n35144_));
  AOI21_X1   g31840(.A1(new_n35144_), .A2(new_n35139_), .B(pi0793), .ZN(po0442));
  INV_X1     g31841(.I(new_n35134_), .ZN(new_n35146_));
  NOR3_X1    g31842(.A1(new_n35146_), .A2(new_n6663_), .A3(new_n6664_), .ZN(new_n35147_));
  AOI21_X1   g31843(.A1(pi0286), .A2(pi0288), .B(new_n35134_), .ZN(new_n35148_));
  OAI21_X1   g31844(.A1(new_n35147_), .A2(new_n35148_), .B(new_n9863_), .ZN(new_n35149_));
  NOR2_X1    g31845(.A1(pi0285), .A2(pi0288), .ZN(new_n35150_));
  AOI21_X1   g31846(.A1(new_n35150_), .A2(new_n6665_), .B(new_n6663_), .ZN(new_n35151_));
  NAND2_X1   g31847(.A1(new_n35151_), .A2(pi0286), .ZN(new_n35152_));
  XOR2_X1    g31848(.A1(new_n6407_), .A2(new_n35152_), .Z(new_n35153_));
  AOI21_X1   g31849(.A1(new_n35146_), .A2(new_n35153_), .B(po1038), .ZN(new_n35154_));
  INV_X1     g31850(.I(pi0793), .ZN(new_n35155_));
  NAND2_X1   g31851(.A1(po1038), .A2(pi0286), .ZN(new_n35156_));
  XOR2_X1    g31852(.A1(new_n35156_), .A2(new_n35151_), .Z(new_n35157_));
  OAI21_X1   g31853(.A1(new_n35157_), .A2(new_n6407_), .B(new_n35155_), .ZN(new_n35158_));
  AOI21_X1   g31854(.A1(new_n35149_), .A2(new_n35154_), .B(new_n35158_), .ZN(po0443));
  AOI21_X1   g31855(.A1(new_n5401_), .A2(pi0457), .B(pi0332), .ZN(po0444));
  NAND2_X1   g31856(.A1(new_n6407_), .A2(new_n6664_), .ZN(new_n35161_));
  OAI21_X1   g31857(.A1(new_n6407_), .A2(new_n35151_), .B(new_n35161_), .ZN(new_n35162_));
  NOR2_X1    g31858(.A1(new_n35134_), .A2(po1038), .ZN(po0637));
  XOR2_X1    g31859(.A1(po0637), .A2(new_n35162_), .Z(new_n35164_));
  NOR2_X1    g31860(.A1(new_n35164_), .A2(pi0793), .ZN(po0445));
  NAND2_X1   g31861(.A1(new_n9863_), .A2(new_n6663_), .ZN(new_n35166_));
  NOR2_X1    g31862(.A1(new_n6665_), .A2(pi0288), .ZN(new_n35167_));
  NOR4_X1    g31863(.A1(new_n35146_), .A2(new_n6662_), .A3(new_n35166_), .A4(new_n35167_), .ZN(new_n35168_));
  OR2_X2     g31864(.A1(new_n35168_), .A2(new_n6665_), .Z(new_n35169_));
  AOI21_X1   g31865(.A1(new_n35168_), .A2(new_n6665_), .B(new_n35135_), .ZN(new_n35170_));
  OAI21_X1   g31866(.A1(pi0289), .A2(new_n7240_), .B(new_n35137_), .ZN(new_n35171_));
  OAI21_X1   g31867(.A1(new_n35171_), .A2(new_n6662_), .B(new_n35155_), .ZN(new_n35172_));
  NAND3_X1   g31868(.A1(new_n35172_), .A2(pi0288), .A3(po1038), .ZN(new_n35173_));
  AOI21_X1   g31869(.A1(new_n35169_), .A2(new_n35170_), .B(new_n35173_), .ZN(po0446));
  INV_X1     g31870(.I(pi1048), .ZN(new_n35175_));
  NAND2_X1   g31871(.A1(pi0290), .A2(pi0476), .ZN(new_n35176_));
  OAI21_X1   g31872(.A1(pi0476), .A2(new_n35175_), .B(new_n35176_), .ZN(po0447));
  INV_X1     g31873(.I(pi1049), .ZN(new_n35178_));
  NAND2_X1   g31874(.A1(pi0291), .A2(pi0476), .ZN(new_n35179_));
  OAI21_X1   g31875(.A1(pi0476), .A2(new_n35178_), .B(new_n35179_), .ZN(po0448));
  INV_X1     g31876(.I(pi1084), .ZN(new_n35181_));
  NAND2_X1   g31877(.A1(pi0292), .A2(pi0476), .ZN(new_n35182_));
  OAI21_X1   g31878(.A1(pi0476), .A2(new_n35181_), .B(new_n35182_), .ZN(po0449));
  INV_X1     g31879(.I(pi1059), .ZN(new_n35184_));
  NAND2_X1   g31880(.A1(pi0293), .A2(pi0476), .ZN(new_n35185_));
  OAI21_X1   g31881(.A1(pi0476), .A2(new_n35184_), .B(new_n35185_), .ZN(po0450));
  INV_X1     g31882(.I(pi1072), .ZN(new_n35187_));
  NAND2_X1   g31883(.A1(pi0294), .A2(pi0476), .ZN(new_n35188_));
  OAI21_X1   g31884(.A1(pi0476), .A2(new_n35187_), .B(new_n35188_), .ZN(po0451));
  NAND2_X1   g31885(.A1(pi0295), .A2(pi0476), .ZN(new_n35190_));
  OAI21_X1   g31886(.A1(pi0476), .A2(new_n33607_), .B(new_n35190_), .ZN(po0452));
  NAND2_X1   g31887(.A1(pi0296), .A2(pi0476), .ZN(new_n35192_));
  OAI21_X1   g31888(.A1(pi0476), .A2(new_n34021_), .B(new_n35192_), .ZN(po0453));
  NAND2_X1   g31889(.A1(pi0297), .A2(pi0476), .ZN(new_n35194_));
  OAI21_X1   g31890(.A1(pi0476), .A2(new_n34014_), .B(new_n35194_), .ZN(po0454));
  NAND2_X1   g31891(.A1(pi0298), .A2(pi0478), .ZN(new_n35196_));
  OAI21_X1   g31892(.A1(pi0478), .A2(new_n34014_), .B(new_n35196_), .ZN(po0455));
  NOR2_X1    g31893(.A1(new_n10472_), .A2(new_n3115_), .ZN(new_n35198_));
  NAND4_X1   g31894(.A1(new_n8529_), .A2(pi0054), .A3(new_n2902_), .A4(new_n3160_), .ZN(new_n35199_));
  XOR2_X1    g31895(.A1(new_n35198_), .A2(new_n35199_), .Z(new_n35200_));
  AOI22_X1   g31896(.A1(new_n7330_), .A2(new_n9135_), .B1(pi0039), .B2(new_n9129_), .ZN(new_n35201_));
  NOR2_X1    g31897(.A1(new_n35200_), .A2(new_n35201_), .ZN(po0456));
  NAND3_X1   g31898(.A1(new_n8224_), .A2(pi0312), .A3(new_n5546_), .ZN(new_n35203_));
  XOR2_X1    g31899(.A1(new_n35203_), .A2(pi0300), .Z(new_n35204_));
  NAND2_X1   g31900(.A1(new_n35204_), .A2(new_n3258_), .ZN(po0457));
  NOR2_X1    g31901(.A1(new_n35203_), .A2(pi0300), .ZN(new_n35206_));
  XOR2_X1    g31902(.A1(new_n35206_), .A2(pi0301), .Z(new_n35207_));
  NOR2_X1    g31903(.A1(new_n35207_), .A2(pi0055), .ZN(po0458));
  NOR2_X1    g31904(.A1(new_n12654_), .A2(new_n3368_), .ZN(new_n35209_));
  OAI21_X1   g31905(.A1(pi0222), .A2(pi0223), .B(pi0937), .ZN(new_n35210_));
  NAND2_X1   g31906(.A1(new_n7240_), .A2(new_n5296_), .ZN(new_n35211_));
  NAND2_X1   g31907(.A1(new_n3386_), .A2(pi0273), .ZN(new_n35212_));
  AOI21_X1   g31908(.A1(new_n35211_), .A2(new_n35210_), .B(new_n35212_), .ZN(new_n35213_));
  OAI21_X1   g31909(.A1(new_n35213_), .A2(new_n35209_), .B(pi0237), .ZN(new_n35214_));
  NOR2_X1    g31910(.A1(new_n6453_), .A2(new_n3058_), .ZN(new_n35215_));
  NAND2_X1   g31911(.A1(new_n35215_), .A2(pi0273), .ZN(new_n35216_));
  NOR2_X1    g31912(.A1(new_n3536_), .A2(new_n3011_), .ZN(new_n35217_));
  NAND2_X1   g31913(.A1(new_n35217_), .A2(pi0937), .ZN(new_n35218_));
  NAND2_X1   g31914(.A1(new_n35216_), .A2(new_n35218_), .ZN(new_n35219_));
  AOI22_X1   g31915(.A1(new_n35219_), .A2(new_n35213_), .B1(new_n3091_), .B2(new_n12654_), .ZN(new_n35220_));
  INV_X1     g31916(.I(new_n35211_), .ZN(new_n35221_));
  NOR2_X1    g31917(.A1(new_n12654_), .A2(new_n5281_), .ZN(new_n35222_));
  NOR2_X1    g31918(.A1(new_n35221_), .A2(new_n35222_), .ZN(new_n35223_));
  NAND2_X1   g31919(.A1(new_n35223_), .A2(pi1148), .ZN(new_n35224_));
  AOI21_X1   g31920(.A1(new_n35220_), .A2(new_n35214_), .B(new_n35224_), .ZN(po0459));
  NAND2_X1   g31921(.A1(pi0303), .A2(pi0478), .ZN(new_n35226_));
  OAI21_X1   g31922(.A1(pi0478), .A2(new_n35178_), .B(new_n35226_), .ZN(po0460));
  NAND2_X1   g31923(.A1(pi0304), .A2(pi0478), .ZN(new_n35228_));
  OAI21_X1   g31924(.A1(pi0478), .A2(new_n35175_), .B(new_n35228_), .ZN(po0461));
  NAND2_X1   g31925(.A1(pi0305), .A2(pi0478), .ZN(new_n35230_));
  OAI21_X1   g31926(.A1(pi0478), .A2(new_n35181_), .B(new_n35230_), .ZN(po0462));
  NAND2_X1   g31927(.A1(pi0306), .A2(pi0478), .ZN(new_n35232_));
  OAI21_X1   g31928(.A1(pi0478), .A2(new_n35184_), .B(new_n35232_), .ZN(po0463));
  NAND2_X1   g31929(.A1(pi0307), .A2(pi0478), .ZN(new_n35234_));
  OAI21_X1   g31930(.A1(pi0478), .A2(new_n33607_), .B(new_n35234_), .ZN(po0464));
  NAND2_X1   g31931(.A1(pi0308), .A2(pi0478), .ZN(new_n35236_));
  OAI21_X1   g31932(.A1(pi0478), .A2(new_n34021_), .B(new_n35236_), .ZN(po0465));
  NAND2_X1   g31933(.A1(pi0309), .A2(pi0478), .ZN(new_n35238_));
  OAI21_X1   g31934(.A1(pi0478), .A2(new_n35187_), .B(new_n35238_), .ZN(po0466));
  NAND4_X1   g31935(.A1(new_n3121_), .A2(pi0216), .A3(pi0271), .A4(pi0934), .ZN(new_n35240_));
  AOI21_X1   g31936(.A1(new_n35240_), .A2(new_n3121_), .B(new_n3111_), .ZN(new_n35241_));
  NOR4_X1    g31937(.A1(new_n12654_), .A2(new_n3312_), .A3(new_n5281_), .A4(new_n35241_), .ZN(new_n35242_));
  NOR2_X1    g31938(.A1(new_n3099_), .A2(pi0271), .ZN(new_n35243_));
  NAND2_X1   g31939(.A1(new_n3101_), .A2(pi0934), .ZN(new_n35244_));
  XOR2_X1    g31940(.A1(new_n35244_), .A2(new_n35243_), .Z(new_n35245_));
  NOR2_X1    g31941(.A1(new_n35211_), .A2(new_n35245_), .ZN(new_n35246_));
  OAI21_X1   g31942(.A1(new_n35242_), .A2(new_n35209_), .B(new_n35246_), .ZN(new_n35247_));
  NAND2_X1   g31943(.A1(new_n35222_), .A2(new_n35241_), .ZN(new_n35248_));
  NAND2_X1   g31944(.A1(new_n12654_), .A2(new_n3128_), .ZN(new_n35249_));
  NAND2_X1   g31945(.A1(new_n35221_), .A2(new_n35245_), .ZN(new_n35250_));
  NAND4_X1   g31946(.A1(new_n35250_), .A2(pi1147), .A3(new_n35248_), .A4(new_n35249_), .ZN(new_n35251_));
  AOI22_X1   g31947(.A1(new_n35221_), .A2(new_n3312_), .B1(new_n3091_), .B2(new_n35222_), .ZN(new_n35252_));
  INV_X1     g31948(.I(new_n35252_), .ZN(new_n35253_));
  NOR2_X1    g31949(.A1(new_n35253_), .A2(pi1147), .ZN(new_n35254_));
  AOI21_X1   g31950(.A1(new_n35254_), .A2(new_n35251_), .B(new_n35247_), .ZN(new_n35255_));
  NOR3_X1    g31951(.A1(new_n35221_), .A2(new_n31940_), .A3(new_n35222_), .ZN(new_n35256_));
  OAI21_X1   g31952(.A1(new_n35247_), .A2(new_n35256_), .B(new_n27639_), .ZN(new_n35257_));
  OAI21_X1   g31953(.A1(new_n35255_), .A2(new_n27639_), .B(new_n35257_), .ZN(po0467));
  NAND2_X1   g31954(.A1(pi0055), .A2(pi0311), .ZN(new_n35259_));
  XOR2_X1    g31955(.A1(new_n35259_), .A2(pi0301), .Z(new_n35260_));
  NOR3_X1    g31956(.A1(new_n35203_), .A2(pi0300), .A3(new_n35260_), .ZN(po0468));
  NAND3_X1   g31957(.A1(new_n8224_), .A2(pi0057), .A3(pi0312), .ZN(new_n35262_));
  OAI21_X1   g31958(.A1(new_n35262_), .A2(pi0059), .B(new_n3258_), .ZN(new_n35263_));
  AOI21_X1   g31959(.A1(pi0059), .A2(new_n35262_), .B(new_n35263_), .ZN(po0469));
  NAND2_X1   g31960(.A1(new_n8464_), .A2(new_n10494_), .ZN(new_n35265_));
  AOI21_X1   g31961(.A1(new_n10500_), .A2(po0740), .B(new_n8292_), .ZN(new_n35266_));
  NAND3_X1   g31962(.A1(new_n35265_), .A2(new_n35266_), .A3(po1110), .ZN(new_n35267_));
  OAI21_X1   g31963(.A1(pi0313), .A2(po1110), .B(new_n35267_), .ZN(po0470));
  NOR2_X1    g31964(.A1(new_n11208_), .A2(new_n3133_), .ZN(new_n35269_));
  XNOR2_X1   g31965(.A1(new_n35269_), .A2(new_n3417_), .ZN(new_n35270_));
  AOI21_X1   g31966(.A1(new_n5765_), .A2(new_n7330_), .B(new_n11417_), .ZN(new_n35271_));
  NAND2_X1   g31967(.A1(new_n10299_), .A2(new_n3206_), .ZN(new_n35272_));
  NAND2_X1   g31968(.A1(new_n11315_), .A2(new_n11557_), .ZN(new_n35273_));
  AOI21_X1   g31969(.A1(new_n3133_), .A2(new_n11175_), .B(new_n35273_), .ZN(new_n35274_));
  OAI21_X1   g31970(.A1(new_n35271_), .A2(new_n35272_), .B(new_n35274_), .ZN(new_n35275_));
  AOI21_X1   g31971(.A1(new_n35270_), .A2(new_n12340_), .B(new_n35275_), .ZN(po0471));
  INV_X1     g31972(.I(pi1080), .ZN(new_n35277_));
  INV_X1     g31973(.I(pi0340), .ZN(new_n35278_));
  NAND3_X1   g31974(.A1(new_n35146_), .A2(new_n35278_), .A3(new_n7240_), .ZN(new_n35279_));
  NAND2_X1   g31975(.A1(new_n35279_), .A2(pi0315), .ZN(new_n35280_));
  OAI21_X1   g31976(.A1(new_n35277_), .A2(new_n35279_), .B(new_n35280_), .ZN(po0472));
  INV_X1     g31977(.I(pi1047), .ZN(new_n35282_));
  NAND2_X1   g31978(.A1(new_n35279_), .A2(pi0316), .ZN(new_n35283_));
  OAI21_X1   g31979(.A1(new_n35282_), .A2(new_n35279_), .B(new_n35283_), .ZN(po0473));
  INV_X1     g31980(.I(po0637), .ZN(new_n35285_));
  NOR2_X1    g31981(.A1(new_n35285_), .A2(pi0330), .ZN(new_n35286_));
  NAND2_X1   g31982(.A1(new_n35286_), .A2(pi1078), .ZN(new_n35287_));
  OAI21_X1   g31983(.A1(new_n6679_), .A2(new_n35286_), .B(new_n35287_), .ZN(po0474));
  INV_X1     g31984(.I(pi1074), .ZN(new_n35289_));
  INV_X1     g31985(.I(pi0341), .ZN(new_n35290_));
  NAND3_X1   g31986(.A1(new_n35146_), .A2(new_n35290_), .A3(new_n7240_), .ZN(new_n35291_));
  NAND2_X1   g31987(.A1(new_n35291_), .A2(pi0318), .ZN(new_n35292_));
  OAI21_X1   g31988(.A1(new_n35289_), .A2(new_n35291_), .B(new_n35292_), .ZN(po0475));
  NAND2_X1   g31989(.A1(new_n35291_), .A2(pi0319), .ZN(new_n35294_));
  OAI21_X1   g31990(.A1(new_n35187_), .A2(new_n35291_), .B(new_n35294_), .ZN(po0476));
  NAND2_X1   g31991(.A1(new_n35279_), .A2(pi0320), .ZN(new_n35296_));
  OAI21_X1   g31992(.A1(new_n35175_), .A2(new_n35279_), .B(new_n35296_), .ZN(po0477));
  INV_X1     g31993(.I(pi1058), .ZN(new_n35298_));
  NAND2_X1   g31994(.A1(new_n35279_), .A2(pi0321), .ZN(new_n35299_));
  OAI21_X1   g31995(.A1(new_n35298_), .A2(new_n35279_), .B(new_n35299_), .ZN(po0478));
  INV_X1     g31996(.I(pi1051), .ZN(new_n35301_));
  NAND2_X1   g31997(.A1(new_n35279_), .A2(pi0322), .ZN(new_n35302_));
  OAI21_X1   g31998(.A1(new_n35301_), .A2(new_n35279_), .B(new_n35302_), .ZN(po0479));
  NAND2_X1   g31999(.A1(new_n35279_), .A2(pi0323), .ZN(new_n35304_));
  OAI21_X1   g32000(.A1(new_n33997_), .A2(new_n35279_), .B(new_n35304_), .ZN(po0480));
  INV_X1     g32001(.I(pi1086), .ZN(new_n35306_));
  NAND2_X1   g32002(.A1(new_n35291_), .A2(pi0324), .ZN(new_n35307_));
  OAI21_X1   g32003(.A1(new_n35306_), .A2(new_n35291_), .B(new_n35307_), .ZN(po0481));
  INV_X1     g32004(.I(pi1063), .ZN(new_n35309_));
  NAND2_X1   g32005(.A1(new_n35291_), .A2(pi0325), .ZN(new_n35310_));
  OAI21_X1   g32006(.A1(new_n35309_), .A2(new_n35291_), .B(new_n35310_), .ZN(po0482));
  INV_X1     g32007(.I(pi1057), .ZN(new_n35312_));
  NAND2_X1   g32008(.A1(new_n35291_), .A2(pi0326), .ZN(new_n35313_));
  OAI21_X1   g32009(.A1(new_n35312_), .A2(new_n35291_), .B(new_n35313_), .ZN(po0483));
  NAND2_X1   g32010(.A1(new_n35279_), .A2(pi0327), .ZN(new_n35315_));
  OAI21_X1   g32011(.A1(new_n34023_), .A2(new_n35279_), .B(new_n35315_), .ZN(po0484));
  NAND2_X1   g32012(.A1(new_n35291_), .A2(pi0328), .ZN(new_n35317_));
  OAI21_X1   g32013(.A1(new_n35298_), .A2(new_n35291_), .B(new_n35317_), .ZN(po0485));
  INV_X1     g32014(.I(pi1043), .ZN(new_n35319_));
  NAND2_X1   g32015(.A1(new_n35291_), .A2(pi0329), .ZN(new_n35320_));
  OAI21_X1   g32016(.A1(new_n35319_), .A2(new_n35291_), .B(new_n35320_), .ZN(po0486));
  INV_X1     g32017(.I(pi0330), .ZN(new_n35322_));
  NOR2_X1    g32018(.A1(new_n2985_), .A2(new_n2979_), .ZN(new_n35323_));
  OAI21_X1   g32019(.A1(new_n35146_), .A2(new_n35322_), .B(new_n35323_), .ZN(new_n35324_));
  AOI21_X1   g32020(.A1(pi0340), .A2(new_n35146_), .B(new_n35324_), .ZN(new_n35325_));
  INV_X1     g32021(.I(new_n35323_), .ZN(new_n35326_));
  NOR2_X1    g32022(.A1(new_n7240_), .A2(new_n35326_), .ZN(new_n35327_));
  XNOR2_X1   g32023(.A1(new_n35325_), .A2(new_n35327_), .ZN(new_n35328_));
  NOR2_X1    g32024(.A1(new_n35328_), .A2(new_n35322_), .ZN(po0487));
  INV_X1     g32025(.I(pi0331), .ZN(new_n35330_));
  OAI21_X1   g32026(.A1(new_n35146_), .A2(new_n35330_), .B(new_n35323_), .ZN(new_n35331_));
  AOI21_X1   g32027(.A1(pi0341), .A2(new_n35146_), .B(new_n35331_), .ZN(new_n35332_));
  XNOR2_X1   g32028(.A1(new_n35332_), .A2(new_n35327_), .ZN(new_n35333_));
  NOR2_X1    g32029(.A1(new_n35333_), .A2(new_n35330_), .ZN(po0488));
  NOR3_X1    g32030(.A1(new_n8946_), .A2(pi0332), .A3(new_n8290_), .ZN(new_n35335_));
  NAND2_X1   g32031(.A1(new_n7350_), .A2(new_n2955_), .ZN(new_n35336_));
  NAND2_X1   g32032(.A1(new_n6367_), .A2(pi0070), .ZN(new_n35337_));
  AOI21_X1   g32033(.A1(new_n8946_), .A2(new_n35337_), .B(new_n10280_), .ZN(new_n35338_));
  OAI21_X1   g32034(.A1(new_n35336_), .A2(new_n35335_), .B(new_n35338_), .ZN(new_n35339_));
  NAND2_X1   g32035(.A1(new_n35339_), .A2(pi0039), .ZN(new_n35340_));
  XOR2_X1    g32036(.A1(new_n35340_), .A2(new_n4368_), .Z(new_n35341_));
  NAND2_X1   g32037(.A1(new_n35341_), .A2(new_n8447_), .ZN(new_n35342_));
  AOI21_X1   g32038(.A1(new_n35342_), .A2(new_n8345_), .B(new_n6281_), .ZN(po0489));
  NAND2_X1   g32039(.A1(new_n35291_), .A2(pi0333), .ZN(new_n35344_));
  OAI21_X1   g32040(.A1(new_n34023_), .A2(new_n35291_), .B(new_n35344_), .ZN(po0490));
  NAND2_X1   g32041(.A1(new_n35291_), .A2(pi0334), .ZN(new_n35346_));
  OAI21_X1   g32042(.A1(new_n33997_), .A2(new_n35291_), .B(new_n35346_), .ZN(po0491));
  NAND2_X1   g32043(.A1(new_n35291_), .A2(pi0335), .ZN(new_n35348_));
  OAI21_X1   g32044(.A1(new_n34009_), .A2(new_n35291_), .B(new_n35348_), .ZN(po0492));
  INV_X1     g32045(.I(pi0336), .ZN(new_n35350_));
  NAND2_X1   g32046(.A1(new_n35286_), .A2(pi1070), .ZN(new_n35351_));
  OAI21_X1   g32047(.A1(new_n35350_), .A2(new_n35286_), .B(new_n35351_), .ZN(po0493));
  INV_X1     g32048(.I(pi0337), .ZN(new_n35353_));
  NAND2_X1   g32049(.A1(new_n35286_), .A2(pi1044), .ZN(new_n35354_));
  OAI21_X1   g32050(.A1(new_n35353_), .A2(new_n35286_), .B(new_n35354_), .ZN(po0494));
  INV_X1     g32051(.I(pi0338), .ZN(new_n35356_));
  NAND2_X1   g32052(.A1(new_n35286_), .A2(pi1072), .ZN(new_n35357_));
  OAI21_X1   g32053(.A1(new_n35356_), .A2(new_n35286_), .B(new_n35357_), .ZN(po0495));
  NAND2_X1   g32054(.A1(new_n35286_), .A2(pi1086), .ZN(new_n35359_));
  OAI21_X1   g32055(.A1(new_n6701_), .A2(new_n35286_), .B(new_n35359_), .ZN(po0496));
  AOI21_X1   g32056(.A1(new_n35278_), .A2(new_n35326_), .B(new_n7240_), .ZN(po0497));
  NAND3_X1   g32057(.A1(po0637), .A2(pi0330), .A3(new_n35323_), .ZN(new_n35364_));
  NAND3_X1   g32058(.A1(new_n35285_), .A2(new_n35322_), .A3(new_n35323_), .ZN(new_n35365_));
  AOI21_X1   g32059(.A1(new_n35365_), .A2(new_n35364_), .B(new_n35290_), .ZN(po0498));
  NAND2_X1   g32060(.A1(new_n35279_), .A2(pi0342), .ZN(new_n35367_));
  OAI21_X1   g32061(.A1(new_n35178_), .A2(new_n35279_), .B(new_n35367_), .ZN(po0499));
  NAND2_X1   g32062(.A1(new_n35279_), .A2(pi0343), .ZN(new_n35369_));
  OAI21_X1   g32063(.A1(new_n34003_), .A2(new_n35279_), .B(new_n35369_), .ZN(po0500));
  NAND2_X1   g32064(.A1(new_n35279_), .A2(pi0344), .ZN(new_n35371_));
  OAI21_X1   g32065(.A1(new_n34009_), .A2(new_n35279_), .B(new_n35371_), .ZN(po0501));
  NAND2_X1   g32066(.A1(new_n35279_), .A2(pi0345), .ZN(new_n35373_));
  OAI21_X1   g32067(.A1(new_n33609_), .A2(new_n35279_), .B(new_n35373_), .ZN(po0502));
  NAND2_X1   g32068(.A1(new_n35279_), .A2(pi0346), .ZN(new_n35375_));
  OAI21_X1   g32069(.A1(new_n34016_), .A2(new_n35279_), .B(new_n35375_), .ZN(po0503));
  INV_X1     g32070(.I(pi1055), .ZN(new_n35377_));
  NAND2_X1   g32071(.A1(new_n35279_), .A2(pi0347), .ZN(new_n35378_));
  OAI21_X1   g32072(.A1(new_n35377_), .A2(new_n35279_), .B(new_n35378_), .ZN(po0504));
  INV_X1     g32073(.I(pi1087), .ZN(new_n35380_));
  NAND2_X1   g32074(.A1(new_n35279_), .A2(pi0348), .ZN(new_n35381_));
  OAI21_X1   g32075(.A1(new_n35380_), .A2(new_n35279_), .B(new_n35381_), .ZN(po0505));
  NAND2_X1   g32076(.A1(new_n35279_), .A2(pi0349), .ZN(new_n35383_));
  OAI21_X1   g32077(.A1(new_n35319_), .A2(new_n35279_), .B(new_n35383_), .ZN(po0506));
  INV_X1     g32078(.I(pi1035), .ZN(new_n35385_));
  NAND2_X1   g32079(.A1(new_n35279_), .A2(pi0350), .ZN(new_n35386_));
  OAI21_X1   g32080(.A1(new_n35385_), .A2(new_n35279_), .B(new_n35386_), .ZN(po0507));
  INV_X1     g32081(.I(pi1079), .ZN(new_n35388_));
  NAND2_X1   g32082(.A1(new_n35279_), .A2(pi0351), .ZN(new_n35389_));
  OAI21_X1   g32083(.A1(new_n35388_), .A2(new_n35279_), .B(new_n35389_), .ZN(po0508));
  INV_X1     g32084(.I(pi1078), .ZN(new_n35391_));
  NAND2_X1   g32085(.A1(new_n35279_), .A2(pi0352), .ZN(new_n35392_));
  OAI21_X1   g32086(.A1(new_n35391_), .A2(new_n35279_), .B(new_n35392_), .ZN(po0509));
  NAND2_X1   g32087(.A1(new_n35279_), .A2(pi0353), .ZN(new_n35394_));
  OAI21_X1   g32088(.A1(new_n35309_), .A2(new_n35279_), .B(new_n35394_), .ZN(po0510));
  INV_X1     g32089(.I(pi1045), .ZN(new_n35396_));
  NAND2_X1   g32090(.A1(new_n35279_), .A2(pi0354), .ZN(new_n35397_));
  OAI21_X1   g32091(.A1(new_n35396_), .A2(new_n35279_), .B(new_n35397_), .ZN(po0511));
  NAND2_X1   g32092(.A1(new_n35279_), .A2(pi0355), .ZN(new_n35399_));
  OAI21_X1   g32093(.A1(new_n35181_), .A2(new_n35279_), .B(new_n35399_), .ZN(po0512));
  INV_X1     g32094(.I(pi1081), .ZN(new_n35401_));
  NAND2_X1   g32095(.A1(new_n35279_), .A2(pi0356), .ZN(new_n35402_));
  OAI21_X1   g32096(.A1(new_n35401_), .A2(new_n35279_), .B(new_n35402_), .ZN(po0513));
  INV_X1     g32097(.I(pi1076), .ZN(new_n35404_));
  NAND2_X1   g32098(.A1(new_n35279_), .A2(pi0357), .ZN(new_n35405_));
  OAI21_X1   g32099(.A1(new_n35404_), .A2(new_n35279_), .B(new_n35405_), .ZN(po0514));
  INV_X1     g32100(.I(pi1071), .ZN(new_n35407_));
  NAND2_X1   g32101(.A1(new_n35279_), .A2(pi0358), .ZN(new_n35408_));
  OAI21_X1   g32102(.A1(new_n35407_), .A2(new_n35279_), .B(new_n35408_), .ZN(po0515));
  INV_X1     g32103(.I(pi1068), .ZN(new_n35410_));
  NAND2_X1   g32104(.A1(new_n35279_), .A2(pi0359), .ZN(new_n35411_));
  OAI21_X1   g32105(.A1(new_n35410_), .A2(new_n35279_), .B(new_n35411_), .ZN(po0516));
  INV_X1     g32106(.I(pi1042), .ZN(new_n35413_));
  NAND2_X1   g32107(.A1(new_n35279_), .A2(pi0360), .ZN(new_n35414_));
  OAI21_X1   g32108(.A1(new_n35413_), .A2(new_n35279_), .B(new_n35414_), .ZN(po0517));
  NAND2_X1   g32109(.A1(new_n35279_), .A2(pi0361), .ZN(new_n35416_));
  OAI21_X1   g32110(.A1(new_n35184_), .A2(new_n35279_), .B(new_n35416_), .ZN(po0518));
  NAND2_X1   g32111(.A1(new_n35279_), .A2(pi0362), .ZN(new_n35418_));
  OAI21_X1   g32112(.A1(new_n33991_), .A2(new_n35279_), .B(new_n35418_), .ZN(po0519));
  NAND2_X1   g32113(.A1(new_n35286_), .A2(pi1049), .ZN(new_n35420_));
  OAI21_X1   g32114(.A1(new_n6705_), .A2(new_n35286_), .B(new_n35420_), .ZN(po0520));
  NAND2_X1   g32115(.A1(new_n35286_), .A2(pi1062), .ZN(new_n35422_));
  OAI21_X1   g32116(.A1(new_n6722_), .A2(new_n35286_), .B(new_n35422_), .ZN(po0521));
  INV_X1     g32117(.I(pi0365), .ZN(new_n35424_));
  NAND2_X1   g32118(.A1(new_n35286_), .A2(pi1065), .ZN(new_n35425_));
  OAI21_X1   g32119(.A1(new_n35424_), .A2(new_n35286_), .B(new_n35425_), .ZN(po0522));
  INV_X1     g32120(.I(pi0366), .ZN(new_n35427_));
  NAND2_X1   g32121(.A1(new_n35286_), .A2(pi1069), .ZN(new_n35428_));
  OAI21_X1   g32122(.A1(new_n35427_), .A2(new_n35286_), .B(new_n35428_), .ZN(po0523));
  NAND2_X1   g32123(.A1(new_n35286_), .A2(pi1039), .ZN(new_n35430_));
  OAI21_X1   g32124(.A1(new_n6729_), .A2(new_n35286_), .B(new_n35430_), .ZN(po0524));
  INV_X1     g32125(.I(pi0368), .ZN(new_n35432_));
  NAND2_X1   g32126(.A1(new_n35286_), .A2(pi1067), .ZN(new_n35433_));
  OAI21_X1   g32127(.A1(new_n35432_), .A2(new_n35286_), .B(new_n35433_), .ZN(po0525));
  NAND2_X1   g32128(.A1(new_n35286_), .A2(pi1080), .ZN(new_n35435_));
  OAI21_X1   g32129(.A1(new_n10140_), .A2(new_n35286_), .B(new_n35435_), .ZN(po0526));
  NAND2_X1   g32130(.A1(new_n35286_), .A2(pi1055), .ZN(new_n35437_));
  OAI21_X1   g32131(.A1(new_n7179_), .A2(new_n35286_), .B(new_n35437_), .ZN(po0527));
  NAND2_X1   g32132(.A1(new_n35286_), .A2(pi1051), .ZN(new_n35439_));
  OAI21_X1   g32133(.A1(new_n6671_), .A2(new_n35286_), .B(new_n35439_), .ZN(po0528));
  NAND2_X1   g32134(.A1(new_n35286_), .A2(pi1048), .ZN(new_n35441_));
  OAI21_X1   g32135(.A1(new_n6707_), .A2(new_n35286_), .B(new_n35441_), .ZN(po0529));
  INV_X1     g32136(.I(pi0373), .ZN(new_n35443_));
  NAND2_X1   g32137(.A1(new_n35286_), .A2(pi1087), .ZN(new_n35444_));
  OAI21_X1   g32138(.A1(new_n35443_), .A2(new_n35286_), .B(new_n35444_), .ZN(po0530));
  NAND2_X1   g32139(.A1(new_n35286_), .A2(pi1035), .ZN(new_n35446_));
  OAI21_X1   g32140(.A1(new_n7178_), .A2(new_n35286_), .B(new_n35446_), .ZN(po0531));
  NAND2_X1   g32141(.A1(new_n35286_), .A2(pi1047), .ZN(new_n35448_));
  OAI21_X1   g32142(.A1(new_n7177_), .A2(new_n35286_), .B(new_n35448_), .ZN(po0532));
  INV_X1     g32143(.I(pi0376), .ZN(new_n35450_));
  NAND2_X1   g32144(.A1(new_n35286_), .A2(pi1079), .ZN(new_n35451_));
  OAI21_X1   g32145(.A1(new_n35450_), .A2(new_n35286_), .B(new_n35451_), .ZN(po0533));
  NAND2_X1   g32146(.A1(new_n35286_), .A2(pi1074), .ZN(new_n35453_));
  OAI21_X1   g32147(.A1(new_n6677_), .A2(new_n35286_), .B(new_n35453_), .ZN(po0534));
  NAND2_X1   g32148(.A1(new_n35286_), .A2(pi1063), .ZN(new_n35455_));
  OAI21_X1   g32149(.A1(new_n6681_), .A2(new_n35286_), .B(new_n35455_), .ZN(po0535));
  INV_X1     g32150(.I(pi0379), .ZN(new_n35457_));
  NAND2_X1   g32151(.A1(new_n35286_), .A2(pi1045), .ZN(new_n35458_));
  OAI21_X1   g32152(.A1(new_n35457_), .A2(new_n35286_), .B(new_n35458_), .ZN(po0536));
  INV_X1     g32153(.I(pi0380), .ZN(new_n35460_));
  NAND2_X1   g32154(.A1(new_n35286_), .A2(pi1084), .ZN(new_n35461_));
  OAI21_X1   g32155(.A1(new_n35460_), .A2(new_n35286_), .B(new_n35461_), .ZN(po0537));
  NAND2_X1   g32156(.A1(new_n35286_), .A2(pi1081), .ZN(new_n35463_));
  OAI21_X1   g32157(.A1(new_n6678_), .A2(new_n35286_), .B(new_n35463_), .ZN(po0538));
  INV_X1     g32158(.I(pi0382), .ZN(new_n35465_));
  NAND2_X1   g32159(.A1(new_n35286_), .A2(pi1076), .ZN(new_n35466_));
  OAI21_X1   g32160(.A1(new_n35465_), .A2(new_n35286_), .B(new_n35466_), .ZN(po0539));
  INV_X1     g32161(.I(pi0383), .ZN(new_n35468_));
  NAND2_X1   g32162(.A1(new_n35286_), .A2(pi1071), .ZN(new_n35469_));
  OAI21_X1   g32163(.A1(new_n35468_), .A2(new_n35286_), .B(new_n35469_), .ZN(po0540));
  NAND2_X1   g32164(.A1(new_n35286_), .A2(pi1068), .ZN(new_n35471_));
  OAI21_X1   g32165(.A1(new_n6743_), .A2(new_n35286_), .B(new_n35471_), .ZN(po0541));
  NAND2_X1   g32166(.A1(new_n35286_), .A2(pi1042), .ZN(new_n35473_));
  OAI21_X1   g32167(.A1(new_n6682_), .A2(new_n35286_), .B(new_n35473_), .ZN(po0542));
  NAND2_X1   g32168(.A1(new_n35286_), .A2(pi1059), .ZN(new_n35475_));
  OAI21_X1   g32169(.A1(new_n6708_), .A2(new_n35286_), .B(new_n35475_), .ZN(po0543));
  NAND2_X1   g32170(.A1(new_n35286_), .A2(pi1053), .ZN(new_n35477_));
  OAI21_X1   g32171(.A1(new_n6700_), .A2(new_n35286_), .B(new_n35477_), .ZN(po0544));
  NAND2_X1   g32172(.A1(new_n35286_), .A2(pi1037), .ZN(new_n35479_));
  OAI21_X1   g32173(.A1(new_n6699_), .A2(new_n35286_), .B(new_n35479_), .ZN(po0545));
  INV_X1     g32174(.I(pi0389), .ZN(new_n35481_));
  NAND2_X1   g32175(.A1(new_n35286_), .A2(pi1036), .ZN(new_n35482_));
  OAI21_X1   g32176(.A1(new_n35481_), .A2(new_n35286_), .B(new_n35482_), .ZN(po0546));
  NAND2_X1   g32177(.A1(new_n35291_), .A2(pi0390), .ZN(new_n35484_));
  OAI21_X1   g32178(.A1(new_n35178_), .A2(new_n35291_), .B(new_n35484_), .ZN(po0547));
  NAND2_X1   g32179(.A1(new_n35291_), .A2(pi0391), .ZN(new_n35486_));
  OAI21_X1   g32180(.A1(new_n34003_), .A2(new_n35291_), .B(new_n35486_), .ZN(po0548));
  NAND2_X1   g32181(.A1(new_n35291_), .A2(pi0392), .ZN(new_n35488_));
  OAI21_X1   g32182(.A1(new_n33609_), .A2(new_n35291_), .B(new_n35488_), .ZN(po0549));
  NAND2_X1   g32183(.A1(new_n35291_), .A2(pi0393), .ZN(new_n35490_));
  OAI21_X1   g32184(.A1(new_n34016_), .A2(new_n35291_), .B(new_n35490_), .ZN(po0550));
  NAND2_X1   g32185(.A1(new_n35291_), .A2(pi0394), .ZN(new_n35492_));
  OAI21_X1   g32186(.A1(new_n35277_), .A2(new_n35291_), .B(new_n35492_), .ZN(po0551));
  NAND2_X1   g32187(.A1(new_n35291_), .A2(pi0395), .ZN(new_n35494_));
  OAI21_X1   g32188(.A1(new_n35377_), .A2(new_n35291_), .B(new_n35494_), .ZN(po0552));
  NAND2_X1   g32189(.A1(new_n35291_), .A2(pi0396), .ZN(new_n35496_));
  OAI21_X1   g32190(.A1(new_n35301_), .A2(new_n35291_), .B(new_n35496_), .ZN(po0553));
  NAND2_X1   g32191(.A1(new_n35291_), .A2(pi0397), .ZN(new_n35498_));
  OAI21_X1   g32192(.A1(new_n35175_), .A2(new_n35291_), .B(new_n35498_), .ZN(po0554));
  NAND2_X1   g32193(.A1(new_n35291_), .A2(pi0398), .ZN(new_n35500_));
  OAI21_X1   g32194(.A1(new_n35380_), .A2(new_n35291_), .B(new_n35500_), .ZN(po0555));
  NAND2_X1   g32195(.A1(new_n35291_), .A2(pi0399), .ZN(new_n35502_));
  OAI21_X1   g32196(.A1(new_n35282_), .A2(new_n35291_), .B(new_n35502_), .ZN(po0556));
  NAND2_X1   g32197(.A1(new_n35291_), .A2(pi0400), .ZN(new_n35504_));
  OAI21_X1   g32198(.A1(new_n35385_), .A2(new_n35291_), .B(new_n35504_), .ZN(po0557));
  NAND2_X1   g32199(.A1(new_n35291_), .A2(pi0401), .ZN(new_n35506_));
  OAI21_X1   g32200(.A1(new_n35388_), .A2(new_n35291_), .B(new_n35506_), .ZN(po0558));
  NAND2_X1   g32201(.A1(new_n35291_), .A2(pi0402), .ZN(new_n35508_));
  OAI21_X1   g32202(.A1(new_n35391_), .A2(new_n35291_), .B(new_n35508_), .ZN(po0559));
  NAND2_X1   g32203(.A1(new_n35291_), .A2(pi0403), .ZN(new_n35510_));
  OAI21_X1   g32204(.A1(new_n35396_), .A2(new_n35291_), .B(new_n35510_), .ZN(po0560));
  NAND2_X1   g32205(.A1(new_n35291_), .A2(pi0404), .ZN(new_n35512_));
  OAI21_X1   g32206(.A1(new_n35181_), .A2(new_n35291_), .B(new_n35512_), .ZN(po0561));
  NAND2_X1   g32207(.A1(new_n35291_), .A2(pi0405), .ZN(new_n35514_));
  OAI21_X1   g32208(.A1(new_n35401_), .A2(new_n35291_), .B(new_n35514_), .ZN(po0562));
  NAND2_X1   g32209(.A1(new_n35291_), .A2(pi0406), .ZN(new_n35516_));
  OAI21_X1   g32210(.A1(new_n35404_), .A2(new_n35291_), .B(new_n35516_), .ZN(po0563));
  NAND2_X1   g32211(.A1(new_n35291_), .A2(pi0407), .ZN(new_n35518_));
  OAI21_X1   g32212(.A1(new_n35407_), .A2(new_n35291_), .B(new_n35518_), .ZN(po0564));
  NAND2_X1   g32213(.A1(new_n35291_), .A2(pi0408), .ZN(new_n35520_));
  OAI21_X1   g32214(.A1(new_n35410_), .A2(new_n35291_), .B(new_n35520_), .ZN(po0565));
  NAND2_X1   g32215(.A1(new_n35291_), .A2(pi0409), .ZN(new_n35522_));
  OAI21_X1   g32216(.A1(new_n35413_), .A2(new_n35291_), .B(new_n35522_), .ZN(po0566));
  NAND2_X1   g32217(.A1(new_n35291_), .A2(pi0410), .ZN(new_n35524_));
  OAI21_X1   g32218(.A1(new_n35184_), .A2(new_n35291_), .B(new_n35524_), .ZN(po0567));
  NAND2_X1   g32219(.A1(new_n35291_), .A2(pi0411), .ZN(new_n35526_));
  OAI21_X1   g32220(.A1(new_n33607_), .A2(new_n35291_), .B(new_n35526_), .ZN(po0568));
  NAND2_X1   g32221(.A1(new_n35291_), .A2(pi0412), .ZN(new_n35528_));
  OAI21_X1   g32222(.A1(new_n34021_), .A2(new_n35291_), .B(new_n35528_), .ZN(po0569));
  NAND2_X1   g32223(.A1(new_n35291_), .A2(pi0413), .ZN(new_n35530_));
  OAI21_X1   g32224(.A1(new_n33985_), .A2(new_n35291_), .B(new_n35530_), .ZN(po0570));
  NAND3_X1   g32225(.A1(new_n35146_), .A2(new_n35330_), .A3(new_n7240_), .ZN(new_n35532_));
  NAND2_X1   g32226(.A1(new_n35532_), .A2(pi0414), .ZN(new_n35533_));
  OAI21_X1   g32227(.A1(new_n35178_), .A2(new_n35532_), .B(new_n35533_), .ZN(po0571));
  NAND2_X1   g32228(.A1(new_n35532_), .A2(pi0415), .ZN(new_n35535_));
  OAI21_X1   g32229(.A1(new_n34003_), .A2(new_n35532_), .B(new_n35535_), .ZN(po0572));
  NAND2_X1   g32230(.A1(new_n35532_), .A2(pi0416), .ZN(new_n35537_));
  OAI21_X1   g32231(.A1(new_n34009_), .A2(new_n35532_), .B(new_n35537_), .ZN(po0573));
  NAND2_X1   g32232(.A1(new_n35532_), .A2(pi0417), .ZN(new_n35539_));
  OAI21_X1   g32233(.A1(new_n33609_), .A2(new_n35532_), .B(new_n35539_), .ZN(po0574));
  NAND2_X1   g32234(.A1(new_n35532_), .A2(pi0418), .ZN(new_n35541_));
  OAI21_X1   g32235(.A1(new_n34016_), .A2(new_n35532_), .B(new_n35541_), .ZN(po0575));
  NAND2_X1   g32236(.A1(new_n35532_), .A2(pi0419), .ZN(new_n35543_));
  OAI21_X1   g32237(.A1(new_n35277_), .A2(new_n35532_), .B(new_n35543_), .ZN(po0576));
  NAND2_X1   g32238(.A1(new_n35532_), .A2(pi0420), .ZN(new_n35545_));
  OAI21_X1   g32239(.A1(new_n35377_), .A2(new_n35532_), .B(new_n35545_), .ZN(po0577));
  NAND2_X1   g32240(.A1(new_n35532_), .A2(pi0421), .ZN(new_n35547_));
  OAI21_X1   g32241(.A1(new_n35301_), .A2(new_n35532_), .B(new_n35547_), .ZN(po0578));
  NAND2_X1   g32242(.A1(new_n35532_), .A2(pi0422), .ZN(new_n35549_));
  OAI21_X1   g32243(.A1(new_n35175_), .A2(new_n35532_), .B(new_n35549_), .ZN(po0579));
  NAND2_X1   g32244(.A1(new_n35532_), .A2(pi0423), .ZN(new_n35551_));
  OAI21_X1   g32245(.A1(new_n35380_), .A2(new_n35532_), .B(new_n35551_), .ZN(po0580));
  NAND2_X1   g32246(.A1(new_n35532_), .A2(pi0424), .ZN(new_n35553_));
  OAI21_X1   g32247(.A1(new_n35282_), .A2(new_n35532_), .B(new_n35553_), .ZN(po0581));
  NAND2_X1   g32248(.A1(new_n35532_), .A2(pi0425), .ZN(new_n35555_));
  OAI21_X1   g32249(.A1(new_n35385_), .A2(new_n35532_), .B(new_n35555_), .ZN(po0582));
  NAND2_X1   g32250(.A1(new_n35532_), .A2(pi0426), .ZN(new_n35557_));
  OAI21_X1   g32251(.A1(new_n35388_), .A2(new_n35532_), .B(new_n35557_), .ZN(po0583));
  NAND2_X1   g32252(.A1(new_n35532_), .A2(pi0427), .ZN(new_n35559_));
  OAI21_X1   g32253(.A1(new_n35391_), .A2(new_n35532_), .B(new_n35559_), .ZN(po0584));
  NAND2_X1   g32254(.A1(new_n35532_), .A2(pi0428), .ZN(new_n35561_));
  OAI21_X1   g32255(.A1(new_n35396_), .A2(new_n35532_), .B(new_n35561_), .ZN(po0585));
  NAND2_X1   g32256(.A1(new_n35532_), .A2(pi0429), .ZN(new_n35563_));
  OAI21_X1   g32257(.A1(new_n35181_), .A2(new_n35532_), .B(new_n35563_), .ZN(po0586));
  NAND2_X1   g32258(.A1(new_n35532_), .A2(pi0430), .ZN(new_n35565_));
  OAI21_X1   g32259(.A1(new_n35404_), .A2(new_n35532_), .B(new_n35565_), .ZN(po0587));
  NAND2_X1   g32260(.A1(new_n35532_), .A2(pi0431), .ZN(new_n35567_));
  OAI21_X1   g32261(.A1(new_n35407_), .A2(new_n35532_), .B(new_n35567_), .ZN(po0588));
  NAND2_X1   g32262(.A1(new_n35532_), .A2(pi0432), .ZN(new_n35569_));
  OAI21_X1   g32263(.A1(new_n35410_), .A2(new_n35532_), .B(new_n35569_), .ZN(po0589));
  NAND2_X1   g32264(.A1(new_n35532_), .A2(pi0433), .ZN(new_n35571_));
  OAI21_X1   g32265(.A1(new_n35413_), .A2(new_n35532_), .B(new_n35571_), .ZN(po0590));
  NAND2_X1   g32266(.A1(new_n35532_), .A2(pi0434), .ZN(new_n35573_));
  OAI21_X1   g32267(.A1(new_n35184_), .A2(new_n35532_), .B(new_n35573_), .ZN(po0591));
  NAND2_X1   g32268(.A1(new_n35532_), .A2(pi0435), .ZN(new_n35575_));
  OAI21_X1   g32269(.A1(new_n33607_), .A2(new_n35532_), .B(new_n35575_), .ZN(po0592));
  NAND2_X1   g32270(.A1(new_n35532_), .A2(pi0436), .ZN(new_n35577_));
  OAI21_X1   g32271(.A1(new_n34021_), .A2(new_n35532_), .B(new_n35577_), .ZN(po0593));
  NAND2_X1   g32272(.A1(new_n35532_), .A2(pi0437), .ZN(new_n35579_));
  OAI21_X1   g32273(.A1(new_n33991_), .A2(new_n35532_), .B(new_n35579_), .ZN(po0594));
  NAND2_X1   g32274(.A1(new_n35532_), .A2(pi0438), .ZN(new_n35581_));
  OAI21_X1   g32275(.A1(new_n33985_), .A2(new_n35532_), .B(new_n35581_), .ZN(po0595));
  INV_X1     g32276(.I(pi0439), .ZN(new_n35583_));
  NAND2_X1   g32277(.A1(new_n35286_), .A2(pi1057), .ZN(new_n35584_));
  OAI21_X1   g32278(.A1(new_n35583_), .A2(new_n35286_), .B(new_n35584_), .ZN(po0596));
  NAND2_X1   g32279(.A1(new_n35286_), .A2(pi1043), .ZN(new_n35586_));
  OAI21_X1   g32280(.A1(new_n6744_), .A2(new_n35286_), .B(new_n35586_), .ZN(po0597));
  NAND2_X1   g32281(.A1(new_n35279_), .A2(pi0441), .ZN(new_n35588_));
  OAI21_X1   g32282(.A1(new_n34014_), .A2(new_n35279_), .B(new_n35588_), .ZN(po0598));
  NAND2_X1   g32283(.A1(new_n35286_), .A2(pi1058), .ZN(new_n35590_));
  OAI21_X1   g32284(.A1(new_n6746_), .A2(new_n35286_), .B(new_n35590_), .ZN(po0599));
  NAND2_X1   g32285(.A1(new_n35532_), .A2(pi0443), .ZN(new_n35592_));
  OAI21_X1   g32286(.A1(new_n34014_), .A2(new_n35532_), .B(new_n35592_), .ZN(po0600));
  NAND2_X1   g32287(.A1(new_n35532_), .A2(pi0444), .ZN(new_n35594_));
  OAI21_X1   g32288(.A1(new_n35187_), .A2(new_n35532_), .B(new_n35594_), .ZN(po0601));
  NAND2_X1   g32289(.A1(new_n35532_), .A2(pi0445), .ZN(new_n35596_));
  OAI21_X1   g32290(.A1(new_n35401_), .A2(new_n35532_), .B(new_n35596_), .ZN(po0602));
  NAND2_X1   g32291(.A1(new_n35532_), .A2(pi0446), .ZN(new_n35598_));
  OAI21_X1   g32292(.A1(new_n35306_), .A2(new_n35532_), .B(new_n35598_), .ZN(po0603));
  INV_X1     g32293(.I(pi0447), .ZN(new_n35600_));
  NAND2_X1   g32294(.A1(new_n35286_), .A2(pi1040), .ZN(new_n35601_));
  OAI21_X1   g32295(.A1(new_n35600_), .A2(new_n35286_), .B(new_n35601_), .ZN(po0604));
  NAND2_X1   g32296(.A1(new_n35532_), .A2(pi0448), .ZN(new_n35603_));
  OAI21_X1   g32297(.A1(new_n35289_), .A2(new_n35532_), .B(new_n35603_), .ZN(po0605));
  NAND2_X1   g32298(.A1(new_n35532_), .A2(pi0449), .ZN(new_n35605_));
  OAI21_X1   g32299(.A1(new_n35312_), .A2(new_n35532_), .B(new_n35605_), .ZN(po0606));
  NAND2_X1   g32300(.A1(new_n35279_), .A2(pi0450), .ZN(new_n35607_));
  OAI21_X1   g32301(.A1(new_n33985_), .A2(new_n35279_), .B(new_n35607_), .ZN(po0607));
  NAND2_X1   g32302(.A1(new_n35532_), .A2(pi0451), .ZN(new_n35609_));
  OAI21_X1   g32303(.A1(new_n35309_), .A2(new_n35532_), .B(new_n35609_), .ZN(po0608));
  NAND2_X1   g32304(.A1(new_n35279_), .A2(pi0452), .ZN(new_n35611_));
  OAI21_X1   g32305(.A1(new_n33607_), .A2(new_n35279_), .B(new_n35611_), .ZN(po0609));
  NAND2_X1   g32306(.A1(new_n35532_), .A2(pi0453), .ZN(new_n35613_));
  OAI21_X1   g32307(.A1(new_n34023_), .A2(new_n35532_), .B(new_n35613_), .ZN(po0610));
  NAND2_X1   g32308(.A1(new_n35532_), .A2(pi0454), .ZN(new_n35615_));
  OAI21_X1   g32309(.A1(new_n35319_), .A2(new_n35532_), .B(new_n35615_), .ZN(po0611));
  NAND2_X1   g32310(.A1(new_n35279_), .A2(pi0455), .ZN(new_n35617_));
  OAI21_X1   g32311(.A1(new_n34021_), .A2(new_n35279_), .B(new_n35617_), .ZN(po0612));
  NAND2_X1   g32312(.A1(new_n35291_), .A2(pi0456), .ZN(new_n35619_));
  OAI21_X1   g32313(.A1(new_n34014_), .A2(new_n35291_), .B(new_n35619_), .ZN(po0613));
  INV_X1     g32314(.I(pi0804), .ZN(new_n35621_));
  INV_X1     g32315(.I(pi0810), .ZN(new_n35622_));
  AOI21_X1   g32316(.A1(pi0600), .A2(new_n35622_), .B(new_n35621_), .ZN(new_n35623_));
  INV_X1     g32317(.I(pi0594), .ZN(new_n35624_));
  INV_X1     g32318(.I(pi0597), .ZN(new_n35625_));
  INV_X1     g32319(.I(pi0600), .ZN(new_n35626_));
  INV_X1     g32320(.I(pi0601), .ZN(new_n35627_));
  NOR4_X1    g32321(.A1(new_n35624_), .A2(new_n35625_), .A3(new_n35626_), .A4(new_n35627_), .ZN(new_n35628_));
  INV_X1     g32322(.I(pi0599), .ZN(new_n35629_));
  AOI21_X1   g32323(.A1(pi0596), .A2(pi0804), .B(pi0810), .ZN(new_n35630_));
  OAI21_X1   g32324(.A1(new_n35630_), .A2(new_n35629_), .B(pi0595), .ZN(new_n35631_));
  INV_X1     g32325(.I(pi0595), .ZN(new_n35632_));
  INV_X1     g32326(.I(pi0815), .ZN(new_n35633_));
  NAND2_X1   g32327(.A1(new_n35621_), .A2(new_n35622_), .ZN(new_n35634_));
  NOR3_X1    g32328(.A1(new_n35634_), .A2(new_n35632_), .A3(new_n35633_), .ZN(new_n35635_));
  XNOR2_X1   g32329(.A1(new_n35635_), .A2(new_n35631_), .ZN(new_n35636_));
  AOI21_X1   g32330(.A1(new_n35634_), .A2(new_n35627_), .B(pi0815), .ZN(new_n35637_));
  AOI22_X1   g32331(.A1(new_n35636_), .A2(new_n35637_), .B1(new_n35623_), .B2(new_n35628_), .ZN(new_n35638_));
  INV_X1     g32332(.I(pi0990), .ZN(new_n35639_));
  NOR3_X1    g32333(.A1(new_n35624_), .A2(new_n35626_), .A3(new_n35639_), .ZN(new_n35640_));
  AND3_X2    g32334(.A1(new_n35623_), .A2(new_n35633_), .A3(pi0821), .Z(new_n35641_));
  AOI21_X1   g32335(.A1(new_n35641_), .A2(new_n35640_), .B(pi0605), .ZN(new_n35642_));
  NOR2_X1    g32336(.A1(new_n35638_), .A2(new_n35642_), .ZN(po0614));
  NAND2_X1   g32337(.A1(new_n35279_), .A2(pi0458), .ZN(new_n35644_));
  OAI21_X1   g32338(.A1(new_n35187_), .A2(new_n35279_), .B(new_n35644_), .ZN(po0615));
  NAND2_X1   g32339(.A1(new_n35532_), .A2(pi0459), .ZN(new_n35646_));
  OAI21_X1   g32340(.A1(new_n35298_), .A2(new_n35532_), .B(new_n35646_), .ZN(po0616));
  NAND2_X1   g32341(.A1(new_n35279_), .A2(pi0460), .ZN(new_n35648_));
  OAI21_X1   g32342(.A1(new_n35306_), .A2(new_n35279_), .B(new_n35648_), .ZN(po0617));
  NAND2_X1   g32343(.A1(new_n35279_), .A2(pi0461), .ZN(new_n35650_));
  OAI21_X1   g32344(.A1(new_n35312_), .A2(new_n35279_), .B(new_n35650_), .ZN(po0618));
  NAND2_X1   g32345(.A1(new_n35279_), .A2(pi0462), .ZN(new_n35652_));
  OAI21_X1   g32346(.A1(new_n35289_), .A2(new_n35279_), .B(new_n35652_), .ZN(po0619));
  NAND2_X1   g32347(.A1(new_n35291_), .A2(pi0463), .ZN(new_n35654_));
  OAI21_X1   g32348(.A1(new_n33991_), .A2(new_n35291_), .B(new_n35654_), .ZN(po0620));
  NAND2_X1   g32349(.A1(new_n35532_), .A2(pi0464), .ZN(new_n35656_));
  OAI21_X1   g32350(.A1(new_n33997_), .A2(new_n35532_), .B(new_n35656_), .ZN(po0621));
  AOI21_X1   g32351(.A1(new_n32579_), .A2(new_n35217_), .B(new_n7240_), .ZN(new_n35658_));
  NOR2_X1    g32352(.A1(new_n5294_), .A2(new_n5296_), .ZN(new_n35659_));
  INV_X1     g32353(.I(new_n9225_), .ZN(new_n35660_));
  NOR2_X1    g32354(.A1(new_n9223_), .A2(new_n35660_), .ZN(new_n35661_));
  INV_X1     g32355(.I(new_n35661_), .ZN(new_n35662_));
  NAND4_X1   g32356(.A1(new_n35662_), .A2(new_n32579_), .A3(pi1157), .A4(new_n35659_), .ZN(new_n35663_));
  NAND2_X1   g32357(.A1(new_n35662_), .A2(new_n32579_), .ZN(new_n35664_));
  NAND3_X1   g32358(.A1(new_n35664_), .A2(new_n35659_), .A3(new_n14006_), .ZN(new_n35665_));
  NAND2_X1   g32359(.A1(new_n35665_), .A2(new_n35663_), .ZN(new_n35666_));
  NOR4_X1    g32360(.A1(new_n3121_), .A2(new_n3098_), .A3(pi0222), .A4(pi0223), .ZN(new_n35667_));
  XOR2_X1    g32361(.A1(new_n35667_), .A2(new_n5190_), .Z(new_n35668_));
  NAND2_X1   g32362(.A1(new_n35668_), .A2(pi0243), .ZN(new_n35669_));
  NAND2_X1   g32363(.A1(new_n35669_), .A2(new_n35662_), .ZN(new_n35670_));
  AOI22_X1   g32364(.A1(new_n35666_), .A2(pi0926), .B1(pi1157), .B2(new_n35670_), .ZN(new_n35671_));
  AOI22_X1   g32365(.A1(new_n35215_), .A2(pi1157), .B1(pi0926), .B2(new_n5280_), .ZN(new_n35672_));
  NAND2_X1   g32366(.A1(new_n5293_), .A2(new_n3121_), .ZN(new_n35673_));
  OAI21_X1   g32367(.A1(new_n35673_), .A2(new_n3383_), .B(pi0216), .ZN(new_n35674_));
  NAND4_X1   g32368(.A1(po1038), .A2(new_n32579_), .A3(pi0926), .A4(pi1157), .ZN(new_n35675_));
  NOR4_X1    g32369(.A1(new_n35671_), .A2(new_n35672_), .A3(new_n35674_), .A4(new_n35675_), .ZN(new_n35676_));
  XOR2_X1    g32370(.A1(new_n35676_), .A2(new_n35658_), .Z(po0622));
  NOR2_X1    g32371(.A1(new_n35661_), .A2(po1038), .ZN(new_n35678_));
  AOI21_X1   g32372(.A1(po1038), .A2(new_n35217_), .B(new_n35678_), .ZN(new_n35679_));
  NAND3_X1   g32373(.A1(new_n35253_), .A2(pi0943), .A3(pi1151), .ZN(new_n35680_));
  NAND3_X1   g32374(.A1(new_n35252_), .A2(pi0943), .A3(new_n31670_), .ZN(new_n35681_));
  AOI21_X1   g32375(.A1(new_n35680_), .A2(new_n35681_), .B(new_n35679_), .ZN(new_n35682_));
  INV_X1     g32376(.I(pi0943), .ZN(new_n35683_));
  NOR2_X1    g32377(.A1(new_n35683_), .A2(new_n31670_), .ZN(new_n35684_));
  INV_X1     g32378(.I(new_n35679_), .ZN(new_n35685_));
  NOR2_X1    g32379(.A1(new_n35685_), .A2(new_n35223_), .ZN(new_n35686_));
  NOR2_X1    g32380(.A1(new_n12654_), .A2(new_n3314_), .ZN(new_n35687_));
  AOI21_X1   g32381(.A1(new_n3136_), .A2(new_n12654_), .B(new_n35687_), .ZN(new_n35688_));
  AOI22_X1   g32382(.A1(new_n35686_), .A2(new_n35683_), .B1(new_n35688_), .B2(new_n35684_), .ZN(new_n35689_));
  NOR2_X1    g32383(.A1(new_n7240_), .A2(pi0215), .ZN(new_n35690_));
  NAND3_X1   g32384(.A1(new_n35668_), .A2(po1038), .A3(pi0221), .ZN(new_n35691_));
  XOR2_X1    g32385(.A1(new_n35691_), .A2(new_n35690_), .Z(new_n35692_));
  NOR4_X1    g32386(.A1(new_n35682_), .A2(new_n32770_), .A3(new_n35689_), .A4(new_n35692_), .ZN(po0623));
  NAND2_X1   g32387(.A1(new_n7269_), .A2(new_n13017_), .ZN(new_n35694_));
  OAI21_X1   g32388(.A1(new_n8290_), .A2(new_n35694_), .B(new_n13002_), .ZN(new_n35695_));
  NOR2_X1    g32389(.A1(new_n10455_), .A2(new_n2454_), .ZN(new_n35696_));
  NAND2_X1   g32390(.A1(new_n35696_), .A2(new_n35695_), .ZN(new_n35697_));
  NAND3_X1   g32391(.A1(new_n33614_), .A2(pi0040), .A3(new_n5401_), .ZN(new_n35698_));
  OAI21_X1   g32392(.A1(new_n5532_), .A2(new_n35698_), .B(new_n35697_), .ZN(new_n35699_));
  INV_X1     g32393(.I(new_n35698_), .ZN(new_n35700_));
  NAND3_X1   g32394(.A1(new_n35696_), .A2(new_n35695_), .A3(new_n35700_), .ZN(new_n35701_));
  OAI21_X1   g32395(.A1(new_n5532_), .A2(new_n35701_), .B(new_n35699_), .ZN(new_n35702_));
  NAND2_X1   g32396(.A1(new_n35697_), .A2(new_n35698_), .ZN(new_n35703_));
  NAND3_X1   g32397(.A1(new_n35703_), .A2(pi1091), .A3(new_n35701_), .ZN(new_n35704_));
  NAND2_X1   g32398(.A1(new_n6474_), .A2(pi1091), .ZN(new_n35705_));
  XOR2_X1    g32399(.A1(new_n35704_), .A2(new_n35705_), .Z(new_n35706_));
  INV_X1     g32400(.I(new_n30541_), .ZN(po0950));
  NAND4_X1   g32401(.A1(new_n8288_), .A2(new_n3193_), .A3(new_n5765_), .A4(new_n7330_), .ZN(new_n35708_));
  AOI21_X1   g32402(.A1(po0950), .A2(new_n35700_), .B(new_n35708_), .ZN(new_n35709_));
  AOI21_X1   g32403(.A1(new_n35706_), .A2(new_n35702_), .B(new_n35709_), .ZN(new_n35710_));
  OAI21_X1   g32404(.A1(new_n6402_), .A2(new_n35698_), .B(new_n35697_), .ZN(new_n35711_));
  OAI21_X1   g32405(.A1(new_n6402_), .A2(new_n35701_), .B(new_n35711_), .ZN(new_n35712_));
  NOR2_X1    g32406(.A1(new_n35702_), .A2(new_n2984_), .ZN(new_n35713_));
  XOR2_X1    g32407(.A1(new_n35713_), .A2(new_n2985_), .Z(new_n35714_));
  NAND2_X1   g32408(.A1(new_n35714_), .A2(new_n35712_), .ZN(new_n35715_));
  NOR2_X1    g32409(.A1(new_n35715_), .A2(new_n35710_), .ZN(po0624));
  NAND3_X1   g32410(.A1(new_n8297_), .A2(new_n3259_), .A3(new_n3262_), .ZN(new_n35717_));
  OAI22_X1   g32411(.A1(new_n7325_), .A2(new_n35717_), .B1(new_n9180_), .B2(new_n9439_), .ZN(po0625));
  AOI21_X1   g32412(.A1(new_n34074_), .A2(new_n35217_), .B(new_n7240_), .ZN(new_n35719_));
  NAND4_X1   g32413(.A1(new_n35662_), .A2(new_n34074_), .A3(pi1156), .A4(new_n35659_), .ZN(new_n35720_));
  NAND2_X1   g32414(.A1(new_n35662_), .A2(new_n34074_), .ZN(new_n35721_));
  NAND3_X1   g32415(.A1(new_n35721_), .A2(new_n35659_), .A3(new_n13969_), .ZN(new_n35722_));
  NAND2_X1   g32416(.A1(new_n35722_), .A2(new_n35720_), .ZN(new_n35723_));
  NAND2_X1   g32417(.A1(new_n35668_), .A2(pi0263), .ZN(new_n35724_));
  NAND2_X1   g32418(.A1(new_n35724_), .A2(new_n35662_), .ZN(new_n35725_));
  AOI22_X1   g32419(.A1(new_n35723_), .A2(pi0942), .B1(pi1156), .B2(new_n35725_), .ZN(new_n35726_));
  AOI22_X1   g32420(.A1(new_n35215_), .A2(pi1156), .B1(pi0942), .B2(new_n5280_), .ZN(new_n35727_));
  NAND4_X1   g32421(.A1(po1038), .A2(new_n34074_), .A3(pi0942), .A4(pi1156), .ZN(new_n35728_));
  NOR4_X1    g32422(.A1(new_n35726_), .A2(new_n35674_), .A3(new_n35727_), .A4(new_n35728_), .ZN(new_n35729_));
  XOR2_X1    g32423(.A1(new_n35729_), .A2(new_n35719_), .Z(po0626));
  AOI21_X1   g32424(.A1(pi0267), .A2(new_n35217_), .B(new_n7240_), .ZN(new_n35731_));
  NAND4_X1   g32425(.A1(new_n35662_), .A2(pi0267), .A3(pi1155), .A4(new_n35659_), .ZN(new_n35732_));
  NAND2_X1   g32426(.A1(new_n35662_), .A2(pi0267), .ZN(new_n35733_));
  NAND3_X1   g32427(.A1(new_n35733_), .A2(new_n35659_), .A3(new_n13778_), .ZN(new_n35734_));
  NAND2_X1   g32428(.A1(new_n35734_), .A2(new_n35732_), .ZN(new_n35735_));
  NAND2_X1   g32429(.A1(new_n35668_), .A2(pi0267), .ZN(new_n35736_));
  NAND2_X1   g32430(.A1(new_n35736_), .A2(new_n35662_), .ZN(new_n35737_));
  AOI22_X1   g32431(.A1(new_n35735_), .A2(pi0925), .B1(pi1155), .B2(new_n35737_), .ZN(new_n35738_));
  AOI22_X1   g32432(.A1(new_n35215_), .A2(pi1155), .B1(pi0925), .B2(new_n5280_), .ZN(new_n35739_));
  NAND4_X1   g32433(.A1(po1038), .A2(pi0267), .A3(pi0925), .A4(pi1155), .ZN(new_n35740_));
  NOR4_X1    g32434(.A1(new_n35738_), .A2(new_n35674_), .A3(new_n35739_), .A4(new_n35740_), .ZN(new_n35741_));
  XOR2_X1    g32435(.A1(new_n35741_), .A2(new_n35731_), .Z(po0627));
  AOI21_X1   g32436(.A1(pi0253), .A2(new_n35217_), .B(new_n7240_), .ZN(new_n35743_));
  NAND4_X1   g32437(.A1(new_n35662_), .A2(pi0253), .A3(pi1153), .A4(new_n35659_), .ZN(new_n35744_));
  NAND2_X1   g32438(.A1(new_n35662_), .A2(pi0253), .ZN(new_n35745_));
  NAND3_X1   g32439(.A1(new_n35745_), .A2(new_n35659_), .A3(new_n13614_), .ZN(new_n35746_));
  NAND2_X1   g32440(.A1(new_n35746_), .A2(new_n35744_), .ZN(new_n35747_));
  NAND2_X1   g32441(.A1(new_n35668_), .A2(pi0253), .ZN(new_n35748_));
  NAND2_X1   g32442(.A1(new_n35748_), .A2(new_n35662_), .ZN(new_n35749_));
  AOI22_X1   g32443(.A1(new_n35747_), .A2(pi0941), .B1(pi1153), .B2(new_n35749_), .ZN(new_n35750_));
  AOI22_X1   g32444(.A1(new_n35215_), .A2(pi1153), .B1(pi0941), .B2(new_n5280_), .ZN(new_n35751_));
  NAND4_X1   g32445(.A1(po1038), .A2(pi0253), .A3(pi0941), .A4(pi1153), .ZN(new_n35752_));
  NOR4_X1    g32446(.A1(new_n35750_), .A2(new_n35674_), .A3(new_n35751_), .A4(new_n35752_), .ZN(new_n35753_));
  XOR2_X1    g32447(.A1(new_n35753_), .A2(new_n35743_), .Z(po0628));
  AOI21_X1   g32448(.A1(pi0254), .A2(new_n35217_), .B(new_n7240_), .ZN(new_n35755_));
  NAND4_X1   g32449(.A1(new_n35662_), .A2(pi0254), .A3(pi1154), .A4(new_n35659_), .ZN(new_n35756_));
  NAND2_X1   g32450(.A1(new_n35662_), .A2(pi0254), .ZN(new_n35757_));
  NAND3_X1   g32451(.A1(new_n35757_), .A2(new_n35659_), .A3(new_n13817_), .ZN(new_n35758_));
  NAND2_X1   g32452(.A1(new_n35758_), .A2(new_n35756_), .ZN(new_n35759_));
  NAND2_X1   g32453(.A1(new_n35668_), .A2(pi0254), .ZN(new_n35760_));
  NAND2_X1   g32454(.A1(new_n35760_), .A2(new_n35662_), .ZN(new_n35761_));
  AOI22_X1   g32455(.A1(new_n35759_), .A2(pi0923), .B1(pi1154), .B2(new_n35761_), .ZN(new_n35762_));
  AOI22_X1   g32456(.A1(new_n35215_), .A2(pi1154), .B1(pi0923), .B2(new_n5280_), .ZN(new_n35763_));
  NAND4_X1   g32457(.A1(po1038), .A2(pi0254), .A3(pi0923), .A4(pi1154), .ZN(new_n35764_));
  NOR4_X1    g32458(.A1(new_n35762_), .A2(new_n35674_), .A3(new_n35763_), .A4(new_n35764_), .ZN(new_n35765_));
  XOR2_X1    g32459(.A1(new_n35765_), .A2(new_n35755_), .Z(po0629));
  NAND3_X1   g32460(.A1(new_n35253_), .A2(pi0922), .A3(pi1152), .ZN(new_n35767_));
  NAND3_X1   g32461(.A1(new_n35252_), .A2(pi0922), .A3(new_n31002_), .ZN(new_n35768_));
  AOI21_X1   g32462(.A1(new_n35767_), .A2(new_n35768_), .B(new_n35679_), .ZN(new_n35769_));
  INV_X1     g32463(.I(pi0922), .ZN(new_n35770_));
  NOR2_X1    g32464(.A1(new_n35770_), .A2(new_n31002_), .ZN(new_n35771_));
  AOI22_X1   g32465(.A1(new_n35686_), .A2(new_n35770_), .B1(new_n35688_), .B2(new_n35771_), .ZN(new_n35772_));
  NOR4_X1    g32466(.A1(new_n35769_), .A2(new_n34534_), .A3(new_n35692_), .A4(new_n35772_), .ZN(po0630));
  NAND3_X1   g32467(.A1(new_n35253_), .A2(pi0931), .A3(pi1150), .ZN(new_n35774_));
  NAND3_X1   g32468(.A1(new_n35252_), .A2(pi0931), .A3(new_n32242_), .ZN(new_n35775_));
  AOI21_X1   g32469(.A1(new_n35774_), .A2(new_n35775_), .B(new_n35679_), .ZN(new_n35776_));
  INV_X1     g32470(.I(pi0931), .ZN(new_n35777_));
  NOR2_X1    g32471(.A1(new_n35777_), .A2(new_n32242_), .ZN(new_n35778_));
  AOI22_X1   g32472(.A1(new_n35686_), .A2(new_n35777_), .B1(new_n35688_), .B2(new_n35778_), .ZN(new_n35779_));
  NOR4_X1    g32473(.A1(new_n35776_), .A2(new_n32769_), .A3(new_n35692_), .A4(new_n35779_), .ZN(po0631));
  NAND3_X1   g32474(.A1(new_n35253_), .A2(pi0936), .A3(pi1149), .ZN(new_n35781_));
  NAND3_X1   g32475(.A1(new_n35252_), .A2(pi0936), .A3(new_n31941_), .ZN(new_n35782_));
  AOI21_X1   g32476(.A1(new_n35781_), .A2(new_n35782_), .B(new_n35679_), .ZN(new_n35783_));
  INV_X1     g32477(.I(pi0936), .ZN(new_n35784_));
  NOR2_X1    g32478(.A1(new_n35784_), .A2(new_n31941_), .ZN(new_n35785_));
  AOI22_X1   g32479(.A1(new_n35686_), .A2(new_n35784_), .B1(new_n35688_), .B2(new_n35785_), .ZN(new_n35786_));
  NOR4_X1    g32480(.A1(new_n35783_), .A2(new_n32771_), .A3(new_n35692_), .A4(new_n35786_), .ZN(po0632));
  NOR3_X1    g32481(.A1(new_n10244_), .A2(new_n8276_), .A3(new_n9263_), .ZN(new_n35788_));
  NOR3_X1    g32482(.A1(new_n35788_), .A2(new_n8282_), .A3(new_n9263_), .ZN(new_n35789_));
  NOR4_X1    g32483(.A1(new_n10244_), .A2(new_n8276_), .A3(new_n8283_), .A4(new_n9263_), .ZN(new_n35790_));
  NAND4_X1   g32484(.A1(new_n10246_), .A2(new_n2446_), .A3(new_n3291_), .A4(new_n8529_), .ZN(new_n35791_));
  NOR3_X1    g32485(.A1(new_n35789_), .A2(new_n35791_), .A3(new_n35790_), .ZN(new_n35792_));
  NOR4_X1    g32486(.A1(new_n35792_), .A2(new_n2450_), .A3(new_n7240_), .A4(new_n9263_), .ZN(new_n35793_));
  XOR2_X1    g32487(.A1(new_n35793_), .A2(new_n34560_), .Z(po0633));
  NAND2_X1   g32488(.A1(new_n35265_), .A2(new_n35266_), .ZN(po0634));
  NOR2_X1    g32489(.A1(new_n34817_), .A2(new_n2450_), .ZN(po0635));
  INV_X1     g32490(.I(pi0481), .ZN(new_n35797_));
  NAND2_X1   g32491(.A1(new_n27674_), .A2(pi0248), .ZN(new_n35798_));
  OAI21_X1   g32492(.A1(new_n35797_), .A2(new_n27674_), .B(new_n35798_), .ZN(po0638));
  INV_X1     g32493(.I(new_n27683_), .ZN(new_n35800_));
  NAND2_X1   g32494(.A1(new_n35800_), .A2(pi0482), .ZN(new_n35801_));
  OAI21_X1   g32495(.A1(new_n3810_), .A2(new_n35800_), .B(new_n35801_), .ZN(po0639));
  NAND2_X1   g32496(.A1(new_n27763_), .A2(new_n27766_), .ZN(new_n35803_));
  NAND2_X1   g32497(.A1(new_n35803_), .A2(pi0483), .ZN(new_n35804_));
  OAI21_X1   g32498(.A1(new_n5364_), .A2(new_n35803_), .B(new_n35804_), .ZN(po0640));
  NAND2_X1   g32499(.A1(new_n35803_), .A2(pi0484), .ZN(new_n35806_));
  OAI21_X1   g32500(.A1(new_n3810_), .A2(new_n35803_), .B(new_n35806_), .ZN(po0641));
  INV_X1     g32501(.I(pi0485), .ZN(new_n35808_));
  NAND2_X1   g32502(.A1(new_n28698_), .A2(pi0234), .ZN(new_n35809_));
  OAI21_X1   g32503(.A1(new_n35808_), .A2(new_n28698_), .B(new_n35809_), .ZN(po0642));
  INV_X1     g32504(.I(pi0486), .ZN(new_n35811_));
  NAND2_X1   g32505(.A1(new_n28698_), .A2(pi0244), .ZN(new_n35812_));
  OAI21_X1   g32506(.A1(new_n35811_), .A2(new_n28698_), .B(new_n35812_), .ZN(po0643));
  INV_X1     g32507(.I(pi0487), .ZN(new_n35814_));
  NAND2_X1   g32508(.A1(new_n27674_), .A2(pi0246), .ZN(new_n35815_));
  OAI21_X1   g32509(.A1(new_n35814_), .A2(new_n27674_), .B(new_n35815_), .ZN(po0644));
  NAND2_X1   g32510(.A1(new_n27674_), .A2(pi0239), .ZN(new_n35817_));
  OAI21_X1   g32511(.A1(pi0488), .A2(new_n27674_), .B(new_n35817_), .ZN(po0645));
  INV_X1     g32512(.I(pi0489), .ZN(new_n35819_));
  NAND2_X1   g32513(.A1(new_n28698_), .A2(pi0242), .ZN(new_n35820_));
  OAI21_X1   g32514(.A1(new_n35819_), .A2(new_n28698_), .B(new_n35820_), .ZN(po0646));
  NAND2_X1   g32515(.A1(new_n35803_), .A2(pi0490), .ZN(new_n35822_));
  OAI21_X1   g32516(.A1(new_n4064_), .A2(new_n35803_), .B(new_n35822_), .ZN(po0647));
  NAND2_X1   g32517(.A1(new_n35803_), .A2(pi0491), .ZN(new_n35824_));
  OAI21_X1   g32518(.A1(new_n3743_), .A2(new_n35803_), .B(new_n35824_), .ZN(po0648));
  NAND2_X1   g32519(.A1(new_n35803_), .A2(pi0492), .ZN(new_n35826_));
  OAI21_X1   g32520(.A1(new_n4710_), .A2(new_n35803_), .B(new_n35826_), .ZN(po0649));
  INV_X1     g32521(.I(pi0244), .ZN(new_n35828_));
  NAND2_X1   g32522(.A1(new_n35803_), .A2(pi0493), .ZN(new_n35829_));
  OAI21_X1   g32523(.A1(new_n35828_), .A2(new_n35803_), .B(new_n35829_), .ZN(po0650));
  INV_X1     g32524(.I(pi0239), .ZN(new_n35831_));
  INV_X1     g32525(.I(pi0494), .ZN(new_n35832_));
  NAND2_X1   g32526(.A1(new_n35803_), .A2(new_n35832_), .ZN(new_n35833_));
  OAI21_X1   g32527(.A1(new_n35831_), .A2(new_n35803_), .B(new_n35833_), .ZN(po0651));
  NAND2_X1   g32528(.A1(new_n35803_), .A2(pi0495), .ZN(new_n35835_));
  OAI21_X1   g32529(.A1(new_n3611_), .A2(new_n35803_), .B(new_n35835_), .ZN(po0652));
  NAND2_X1   g32530(.A1(new_n27763_), .A2(new_n27678_), .ZN(new_n35837_));
  NAND2_X1   g32531(.A1(new_n35837_), .A2(pi0496), .ZN(new_n35838_));
  OAI21_X1   g32532(.A1(new_n3810_), .A2(new_n35837_), .B(new_n35838_), .ZN(po0653));
  INV_X1     g32533(.I(pi0497), .ZN(new_n35840_));
  NAND2_X1   g32534(.A1(new_n35837_), .A2(new_n35840_), .ZN(new_n35841_));
  OAI21_X1   g32535(.A1(new_n35831_), .A2(new_n35837_), .B(new_n35841_), .ZN(po0654));
  INV_X1     g32536(.I(pi0498), .ZN(new_n35843_));
  NAND2_X1   g32537(.A1(new_n27683_), .A2(pi0238), .ZN(new_n35844_));
  OAI21_X1   g32538(.A1(new_n35843_), .A2(new_n27683_), .B(new_n35844_), .ZN(po0655));
  NAND2_X1   g32539(.A1(new_n35837_), .A2(pi0499), .ZN(new_n35846_));
  OAI21_X1   g32540(.A1(new_n4549_), .A2(new_n35837_), .B(new_n35846_), .ZN(po0656));
  NAND2_X1   g32541(.A1(new_n35837_), .A2(pi0500), .ZN(new_n35848_));
  OAI21_X1   g32542(.A1(new_n4064_), .A2(new_n35837_), .B(new_n35848_), .ZN(po0657));
  NAND2_X1   g32543(.A1(new_n35837_), .A2(pi0501), .ZN(new_n35850_));
  OAI21_X1   g32544(.A1(new_n4225_), .A2(new_n35837_), .B(new_n35850_), .ZN(po0658));
  NAND2_X1   g32545(.A1(new_n35837_), .A2(pi0502), .ZN(new_n35852_));
  OAI21_X1   g32546(.A1(new_n4459_), .A2(new_n35837_), .B(new_n35852_), .ZN(po0659));
  NAND2_X1   g32547(.A1(new_n35837_), .A2(pi0503), .ZN(new_n35854_));
  OAI21_X1   g32548(.A1(new_n4955_), .A2(new_n35837_), .B(new_n35854_), .ZN(po0660));
  INV_X1     g32549(.I(pi0504), .ZN(new_n35856_));
  NAND2_X1   g32550(.A1(new_n27760_), .A2(pi0242), .ZN(new_n35857_));
  OAI21_X1   g32551(.A1(new_n35856_), .A2(new_n27760_), .B(new_n35857_), .ZN(po0661));
  NAND3_X1   g32552(.A1(new_n32522_), .A2(new_n5555_), .A3(new_n5656_), .ZN(new_n35859_));
  NAND3_X1   g32553(.A1(new_n5638_), .A2(new_n5652_), .A3(new_n32522_), .ZN(new_n35860_));
  NAND2_X1   g32554(.A1(new_n35860_), .A2(new_n35859_), .ZN(new_n35861_));
  NAND2_X1   g32555(.A1(new_n35861_), .A2(new_n2768_), .ZN(new_n35862_));
  NOR2_X1    g32556(.A1(new_n27759_), .A2(new_n2768_), .ZN(new_n35863_));
  NAND3_X1   g32557(.A1(new_n35863_), .A2(pi0505), .A3(new_n27641_), .ZN(new_n35864_));
  AOI21_X1   g32558(.A1(new_n35864_), .A2(new_n35862_), .B(new_n35837_), .ZN(po0662));
  INV_X1     g32559(.I(pi0506), .ZN(new_n35866_));
  NAND2_X1   g32560(.A1(new_n27760_), .A2(pi0241), .ZN(new_n35867_));
  OAI21_X1   g32561(.A1(new_n35866_), .A2(new_n27760_), .B(new_n35867_), .ZN(po0663));
  INV_X1     g32562(.I(new_n27760_), .ZN(new_n35869_));
  NAND2_X1   g32563(.A1(new_n35869_), .A2(pi0507), .ZN(new_n35870_));
  OAI21_X1   g32564(.A1(new_n3743_), .A2(new_n35869_), .B(new_n35870_), .ZN(po0664));
  INV_X1     g32565(.I(pi0508), .ZN(new_n35872_));
  NAND2_X1   g32566(.A1(new_n27760_), .A2(pi0247), .ZN(new_n35873_));
  OAI21_X1   g32567(.A1(new_n35872_), .A2(new_n27760_), .B(new_n35873_), .ZN(po0665));
  INV_X1     g32568(.I(pi0509), .ZN(new_n35875_));
  NAND2_X1   g32569(.A1(new_n27760_), .A2(pi0245), .ZN(new_n35876_));
  OAI21_X1   g32570(.A1(new_n35875_), .A2(new_n27760_), .B(new_n35876_), .ZN(po0666));
  INV_X1     g32571(.I(pi0510), .ZN(new_n35878_));
  NAND2_X1   g32572(.A1(new_n27674_), .A2(pi0242), .ZN(new_n35879_));
  OAI21_X1   g32573(.A1(new_n35878_), .A2(new_n27674_), .B(new_n35879_), .ZN(po0667));
  INV_X1     g32574(.I(pi0511), .ZN(new_n35881_));
  NOR3_X1    g32575(.A1(new_n5798_), .A2(new_n5807_), .A3(new_n32521_), .ZN(new_n35882_));
  NOR3_X1    g32576(.A1(new_n5802_), .A2(new_n5809_), .A3(new_n32521_), .ZN(new_n35883_));
  NOR2_X1    g32577(.A1(new_n35883_), .A2(new_n35882_), .ZN(new_n35884_));
  NOR2_X1    g32578(.A1(new_n35884_), .A2(pi0234), .ZN(new_n35885_));
  INV_X1     g32579(.I(new_n35885_), .ZN(new_n35886_));
  NAND2_X1   g32580(.A1(new_n35886_), .A2(new_n27674_), .ZN(new_n35887_));
  OAI21_X1   g32581(.A1(new_n35881_), .A2(new_n27674_), .B(new_n35887_), .ZN(po0668));
  INV_X1     g32582(.I(pi0512), .ZN(new_n35889_));
  NAND2_X1   g32583(.A1(new_n27674_), .A2(pi0235), .ZN(new_n35890_));
  OAI21_X1   g32584(.A1(new_n35889_), .A2(new_n27674_), .B(new_n35890_), .ZN(po0669));
  INV_X1     g32585(.I(pi0513), .ZN(new_n35892_));
  NAND2_X1   g32586(.A1(new_n27674_), .A2(pi0244), .ZN(new_n35893_));
  OAI21_X1   g32587(.A1(new_n35892_), .A2(new_n27674_), .B(new_n35893_), .ZN(po0670));
  INV_X1     g32588(.I(pi0514), .ZN(new_n35895_));
  NAND2_X1   g32589(.A1(new_n27674_), .A2(pi0245), .ZN(new_n35896_));
  OAI21_X1   g32590(.A1(new_n35895_), .A2(new_n27674_), .B(new_n35896_), .ZN(po0671));
  INV_X1     g32591(.I(pi0515), .ZN(new_n35898_));
  NAND2_X1   g32592(.A1(new_n27674_), .A2(pi0240), .ZN(new_n35899_));
  OAI21_X1   g32593(.A1(new_n35898_), .A2(new_n27674_), .B(new_n35899_), .ZN(po0672));
  INV_X1     g32594(.I(pi0516), .ZN(new_n35901_));
  NAND2_X1   g32595(.A1(new_n27674_), .A2(pi0247), .ZN(new_n35902_));
  OAI21_X1   g32596(.A1(new_n35901_), .A2(new_n27674_), .B(new_n35902_), .ZN(po0673));
  INV_X1     g32597(.I(pi0517), .ZN(new_n35904_));
  NAND2_X1   g32598(.A1(new_n27674_), .A2(pi0238), .ZN(new_n35905_));
  OAI21_X1   g32599(.A1(new_n35904_), .A2(new_n27674_), .B(new_n35905_), .ZN(po0674));
  NOR2_X1    g32600(.A1(new_n27673_), .A2(new_n2768_), .ZN(new_n35907_));
  NAND3_X1   g32601(.A1(new_n35907_), .A2(pi0518), .A3(new_n27641_), .ZN(new_n35908_));
  AOI21_X1   g32602(.A1(new_n35908_), .A2(new_n35886_), .B(new_n27679_), .ZN(po0675));
  NAND2_X1   g32603(.A1(new_n27680_), .A2(pi0239), .ZN(new_n35910_));
  OAI21_X1   g32604(.A1(pi0519), .A2(new_n27680_), .B(new_n35910_), .ZN(po0676));
  NAND2_X1   g32605(.A1(new_n27679_), .A2(pi0520), .ZN(new_n35912_));
  OAI21_X1   g32606(.A1(new_n4549_), .A2(new_n27679_), .B(new_n35912_), .ZN(po0677));
  NAND2_X1   g32607(.A1(new_n27679_), .A2(pi0521), .ZN(new_n35914_));
  OAI21_X1   g32608(.A1(new_n4225_), .A2(new_n27679_), .B(new_n35914_), .ZN(po0678));
  NAND2_X1   g32609(.A1(new_n27679_), .A2(pi0522), .ZN(new_n35916_));
  OAI21_X1   g32610(.A1(new_n3743_), .A2(new_n27679_), .B(new_n35916_), .ZN(po0679));
  NAND2_X1   g32611(.A1(new_n27677_), .A2(new_n27766_), .ZN(new_n35918_));
  NAND3_X1   g32612(.A1(new_n35907_), .A2(pi0523), .A3(new_n27641_), .ZN(new_n35919_));
  AOI21_X1   g32613(.A1(new_n35919_), .A2(new_n35886_), .B(new_n35918_), .ZN(po0680));
  INV_X1     g32614(.I(pi0524), .ZN(new_n35921_));
  NAND2_X1   g32615(.A1(new_n35918_), .A2(new_n35921_), .ZN(new_n35922_));
  OAI21_X1   g32616(.A1(new_n35831_), .A2(new_n35918_), .B(new_n35922_), .ZN(po0681));
  NAND2_X1   g32617(.A1(new_n35918_), .A2(pi0525), .ZN(new_n35924_));
  OAI21_X1   g32618(.A1(new_n4955_), .A2(new_n35918_), .B(new_n35924_), .ZN(po0682));
  NAND2_X1   g32619(.A1(new_n35918_), .A2(pi0526), .ZN(new_n35926_));
  OAI21_X1   g32620(.A1(new_n4549_), .A2(new_n35918_), .B(new_n35926_), .ZN(po0683));
  NAND2_X1   g32621(.A1(new_n35918_), .A2(pi0527), .ZN(new_n35928_));
  OAI21_X1   g32622(.A1(new_n4459_), .A2(new_n35918_), .B(new_n35928_), .ZN(po0684));
  NAND2_X1   g32623(.A1(new_n35918_), .A2(pi0528), .ZN(new_n35930_));
  OAI21_X1   g32624(.A1(new_n3810_), .A2(new_n35918_), .B(new_n35930_), .ZN(po0685));
  NAND2_X1   g32625(.A1(new_n35918_), .A2(pi0529), .ZN(new_n35932_));
  OAI21_X1   g32626(.A1(new_n3743_), .A2(new_n35918_), .B(new_n35932_), .ZN(po0686));
  NAND2_X1   g32627(.A1(new_n35918_), .A2(pi0530), .ZN(new_n35934_));
  OAI21_X1   g32628(.A1(new_n4710_), .A2(new_n35918_), .B(new_n35934_), .ZN(po0687));
  INV_X1     g32629(.I(pi0531), .ZN(new_n35936_));
  NAND2_X1   g32630(.A1(new_n27683_), .A2(pi0235), .ZN(new_n35937_));
  OAI21_X1   g32631(.A1(new_n35936_), .A2(new_n27683_), .B(new_n35937_), .ZN(po0688));
  INV_X1     g32632(.I(pi0532), .ZN(new_n35939_));
  NAND2_X1   g32633(.A1(new_n27683_), .A2(pi0247), .ZN(new_n35940_));
  OAI21_X1   g32634(.A1(new_n35939_), .A2(new_n27683_), .B(new_n35940_), .ZN(po0689));
  INV_X1     g32635(.I(pi0533), .ZN(new_n35942_));
  NAND2_X1   g32636(.A1(new_n27760_), .A2(pi0235), .ZN(new_n35943_));
  OAI21_X1   g32637(.A1(new_n35942_), .A2(new_n27760_), .B(new_n35943_), .ZN(po0690));
  NAND2_X1   g32638(.A1(new_n27760_), .A2(pi0239), .ZN(new_n35945_));
  OAI21_X1   g32639(.A1(pi0534), .A2(new_n27760_), .B(new_n35945_), .ZN(po0691));
  INV_X1     g32640(.I(pi0535), .ZN(new_n35947_));
  NAND2_X1   g32641(.A1(new_n27760_), .A2(pi0240), .ZN(new_n35948_));
  OAI21_X1   g32642(.A1(new_n35947_), .A2(new_n27760_), .B(new_n35948_), .ZN(po0692));
  INV_X1     g32643(.I(pi0536), .ZN(new_n35950_));
  NAND2_X1   g32644(.A1(new_n27760_), .A2(pi0246), .ZN(new_n35951_));
  OAI21_X1   g32645(.A1(new_n35950_), .A2(new_n27760_), .B(new_n35951_), .ZN(po0693));
  INV_X1     g32646(.I(pi0537), .ZN(new_n35953_));
  NAND2_X1   g32647(.A1(new_n27760_), .A2(pi0248), .ZN(new_n35954_));
  OAI21_X1   g32648(.A1(new_n35953_), .A2(new_n27760_), .B(new_n35954_), .ZN(po0694));
  INV_X1     g32649(.I(pi0538), .ZN(new_n35956_));
  NAND2_X1   g32650(.A1(new_n27760_), .A2(pi0249), .ZN(new_n35957_));
  OAI21_X1   g32651(.A1(new_n35956_), .A2(new_n27760_), .B(new_n35957_), .ZN(po0695));
  NAND2_X1   g32652(.A1(new_n35837_), .A2(pi0539), .ZN(new_n35959_));
  OAI21_X1   g32653(.A1(new_n5364_), .A2(new_n35837_), .B(new_n35959_), .ZN(po0696));
  NAND2_X1   g32654(.A1(new_n35837_), .A2(pi0540), .ZN(new_n35961_));
  OAI21_X1   g32655(.A1(new_n3611_), .A2(new_n35837_), .B(new_n35961_), .ZN(po0697));
  NAND2_X1   g32656(.A1(new_n35837_), .A2(pi0541), .ZN(new_n35963_));
  OAI21_X1   g32657(.A1(new_n35828_), .A2(new_n35837_), .B(new_n35963_), .ZN(po0698));
  NAND2_X1   g32658(.A1(new_n35837_), .A2(pi0542), .ZN(new_n35965_));
  OAI21_X1   g32659(.A1(new_n4710_), .A2(new_n35837_), .B(new_n35965_), .ZN(po0699));
  NAND2_X1   g32660(.A1(new_n35837_), .A2(pi0543), .ZN(new_n35967_));
  OAI21_X1   g32661(.A1(new_n3743_), .A2(new_n35837_), .B(new_n35967_), .ZN(po0700));
  NAND3_X1   g32662(.A1(new_n35863_), .A2(pi0544), .A3(new_n27641_), .ZN(new_n35969_));
  AOI21_X1   g32663(.A1(new_n35969_), .A2(new_n35862_), .B(new_n35803_), .ZN(po0701));
  NAND2_X1   g32664(.A1(new_n35803_), .A2(pi0545), .ZN(new_n35971_));
  OAI21_X1   g32665(.A1(new_n4955_), .A2(new_n35803_), .B(new_n35971_), .ZN(po0702));
  NAND2_X1   g32666(.A1(new_n35803_), .A2(pi0546), .ZN(new_n35973_));
  OAI21_X1   g32667(.A1(new_n4549_), .A2(new_n35803_), .B(new_n35973_), .ZN(po0703));
  NAND2_X1   g32668(.A1(new_n35803_), .A2(pi0547), .ZN(new_n35975_));
  OAI21_X1   g32669(.A1(new_n4459_), .A2(new_n35803_), .B(new_n35975_), .ZN(po0704));
  NAND2_X1   g32670(.A1(new_n35803_), .A2(pi0548), .ZN(new_n35977_));
  OAI21_X1   g32671(.A1(new_n4225_), .A2(new_n35803_), .B(new_n35977_), .ZN(po0705));
  INV_X1     g32672(.I(pi0549), .ZN(new_n35979_));
  NAND2_X1   g32673(.A1(new_n28698_), .A2(pi0235), .ZN(new_n35980_));
  OAI21_X1   g32674(.A1(new_n35979_), .A2(new_n28698_), .B(new_n35980_), .ZN(po0706));
  NAND2_X1   g32675(.A1(new_n28698_), .A2(pi0239), .ZN(new_n35982_));
  OAI21_X1   g32676(.A1(pi0550), .A2(new_n28698_), .B(new_n35982_), .ZN(po0707));
  INV_X1     g32677(.I(pi0551), .ZN(new_n35984_));
  NAND2_X1   g32678(.A1(new_n28698_), .A2(pi0240), .ZN(new_n35985_));
  OAI21_X1   g32679(.A1(new_n35984_), .A2(new_n28698_), .B(new_n35985_), .ZN(po0708));
  INV_X1     g32680(.I(pi0552), .ZN(new_n35987_));
  NAND2_X1   g32681(.A1(new_n28698_), .A2(pi0247), .ZN(new_n35988_));
  OAI21_X1   g32682(.A1(new_n35987_), .A2(new_n28698_), .B(new_n35988_), .ZN(po0709));
  INV_X1     g32683(.I(pi0553), .ZN(new_n35990_));
  NAND2_X1   g32684(.A1(new_n28698_), .A2(pi0241), .ZN(new_n35991_));
  OAI21_X1   g32685(.A1(new_n35990_), .A2(new_n28698_), .B(new_n35991_), .ZN(po0710));
  INV_X1     g32686(.I(pi0554), .ZN(new_n35993_));
  NAND2_X1   g32687(.A1(new_n28698_), .A2(pi0248), .ZN(new_n35994_));
  OAI21_X1   g32688(.A1(new_n35993_), .A2(new_n28698_), .B(new_n35994_), .ZN(po0711));
  INV_X1     g32689(.I(pi0555), .ZN(new_n35996_));
  NAND2_X1   g32690(.A1(new_n28698_), .A2(pi0249), .ZN(new_n35997_));
  OAI21_X1   g32691(.A1(new_n35996_), .A2(new_n28698_), .B(new_n35997_), .ZN(po0712));
  INV_X1     g32692(.I(pi0556), .ZN(new_n35999_));
  NAND2_X1   g32693(.A1(new_n27683_), .A2(pi0242), .ZN(new_n36000_));
  OAI21_X1   g32694(.A1(new_n35999_), .A2(new_n27683_), .B(new_n36000_), .ZN(po0713));
  NAND3_X1   g32695(.A1(new_n35863_), .A2(pi0557), .A3(new_n27641_), .ZN(new_n36002_));
  AOI21_X1   g32696(.A1(new_n36002_), .A2(new_n35862_), .B(new_n35869_), .ZN(po0714));
  INV_X1     g32697(.I(pi0558), .ZN(new_n36004_));
  NAND2_X1   g32698(.A1(new_n27760_), .A2(pi0244), .ZN(new_n36005_));
  OAI21_X1   g32699(.A1(new_n36004_), .A2(new_n27760_), .B(new_n36005_), .ZN(po0715));
  INV_X1     g32700(.I(pi0559), .ZN(new_n36007_));
  NAND2_X1   g32701(.A1(new_n27674_), .A2(pi0241), .ZN(new_n36008_));
  OAI21_X1   g32702(.A1(new_n36007_), .A2(new_n27674_), .B(new_n36008_), .ZN(po0716));
  INV_X1     g32703(.I(pi0560), .ZN(new_n36010_));
  NAND2_X1   g32704(.A1(new_n27683_), .A2(pi0240), .ZN(new_n36011_));
  OAI21_X1   g32705(.A1(new_n36010_), .A2(new_n27683_), .B(new_n36011_), .ZN(po0717));
  NAND2_X1   g32706(.A1(new_n27679_), .A2(pi0561), .ZN(new_n36013_));
  OAI21_X1   g32707(.A1(new_n4459_), .A2(new_n27679_), .B(new_n36013_), .ZN(po0718));
  NAND2_X1   g32708(.A1(new_n35800_), .A2(pi0562), .ZN(new_n36015_));
  OAI21_X1   g32709(.A1(new_n4064_), .A2(new_n35800_), .B(new_n36015_), .ZN(po0719));
  INV_X1     g32710(.I(pi0563), .ZN(new_n36017_));
  NAND2_X1   g32711(.A1(new_n28698_), .A2(pi0246), .ZN(new_n36018_));
  OAI21_X1   g32712(.A1(new_n36017_), .A2(new_n28698_), .B(new_n36018_), .ZN(po0720));
  NAND2_X1   g32713(.A1(new_n35800_), .A2(pi0564), .ZN(new_n36020_));
  OAI21_X1   g32714(.A1(new_n4549_), .A2(new_n35800_), .B(new_n36020_), .ZN(po0721));
  NAND2_X1   g32715(.A1(new_n35800_), .A2(pi0565), .ZN(new_n36022_));
  OAI21_X1   g32716(.A1(new_n4225_), .A2(new_n35800_), .B(new_n36022_), .ZN(po0722));
  INV_X1     g32717(.I(pi0566), .ZN(new_n36024_));
  NAND2_X1   g32718(.A1(new_n27683_), .A2(pi0244), .ZN(new_n36025_));
  OAI21_X1   g32719(.A1(new_n36024_), .A2(new_n27683_), .B(new_n36025_), .ZN(po0723));
  NAND2_X1   g32720(.A1(new_n6514_), .A2(pi0230), .ZN(new_n36027_));
  NOR3_X1    g32721(.A1(new_n2979_), .A2(pi0567), .A3(pi1093), .ZN(new_n36028_));
  INV_X1     g32722(.I(new_n15392_), .ZN(new_n36029_));
  NOR2_X1    g32723(.A1(new_n36028_), .A2(pi0680), .ZN(new_n36030_));
  AOI21_X1   g32724(.A1(new_n13680_), .A2(new_n36030_), .B(new_n36029_), .ZN(new_n36031_));
  NOR2_X1    g32725(.A1(new_n15396_), .A2(new_n36031_), .ZN(new_n36032_));
  NAND2_X1   g32726(.A1(new_n36032_), .A2(new_n14059_), .ZN(new_n36033_));
  NOR2_X1    g32727(.A1(new_n36033_), .A2(new_n15401_), .ZN(new_n36034_));
  NOR2_X1    g32728(.A1(new_n36034_), .A2(new_n36028_), .ZN(new_n36035_));
  NOR4_X1    g32729(.A1(new_n16384_), .A2(new_n5794_), .A3(new_n14304_), .A4(new_n16375_), .ZN(new_n36036_));
  INV_X1     g32730(.I(new_n36028_), .ZN(new_n36037_));
  NAND2_X1   g32731(.A1(new_n36036_), .A2(new_n13860_), .ZN(new_n36038_));
  AOI21_X1   g32732(.A1(new_n36038_), .A2(new_n36037_), .B(new_n13896_), .ZN(new_n36039_));
  NOR2_X1    g32733(.A1(new_n13896_), .A2(new_n13868_), .ZN(new_n36040_));
  XOR2_X1    g32734(.A1(new_n36039_), .A2(new_n36040_), .Z(new_n36041_));
  AOI21_X1   g32735(.A1(new_n36036_), .A2(pi0619), .B(new_n36028_), .ZN(new_n36042_));
  NAND2_X1   g32736(.A1(new_n36041_), .A2(new_n36042_), .ZN(new_n36043_));
  NAND3_X1   g32737(.A1(new_n36043_), .A2(new_n13896_), .A3(new_n36037_), .ZN(new_n36044_));
  NAND2_X1   g32738(.A1(new_n36044_), .A2(new_n36036_), .ZN(new_n36045_));
  NOR2_X1    g32739(.A1(new_n16372_), .A2(new_n36028_), .ZN(new_n36046_));
  AOI21_X1   g32740(.A1(new_n36045_), .A2(new_n16372_), .B(new_n36046_), .ZN(new_n36047_));
  OAI22_X1   g32741(.A1(new_n36045_), .A2(new_n15479_), .B1(new_n27904_), .B2(new_n36031_), .ZN(new_n36048_));
  NAND4_X1   g32742(.A1(new_n36048_), .A2(new_n27914_), .A3(new_n36041_), .A4(new_n36042_), .ZN(new_n36049_));
  XOR2_X1    g32743(.A1(new_n36045_), .A2(pi1158), .Z(new_n36050_));
  NOR3_X1    g32744(.A1(new_n36050_), .A2(new_n13901_), .A3(new_n13964_), .ZN(new_n36051_));
  OR3_X2     g32745(.A1(new_n36031_), .A2(new_n13918_), .A3(new_n27904_), .Z(new_n36052_));
  OAI21_X1   g32746(.A1(new_n28070_), .A2(new_n36037_), .B(new_n36052_), .ZN(new_n36053_));
  NAND2_X1   g32747(.A1(new_n36053_), .A2(pi0641), .ZN(new_n36054_));
  NAND2_X1   g32748(.A1(new_n36054_), .A2(new_n13937_), .ZN(new_n36055_));
  AOI21_X1   g32749(.A1(new_n36028_), .A2(new_n14139_), .B(pi0641), .ZN(new_n36056_));
  NOR2_X1    g32750(.A1(new_n36052_), .A2(new_n36056_), .ZN(new_n36057_));
  OAI21_X1   g32751(.A1(new_n36051_), .A2(new_n36055_), .B(new_n36057_), .ZN(new_n36058_));
  NAND2_X1   g32752(.A1(new_n36058_), .A2(new_n36049_), .ZN(new_n36059_));
  NAND3_X1   g32753(.A1(new_n13942_), .A2(pi0629), .A3(pi1156), .ZN(new_n36060_));
  OAI21_X1   g32754(.A1(new_n36047_), .A2(new_n36060_), .B(new_n12777_), .ZN(new_n36061_));
  AOI21_X1   g32755(.A1(new_n36059_), .A2(new_n16424_), .B(new_n36061_), .ZN(new_n36062_));
  OAI21_X1   g32756(.A1(new_n36037_), .A2(new_n13969_), .B(new_n13942_), .ZN(new_n36063_));
  AOI21_X1   g32757(.A1(new_n36032_), .A2(new_n36063_), .B(pi0629), .ZN(new_n36064_));
  NOR4_X1    g32758(.A1(new_n36062_), .A2(new_n16567_), .A3(new_n36047_), .A4(new_n36064_), .ZN(new_n36065_));
  NAND2_X1   g32759(.A1(new_n36065_), .A2(new_n12776_), .ZN(new_n36066_));
  INV_X1     g32760(.I(new_n36047_), .ZN(new_n36067_));
  NOR2_X1    g32761(.A1(new_n13994_), .A2(new_n36028_), .ZN(new_n36068_));
  AOI21_X1   g32762(.A1(new_n36067_), .A2(new_n13994_), .B(new_n36068_), .ZN(new_n36069_));
  OAI21_X1   g32763(.A1(new_n36028_), .A2(pi1157), .B(pi0647), .ZN(new_n36070_));
  NOR2_X1    g32764(.A1(new_n36033_), .A2(new_n36070_), .ZN(new_n36071_));
  NOR2_X1    g32765(.A1(new_n36065_), .A2(new_n14006_), .ZN(new_n36072_));
  XOR2_X1    g32766(.A1(new_n36072_), .A2(new_n14008_), .Z(new_n36073_));
  NOR2_X1    g32767(.A1(new_n36073_), .A2(new_n36069_), .ZN(new_n36074_));
  NOR3_X1    g32768(.A1(new_n36074_), .A2(new_n14010_), .A3(new_n36071_), .ZN(new_n36075_));
  NOR3_X1    g32769(.A1(new_n36075_), .A2(pi0630), .A3(new_n36071_), .ZN(new_n36076_));
  NOR2_X1    g32770(.A1(new_n36065_), .A2(new_n14005_), .ZN(new_n36077_));
  XOR2_X1    g32771(.A1(new_n36077_), .A2(new_n14008_), .Z(new_n36078_));
  OR4_X2     g32772(.A1(new_n12776_), .A2(new_n36076_), .A3(new_n36069_), .A4(new_n36078_), .Z(new_n36079_));
  NAND2_X1   g32773(.A1(new_n36079_), .A2(new_n36066_), .ZN(new_n36080_));
  NOR2_X1    g32774(.A1(new_n36080_), .A2(new_n14200_), .ZN(new_n36081_));
  XOR2_X1    g32775(.A1(new_n36081_), .A2(new_n14205_), .Z(new_n36082_));
  NAND2_X1   g32776(.A1(new_n36082_), .A2(new_n36035_), .ZN(new_n36083_));
  NOR3_X1    g32777(.A1(new_n36067_), .A2(new_n13993_), .A3(new_n14210_), .ZN(new_n36084_));
  OAI21_X1   g32778(.A1(new_n36037_), .A2(new_n14200_), .B(new_n14204_), .ZN(new_n36085_));
  AOI21_X1   g32779(.A1(new_n36084_), .A2(new_n36085_), .B(new_n14203_), .ZN(new_n36086_));
  AOI21_X1   g32780(.A1(new_n36083_), .A2(new_n36086_), .B(new_n12775_), .ZN(new_n36087_));
  AOI21_X1   g32781(.A1(new_n36037_), .A2(new_n14200_), .B(new_n14204_), .ZN(new_n36088_));
  NOR2_X1    g32782(.A1(new_n36080_), .A2(new_n14204_), .ZN(new_n36089_));
  XOR2_X1    g32783(.A1(new_n36089_), .A2(new_n14205_), .Z(new_n36090_));
  AOI22_X1   g32784(.A1(new_n36090_), .A2(new_n36035_), .B1(new_n36084_), .B2(new_n36088_), .ZN(new_n36091_));
  NAND2_X1   g32785(.A1(new_n36080_), .A2(new_n19043_), .ZN(new_n36092_));
  NOR2_X1    g32786(.A1(new_n36091_), .A2(new_n36092_), .ZN(new_n36093_));
  XOR2_X1    g32787(.A1(new_n36093_), .A2(new_n36087_), .Z(new_n36094_));
  NAND3_X1   g32788(.A1(new_n36094_), .A2(pi0230), .A3(pi1092), .ZN(new_n36095_));
  XOR2_X1    g32789(.A1(new_n36095_), .A2(new_n36027_), .Z(po0724));
  INV_X1     g32790(.I(pi0568), .ZN(new_n36097_));
  NAND2_X1   g32791(.A1(new_n27683_), .A2(pi0245), .ZN(new_n36098_));
  OAI21_X1   g32792(.A1(new_n36097_), .A2(new_n27683_), .B(new_n36098_), .ZN(po0725));
  NAND2_X1   g32793(.A1(new_n27683_), .A2(pi0239), .ZN(new_n36100_));
  OAI21_X1   g32794(.A1(pi0569), .A2(new_n27683_), .B(new_n36100_), .ZN(po0726));
  NAND3_X1   g32795(.A1(new_n35907_), .A2(pi0570), .A3(new_n27641_), .ZN(new_n36102_));
  AOI21_X1   g32796(.A1(new_n36102_), .A2(new_n35886_), .B(new_n35800_), .ZN(po0727));
  NAND2_X1   g32797(.A1(new_n35918_), .A2(pi0571), .ZN(new_n36104_));
  OAI21_X1   g32798(.A1(new_n4064_), .A2(new_n35918_), .B(new_n36104_), .ZN(po0728));
  NAND2_X1   g32799(.A1(new_n35918_), .A2(pi0572), .ZN(new_n36106_));
  OAI21_X1   g32800(.A1(new_n35828_), .A2(new_n35918_), .B(new_n36106_), .ZN(po0729));
  NAND2_X1   g32801(.A1(new_n35918_), .A2(pi0573), .ZN(new_n36108_));
  OAI21_X1   g32802(.A1(new_n5364_), .A2(new_n35918_), .B(new_n36108_), .ZN(po0730));
  NAND2_X1   g32803(.A1(new_n27679_), .A2(pi0574), .ZN(new_n36110_));
  OAI21_X1   g32804(.A1(new_n4064_), .A2(new_n27679_), .B(new_n36110_), .ZN(po0731));
  NAND2_X1   g32805(.A1(new_n35918_), .A2(pi0575), .ZN(new_n36112_));
  OAI21_X1   g32806(.A1(new_n3611_), .A2(new_n35918_), .B(new_n36112_), .ZN(po0732));
  NAND2_X1   g32807(.A1(new_n35918_), .A2(pi0576), .ZN(new_n36114_));
  OAI21_X1   g32808(.A1(new_n4225_), .A2(new_n35918_), .B(new_n36114_), .ZN(po0733));
  INV_X1     g32809(.I(pi0577), .ZN(new_n36116_));
  NAND2_X1   g32810(.A1(new_n28698_), .A2(pi0238), .ZN(new_n36117_));
  OAI21_X1   g32811(.A1(new_n36116_), .A2(new_n28698_), .B(new_n36117_), .ZN(po0734));
  NAND2_X1   g32812(.A1(new_n27679_), .A2(pi0578), .ZN(new_n36119_));
  OAI21_X1   g32813(.A1(new_n3810_), .A2(new_n27679_), .B(new_n36119_), .ZN(po0735));
  INV_X1     g32814(.I(pi0579), .ZN(new_n36121_));
  NAND2_X1   g32815(.A1(new_n27674_), .A2(pi0249), .ZN(new_n36122_));
  OAI21_X1   g32816(.A1(new_n36121_), .A2(new_n27674_), .B(new_n36122_), .ZN(po0736));
  INV_X1     g32817(.I(pi0580), .ZN(new_n36124_));
  NAND2_X1   g32818(.A1(new_n28698_), .A2(pi0245), .ZN(new_n36125_));
  OAI21_X1   g32819(.A1(new_n36124_), .A2(new_n28698_), .B(new_n36125_), .ZN(po0737));
  NAND2_X1   g32820(.A1(new_n27679_), .A2(pi0581), .ZN(new_n36127_));
  OAI21_X1   g32821(.A1(new_n3611_), .A2(new_n27679_), .B(new_n36127_), .ZN(po0738));
  NAND2_X1   g32822(.A1(new_n27679_), .A2(pi0582), .ZN(new_n36129_));
  OAI21_X1   g32823(.A1(new_n4710_), .A2(new_n27679_), .B(new_n36129_), .ZN(po0739));
  NAND2_X1   g32824(.A1(new_n27679_), .A2(pi0584), .ZN(new_n36131_));
  OAI21_X1   g32825(.A1(new_n4955_), .A2(new_n27679_), .B(new_n36131_), .ZN(po0741));
  NAND2_X1   g32826(.A1(new_n27679_), .A2(pi0585), .ZN(new_n36133_));
  OAI21_X1   g32827(.A1(new_n35828_), .A2(new_n27679_), .B(new_n36133_), .ZN(po0742));
  NAND2_X1   g32828(.A1(new_n27679_), .A2(pi0586), .ZN(new_n36135_));
  OAI21_X1   g32829(.A1(new_n5364_), .A2(new_n27679_), .B(new_n36135_), .ZN(po0743));
  NOR3_X1    g32830(.A1(new_n16375_), .A2(new_n30557_), .A3(new_n13103_), .ZN(new_n36137_));
  NAND4_X1   g32831(.A1(new_n18967_), .A2(new_n14142_), .A3(new_n28375_), .A4(new_n36137_), .ZN(new_n36138_));
  OAI22_X1   g32832(.A1(new_n16388_), .A2(new_n36138_), .B1(pi0230), .B2(new_n5392_), .ZN(po0744));
  NOR4_X1    g32833(.A1(new_n35326_), .A2(pi0123), .A3(new_n5683_), .A4(new_n2722_), .ZN(new_n36140_));
  OAI21_X1   g32834(.A1(pi0591), .A2(new_n35326_), .B(new_n36140_), .ZN(new_n36141_));
  INV_X1     g32835(.I(new_n36140_), .ZN(new_n36142_));
  NAND3_X1   g32836(.A1(new_n36142_), .A2(new_n6350_), .A3(new_n35323_), .ZN(new_n36143_));
  AOI21_X1   g32837(.A1(new_n36143_), .A2(new_n36141_), .B(new_n9787_), .ZN(po0745));
  NOR3_X1    g32838(.A1(new_n5638_), .A2(new_n5652_), .A3(new_n32521_), .ZN(new_n36145_));
  NOR3_X1    g32839(.A1(new_n5555_), .A2(new_n5656_), .A3(new_n32521_), .ZN(new_n36146_));
  NOR2_X1    g32840(.A1(new_n36145_), .A2(new_n36146_), .ZN(new_n36147_));
  NAND2_X1   g32841(.A1(new_n27640_), .A2(pi0206), .ZN(new_n36148_));
  NAND2_X1   g32842(.A1(pi0204), .A2(pi0237), .ZN(new_n36149_));
  AOI21_X1   g32843(.A1(new_n36148_), .A2(new_n36149_), .B(new_n36147_), .ZN(po0746));
  OAI21_X1   g32844(.A1(pi0588), .A2(new_n35326_), .B(new_n36140_), .ZN(new_n36151_));
  NAND3_X1   g32845(.A1(new_n36142_), .A2(new_n9787_), .A3(new_n35323_), .ZN(new_n36152_));
  AOI21_X1   g32846(.A1(new_n36152_), .A2(new_n36151_), .B(new_n6933_), .ZN(po0747));
  OAI21_X1   g32847(.A1(pi0592), .A2(new_n35326_), .B(new_n36140_), .ZN(new_n36154_));
  NAND3_X1   g32848(.A1(new_n36142_), .A2(new_n6358_), .A3(new_n35323_), .ZN(new_n36155_));
  AOI21_X1   g32849(.A1(new_n36155_), .A2(new_n36154_), .B(new_n6350_), .ZN(po0748));
  OAI21_X1   g32850(.A1(pi0590), .A2(new_n35326_), .B(new_n36140_), .ZN(new_n36157_));
  NAND3_X1   g32851(.A1(new_n36142_), .A2(new_n6933_), .A3(new_n35323_), .ZN(new_n36158_));
  AOI21_X1   g32852(.A1(new_n36158_), .A2(new_n36157_), .B(new_n6358_), .ZN(po0749));
  INV_X1     g32853(.I(pi0534), .ZN(new_n36160_));
  NOR2_X1    g32854(.A1(new_n35884_), .A2(pi0511), .ZN(new_n36161_));
  NOR3_X1    g32855(.A1(new_n35883_), .A2(new_n35882_), .A3(new_n35881_), .ZN(new_n36162_));
  NAND2_X1   g32856(.A1(new_n4549_), .A2(pi0487), .ZN(new_n36163_));
  NAND2_X1   g32857(.A1(new_n35814_), .A2(pi0246), .ZN(new_n36164_));
  AOI21_X1   g32858(.A1(new_n36163_), .A2(new_n36164_), .B(new_n2768_), .ZN(new_n36165_));
  OAI21_X1   g32859(.A1(new_n36161_), .A2(new_n36162_), .B(new_n36165_), .ZN(new_n36166_));
  XOR2_X1    g32860(.A1(pi0249), .A2(pi0579), .Z(new_n36167_));
  NOR2_X1    g32861(.A1(new_n36166_), .A2(new_n36167_), .ZN(new_n36168_));
  NOR2_X1    g32862(.A1(new_n36147_), .A2(pi0557), .ZN(new_n36169_));
  INV_X1     g32863(.I(pi0557), .ZN(new_n36170_));
  NOR2_X1    g32864(.A1(new_n35861_), .A2(new_n36170_), .ZN(new_n36171_));
  NOR2_X1    g32865(.A1(new_n35950_), .A2(pi0246), .ZN(new_n36172_));
  NOR2_X1    g32866(.A1(new_n4549_), .A2(pi0536), .ZN(new_n36173_));
  OAI21_X1   g32867(.A1(new_n36172_), .A2(new_n36173_), .B(pi0234), .ZN(new_n36174_));
  INV_X1     g32868(.I(new_n36174_), .ZN(new_n36175_));
  OAI21_X1   g32869(.A1(new_n36169_), .A2(new_n36171_), .B(new_n36175_), .ZN(new_n36176_));
  XOR2_X1    g32870(.A1(pi0249), .A2(pi0538), .Z(new_n36177_));
  NOR2_X1    g32871(.A1(new_n36176_), .A2(new_n36177_), .ZN(new_n36178_));
  NAND3_X1   g32872(.A1(new_n36178_), .A2(pi0579), .A3(new_n36168_), .ZN(new_n36179_));
  XOR2_X1    g32873(.A1(new_n35884_), .A2(new_n35881_), .Z(new_n36180_));
  INV_X1     g32874(.I(new_n36167_), .ZN(new_n36181_));
  NAND3_X1   g32875(.A1(new_n36180_), .A2(new_n36165_), .A3(new_n36181_), .ZN(new_n36182_));
  NAND2_X1   g32876(.A1(new_n35861_), .A2(new_n36170_), .ZN(new_n36183_));
  NAND2_X1   g32877(.A1(new_n36147_), .A2(pi0557), .ZN(new_n36184_));
  AOI21_X1   g32878(.A1(new_n36184_), .A2(new_n36183_), .B(new_n36174_), .ZN(new_n36185_));
  INV_X1     g32879(.I(new_n36177_), .ZN(new_n36186_));
  NAND2_X1   g32880(.A1(new_n36185_), .A2(new_n36186_), .ZN(new_n36187_));
  NAND3_X1   g32881(.A1(new_n36187_), .A2(pi0579), .A3(new_n36182_), .ZN(new_n36188_));
  NOR2_X1    g32882(.A1(new_n36166_), .A2(new_n3810_), .ZN(new_n36189_));
  OAI21_X1   g32883(.A1(new_n36189_), .A2(new_n36185_), .B(pi0538), .ZN(new_n36190_));
  AOI21_X1   g32884(.A1(new_n36179_), .A2(new_n36188_), .B(new_n36190_), .ZN(new_n36191_));
  NAND4_X1   g32885(.A1(new_n36191_), .A2(pi0248), .A3(pi0537), .A4(new_n36168_), .ZN(new_n36192_));
  NOR2_X1    g32886(.A1(new_n36187_), .A2(pi0481), .ZN(new_n36193_));
  INV_X1     g32887(.I(new_n36193_), .ZN(new_n36194_));
  AOI21_X1   g32888(.A1(new_n36192_), .A2(new_n35953_), .B(new_n36194_), .ZN(new_n36195_));
  INV_X1     g32889(.I(new_n36195_), .ZN(new_n36196_));
  NAND2_X1   g32890(.A1(new_n36168_), .A2(pi0248), .ZN(new_n36197_));
  NAND3_X1   g32891(.A1(new_n36191_), .A2(pi0248), .A3(pi0537), .ZN(new_n36198_));
  NOR3_X1    g32892(.A1(new_n36187_), .A2(new_n36121_), .A3(new_n36182_), .ZN(new_n36199_));
  NOR3_X1    g32893(.A1(new_n36178_), .A2(new_n36121_), .A3(new_n36168_), .ZN(new_n36200_));
  INV_X1     g32894(.I(new_n36190_), .ZN(new_n36201_));
  OAI21_X1   g32895(.A1(new_n36200_), .A2(new_n36199_), .B(new_n36201_), .ZN(new_n36202_));
  NAND3_X1   g32896(.A1(new_n36202_), .A2(pi0248), .A3(new_n35953_), .ZN(new_n36203_));
  AOI21_X1   g32897(.A1(new_n36203_), .A2(new_n36198_), .B(new_n36197_), .ZN(new_n36204_));
  NOR2_X1    g32898(.A1(new_n35797_), .A2(new_n35953_), .ZN(new_n36205_));
  OAI21_X1   g32899(.A1(new_n36204_), .A2(new_n36178_), .B(new_n36205_), .ZN(new_n36206_));
  NAND2_X1   g32900(.A1(new_n36206_), .A2(new_n36196_), .ZN(new_n36207_));
  XOR2_X1    g32901(.A1(pi0248), .A2(pi0537), .Z(new_n36208_));
  NOR2_X1    g32902(.A1(new_n36187_), .A2(new_n36208_), .ZN(new_n36209_));
  NAND4_X1   g32903(.A1(new_n36207_), .A2(pi0241), .A3(pi0559), .A4(new_n36209_), .ZN(new_n36210_));
  XNOR2_X1   g32904(.A1(pi0248), .A2(pi0481), .ZN(new_n36211_));
  NAND2_X1   g32905(.A1(new_n36168_), .A2(new_n36211_), .ZN(new_n36212_));
  NOR2_X1    g32906(.A1(new_n36212_), .A2(pi0506), .ZN(new_n36213_));
  INV_X1     g32907(.I(new_n36213_), .ZN(new_n36214_));
  AOI21_X1   g32908(.A1(new_n36210_), .A2(new_n36007_), .B(new_n36214_), .ZN(new_n36215_));
  INV_X1     g32909(.I(new_n36215_), .ZN(new_n36216_));
  INV_X1     g32910(.I(new_n36209_), .ZN(new_n36217_));
  NOR2_X1    g32911(.A1(new_n36217_), .A2(new_n4064_), .ZN(new_n36218_));
  INV_X1     g32912(.I(new_n36212_), .ZN(new_n36219_));
  NAND3_X1   g32913(.A1(new_n36207_), .A2(pi0241), .A3(pi0559), .ZN(new_n36220_));
  NOR3_X1    g32914(.A1(new_n36202_), .A2(new_n4225_), .A3(new_n35953_), .ZN(new_n36221_));
  NOR3_X1    g32915(.A1(new_n36191_), .A2(new_n4225_), .A3(pi0537), .ZN(new_n36222_));
  NOR2_X1    g32916(.A1(new_n36221_), .A2(new_n36222_), .ZN(new_n36223_));
  OAI21_X1   g32917(.A1(new_n36223_), .A2(new_n36197_), .B(new_n36187_), .ZN(new_n36224_));
  AOI21_X1   g32918(.A1(new_n36224_), .A2(new_n36205_), .B(new_n36195_), .ZN(new_n36225_));
  NAND3_X1   g32919(.A1(new_n36225_), .A2(pi0241), .A3(new_n36007_), .ZN(new_n36226_));
  NAND2_X1   g32920(.A1(new_n36226_), .A2(new_n36220_), .ZN(new_n36227_));
  AOI21_X1   g32921(.A1(new_n36227_), .A2(new_n36218_), .B(new_n36219_), .ZN(new_n36228_));
  NOR2_X1    g32922(.A1(new_n35866_), .A2(new_n36007_), .ZN(new_n36229_));
  INV_X1     g32923(.I(new_n36229_), .ZN(new_n36230_));
  OAI21_X1   g32924(.A1(new_n36228_), .A2(new_n36230_), .B(new_n36216_), .ZN(new_n36231_));
  XOR2_X1    g32925(.A1(pi0241), .A2(pi0506), .Z(new_n36232_));
  NOR2_X1    g32926(.A1(new_n36217_), .A2(new_n36232_), .ZN(new_n36233_));
  NAND4_X1   g32927(.A1(new_n36231_), .A2(pi0240), .A3(pi0515), .A4(new_n36233_), .ZN(new_n36234_));
  XOR2_X1    g32928(.A1(pi0241), .A2(pi0559), .Z(new_n36235_));
  NOR2_X1    g32929(.A1(new_n36212_), .A2(new_n36235_), .ZN(new_n36236_));
  INV_X1     g32930(.I(new_n36236_), .ZN(new_n36237_));
  NOR2_X1    g32931(.A1(new_n36237_), .A2(pi0535), .ZN(new_n36238_));
  INV_X1     g32932(.I(new_n36238_), .ZN(new_n36239_));
  AOI21_X1   g32933(.A1(new_n36234_), .A2(new_n35898_), .B(new_n36239_), .ZN(new_n36240_));
  INV_X1     g32934(.I(new_n36233_), .ZN(new_n36241_));
  NOR2_X1    g32935(.A1(new_n36241_), .A2(new_n4710_), .ZN(new_n36242_));
  NOR3_X1    g32936(.A1(new_n36225_), .A2(new_n4064_), .A3(new_n36007_), .ZN(new_n36243_));
  NOR3_X1    g32937(.A1(new_n36207_), .A2(new_n4064_), .A3(pi0559), .ZN(new_n36244_));
  OAI21_X1   g32938(.A1(new_n36243_), .A2(new_n36244_), .B(new_n36218_), .ZN(new_n36245_));
  AOI21_X1   g32939(.A1(new_n36245_), .A2(new_n36212_), .B(new_n36230_), .ZN(new_n36246_));
  NOR2_X1    g32940(.A1(new_n36246_), .A2(new_n36215_), .ZN(new_n36247_));
  NOR3_X1    g32941(.A1(new_n36247_), .A2(new_n4710_), .A3(new_n35898_), .ZN(new_n36248_));
  NOR4_X1    g32942(.A1(new_n36246_), .A2(new_n4710_), .A3(pi0515), .A4(new_n36215_), .ZN(new_n36249_));
  OAI21_X1   g32943(.A1(new_n36248_), .A2(new_n36249_), .B(new_n36242_), .ZN(new_n36250_));
  NAND2_X1   g32944(.A1(new_n36250_), .A2(new_n36237_), .ZN(new_n36251_));
  NOR2_X1    g32945(.A1(new_n35898_), .A2(new_n35947_), .ZN(new_n36252_));
  AOI21_X1   g32946(.A1(new_n36251_), .A2(new_n36252_), .B(new_n36240_), .ZN(new_n36253_));
  NOR3_X1    g32947(.A1(new_n36253_), .A2(new_n35831_), .A3(new_n36160_), .ZN(new_n36254_));
  INV_X1     g32948(.I(new_n36252_), .ZN(new_n36255_));
  AOI21_X1   g32949(.A1(new_n36250_), .A2(new_n36237_), .B(new_n36255_), .ZN(new_n36256_));
  NOR4_X1    g32950(.A1(new_n36256_), .A2(new_n35831_), .A3(pi0534), .A4(new_n36240_), .ZN(new_n36257_));
  XOR2_X1    g32951(.A1(pi0240), .A2(pi0515), .Z(new_n36258_));
  NOR2_X1    g32952(.A1(new_n36237_), .A2(new_n36258_), .ZN(new_n36259_));
  INV_X1     g32953(.I(new_n36259_), .ZN(new_n36260_));
  NOR2_X1    g32954(.A1(new_n36260_), .A2(new_n35831_), .ZN(new_n36261_));
  OAI21_X1   g32955(.A1(new_n36254_), .A2(new_n36257_), .B(new_n36261_), .ZN(new_n36262_));
  XOR2_X1    g32956(.A1(pi0240), .A2(pi0535), .Z(new_n36263_));
  NOR2_X1    g32957(.A1(new_n36241_), .A2(new_n36263_), .ZN(new_n36264_));
  INV_X1     g32958(.I(new_n36264_), .ZN(new_n36265_));
  NOR2_X1    g32959(.A1(new_n36265_), .A2(pi0488), .ZN(new_n36266_));
  INV_X1     g32960(.I(new_n36266_), .ZN(new_n36267_));
  AOI21_X1   g32961(.A1(new_n36262_), .A2(new_n36160_), .B(new_n36267_), .ZN(new_n36268_));
  NOR4_X1    g32962(.A1(new_n36253_), .A2(new_n35831_), .A3(new_n36160_), .A4(new_n36260_), .ZN(new_n36269_));
  NAND2_X1   g32963(.A1(pi0488), .A2(pi0534), .ZN(new_n36270_));
  INV_X1     g32964(.I(new_n36270_), .ZN(new_n36271_));
  OAI21_X1   g32965(.A1(new_n36269_), .A2(new_n36264_), .B(new_n36271_), .ZN(new_n36272_));
  INV_X1     g32966(.I(new_n36272_), .ZN(new_n36273_));
  NOR2_X1    g32967(.A1(new_n36268_), .A2(new_n36273_), .ZN(new_n36274_));
  XOR2_X1    g32968(.A1(pi0239), .A2(pi0488), .Z(new_n36275_));
  NAND2_X1   g32969(.A1(new_n36259_), .A2(new_n36275_), .ZN(new_n36276_));
  NOR4_X1    g32970(.A1(new_n36274_), .A2(new_n5364_), .A3(new_n35856_), .A4(new_n36276_), .ZN(new_n36277_));
  XNOR2_X1   g32971(.A1(pi0239), .A2(pi0534), .ZN(new_n36278_));
  NOR2_X1    g32972(.A1(new_n36265_), .A2(new_n36278_), .ZN(new_n36279_));
  INV_X1     g32973(.I(new_n36279_), .ZN(new_n36280_));
  NOR2_X1    g32974(.A1(new_n36280_), .A2(pi0510), .ZN(new_n36281_));
  OAI21_X1   g32975(.A1(new_n36277_), .A2(pi0504), .B(new_n36281_), .ZN(new_n36282_));
  NOR2_X1    g32976(.A1(new_n36276_), .A2(new_n5364_), .ZN(new_n36283_));
  INV_X1     g32977(.I(new_n36283_), .ZN(new_n36284_));
  INV_X1     g32978(.I(new_n36240_), .ZN(new_n36285_));
  INV_X1     g32979(.I(new_n36242_), .ZN(new_n36286_));
  NAND3_X1   g32980(.A1(new_n36231_), .A2(pi0240), .A3(pi0515), .ZN(new_n36287_));
  INV_X1     g32981(.I(new_n36249_), .ZN(new_n36288_));
  AOI21_X1   g32982(.A1(new_n36288_), .A2(new_n36287_), .B(new_n36286_), .ZN(new_n36289_));
  OAI21_X1   g32983(.A1(new_n36289_), .A2(new_n36236_), .B(new_n36252_), .ZN(new_n36290_));
  NAND2_X1   g32984(.A1(new_n36290_), .A2(new_n36285_), .ZN(new_n36291_));
  NAND3_X1   g32985(.A1(new_n36291_), .A2(pi0239), .A3(pi0534), .ZN(new_n36292_));
  NAND3_X1   g32986(.A1(new_n36253_), .A2(pi0239), .A3(new_n36160_), .ZN(new_n36293_));
  INV_X1     g32987(.I(new_n36261_), .ZN(new_n36294_));
  AOI21_X1   g32988(.A1(new_n36292_), .A2(new_n36293_), .B(new_n36294_), .ZN(new_n36295_));
  OAI21_X1   g32989(.A1(new_n36295_), .A2(pi0534), .B(new_n36266_), .ZN(new_n36296_));
  NAND2_X1   g32990(.A1(new_n36296_), .A2(new_n36272_), .ZN(new_n36297_));
  NAND3_X1   g32991(.A1(new_n36297_), .A2(pi0242), .A3(pi0504), .ZN(new_n36298_));
  NAND4_X1   g32992(.A1(new_n36296_), .A2(pi0242), .A3(new_n35856_), .A4(new_n36272_), .ZN(new_n36299_));
  AOI21_X1   g32993(.A1(new_n36298_), .A2(new_n36299_), .B(new_n36284_), .ZN(new_n36300_));
  NOR2_X1    g32994(.A1(new_n35856_), .A2(new_n35878_), .ZN(new_n36301_));
  OAI21_X1   g32995(.A1(new_n36300_), .A2(new_n36279_), .B(new_n36301_), .ZN(new_n36302_));
  NAND2_X1   g32996(.A1(new_n36302_), .A2(new_n36282_), .ZN(new_n36303_));
  XOR2_X1    g32997(.A1(pi0242), .A2(pi0510), .Z(new_n36304_));
  NOR2_X1    g32998(.A1(new_n36276_), .A2(new_n36304_), .ZN(new_n36305_));
  NAND4_X1   g32999(.A1(new_n36303_), .A2(pi0235), .A3(pi0533), .A4(new_n36305_), .ZN(new_n36306_));
  XOR2_X1    g33000(.A1(pi0242), .A2(pi0504), .Z(new_n36307_));
  NOR2_X1    g33001(.A1(new_n36280_), .A2(new_n36307_), .ZN(new_n36308_));
  INV_X1     g33002(.I(new_n36308_), .ZN(new_n36309_));
  NOR2_X1    g33003(.A1(new_n36309_), .A2(pi0512), .ZN(new_n36310_));
  INV_X1     g33004(.I(new_n36310_), .ZN(new_n36311_));
  AOI21_X1   g33005(.A1(new_n36306_), .A2(new_n35942_), .B(new_n36311_), .ZN(new_n36312_));
  INV_X1     g33006(.I(new_n36312_), .ZN(new_n36313_));
  INV_X1     g33007(.I(new_n36305_), .ZN(new_n36314_));
  NOR2_X1    g33008(.A1(new_n36314_), .A2(new_n3611_), .ZN(new_n36315_));
  INV_X1     g33009(.I(new_n36315_), .ZN(new_n36316_));
  NAND3_X1   g33010(.A1(new_n36303_), .A2(pi0235), .A3(pi0533), .ZN(new_n36317_));
  NAND4_X1   g33011(.A1(new_n36302_), .A2(pi0235), .A3(new_n35942_), .A4(new_n36282_), .ZN(new_n36318_));
  AOI21_X1   g33012(.A1(new_n36317_), .A2(new_n36318_), .B(new_n36316_), .ZN(new_n36319_));
  NOR2_X1    g33013(.A1(new_n35889_), .A2(new_n35942_), .ZN(new_n36320_));
  OAI21_X1   g33014(.A1(new_n36319_), .A2(new_n36308_), .B(new_n36320_), .ZN(new_n36321_));
  NAND2_X1   g33015(.A1(new_n36321_), .A2(new_n36313_), .ZN(new_n36322_));
  XOR2_X1    g33016(.A1(pi0235), .A2(pi0512), .Z(new_n36323_));
  NOR2_X1    g33017(.A1(new_n36314_), .A2(new_n36323_), .ZN(new_n36324_));
  NAND4_X1   g33018(.A1(new_n36322_), .A2(pi0244), .A3(pi0558), .A4(new_n36324_), .ZN(new_n36325_));
  XOR2_X1    g33019(.A1(pi0235), .A2(pi0533), .Z(new_n36326_));
  NOR2_X1    g33020(.A1(new_n36309_), .A2(new_n36326_), .ZN(new_n36327_));
  INV_X1     g33021(.I(new_n36327_), .ZN(new_n36328_));
  NOR2_X1    g33022(.A1(new_n36328_), .A2(pi0513), .ZN(new_n36329_));
  INV_X1     g33023(.I(new_n36329_), .ZN(new_n36330_));
  AOI21_X1   g33024(.A1(new_n36325_), .A2(new_n36004_), .B(new_n36330_), .ZN(new_n36331_));
  INV_X1     g33025(.I(new_n36331_), .ZN(new_n36332_));
  INV_X1     g33026(.I(new_n36324_), .ZN(new_n36333_));
  NOR2_X1    g33027(.A1(new_n36333_), .A2(new_n35828_), .ZN(new_n36334_));
  INV_X1     g33028(.I(new_n36334_), .ZN(new_n36335_));
  NAND3_X1   g33029(.A1(new_n36322_), .A2(pi0244), .A3(pi0558), .ZN(new_n36336_));
  NAND4_X1   g33030(.A1(new_n36321_), .A2(new_n36313_), .A3(pi0244), .A4(new_n36004_), .ZN(new_n36337_));
  AOI21_X1   g33031(.A1(new_n36336_), .A2(new_n36337_), .B(new_n36335_), .ZN(new_n36338_));
  NOR2_X1    g33032(.A1(new_n35892_), .A2(new_n36004_), .ZN(new_n36339_));
  OAI21_X1   g33033(.A1(new_n36338_), .A2(new_n36327_), .B(new_n36339_), .ZN(new_n36340_));
  NAND2_X1   g33034(.A1(new_n36340_), .A2(new_n36332_), .ZN(new_n36341_));
  XOR2_X1    g33035(.A1(pi0244), .A2(pi0513), .Z(new_n36342_));
  NOR2_X1    g33036(.A1(new_n36333_), .A2(new_n36342_), .ZN(new_n36343_));
  NAND4_X1   g33037(.A1(new_n36341_), .A2(pi0245), .A3(pi0509), .A4(new_n36343_), .ZN(new_n36344_));
  XOR2_X1    g33038(.A1(pi0244), .A2(pi0558), .Z(new_n36345_));
  NOR2_X1    g33039(.A1(new_n36328_), .A2(new_n36345_), .ZN(new_n36346_));
  INV_X1     g33040(.I(new_n36346_), .ZN(new_n36347_));
  NOR2_X1    g33041(.A1(new_n36347_), .A2(pi0514), .ZN(new_n36348_));
  INV_X1     g33042(.I(new_n36348_), .ZN(new_n36349_));
  AOI21_X1   g33043(.A1(new_n36344_), .A2(new_n35875_), .B(new_n36349_), .ZN(new_n36350_));
  INV_X1     g33044(.I(new_n36343_), .ZN(new_n36351_));
  NOR2_X1    g33045(.A1(new_n36351_), .A2(new_n4955_), .ZN(new_n36352_));
  INV_X1     g33046(.I(new_n36282_), .ZN(new_n36353_));
  NOR3_X1    g33047(.A1(new_n36274_), .A2(new_n5364_), .A3(new_n35856_), .ZN(new_n36354_));
  NOR4_X1    g33048(.A1(new_n36268_), .A2(new_n36273_), .A3(new_n5364_), .A4(pi0504), .ZN(new_n36355_));
  OAI21_X1   g33049(.A1(new_n36354_), .A2(new_n36355_), .B(new_n36283_), .ZN(new_n36356_));
  INV_X1     g33050(.I(new_n36301_), .ZN(new_n36357_));
  AOI21_X1   g33051(.A1(new_n36356_), .A2(new_n36280_), .B(new_n36357_), .ZN(new_n36358_));
  NOR2_X1    g33052(.A1(new_n36358_), .A2(new_n36353_), .ZN(new_n36359_));
  NOR3_X1    g33053(.A1(new_n36359_), .A2(new_n3611_), .A3(new_n35942_), .ZN(new_n36360_));
  NOR4_X1    g33054(.A1(new_n36358_), .A2(new_n36353_), .A3(new_n3611_), .A4(pi0533), .ZN(new_n36361_));
  OAI21_X1   g33055(.A1(new_n36360_), .A2(new_n36361_), .B(new_n36315_), .ZN(new_n36362_));
  INV_X1     g33056(.I(new_n36320_), .ZN(new_n36363_));
  AOI21_X1   g33057(.A1(new_n36362_), .A2(new_n36309_), .B(new_n36363_), .ZN(new_n36364_));
  NOR2_X1    g33058(.A1(new_n36364_), .A2(new_n36312_), .ZN(new_n36365_));
  NOR3_X1    g33059(.A1(new_n36365_), .A2(new_n35828_), .A3(new_n36004_), .ZN(new_n36366_));
  NOR4_X1    g33060(.A1(new_n36364_), .A2(new_n35828_), .A3(pi0558), .A4(new_n36312_), .ZN(new_n36367_));
  OAI21_X1   g33061(.A1(new_n36366_), .A2(new_n36367_), .B(new_n36334_), .ZN(new_n36368_));
  NAND2_X1   g33062(.A1(new_n36368_), .A2(new_n36328_), .ZN(new_n36369_));
  AOI21_X1   g33063(.A1(new_n36369_), .A2(new_n36339_), .B(new_n36331_), .ZN(new_n36370_));
  NOR3_X1    g33064(.A1(new_n36370_), .A2(new_n4955_), .A3(new_n35875_), .ZN(new_n36371_));
  INV_X1     g33065(.I(new_n36339_), .ZN(new_n36372_));
  AOI21_X1   g33066(.A1(new_n36368_), .A2(new_n36328_), .B(new_n36372_), .ZN(new_n36373_));
  NOR4_X1    g33067(.A1(new_n36373_), .A2(new_n4955_), .A3(pi0509), .A4(new_n36331_), .ZN(new_n36374_));
  OAI21_X1   g33068(.A1(new_n36371_), .A2(new_n36374_), .B(new_n36352_), .ZN(new_n36375_));
  NAND2_X1   g33069(.A1(new_n36375_), .A2(new_n36347_), .ZN(new_n36376_));
  NOR2_X1    g33070(.A1(new_n35875_), .A2(new_n35895_), .ZN(new_n36377_));
  AOI21_X1   g33071(.A1(new_n36376_), .A2(new_n36377_), .B(new_n36350_), .ZN(new_n36378_));
  XOR2_X1    g33072(.A1(pi0245), .A2(pi0514), .Z(new_n36379_));
  NOR2_X1    g33073(.A1(new_n36351_), .A2(new_n36379_), .ZN(new_n36380_));
  INV_X1     g33074(.I(new_n36380_), .ZN(new_n36381_));
  NOR4_X1    g33075(.A1(new_n36378_), .A2(new_n4459_), .A3(new_n35872_), .A4(new_n36381_), .ZN(new_n36382_));
  XOR2_X1    g33076(.A1(pi0245), .A2(pi0509), .Z(new_n36383_));
  NOR2_X1    g33077(.A1(new_n36347_), .A2(new_n36383_), .ZN(new_n36384_));
  INV_X1     g33078(.I(new_n36384_), .ZN(new_n36385_));
  NOR2_X1    g33079(.A1(new_n36385_), .A2(pi0516), .ZN(new_n36386_));
  OAI21_X1   g33080(.A1(new_n36382_), .A2(pi0508), .B(new_n36386_), .ZN(new_n36387_));
  NOR2_X1    g33081(.A1(new_n36381_), .A2(new_n4459_), .ZN(new_n36388_));
  INV_X1     g33082(.I(new_n36350_), .ZN(new_n36389_));
  INV_X1     g33083(.I(new_n36352_), .ZN(new_n36390_));
  NAND3_X1   g33084(.A1(new_n36341_), .A2(pi0245), .A3(pi0509), .ZN(new_n36391_));
  NAND4_X1   g33085(.A1(new_n36340_), .A2(new_n36332_), .A3(pi0245), .A4(new_n35875_), .ZN(new_n36392_));
  AOI21_X1   g33086(.A1(new_n36391_), .A2(new_n36392_), .B(new_n36390_), .ZN(new_n36393_));
  OAI21_X1   g33087(.A1(new_n36393_), .A2(new_n36346_), .B(new_n36377_), .ZN(new_n36394_));
  NAND2_X1   g33088(.A1(new_n36394_), .A2(new_n36389_), .ZN(new_n36395_));
  NAND3_X1   g33089(.A1(new_n36395_), .A2(pi0247), .A3(pi0508), .ZN(new_n36396_));
  NAND4_X1   g33090(.A1(new_n36394_), .A2(new_n36389_), .A3(pi0247), .A4(new_n35872_), .ZN(new_n36397_));
  NAND2_X1   g33091(.A1(new_n36396_), .A2(new_n36397_), .ZN(new_n36398_));
  AOI21_X1   g33092(.A1(new_n36398_), .A2(new_n36388_), .B(new_n36384_), .ZN(new_n36399_));
  NAND2_X1   g33093(.A1(pi0508), .A2(pi0516), .ZN(new_n36400_));
  OAI21_X1   g33094(.A1(new_n36399_), .A2(new_n36400_), .B(new_n36387_), .ZN(new_n36401_));
  AOI21_X1   g33095(.A1(new_n36401_), .A2(pi0238), .B(new_n35904_), .ZN(new_n36402_));
  XOR2_X1    g33096(.A1(pi0247), .A2(pi0516), .Z(new_n36403_));
  NOR2_X1    g33097(.A1(new_n36381_), .A2(new_n36403_), .ZN(new_n36404_));
  XOR2_X1    g33098(.A1(pi0247), .A2(pi0508), .Z(new_n36405_));
  NOR2_X1    g33099(.A1(new_n36385_), .A2(new_n36405_), .ZN(new_n36406_));
  NOR2_X1    g33100(.A1(new_n36406_), .A2(new_n3743_), .ZN(new_n36407_));
  NOR2_X1    g33101(.A1(new_n3743_), .A2(new_n35904_), .ZN(new_n36408_));
  XOR2_X1    g33102(.A1(new_n36407_), .A2(new_n36408_), .Z(new_n36409_));
  NAND2_X1   g33103(.A1(new_n36409_), .A2(new_n36404_), .ZN(new_n36410_));
  NAND2_X1   g33104(.A1(new_n36410_), .A2(pi0507), .ZN(new_n36411_));
  NOR2_X1    g33105(.A1(new_n36406_), .A2(new_n35904_), .ZN(new_n36412_));
  XOR2_X1    g33106(.A1(new_n36412_), .A2(new_n36408_), .Z(new_n36413_));
  AOI21_X1   g33107(.A1(new_n36413_), .A2(new_n36404_), .B(pi0507), .ZN(new_n36414_));
  OAI21_X1   g33108(.A1(new_n36402_), .A2(new_n36411_), .B(new_n36414_), .ZN(new_n36415_));
  AOI21_X1   g33109(.A1(new_n36401_), .A2(new_n3743_), .B(pi0517), .ZN(new_n36416_));
  NAND4_X1   g33110(.A1(new_n36415_), .A2(pi0233), .A3(pi0237), .A4(new_n36416_), .ZN(new_n36417_));
  INV_X1     g33111(.I(new_n36387_), .ZN(new_n36418_));
  NOR3_X1    g33112(.A1(new_n36378_), .A2(new_n4459_), .A3(new_n35872_), .ZN(new_n36419_));
  INV_X1     g33113(.I(new_n36397_), .ZN(new_n36420_));
  OAI21_X1   g33114(.A1(new_n36419_), .A2(new_n36420_), .B(new_n36388_), .ZN(new_n36421_));
  AOI21_X1   g33115(.A1(new_n36421_), .A2(new_n36385_), .B(new_n36400_), .ZN(new_n36422_));
  OAI21_X1   g33116(.A1(new_n36422_), .A2(new_n36418_), .B(pi0238), .ZN(new_n36423_));
  AOI21_X1   g33117(.A1(new_n36423_), .A2(pi0517), .B(new_n36411_), .ZN(new_n36424_));
  INV_X1     g33118(.I(new_n36414_), .ZN(new_n36425_));
  OAI21_X1   g33119(.A1(new_n36424_), .A2(new_n36425_), .B(new_n36416_), .ZN(new_n36426_));
  NAND3_X1   g33120(.A1(new_n36426_), .A2(new_n27639_), .A3(pi0237), .ZN(new_n36427_));
  NAND2_X1   g33121(.A1(new_n36427_), .A2(new_n36417_), .ZN(new_n36428_));
  INV_X1     g33122(.I(pi0585), .ZN(new_n36429_));
  INV_X1     g33123(.I(pi0539), .ZN(new_n36430_));
  INV_X1     g33124(.I(pi0582), .ZN(new_n36431_));
  XOR2_X1    g33125(.A1(pi0248), .A2(pi0501), .Z(new_n36432_));
  XNOR2_X1   g33126(.A1(pi0249), .A2(pi0496), .ZN(new_n36433_));
  XNOR2_X1   g33127(.A1(pi0246), .A2(pi0499), .ZN(new_n36434_));
  NOR3_X1    g33128(.A1(new_n36433_), .A2(new_n36434_), .A3(new_n36432_), .ZN(new_n36435_));
  XOR2_X1    g33129(.A1(new_n35861_), .A2(new_n36435_), .Z(new_n36436_));
  NAND3_X1   g33130(.A1(new_n36436_), .A2(pi0234), .A3(pi0505), .ZN(new_n36437_));
  XOR2_X1    g33131(.A1(pi0241), .A2(pi0500), .Z(new_n36438_));
  OR2_X2     g33132(.A1(new_n36437_), .A2(new_n36438_), .Z(new_n36439_));
  INV_X1     g33133(.I(new_n36439_), .ZN(new_n36440_));
  XNOR2_X1   g33134(.A1(pi0248), .A2(pi0521), .ZN(new_n36441_));
  XNOR2_X1   g33135(.A1(pi0246), .A2(pi0520), .ZN(new_n36442_));
  XNOR2_X1   g33136(.A1(pi0249), .A2(pi0578), .ZN(new_n36443_));
  XNOR2_X1   g33137(.A1(pi0241), .A2(pi0574), .ZN(new_n36444_));
  NOR4_X1    g33138(.A1(new_n36441_), .A2(new_n36442_), .A3(new_n36443_), .A4(new_n36444_), .ZN(new_n36445_));
  XNOR2_X1   g33139(.A1(new_n35884_), .A2(new_n36445_), .ZN(new_n36446_));
  NAND3_X1   g33140(.A1(new_n36446_), .A2(pi0234), .A3(pi0518), .ZN(new_n36447_));
  NAND2_X1   g33141(.A1(new_n36447_), .A2(pi0500), .ZN(new_n36448_));
  NOR2_X1    g33142(.A1(new_n36447_), .A2(pi0500), .ZN(new_n36449_));
  NOR2_X1    g33143(.A1(new_n36449_), .A2(pi0241), .ZN(new_n36450_));
  AOI21_X1   g33144(.A1(new_n36450_), .A2(new_n36448_), .B(new_n36437_), .ZN(new_n36451_));
  NAND4_X1   g33145(.A1(new_n36451_), .A2(new_n36440_), .A3(pi0240), .A4(pi0582), .ZN(new_n36452_));
  NAND2_X1   g33146(.A1(new_n36452_), .A2(new_n36431_), .ZN(new_n36453_));
  NOR2_X1    g33147(.A1(new_n36447_), .A2(pi0542), .ZN(new_n36454_));
  NAND2_X1   g33148(.A1(new_n36453_), .A2(new_n36454_), .ZN(new_n36455_));
  NAND2_X1   g33149(.A1(new_n36451_), .A2(pi0240), .ZN(new_n36456_));
  NOR2_X1    g33150(.A1(new_n4710_), .A2(new_n36431_), .ZN(new_n36457_));
  NAND2_X1   g33151(.A1(new_n36439_), .A2(pi0240), .ZN(new_n36458_));
  XOR2_X1    g33152(.A1(new_n36458_), .A2(new_n36457_), .Z(new_n36459_));
  OAI21_X1   g33153(.A1(new_n36459_), .A2(new_n36456_), .B(new_n36447_), .ZN(new_n36460_));
  AND2_X2    g33154(.A1(pi0542), .A2(pi0582), .Z(new_n36461_));
  NAND2_X1   g33155(.A1(new_n36460_), .A2(new_n36461_), .ZN(new_n36462_));
  NAND2_X1   g33156(.A1(new_n36462_), .A2(new_n36455_), .ZN(new_n36463_));
  NAND3_X1   g33157(.A1(new_n36463_), .A2(pi0239), .A3(pi0497), .ZN(new_n36464_));
  NAND4_X1   g33158(.A1(new_n36462_), .A2(pi0239), .A3(new_n35840_), .A4(new_n36455_), .ZN(new_n36465_));
  NAND2_X1   g33159(.A1(new_n36464_), .A2(new_n36465_), .ZN(new_n36466_));
  NOR2_X1    g33160(.A1(pi0240), .A2(pi0582), .ZN(new_n36467_));
  NOR2_X1    g33161(.A1(new_n36457_), .A2(new_n36467_), .ZN(new_n36468_));
  NOR2_X1    g33162(.A1(new_n36447_), .A2(new_n36468_), .ZN(new_n36469_));
  NAND3_X1   g33163(.A1(new_n36466_), .A2(pi0239), .A3(new_n36469_), .ZN(new_n36470_));
  NAND2_X1   g33164(.A1(new_n36470_), .A2(new_n35840_), .ZN(new_n36471_));
  XOR2_X1    g33165(.A1(pi0240), .A2(pi0542), .Z(new_n36472_));
  NOR2_X1    g33166(.A1(new_n36439_), .A2(new_n36472_), .ZN(new_n36473_));
  INV_X1     g33167(.I(new_n36473_), .ZN(new_n36474_));
  NOR2_X1    g33168(.A1(new_n36474_), .A2(pi0519), .ZN(new_n36475_));
  NAND4_X1   g33169(.A1(new_n36463_), .A2(pi0239), .A3(pi0497), .A4(new_n36469_), .ZN(new_n36476_));
  NAND2_X1   g33170(.A1(pi0497), .A2(pi0519), .ZN(new_n36477_));
  AOI21_X1   g33171(.A1(new_n36476_), .A2(new_n36474_), .B(new_n36477_), .ZN(new_n36478_));
  AOI21_X1   g33172(.A1(new_n36471_), .A2(new_n36475_), .B(new_n36478_), .ZN(new_n36479_));
  XOR2_X1    g33173(.A1(pi0239), .A2(pi0519), .Z(new_n36480_));
  NAND2_X1   g33174(.A1(new_n36469_), .A2(new_n36480_), .ZN(new_n36481_));
  NOR4_X1    g33175(.A1(new_n36479_), .A2(new_n5364_), .A3(new_n36430_), .A4(new_n36481_), .ZN(new_n36482_));
  XNOR2_X1   g33176(.A1(pi0239), .A2(pi0497), .ZN(new_n36483_));
  NOR2_X1    g33177(.A1(new_n36474_), .A2(new_n36483_), .ZN(new_n36484_));
  INV_X1     g33178(.I(new_n36484_), .ZN(new_n36485_));
  NOR2_X1    g33179(.A1(new_n36485_), .A2(pi0586), .ZN(new_n36486_));
  OAI21_X1   g33180(.A1(new_n36482_), .A2(pi0539), .B(new_n36486_), .ZN(new_n36487_));
  NAND3_X1   g33181(.A1(new_n36469_), .A2(pi0242), .A3(new_n36480_), .ZN(new_n36488_));
  NAND2_X1   g33182(.A1(pi0242), .A2(pi0539), .ZN(new_n36489_));
  NAND2_X1   g33183(.A1(new_n36479_), .A2(pi0242), .ZN(new_n36490_));
  XNOR2_X1   g33184(.A1(new_n36490_), .A2(new_n36489_), .ZN(new_n36491_));
  NOR2_X1    g33185(.A1(new_n36491_), .A2(new_n36488_), .ZN(new_n36492_));
  NOR2_X1    g33186(.A1(new_n36492_), .A2(new_n36484_), .ZN(new_n36493_));
  NAND2_X1   g33187(.A1(pi0539), .A2(pi0586), .ZN(new_n36494_));
  OAI21_X1   g33188(.A1(new_n36493_), .A2(new_n36494_), .B(new_n36487_), .ZN(new_n36495_));
  XOR2_X1    g33189(.A1(pi0242), .A2(pi0586), .Z(new_n36496_));
  NOR2_X1    g33190(.A1(new_n36481_), .A2(new_n36496_), .ZN(new_n36497_));
  AND4_X2    g33191(.A1(pi0235), .A2(new_n36495_), .A3(pi0540), .A4(new_n36497_), .Z(new_n36498_));
  NAND2_X1   g33192(.A1(new_n5364_), .A2(new_n36430_), .ZN(new_n36499_));
  AOI21_X1   g33193(.A1(new_n36489_), .A2(new_n36499_), .B(new_n36485_), .ZN(new_n36500_));
  INV_X1     g33194(.I(new_n36500_), .ZN(new_n36501_));
  NOR2_X1    g33195(.A1(new_n36501_), .A2(pi0581), .ZN(new_n36502_));
  OAI21_X1   g33196(.A1(new_n36498_), .A2(pi0540), .B(new_n36502_), .ZN(new_n36503_));
  NAND2_X1   g33197(.A1(new_n36497_), .A2(pi0235), .ZN(new_n36504_));
  NAND2_X1   g33198(.A1(pi0235), .A2(pi0540), .ZN(new_n36505_));
  NOR2_X1    g33199(.A1(new_n36495_), .A2(new_n3611_), .ZN(new_n36506_));
  XOR2_X1    g33200(.A1(new_n36506_), .A2(new_n36505_), .Z(new_n36507_));
  OAI21_X1   g33201(.A1(new_n36507_), .A2(new_n36504_), .B(new_n36501_), .ZN(new_n36508_));
  NAND3_X1   g33202(.A1(new_n36508_), .A2(pi0540), .A3(pi0581), .ZN(new_n36509_));
  NAND2_X1   g33203(.A1(new_n36509_), .A2(new_n36503_), .ZN(new_n36510_));
  XOR2_X1    g33204(.A1(pi0235), .A2(pi0540), .Z(new_n36511_));
  NOR2_X1    g33205(.A1(new_n36501_), .A2(new_n36511_), .ZN(new_n36512_));
  NAND4_X1   g33206(.A1(new_n36510_), .A2(pi0244), .A3(pi0585), .A4(new_n36512_), .ZN(new_n36513_));
  NAND2_X1   g33207(.A1(new_n36513_), .A2(new_n36429_), .ZN(new_n36514_));
  XOR2_X1    g33208(.A1(pi0235), .A2(pi0581), .Z(new_n36515_));
  NOR4_X1    g33209(.A1(new_n36481_), .A2(pi0541), .A3(new_n36496_), .A4(new_n36515_), .ZN(new_n36516_));
  AND2_X2    g33210(.A1(new_n36514_), .A2(new_n36516_), .Z(new_n36517_));
  INV_X1     g33211(.I(new_n36517_), .ZN(new_n36518_));
  INV_X1     g33212(.I(new_n36512_), .ZN(new_n36519_));
  NOR2_X1    g33213(.A1(new_n36519_), .A2(new_n35828_), .ZN(new_n36520_));
  NOR3_X1    g33214(.A1(new_n36481_), .A2(new_n36496_), .A3(new_n36515_), .ZN(new_n36521_));
  NOR2_X1    g33215(.A1(new_n35828_), .A2(new_n36429_), .ZN(new_n36522_));
  NOR2_X1    g33216(.A1(new_n36510_), .A2(new_n35828_), .ZN(new_n36523_));
  XOR2_X1    g33217(.A1(new_n36523_), .A2(new_n36522_), .Z(new_n36524_));
  AOI21_X1   g33218(.A1(new_n36524_), .A2(new_n36520_), .B(new_n36521_), .ZN(new_n36525_));
  NAND2_X1   g33219(.A1(pi0541), .A2(pi0585), .ZN(new_n36526_));
  OAI21_X1   g33220(.A1(new_n36525_), .A2(new_n36526_), .B(new_n36518_), .ZN(new_n36527_));
  XOR2_X1    g33221(.A1(pi0244), .A2(pi0541), .Z(new_n36528_));
  NOR2_X1    g33222(.A1(new_n36519_), .A2(new_n36528_), .ZN(new_n36529_));
  AND4_X2    g33223(.A1(pi0245), .A2(new_n36527_), .A3(pi0584), .A4(new_n36529_), .Z(new_n36530_));
  NOR2_X1    g33224(.A1(pi0244), .A2(pi0585), .ZN(new_n36531_));
  OAI21_X1   g33225(.A1(new_n36522_), .A2(new_n36531_), .B(new_n36521_), .ZN(new_n36532_));
  NOR2_X1    g33226(.A1(new_n36532_), .A2(pi0503), .ZN(new_n36533_));
  OAI21_X1   g33227(.A1(new_n36530_), .A2(pi0584), .B(new_n36533_), .ZN(new_n36534_));
  INV_X1     g33228(.I(new_n36529_), .ZN(new_n36535_));
  NOR2_X1    g33229(.A1(new_n36535_), .A2(new_n4955_), .ZN(new_n36536_));
  INV_X1     g33230(.I(new_n36532_), .ZN(new_n36537_));
  NAND3_X1   g33231(.A1(new_n36527_), .A2(pi0245), .A3(pi0584), .ZN(new_n36538_));
  NOR3_X1    g33232(.A1(new_n36527_), .A2(new_n4955_), .A3(pi0584), .ZN(new_n36539_));
  INV_X1     g33233(.I(new_n36539_), .ZN(new_n36540_));
  NAND2_X1   g33234(.A1(new_n36540_), .A2(new_n36538_), .ZN(new_n36541_));
  AOI21_X1   g33235(.A1(new_n36541_), .A2(new_n36536_), .B(new_n36537_), .ZN(new_n36542_));
  NAND2_X1   g33236(.A1(pi0503), .A2(pi0584), .ZN(new_n36543_));
  OAI21_X1   g33237(.A1(new_n36542_), .A2(new_n36543_), .B(new_n36534_), .ZN(new_n36544_));
  NAND3_X1   g33238(.A1(new_n36544_), .A2(pi0502), .A3(pi0561), .ZN(new_n36545_));
  INV_X1     g33239(.I(pi0502), .ZN(new_n36546_));
  INV_X1     g33240(.I(new_n36544_), .ZN(new_n36547_));
  NAND3_X1   g33241(.A1(new_n36547_), .A2(new_n36546_), .A3(pi0561), .ZN(new_n36548_));
  NAND2_X1   g33242(.A1(new_n36548_), .A2(new_n36545_), .ZN(new_n36549_));
  XOR2_X1    g33243(.A1(pi0245), .A2(pi0503), .Z(new_n36550_));
  NOR2_X1    g33244(.A1(new_n36535_), .A2(new_n36550_), .ZN(new_n36551_));
  NOR3_X1    g33245(.A1(new_n36551_), .A2(pi0247), .A3(pi0561), .ZN(new_n36552_));
  XOR2_X1    g33246(.A1(pi0245), .A2(pi0584), .Z(new_n36553_));
  NOR2_X1    g33247(.A1(new_n36532_), .A2(new_n36553_), .ZN(new_n36554_));
  INV_X1     g33248(.I(new_n36554_), .ZN(new_n36555_));
  NOR3_X1    g33249(.A1(new_n36552_), .A2(new_n36546_), .A3(new_n36555_), .ZN(new_n36556_));
  AND2_X2    g33250(.A1(new_n36549_), .A2(new_n36556_), .Z(new_n36557_));
  INV_X1     g33251(.I(pi0561), .ZN(new_n36558_));
  NOR3_X1    g33252(.A1(new_n36547_), .A2(new_n36546_), .A3(new_n36558_), .ZN(new_n36559_));
  NOR3_X1    g33253(.A1(new_n36544_), .A2(new_n36546_), .A3(pi0561), .ZN(new_n36560_));
  NOR3_X1    g33254(.A1(new_n36551_), .A2(pi0247), .A3(pi0502), .ZN(new_n36561_));
  NOR3_X1    g33255(.A1(new_n36561_), .A2(new_n36558_), .A3(new_n36555_), .ZN(new_n36562_));
  OAI21_X1   g33256(.A1(new_n36559_), .A2(new_n36560_), .B(new_n36562_), .ZN(new_n36563_));
  INV_X1     g33257(.I(new_n36563_), .ZN(new_n36564_));
  NOR2_X1    g33258(.A1(new_n36557_), .A2(new_n36564_), .ZN(new_n36565_));
  OAI21_X1   g33259(.A1(new_n36565_), .A2(new_n3743_), .B(pi0522), .ZN(new_n36566_));
  INV_X1     g33260(.I(pi0543), .ZN(new_n36567_));
  XOR2_X1    g33261(.A1(pi0247), .A2(pi0561), .Z(new_n36568_));
  NOR2_X1    g33262(.A1(new_n36555_), .A2(new_n36568_), .ZN(new_n36569_));
  XNOR2_X1   g33263(.A1(pi0247), .A2(pi0502), .ZN(new_n36570_));
  NAND2_X1   g33264(.A1(new_n36551_), .A2(new_n36570_), .ZN(new_n36571_));
  NAND2_X1   g33265(.A1(new_n36571_), .A2(pi0238), .ZN(new_n36572_));
  NAND2_X1   g33266(.A1(pi0238), .A2(pi0522), .ZN(new_n36573_));
  XOR2_X1    g33267(.A1(new_n36572_), .A2(new_n36573_), .Z(new_n36574_));
  AOI21_X1   g33268(.A1(new_n36574_), .A2(new_n36569_), .B(new_n36567_), .ZN(new_n36575_));
  NAND2_X1   g33269(.A1(new_n36566_), .A2(new_n36575_), .ZN(new_n36576_));
  NAND2_X1   g33270(.A1(new_n36571_), .A2(pi0522), .ZN(new_n36577_));
  XOR2_X1    g33271(.A1(new_n36577_), .A2(new_n36573_), .Z(new_n36578_));
  AOI21_X1   g33272(.A1(new_n36578_), .A2(new_n36569_), .B(pi0543), .ZN(new_n36579_));
  INV_X1     g33273(.I(pi0522), .ZN(new_n36580_));
  OAI21_X1   g33274(.A1(new_n36565_), .A2(pi0238), .B(new_n36580_), .ZN(new_n36581_));
  AOI21_X1   g33275(.A1(new_n36576_), .A2(new_n36579_), .B(new_n36581_), .ZN(new_n36582_));
  INV_X1     g33276(.I(pi0529), .ZN(new_n36583_));
  INV_X1     g33277(.I(pi0547), .ZN(new_n36584_));
  INV_X1     g33278(.I(pi0545), .ZN(new_n36585_));
  INV_X1     g33279(.I(pi0572), .ZN(new_n36586_));
  INV_X1     g33280(.I(pi0495), .ZN(new_n36587_));
  INV_X1     g33281(.I(pi0483), .ZN(new_n36588_));
  INV_X1     g33282(.I(pi0571), .ZN(new_n36589_));
  XOR2_X1    g33283(.A1(pi0249), .A2(pi0528), .Z(new_n36590_));
  XNOR2_X1   g33284(.A1(pi0248), .A2(pi0576), .ZN(new_n36591_));
  XNOR2_X1   g33285(.A1(pi0246), .A2(pi0526), .ZN(new_n36592_));
  NOR3_X1    g33286(.A1(new_n36591_), .A2(new_n36592_), .A3(new_n36590_), .ZN(new_n36593_));
  XNOR2_X1   g33287(.A1(new_n35884_), .A2(new_n36593_), .ZN(new_n36594_));
  NAND3_X1   g33288(.A1(new_n36594_), .A2(pi0234), .A3(pi0523), .ZN(new_n36595_));
  NOR2_X1    g33289(.A1(new_n36595_), .A2(new_n36589_), .ZN(new_n36596_));
  XOR2_X1    g33290(.A1(pi0249), .A2(pi0484), .Z(new_n36597_));
  XNOR2_X1   g33291(.A1(pi0248), .A2(pi0548), .ZN(new_n36598_));
  XNOR2_X1   g33292(.A1(pi0246), .A2(pi0546), .ZN(new_n36599_));
  NOR3_X1    g33293(.A1(new_n36598_), .A2(new_n36599_), .A3(new_n36597_), .ZN(new_n36600_));
  XOR2_X1    g33294(.A1(new_n35861_), .A2(new_n36600_), .Z(new_n36601_));
  NAND3_X1   g33295(.A1(new_n36601_), .A2(pi0234), .A3(pi0544), .ZN(new_n36602_));
  XNOR2_X1   g33296(.A1(pi0241), .A2(pi0571), .ZN(new_n36603_));
  NOR2_X1    g33297(.A1(new_n36602_), .A2(new_n36603_), .ZN(new_n36604_));
  NOR2_X1    g33298(.A1(new_n36604_), .A2(new_n36596_), .ZN(new_n36605_));
  NOR2_X1    g33299(.A1(new_n36605_), .A2(pi0490), .ZN(new_n36606_));
  INV_X1     g33300(.I(pi0490), .ZN(new_n36607_));
  NOR2_X1    g33301(.A1(new_n36605_), .A2(new_n36607_), .ZN(new_n36608_));
  NOR2_X1    g33302(.A1(new_n36606_), .A2(new_n36608_), .ZN(new_n36609_));
  NAND2_X1   g33303(.A1(new_n36609_), .A2(pi0492), .ZN(new_n36610_));
  NAND2_X1   g33304(.A1(pi0492), .A2(pi0530), .ZN(new_n36611_));
  XOR2_X1    g33305(.A1(new_n36610_), .A2(new_n36611_), .Z(new_n36612_));
  XOR2_X1    g33306(.A1(pi0241), .A2(pi0571), .Z(new_n36613_));
  NOR2_X1    g33307(.A1(new_n36595_), .A2(new_n36613_), .ZN(new_n36614_));
  NOR3_X1    g33308(.A1(new_n36614_), .A2(pi0240), .A3(pi0492), .ZN(new_n36615_));
  XOR2_X1    g33309(.A1(pi0241), .A2(pi0490), .Z(new_n36616_));
  NOR2_X1    g33310(.A1(new_n36602_), .A2(new_n36616_), .ZN(new_n36617_));
  NAND2_X1   g33311(.A1(new_n36617_), .A2(pi0530), .ZN(new_n36618_));
  NOR2_X1    g33312(.A1(new_n36618_), .A2(new_n36615_), .ZN(new_n36619_));
  NAND2_X1   g33313(.A1(new_n36612_), .A2(new_n36619_), .ZN(new_n36620_));
  NAND2_X1   g33314(.A1(new_n36609_), .A2(pi0530), .ZN(new_n36621_));
  XOR2_X1    g33315(.A1(new_n36621_), .A2(new_n36611_), .Z(new_n36622_));
  NOR3_X1    g33316(.A1(new_n36614_), .A2(pi0240), .A3(pi0530), .ZN(new_n36623_));
  NAND2_X1   g33317(.A1(new_n36617_), .A2(pi0492), .ZN(new_n36624_));
  NOR2_X1    g33318(.A1(new_n36624_), .A2(new_n36623_), .ZN(new_n36625_));
  NAND2_X1   g33319(.A1(new_n36622_), .A2(new_n36625_), .ZN(new_n36626_));
  NAND2_X1   g33320(.A1(new_n36620_), .A2(new_n36626_), .ZN(new_n36627_));
  NAND3_X1   g33321(.A1(new_n36627_), .A2(pi0239), .A3(pi0494), .ZN(new_n36628_));
  NAND4_X1   g33322(.A1(new_n36620_), .A2(new_n36626_), .A3(pi0239), .A4(new_n35832_), .ZN(new_n36629_));
  NAND2_X1   g33323(.A1(new_n36628_), .A2(new_n36629_), .ZN(new_n36630_));
  XNOR2_X1   g33324(.A1(pi0240), .A2(pi0530), .ZN(new_n36631_));
  NAND2_X1   g33325(.A1(new_n36614_), .A2(new_n36631_), .ZN(new_n36632_));
  INV_X1     g33326(.I(new_n36632_), .ZN(new_n36633_));
  NAND3_X1   g33327(.A1(new_n36630_), .A2(pi0239), .A3(new_n36633_), .ZN(new_n36634_));
  NAND2_X1   g33328(.A1(new_n36634_), .A2(new_n35832_), .ZN(new_n36635_));
  XNOR2_X1   g33329(.A1(pi0240), .A2(pi0492), .ZN(new_n36636_));
  NAND2_X1   g33330(.A1(new_n36617_), .A2(new_n36636_), .ZN(new_n36637_));
  NOR2_X1    g33331(.A1(new_n36637_), .A2(pi0524), .ZN(new_n36638_));
  NAND4_X1   g33332(.A1(new_n36627_), .A2(pi0239), .A3(pi0494), .A4(new_n36633_), .ZN(new_n36639_));
  NAND2_X1   g33333(.A1(new_n36639_), .A2(new_n36637_), .ZN(new_n36640_));
  NOR2_X1    g33334(.A1(new_n35832_), .A2(new_n35921_), .ZN(new_n36641_));
  AOI22_X1   g33335(.A1(new_n36635_), .A2(new_n36638_), .B1(new_n36640_), .B2(new_n36641_), .ZN(new_n36642_));
  XNOR2_X1   g33336(.A1(pi0239), .A2(pi0524), .ZN(new_n36643_));
  NOR2_X1    g33337(.A1(new_n36632_), .A2(new_n36643_), .ZN(new_n36644_));
  INV_X1     g33338(.I(new_n36644_), .ZN(new_n36645_));
  NOR4_X1    g33339(.A1(new_n36642_), .A2(new_n5364_), .A3(new_n36588_), .A4(new_n36645_), .ZN(new_n36646_));
  XNOR2_X1   g33340(.A1(pi0239), .A2(pi0494), .ZN(new_n36647_));
  NOR2_X1    g33341(.A1(new_n36637_), .A2(new_n36647_), .ZN(new_n36648_));
  INV_X1     g33342(.I(new_n36648_), .ZN(new_n36649_));
  NOR2_X1    g33343(.A1(new_n36649_), .A2(pi0573), .ZN(new_n36650_));
  OAI21_X1   g33344(.A1(new_n36646_), .A2(pi0483), .B(new_n36650_), .ZN(new_n36651_));
  NAND2_X1   g33345(.A1(new_n36644_), .A2(pi0242), .ZN(new_n36652_));
  NAND2_X1   g33346(.A1(pi0242), .A2(pi0483), .ZN(new_n36653_));
  NAND2_X1   g33347(.A1(new_n36642_), .A2(pi0242), .ZN(new_n36654_));
  XNOR2_X1   g33348(.A1(new_n36654_), .A2(new_n36653_), .ZN(new_n36655_));
  OAI21_X1   g33349(.A1(new_n36655_), .A2(new_n36652_), .B(new_n36649_), .ZN(new_n36656_));
  NAND3_X1   g33350(.A1(new_n36656_), .A2(pi0483), .A3(pi0573), .ZN(new_n36657_));
  NAND2_X1   g33351(.A1(new_n36657_), .A2(new_n36651_), .ZN(new_n36658_));
  INV_X1     g33352(.I(new_n36658_), .ZN(new_n36659_));
  XOR2_X1    g33353(.A1(pi0242), .A2(pi0573), .Z(new_n36660_));
  NOR2_X1    g33354(.A1(new_n36645_), .A2(new_n36660_), .ZN(new_n36661_));
  INV_X1     g33355(.I(new_n36661_), .ZN(new_n36662_));
  NOR4_X1    g33356(.A1(new_n36659_), .A2(new_n3611_), .A3(new_n36587_), .A4(new_n36662_), .ZN(new_n36663_));
  XOR2_X1    g33357(.A1(pi0242), .A2(pi0483), .Z(new_n36664_));
  NOR2_X1    g33358(.A1(new_n36649_), .A2(new_n36664_), .ZN(new_n36665_));
  INV_X1     g33359(.I(new_n36665_), .ZN(new_n36666_));
  NOR2_X1    g33360(.A1(new_n36666_), .A2(pi0575), .ZN(new_n36667_));
  OAI21_X1   g33361(.A1(new_n36663_), .A2(pi0495), .B(new_n36667_), .ZN(new_n36668_));
  NOR2_X1    g33362(.A1(new_n36662_), .A2(new_n3611_), .ZN(new_n36669_));
  INV_X1     g33363(.I(new_n36669_), .ZN(new_n36670_));
  NAND3_X1   g33364(.A1(new_n36658_), .A2(pi0235), .A3(pi0495), .ZN(new_n36671_));
  NAND3_X1   g33365(.A1(new_n36659_), .A2(pi0235), .A3(new_n36587_), .ZN(new_n36672_));
  AOI21_X1   g33366(.A1(new_n36672_), .A2(new_n36671_), .B(new_n36670_), .ZN(new_n36673_));
  AND2_X2    g33367(.A1(pi0495), .A2(pi0575), .Z(new_n36674_));
  OAI21_X1   g33368(.A1(new_n36673_), .A2(new_n36665_), .B(new_n36674_), .ZN(new_n36675_));
  NAND2_X1   g33369(.A1(new_n36675_), .A2(new_n36668_), .ZN(new_n36676_));
  XOR2_X1    g33370(.A1(pi0235), .A2(pi0495), .Z(new_n36677_));
  NOR2_X1    g33371(.A1(new_n36666_), .A2(new_n36677_), .ZN(new_n36678_));
  NAND4_X1   g33372(.A1(new_n36676_), .A2(pi0244), .A3(pi0572), .A4(new_n36678_), .ZN(new_n36679_));
  NAND2_X1   g33373(.A1(new_n36679_), .A2(new_n36586_), .ZN(new_n36680_));
  XOR2_X1    g33374(.A1(pi0235), .A2(pi0575), .Z(new_n36681_));
  NOR2_X1    g33375(.A1(new_n36662_), .A2(new_n36681_), .ZN(new_n36682_));
  INV_X1     g33376(.I(new_n36682_), .ZN(new_n36683_));
  NOR2_X1    g33377(.A1(new_n36683_), .A2(pi0493), .ZN(new_n36684_));
  NAND2_X1   g33378(.A1(new_n36680_), .A2(new_n36684_), .ZN(new_n36685_));
  INV_X1     g33379(.I(new_n36678_), .ZN(new_n36686_));
  NOR2_X1    g33380(.A1(new_n36686_), .A2(new_n35828_), .ZN(new_n36687_));
  NAND3_X1   g33381(.A1(new_n36676_), .A2(pi0244), .A3(pi0572), .ZN(new_n36688_));
  NOR3_X1    g33382(.A1(new_n36676_), .A2(new_n35828_), .A3(pi0572), .ZN(new_n36689_));
  INV_X1     g33383(.I(new_n36689_), .ZN(new_n36690_));
  NAND2_X1   g33384(.A1(new_n36690_), .A2(new_n36688_), .ZN(new_n36691_));
  AOI21_X1   g33385(.A1(new_n36691_), .A2(new_n36687_), .B(new_n36682_), .ZN(new_n36692_));
  NAND2_X1   g33386(.A1(pi0493), .A2(pi0572), .ZN(new_n36693_));
  OAI21_X1   g33387(.A1(new_n36692_), .A2(new_n36693_), .B(new_n36685_), .ZN(new_n36694_));
  XOR2_X1    g33388(.A1(pi0244), .A2(pi0572), .Z(new_n36695_));
  NOR2_X1    g33389(.A1(new_n36683_), .A2(new_n36695_), .ZN(new_n36696_));
  NAND4_X1   g33390(.A1(new_n36694_), .A2(pi0245), .A3(pi0545), .A4(new_n36696_), .ZN(new_n36697_));
  NAND2_X1   g33391(.A1(new_n36697_), .A2(new_n36585_), .ZN(new_n36698_));
  XOR2_X1    g33392(.A1(pi0244), .A2(pi0493), .Z(new_n36699_));
  NOR2_X1    g33393(.A1(new_n36686_), .A2(new_n36699_), .ZN(new_n36700_));
  INV_X1     g33394(.I(new_n36700_), .ZN(new_n36701_));
  NOR2_X1    g33395(.A1(new_n36701_), .A2(pi0525), .ZN(new_n36702_));
  NAND2_X1   g33396(.A1(new_n36698_), .A2(new_n36702_), .ZN(new_n36703_));
  INV_X1     g33397(.I(new_n36696_), .ZN(new_n36704_));
  NOR2_X1    g33398(.A1(new_n36704_), .A2(new_n4955_), .ZN(new_n36705_));
  NAND3_X1   g33399(.A1(new_n36694_), .A2(pi0245), .A3(pi0545), .ZN(new_n36706_));
  INV_X1     g33400(.I(new_n36688_), .ZN(new_n36707_));
  OAI21_X1   g33401(.A1(new_n36707_), .A2(new_n36689_), .B(new_n36687_), .ZN(new_n36708_));
  NAND2_X1   g33402(.A1(new_n36708_), .A2(new_n36683_), .ZN(new_n36709_));
  INV_X1     g33403(.I(new_n36693_), .ZN(new_n36710_));
  AOI22_X1   g33404(.A1(new_n36709_), .A2(new_n36710_), .B1(new_n36680_), .B2(new_n36684_), .ZN(new_n36711_));
  NAND3_X1   g33405(.A1(new_n36711_), .A2(pi0245), .A3(new_n36585_), .ZN(new_n36712_));
  NAND2_X1   g33406(.A1(new_n36712_), .A2(new_n36706_), .ZN(new_n36713_));
  AOI21_X1   g33407(.A1(new_n36713_), .A2(new_n36705_), .B(new_n36700_), .ZN(new_n36714_));
  NAND2_X1   g33408(.A1(pi0525), .A2(pi0545), .ZN(new_n36715_));
  OAI21_X1   g33409(.A1(new_n36714_), .A2(new_n36715_), .B(new_n36703_), .ZN(new_n36716_));
  XOR2_X1    g33410(.A1(pi0245), .A2(pi0525), .Z(new_n36717_));
  NOR2_X1    g33411(.A1(new_n36704_), .A2(new_n36717_), .ZN(new_n36718_));
  NAND4_X1   g33412(.A1(new_n36716_), .A2(pi0247), .A3(pi0547), .A4(new_n36718_), .ZN(new_n36719_));
  NAND2_X1   g33413(.A1(new_n36719_), .A2(new_n36584_), .ZN(new_n36720_));
  XOR2_X1    g33414(.A1(pi0245), .A2(pi0545), .Z(new_n36721_));
  NOR2_X1    g33415(.A1(new_n36701_), .A2(new_n36721_), .ZN(new_n36722_));
  INV_X1     g33416(.I(new_n36722_), .ZN(new_n36723_));
  NOR2_X1    g33417(.A1(new_n36723_), .A2(pi0527), .ZN(new_n36724_));
  NAND2_X1   g33418(.A1(new_n36720_), .A2(new_n36724_), .ZN(new_n36725_));
  INV_X1     g33419(.I(new_n36718_), .ZN(new_n36726_));
  NOR2_X1    g33420(.A1(new_n36726_), .A2(new_n4459_), .ZN(new_n36727_));
  NAND3_X1   g33421(.A1(new_n36716_), .A2(pi0247), .A3(pi0547), .ZN(new_n36728_));
  NOR3_X1    g33422(.A1(new_n36711_), .A2(new_n4955_), .A3(new_n36585_), .ZN(new_n36729_));
  NOR3_X1    g33423(.A1(new_n36694_), .A2(new_n4955_), .A3(pi0545), .ZN(new_n36730_));
  OAI21_X1   g33424(.A1(new_n36729_), .A2(new_n36730_), .B(new_n36705_), .ZN(new_n36731_));
  NAND2_X1   g33425(.A1(new_n36731_), .A2(new_n36701_), .ZN(new_n36732_));
  INV_X1     g33426(.I(new_n36715_), .ZN(new_n36733_));
  NAND2_X1   g33427(.A1(new_n36732_), .A2(new_n36733_), .ZN(new_n36734_));
  NAND4_X1   g33428(.A1(new_n36734_), .A2(pi0247), .A3(new_n36584_), .A4(new_n36703_), .ZN(new_n36735_));
  NAND2_X1   g33429(.A1(new_n36728_), .A2(new_n36735_), .ZN(new_n36736_));
  AOI21_X1   g33430(.A1(new_n36736_), .A2(new_n36727_), .B(new_n36722_), .ZN(new_n36737_));
  NAND2_X1   g33431(.A1(pi0527), .A2(pi0547), .ZN(new_n36738_));
  OAI21_X1   g33432(.A1(new_n36737_), .A2(new_n36738_), .B(new_n36725_), .ZN(new_n36739_));
  AOI21_X1   g33433(.A1(new_n36739_), .A2(pi0238), .B(new_n36583_), .ZN(new_n36740_));
  XOR2_X1    g33434(.A1(pi0247), .A2(pi0527), .Z(new_n36741_));
  NOR2_X1    g33435(.A1(new_n36726_), .A2(new_n36741_), .ZN(new_n36742_));
  XNOR2_X1   g33436(.A1(pi0247), .A2(pi0547), .ZN(new_n36743_));
  NAND2_X1   g33437(.A1(new_n36722_), .A2(new_n36743_), .ZN(new_n36744_));
  NAND2_X1   g33438(.A1(new_n36744_), .A2(pi0238), .ZN(new_n36745_));
  NAND2_X1   g33439(.A1(pi0238), .A2(pi0529), .ZN(new_n36746_));
  XOR2_X1    g33440(.A1(new_n36745_), .A2(new_n36746_), .Z(new_n36747_));
  NAND2_X1   g33441(.A1(new_n36747_), .A2(new_n36742_), .ZN(new_n36748_));
  NAND2_X1   g33442(.A1(new_n36748_), .A2(pi0491), .ZN(new_n36749_));
  NAND2_X1   g33443(.A1(new_n36744_), .A2(pi0529), .ZN(new_n36750_));
  XOR2_X1    g33444(.A1(new_n36750_), .A2(new_n36746_), .Z(new_n36751_));
  AOI21_X1   g33445(.A1(new_n36751_), .A2(new_n36742_), .B(pi0491), .ZN(new_n36752_));
  OAI21_X1   g33446(.A1(new_n36740_), .A2(new_n36749_), .B(new_n36752_), .ZN(new_n36753_));
  AOI21_X1   g33447(.A1(new_n36739_), .A2(new_n3743_), .B(pi0529), .ZN(new_n36754_));
  NAND4_X1   g33448(.A1(new_n36753_), .A2(pi0233), .A3(pi0237), .A4(new_n36754_), .ZN(new_n36755_));
  INV_X1     g33449(.I(new_n36725_), .ZN(new_n36756_));
  INV_X1     g33450(.I(new_n36728_), .ZN(new_n36757_));
  NOR3_X1    g33451(.A1(new_n36716_), .A2(new_n4459_), .A3(pi0547), .ZN(new_n36758_));
  OAI21_X1   g33452(.A1(new_n36757_), .A2(new_n36758_), .B(new_n36727_), .ZN(new_n36759_));
  AOI21_X1   g33453(.A1(new_n36759_), .A2(new_n36723_), .B(new_n36738_), .ZN(new_n36760_));
  OAI21_X1   g33454(.A1(new_n36760_), .A2(new_n36756_), .B(pi0238), .ZN(new_n36761_));
  AOI21_X1   g33455(.A1(new_n36761_), .A2(pi0529), .B(new_n36749_), .ZN(new_n36762_));
  INV_X1     g33456(.I(new_n36752_), .ZN(new_n36763_));
  OAI21_X1   g33457(.A1(new_n36762_), .A2(new_n36763_), .B(new_n36754_), .ZN(new_n36764_));
  NAND3_X1   g33458(.A1(new_n36764_), .A2(pi0233), .A3(new_n27640_), .ZN(new_n36765_));
  XOR2_X1    g33459(.A1(pi0241), .A2(pi0562), .Z(new_n36766_));
  XNOR2_X1   g33460(.A1(pi0249), .A2(pi0482), .ZN(new_n36767_));
  NOR2_X1    g33461(.A1(pi0246), .A2(pi0564), .ZN(new_n36768_));
  NOR3_X1    g33462(.A1(new_n36767_), .A2(new_n36766_), .A3(new_n36768_), .ZN(new_n36769_));
  XNOR2_X1   g33463(.A1(new_n35884_), .A2(new_n36769_), .ZN(new_n36770_));
  NAND3_X1   g33464(.A1(new_n36770_), .A2(pi0234), .A3(pi0570), .ZN(new_n36771_));
  NAND2_X1   g33465(.A1(new_n36771_), .A2(pi0240), .ZN(new_n36772_));
  NOR2_X1    g33466(.A1(new_n36010_), .A2(pi0240), .ZN(new_n36773_));
  NOR2_X1    g33467(.A1(new_n4710_), .A2(pi0560), .ZN(new_n36774_));
  OAI22_X1   g33468(.A1(new_n36773_), .A2(new_n36774_), .B1(pi0246), .B2(pi0564), .ZN(new_n36775_));
  XOR2_X1    g33469(.A1(new_n36771_), .A2(new_n36775_), .Z(new_n36776_));
  NOR2_X1    g33470(.A1(new_n4549_), .A2(pi0564), .ZN(new_n36777_));
  NOR3_X1    g33471(.A1(new_n36777_), .A2(new_n4710_), .A3(new_n36010_), .ZN(new_n36778_));
  NAND4_X1   g33472(.A1(new_n36776_), .A2(pi0248), .A3(pi0565), .A4(new_n36778_), .ZN(new_n36779_));
  XOR2_X1    g33473(.A1(new_n36779_), .A2(new_n36772_), .Z(new_n36780_));
  XOR2_X1    g33474(.A1(pi0239), .A2(pi0569), .Z(new_n36781_));
  NAND2_X1   g33475(.A1(new_n36780_), .A2(new_n36781_), .ZN(new_n36782_));
  NAND2_X1   g33476(.A1(new_n36782_), .A2(pi0556), .ZN(new_n36783_));
  NAND2_X1   g33477(.A1(pi0489), .A2(pi0556), .ZN(new_n36784_));
  XOR2_X1    g33478(.A1(new_n36783_), .A2(new_n36784_), .Z(new_n36785_));
  NAND2_X1   g33479(.A1(new_n3810_), .A2(pi0555), .ZN(new_n36787_));
  NAND2_X1   g33480(.A1(new_n35996_), .A2(pi0249), .ZN(new_n36788_));
  NAND2_X1   g33481(.A1(new_n4064_), .A2(pi0553), .ZN(new_n36789_));
  NAND2_X1   g33482(.A1(new_n35990_), .A2(pi0241), .ZN(new_n36790_));
  AOI22_X1   g33483(.A1(new_n36787_), .A2(new_n36788_), .B1(new_n36789_), .B2(new_n36790_), .ZN(new_n36791_));
  NAND2_X1   g33484(.A1(new_n35993_), .A2(pi0248), .ZN(new_n36792_));
  NAND2_X1   g33485(.A1(new_n4225_), .A2(pi0554), .ZN(new_n36793_));
  NAND2_X1   g33486(.A1(new_n4549_), .A2(pi0563), .ZN(new_n36794_));
  NAND2_X1   g33487(.A1(new_n36017_), .A2(pi0246), .ZN(new_n36795_));
  AOI22_X1   g33488(.A1(new_n36792_), .A2(new_n36793_), .B1(new_n36794_), .B2(new_n36795_), .ZN(new_n36796_));
  XOR2_X1    g33489(.A1(new_n36791_), .A2(new_n36796_), .Z(new_n36797_));
  NAND3_X1   g33490(.A1(new_n36797_), .A2(pi0240), .A3(pi0551), .ZN(new_n36798_));
  XOR2_X1    g33491(.A1(new_n36147_), .A2(new_n36798_), .Z(new_n36799_));
  NAND3_X1   g33492(.A1(new_n36799_), .A2(pi0234), .A3(pi0485), .ZN(new_n36800_));
  XNOR2_X1   g33493(.A1(pi0239), .A2(pi0550), .ZN(new_n36801_));
  NOR2_X1    g33494(.A1(new_n36800_), .A2(new_n36801_), .ZN(new_n36802_));
  INV_X1     g33495(.I(new_n36802_), .ZN(new_n36803_));
  NOR2_X1    g33496(.A1(new_n36780_), .A2(pi0569), .ZN(new_n36805_));
  OAI21_X1   g33497(.A1(new_n36800_), .A2(pi0550), .B(pi0239), .ZN(new_n36806_));
  NOR2_X1    g33498(.A1(new_n36805_), .A2(new_n36806_), .ZN(new_n36807_));
  NAND3_X1   g33499(.A1(new_n36803_), .A2(new_n5364_), .A3(new_n35999_), .ZN(new_n36808_));
  NAND4_X1   g33500(.A1(new_n36785_), .A2(pi0489), .A3(new_n36807_), .A4(new_n36808_), .ZN(new_n36809_));
  NAND2_X1   g33501(.A1(new_n36782_), .A2(pi0489), .ZN(new_n36810_));
  XOR2_X1    g33502(.A1(new_n36810_), .A2(new_n36784_), .Z(new_n36811_));
  NAND3_X1   g33503(.A1(new_n36803_), .A2(new_n5364_), .A3(new_n35819_), .ZN(new_n36812_));
  NAND4_X1   g33504(.A1(new_n36811_), .A2(pi0556), .A3(new_n36807_), .A4(new_n36812_), .ZN(new_n36813_));
  NAND2_X1   g33505(.A1(new_n36809_), .A2(new_n36813_), .ZN(new_n36814_));
  XOR2_X1    g33506(.A1(pi0242), .A2(pi0556), .Z(new_n36815_));
  NOR2_X1    g33507(.A1(new_n36782_), .A2(new_n36815_), .ZN(new_n36816_));
  NAND4_X1   g33508(.A1(new_n36814_), .A2(pi0235), .A3(pi0549), .A4(new_n36816_), .ZN(new_n36817_));
  NAND2_X1   g33509(.A1(new_n36817_), .A2(new_n35979_), .ZN(new_n36818_));
  XOR2_X1    g33510(.A1(pi0242), .A2(pi0489), .Z(new_n36819_));
  NOR2_X1    g33511(.A1(new_n36803_), .A2(new_n36819_), .ZN(new_n36820_));
  INV_X1     g33512(.I(new_n36820_), .ZN(new_n36821_));
  NOR2_X1    g33513(.A1(new_n36821_), .A2(pi0531), .ZN(new_n36822_));
  NAND2_X1   g33514(.A1(new_n36816_), .A2(pi0235), .ZN(new_n36823_));
  NOR2_X1    g33515(.A1(new_n3611_), .A2(new_n35979_), .ZN(new_n36824_));
  NOR2_X1    g33516(.A1(new_n36814_), .A2(new_n3611_), .ZN(new_n36825_));
  XNOR2_X1   g33517(.A1(new_n36825_), .A2(new_n36824_), .ZN(new_n36826_));
  OAI21_X1   g33518(.A1(new_n36826_), .A2(new_n36823_), .B(new_n36821_), .ZN(new_n36827_));
  NOR2_X1    g33519(.A1(new_n35936_), .A2(new_n35979_), .ZN(new_n36828_));
  AOI22_X1   g33520(.A1(new_n36827_), .A2(new_n36828_), .B1(new_n36818_), .B2(new_n36822_), .ZN(new_n36829_));
  XNOR2_X1   g33521(.A1(pi0235), .A2(pi0531), .ZN(new_n36830_));
  NAND2_X1   g33522(.A1(new_n36816_), .A2(new_n36830_), .ZN(new_n36831_));
  NOR4_X1    g33523(.A1(new_n36829_), .A2(new_n35828_), .A3(new_n35811_), .A4(new_n36831_), .ZN(new_n36832_));
  NOR2_X1    g33524(.A1(pi0235), .A2(pi0549), .ZN(new_n36833_));
  OAI21_X1   g33525(.A1(new_n36824_), .A2(new_n36833_), .B(new_n36820_), .ZN(new_n36834_));
  NOR2_X1    g33526(.A1(new_n36834_), .A2(pi0566), .ZN(new_n36835_));
  OAI21_X1   g33527(.A1(new_n36832_), .A2(pi0486), .B(new_n36835_), .ZN(new_n36836_));
  NAND3_X1   g33528(.A1(new_n36816_), .A2(pi0244), .A3(new_n36830_), .ZN(new_n36837_));
  NAND2_X1   g33529(.A1(pi0244), .A2(pi0486), .ZN(new_n36838_));
  NAND2_X1   g33530(.A1(new_n36829_), .A2(pi0244), .ZN(new_n36839_));
  XNOR2_X1   g33531(.A1(new_n36839_), .A2(new_n36838_), .ZN(new_n36840_));
  OAI21_X1   g33532(.A1(new_n36840_), .A2(new_n36837_), .B(new_n36834_), .ZN(new_n36841_));
  NAND3_X1   g33533(.A1(new_n36841_), .A2(pi0486), .A3(pi0566), .ZN(new_n36842_));
  NAND2_X1   g33534(.A1(new_n36842_), .A2(new_n36836_), .ZN(new_n36843_));
  INV_X1     g33535(.I(new_n36843_), .ZN(new_n36844_));
  XOR2_X1    g33536(.A1(pi0244), .A2(pi0486), .Z(new_n36845_));
  NOR2_X1    g33537(.A1(new_n36834_), .A2(new_n36845_), .ZN(new_n36846_));
  INV_X1     g33538(.I(new_n36846_), .ZN(new_n36847_));
  NOR4_X1    g33539(.A1(new_n36844_), .A2(new_n4955_), .A3(new_n36097_), .A4(new_n36847_), .ZN(new_n36848_));
  XOR2_X1    g33540(.A1(pi0244), .A2(pi0566), .Z(new_n36849_));
  NOR2_X1    g33541(.A1(new_n36831_), .A2(new_n36849_), .ZN(new_n36850_));
  INV_X1     g33542(.I(new_n36850_), .ZN(new_n36851_));
  NOR2_X1    g33543(.A1(new_n36851_), .A2(pi0580), .ZN(new_n36852_));
  OAI21_X1   g33544(.A1(new_n36848_), .A2(pi0568), .B(new_n36852_), .ZN(new_n36853_));
  NAND2_X1   g33545(.A1(new_n36846_), .A2(pi0245), .ZN(new_n36854_));
  NOR2_X1    g33546(.A1(new_n4955_), .A2(new_n36097_), .ZN(new_n36855_));
  NOR2_X1    g33547(.A1(new_n36843_), .A2(new_n4955_), .ZN(new_n36856_));
  XNOR2_X1   g33548(.A1(new_n36856_), .A2(new_n36855_), .ZN(new_n36857_));
  OAI21_X1   g33549(.A1(new_n36857_), .A2(new_n36854_), .B(new_n36851_), .ZN(new_n36858_));
  NAND3_X1   g33550(.A1(new_n36858_), .A2(pi0568), .A3(pi0580), .ZN(new_n36859_));
  NAND2_X1   g33551(.A1(new_n36859_), .A2(new_n36853_), .ZN(new_n36860_));
  INV_X1     g33552(.I(new_n36860_), .ZN(new_n36861_));
  NOR2_X1    g33553(.A1(pi0245), .A2(pi0568), .ZN(new_n36862_));
  OAI21_X1   g33554(.A1(new_n36855_), .A2(new_n36862_), .B(new_n36850_), .ZN(new_n36863_));
  NOR4_X1    g33555(.A1(new_n36861_), .A2(new_n4459_), .A3(new_n35987_), .A4(new_n36863_), .ZN(new_n36864_));
  NOR2_X1    g33556(.A1(new_n36864_), .A2(pi0552), .ZN(new_n36865_));
  XOR2_X1    g33557(.A1(pi0245), .A2(pi0580), .Z(new_n36866_));
  NOR2_X1    g33558(.A1(new_n36847_), .A2(new_n36866_), .ZN(new_n36867_));
  NAND2_X1   g33559(.A1(new_n36867_), .A2(new_n35939_), .ZN(new_n36868_));
  NOR2_X1    g33560(.A1(new_n36863_), .A2(new_n4459_), .ZN(new_n36869_));
  NAND2_X1   g33561(.A1(pi0247), .A2(pi0552), .ZN(new_n36870_));
  NOR2_X1    g33562(.A1(new_n36860_), .A2(new_n4459_), .ZN(new_n36871_));
  XNOR2_X1   g33563(.A1(new_n36871_), .A2(new_n36870_), .ZN(new_n36872_));
  AOI21_X1   g33564(.A1(new_n36872_), .A2(new_n36869_), .B(new_n36867_), .ZN(new_n36873_));
  NAND2_X1   g33565(.A1(pi0532), .A2(pi0552), .ZN(new_n36874_));
  OAI22_X1   g33566(.A1(new_n36873_), .A2(new_n36874_), .B1(new_n36865_), .B2(new_n36868_), .ZN(new_n36875_));
  NAND2_X1   g33567(.A1(new_n36875_), .A2(pi0238), .ZN(new_n36876_));
  INV_X1     g33568(.I(new_n36867_), .ZN(new_n36877_));
  NAND2_X1   g33569(.A1(new_n4459_), .A2(new_n35987_), .ZN(new_n36878_));
  AOI21_X1   g33570(.A1(new_n36870_), .A2(new_n36878_), .B(new_n36877_), .ZN(new_n36879_));
  XOR2_X1    g33571(.A1(pi0247), .A2(pi0532), .Z(new_n36880_));
  NOR2_X1    g33572(.A1(new_n36863_), .A2(new_n36880_), .ZN(new_n36881_));
  NOR2_X1    g33573(.A1(new_n36881_), .A2(new_n3743_), .ZN(new_n36882_));
  NAND2_X1   g33574(.A1(pi0238), .A2(pi0577), .ZN(new_n36883_));
  XNOR2_X1   g33575(.A1(new_n36882_), .A2(new_n36883_), .ZN(new_n36884_));
  NAND2_X1   g33576(.A1(new_n36884_), .A2(new_n36879_), .ZN(new_n36885_));
  NAND2_X1   g33577(.A1(new_n36885_), .A2(pi0498), .ZN(new_n36886_));
  AOI21_X1   g33578(.A1(new_n36876_), .A2(pi0577), .B(new_n36886_), .ZN(new_n36887_));
  NOR2_X1    g33579(.A1(new_n36881_), .A2(new_n36116_), .ZN(new_n36888_));
  XNOR2_X1   g33580(.A1(new_n36888_), .A2(new_n36883_), .ZN(new_n36889_));
  NAND2_X1   g33581(.A1(new_n36889_), .A2(new_n36879_), .ZN(new_n36890_));
  NAND2_X1   g33582(.A1(new_n36890_), .A2(new_n35843_), .ZN(new_n36891_));
  AOI21_X1   g33583(.A1(new_n36875_), .A2(new_n3743_), .B(pi0577), .ZN(new_n36892_));
  OAI21_X1   g33584(.A1(new_n36887_), .A2(new_n36891_), .B(new_n36892_), .ZN(new_n36893_));
  AOI21_X1   g33585(.A1(new_n36765_), .A2(new_n36755_), .B(new_n36893_), .ZN(new_n36894_));
  AOI21_X1   g33586(.A1(new_n36428_), .A2(new_n36582_), .B(new_n36894_), .ZN(po0750));
  NOR2_X1    g33587(.A1(new_n2955_), .A2(new_n35624_), .ZN(po0751));
  INV_X1     g33588(.I(pi0806), .ZN(new_n36897_));
  NAND3_X1   g33589(.A1(new_n35628_), .A2(pi0605), .A3(new_n36897_), .ZN(new_n36898_));
  XOR2_X1    g33590(.A1(new_n36898_), .A2(pi0595), .Z(new_n36899_));
  NOR2_X1    g33591(.A1(new_n36899_), .A2(pi0332), .ZN(po0752));
  NOR2_X1    g33592(.A1(new_n2955_), .A2(new_n35626_), .ZN(new_n36901_));
  NOR3_X1    g33593(.A1(new_n35624_), .A2(new_n36897_), .A3(new_n35639_), .ZN(new_n36902_));
  NOR2_X1    g33594(.A1(new_n35632_), .A2(new_n35625_), .ZN(new_n36903_));
  NAND3_X1   g33595(.A1(new_n36902_), .A2(new_n36901_), .A3(new_n36903_), .ZN(new_n36904_));
  NAND2_X1   g33596(.A1(new_n2955_), .A2(pi0596), .ZN(new_n36905_));
  OAI21_X1   g33597(.A1(new_n36904_), .A2(pi0596), .B(new_n36905_), .ZN(po0753));
  NAND2_X1   g33598(.A1(new_n35640_), .A2(new_n36897_), .ZN(new_n36907_));
  XOR2_X1    g33599(.A1(new_n36907_), .A2(pi0597), .Z(new_n36908_));
  NOR2_X1    g33600(.A1(new_n36908_), .A2(pi0332), .ZN(po0754));
  INV_X1     g33601(.I(pi0598), .ZN(new_n36910_));
  NOR2_X1    g33602(.A1(pi0882), .A2(pi0947), .ZN(new_n36911_));
  NAND2_X1   g33603(.A1(new_n36911_), .A2(new_n36910_), .ZN(new_n36912_));
  NAND2_X1   g33604(.A1(po1038), .A2(new_n36912_), .ZN(new_n36913_));
  NOR2_X1    g33605(.A1(pi0740), .A2(pi0780), .ZN(new_n36914_));
  AOI21_X1   g33606(.A1(new_n36913_), .A2(new_n36914_), .B(new_n5796_), .ZN(po0755));
  NAND2_X1   g33607(.A1(pi0332), .A2(pi0596), .ZN(new_n36916_));
  AOI21_X1   g33608(.A1(new_n36904_), .A2(new_n36916_), .B(pi0599), .ZN(new_n36917_));
  XNOR2_X1   g33609(.A1(new_n36917_), .A2(new_n36916_), .ZN(po0756));
  NAND2_X1   g33610(.A1(new_n36901_), .A2(new_n35639_), .ZN(new_n36919_));
  OAI21_X1   g33611(.A1(new_n2955_), .A2(new_n35626_), .B(pi0990), .ZN(new_n36920_));
  AOI21_X1   g33612(.A1(new_n36919_), .A2(new_n36920_), .B(new_n36897_), .ZN(po0757));
  INV_X1     g33613(.I(pi0989), .ZN(new_n36922_));
  NAND3_X1   g33614(.A1(pi0332), .A2(pi0601), .A3(pi0806), .ZN(new_n36923_));
  NAND3_X1   g33615(.A1(new_n2955_), .A2(new_n35627_), .A3(pi0806), .ZN(new_n36924_));
  AOI21_X1   g33616(.A1(new_n36924_), .A2(new_n36923_), .B(new_n36922_), .ZN(po0758));
  NAND4_X1   g33617(.A1(new_n14058_), .A2(pi0230), .A3(pi0602), .A4(new_n13206_), .ZN(new_n36926_));
  NOR2_X1    g33618(.A1(new_n14200_), .A2(pi1160), .ZN(new_n36927_));
  OAI21_X1   g33619(.A1(new_n14254_), .A2(new_n36927_), .B(pi0790), .ZN(new_n36928_));
  NAND3_X1   g33620(.A1(new_n15402_), .A2(new_n36029_), .A3(new_n36928_), .ZN(new_n36929_));
  OAI22_X1   g33621(.A1(new_n15396_), .A2(new_n30557_), .B1(new_n36926_), .B2(new_n36929_), .ZN(po0759));
  INV_X1     g33622(.I(pi0871), .ZN(new_n36931_));
  INV_X1     g33623(.I(pi0872), .ZN(new_n36932_));
  INV_X1     g33624(.I(pi0952), .ZN(new_n36933_));
  INV_X1     g33625(.I(pi0980), .ZN(new_n36934_));
  NAND3_X1   g33626(.A1(new_n36934_), .A2(pi1038), .A3(pi1060), .ZN(new_n36935_));
  NOR3_X1    g33627(.A1(new_n36935_), .A2(new_n36933_), .A3(pi1061), .ZN(new_n36936_));
  NOR2_X1    g33628(.A1(new_n14799_), .A2(pi1100), .ZN(new_n36937_));
  NAND4_X1   g33629(.A1(new_n36936_), .A2(pi0603), .A3(pi0832), .A4(pi0966), .ZN(new_n36938_));
  AOI21_X1   g33630(.A1(new_n36938_), .A2(new_n36932_), .B(new_n36931_), .ZN(po0760));
  INV_X1     g33631(.I(pi0779), .ZN(new_n36940_));
  NAND3_X1   g33632(.A1(new_n12844_), .A2(new_n36940_), .A3(pi0823), .ZN(new_n36941_));
  INV_X1     g33633(.I(pi0604), .ZN(new_n36942_));
  INV_X1     g33634(.I(pi0983), .ZN(new_n36943_));
  NAND3_X1   g33635(.A1(new_n36942_), .A2(new_n5741_), .A3(new_n36943_), .ZN(new_n36944_));
  NAND4_X1   g33636(.A1(new_n12844_), .A2(pi0299), .A3(pi0823), .A4(new_n36944_), .ZN(new_n36945_));
  XOR2_X1    g33637(.A1(new_n36945_), .A2(new_n36941_), .Z(po0761));
  OR2_X2     g33638(.A1(pi0605), .A2(pi0806), .Z(new_n36947_));
  NAND2_X1   g33639(.A1(pi0605), .A2(pi0806), .ZN(new_n36948_));
  AOI21_X1   g33640(.A1(new_n36947_), .A2(new_n36948_), .B(pi0332), .ZN(po0762));
  NAND2_X1   g33641(.A1(new_n36936_), .A2(pi0832), .ZN(new_n36950_));
  INV_X1     g33642(.I(pi1104), .ZN(new_n36951_));
  NOR2_X1    g33643(.A1(new_n36950_), .A2(new_n36951_), .ZN(new_n36952_));
  AOI21_X1   g33644(.A1(pi0606), .A2(new_n36950_), .B(new_n36952_), .ZN(new_n36953_));
  NAND2_X1   g33645(.A1(pi0837), .A2(pi0966), .ZN(new_n36954_));
  OAI21_X1   g33646(.A1(new_n36953_), .A2(pi0966), .B(new_n36954_), .ZN(po0763));
  INV_X1     g33647(.I(new_n36950_), .ZN(po0897));
  NAND3_X1   g33648(.A1(po0897), .A2(pi0966), .A3(pi1107), .ZN(new_n36957_));
  INV_X1     g33649(.I(pi0966), .ZN(new_n36958_));
  INV_X1     g33650(.I(pi1107), .ZN(new_n36959_));
  NAND3_X1   g33651(.A1(po0897), .A2(new_n36958_), .A3(new_n36959_), .ZN(new_n36960_));
  AOI21_X1   g33652(.A1(new_n36957_), .A2(new_n36960_), .B(new_n28263_), .ZN(po0764));
  NAND3_X1   g33653(.A1(po0897), .A2(pi0966), .A3(pi1116), .ZN(new_n36962_));
  INV_X1     g33654(.I(pi1116), .ZN(new_n36963_));
  NAND3_X1   g33655(.A1(po0897), .A2(new_n36958_), .A3(new_n36963_), .ZN(new_n36964_));
  AOI21_X1   g33656(.A1(new_n36962_), .A2(new_n36964_), .B(new_n14081_), .ZN(po0765));
  NAND3_X1   g33657(.A1(po0897), .A2(pi0966), .A3(pi1118), .ZN(new_n36966_));
  INV_X1     g33658(.I(pi1118), .ZN(new_n36967_));
  NAND3_X1   g33659(.A1(po0897), .A2(new_n36958_), .A3(new_n36967_), .ZN(new_n36968_));
  AOI21_X1   g33660(.A1(new_n36966_), .A2(new_n36968_), .B(new_n13766_), .ZN(po0766));
  INV_X1     g33661(.I(pi0610), .ZN(new_n36970_));
  NAND3_X1   g33662(.A1(po0897), .A2(pi0966), .A3(pi1113), .ZN(new_n36971_));
  INV_X1     g33663(.I(pi1113), .ZN(new_n36972_));
  NAND3_X1   g33664(.A1(po0897), .A2(new_n36958_), .A3(new_n36972_), .ZN(new_n36973_));
  AOI21_X1   g33665(.A1(new_n36971_), .A2(new_n36973_), .B(new_n36970_), .ZN(po0767));
  INV_X1     g33666(.I(pi0611), .ZN(new_n36975_));
  NAND3_X1   g33667(.A1(po0897), .A2(pi0966), .A3(pi1114), .ZN(new_n36976_));
  INV_X1     g33668(.I(pi1114), .ZN(new_n36977_));
  NAND3_X1   g33669(.A1(po0897), .A2(new_n36958_), .A3(new_n36977_), .ZN(new_n36978_));
  AOI21_X1   g33670(.A1(new_n36976_), .A2(new_n36978_), .B(new_n36975_), .ZN(po0768));
  NAND3_X1   g33671(.A1(po0897), .A2(pi0966), .A3(pi1111), .ZN(new_n36980_));
  INV_X1     g33672(.I(pi1111), .ZN(new_n36981_));
  NAND3_X1   g33673(.A1(po0897), .A2(new_n36958_), .A3(new_n36981_), .ZN(new_n36982_));
  AOI21_X1   g33674(.A1(new_n36980_), .A2(new_n36982_), .B(new_n28683_), .ZN(po0769));
  INV_X1     g33675(.I(pi0613), .ZN(new_n36984_));
  NAND3_X1   g33676(.A1(po0897), .A2(pi0966), .A3(pi1115), .ZN(new_n36985_));
  INV_X1     g33677(.I(pi1115), .ZN(new_n36986_));
  NAND3_X1   g33678(.A1(po0897), .A2(new_n36958_), .A3(new_n36986_), .ZN(new_n36987_));
  AOI21_X1   g33679(.A1(new_n36985_), .A2(new_n36987_), .B(new_n36984_), .ZN(po0770));
  NOR2_X1    g33680(.A1(new_n36950_), .A2(new_n36958_), .ZN(new_n36989_));
  NOR2_X1    g33681(.A1(new_n36950_), .A2(pi1102), .ZN(new_n36990_));
  XNOR2_X1   g33682(.A1(new_n36989_), .A2(new_n36990_), .ZN(new_n36991_));
  OAI22_X1   g33683(.A1(new_n36991_), .A2(new_n12868_), .B1(new_n36931_), .B2(new_n36958_), .ZN(po0771));
  INV_X1     g33684(.I(pi0615), .ZN(new_n36993_));
  NOR2_X1    g33685(.A1(pi0882), .A2(pi0907), .ZN(new_n36994_));
  NAND2_X1   g33686(.A1(new_n36994_), .A2(new_n36993_), .ZN(new_n36995_));
  NAND2_X1   g33687(.A1(po1038), .A2(new_n36995_), .ZN(new_n36996_));
  NOR2_X1    g33688(.A1(pi0779), .A2(pi0797), .ZN(new_n36997_));
  AOI21_X1   g33689(.A1(new_n36996_), .A2(new_n36997_), .B(new_n5636_), .ZN(po0772));
  NOR2_X1    g33690(.A1(new_n36950_), .A2(pi1101), .ZN(new_n36999_));
  XNOR2_X1   g33691(.A1(new_n36989_), .A2(new_n36999_), .ZN(new_n37000_));
  OAI22_X1   g33692(.A1(new_n37000_), .A2(new_n12841_), .B1(new_n36932_), .B2(new_n36958_), .ZN(po0773));
  INV_X1     g33693(.I(pi1105), .ZN(new_n37002_));
  NOR2_X1    g33694(.A1(new_n36950_), .A2(new_n37002_), .ZN(new_n37003_));
  AOI21_X1   g33695(.A1(pi0617), .A2(new_n36950_), .B(new_n37003_), .ZN(new_n37004_));
  NAND2_X1   g33696(.A1(pi0850), .A2(pi0966), .ZN(new_n37005_));
  OAI21_X1   g33697(.A1(new_n37004_), .A2(pi0966), .B(new_n37005_), .ZN(po0774));
  NAND3_X1   g33698(.A1(po0897), .A2(pi0966), .A3(pi1117), .ZN(new_n37007_));
  INV_X1     g33699(.I(pi1117), .ZN(new_n37008_));
  NAND3_X1   g33700(.A1(po0897), .A2(new_n36958_), .A3(new_n37008_), .ZN(new_n37009_));
  AOI21_X1   g33701(.A1(new_n37007_), .A2(new_n37009_), .B(new_n13816_), .ZN(po0775));
  NAND3_X1   g33702(.A1(po0897), .A2(pi0966), .A3(pi1122), .ZN(new_n37011_));
  INV_X1     g33703(.I(pi1122), .ZN(new_n37012_));
  NAND3_X1   g33704(.A1(po0897), .A2(new_n36958_), .A3(new_n37012_), .ZN(new_n37013_));
  AOI21_X1   g33705(.A1(new_n37011_), .A2(new_n37013_), .B(new_n13860_), .ZN(po0776));
  INV_X1     g33706(.I(pi0620), .ZN(new_n37015_));
  NAND3_X1   g33707(.A1(po0897), .A2(pi0966), .A3(pi1112), .ZN(new_n37016_));
  INV_X1     g33708(.I(pi1112), .ZN(new_n37017_));
  NAND3_X1   g33709(.A1(po0897), .A2(new_n36958_), .A3(new_n37017_), .ZN(new_n37018_));
  AOI21_X1   g33710(.A1(new_n37016_), .A2(new_n37018_), .B(new_n37015_), .ZN(po0777));
  NAND3_X1   g33711(.A1(po0897), .A2(pi0966), .A3(pi1108), .ZN(new_n37020_));
  INV_X1     g33712(.I(pi1108), .ZN(new_n37021_));
  NAND3_X1   g33713(.A1(po0897), .A2(new_n36958_), .A3(new_n37021_), .ZN(new_n37022_));
  AOI21_X1   g33714(.A1(new_n37020_), .A2(new_n37022_), .B(new_n13142_), .ZN(po0778));
  NAND3_X1   g33715(.A1(po0897), .A2(pi0966), .A3(pi1109), .ZN(new_n37024_));
  INV_X1     g33716(.I(pi1109), .ZN(new_n37025_));
  NAND3_X1   g33717(.A1(po0897), .A2(new_n36958_), .A3(new_n37025_), .ZN(new_n37026_));
  AOI21_X1   g33718(.A1(new_n37024_), .A2(new_n37026_), .B(new_n28296_), .ZN(po0779));
  NAND3_X1   g33719(.A1(po0897), .A2(pi0966), .A3(pi1106), .ZN(new_n37028_));
  INV_X1     g33720(.I(pi1106), .ZN(new_n37029_));
  NAND3_X1   g33721(.A1(po0897), .A2(new_n36958_), .A3(new_n37029_), .ZN(new_n37030_));
  AOI21_X1   g33722(.A1(new_n37028_), .A2(new_n37030_), .B(new_n28200_), .ZN(po0780));
  INV_X1     g33723(.I(pi0780), .ZN(new_n37032_));
  NAND3_X1   g33724(.A1(new_n13336_), .A2(new_n37032_), .A3(pi0831), .ZN(new_n37033_));
  INV_X1     g33725(.I(pi0624), .ZN(new_n37034_));
  NAND3_X1   g33726(.A1(new_n37034_), .A2(new_n5800_), .A3(new_n36943_), .ZN(new_n37035_));
  NAND4_X1   g33727(.A1(new_n13336_), .A2(pi0299), .A3(pi0831), .A4(new_n37035_), .ZN(new_n37036_));
  XOR2_X1    g33728(.A1(new_n37036_), .A2(new_n37033_), .Z(po0781));
  INV_X1     g33729(.I(pi0953), .ZN(new_n37038_));
  INV_X1     g33730(.I(pi1054), .ZN(new_n37039_));
  NAND3_X1   g33731(.A1(new_n37039_), .A2(pi1066), .A3(pi1088), .ZN(new_n37040_));
  NOR3_X1    g33732(.A1(new_n37040_), .A2(new_n14799_), .A3(pi0973), .ZN(new_n37041_));
  NAND2_X1   g33733(.A1(new_n37041_), .A2(new_n37038_), .ZN(new_n37042_));
  INV_X1     g33734(.I(new_n37042_), .ZN(po0954));
  NAND3_X1   g33735(.A1(po0954), .A2(pi0962), .A3(pi1116), .ZN(new_n37044_));
  INV_X1     g33736(.I(pi0962), .ZN(new_n37045_));
  NAND3_X1   g33737(.A1(po0954), .A2(new_n37045_), .A3(new_n36963_), .ZN(new_n37046_));
  AOI21_X1   g33738(.A1(new_n37044_), .A2(new_n37046_), .B(new_n13613_), .ZN(po0782));
  NAND3_X1   g33739(.A1(po0897), .A2(pi0966), .A3(pi1121), .ZN(new_n37048_));
  INV_X1     g33740(.I(pi1121), .ZN(new_n37049_));
  NAND3_X1   g33741(.A1(po0897), .A2(new_n36958_), .A3(new_n37049_), .ZN(new_n37050_));
  AOI21_X1   g33742(.A1(new_n37048_), .A2(new_n37050_), .B(new_n13901_), .ZN(po0783));
  NAND3_X1   g33743(.A1(po0954), .A2(pi0962), .A3(pi1117), .ZN(new_n37052_));
  NAND3_X1   g33744(.A1(po0954), .A2(new_n37045_), .A3(new_n37008_), .ZN(new_n37053_));
  AOI21_X1   g33745(.A1(new_n37052_), .A2(new_n37053_), .B(new_n13823_), .ZN(po0784));
  NAND3_X1   g33746(.A1(po0954), .A2(pi0962), .A3(pi1119), .ZN(new_n37055_));
  INV_X1     g33747(.I(pi1119), .ZN(new_n37056_));
  NAND3_X1   g33748(.A1(po0954), .A2(new_n37045_), .A3(new_n37056_), .ZN(new_n37057_));
  AOI21_X1   g33749(.A1(new_n37055_), .A2(new_n37057_), .B(new_n13942_), .ZN(po0785));
  NAND3_X1   g33750(.A1(po0897), .A2(pi0966), .A3(pi1119), .ZN(new_n37059_));
  NAND3_X1   g33751(.A1(po0897), .A2(new_n36958_), .A3(new_n37056_), .ZN(new_n37060_));
  AOI21_X1   g33752(.A1(new_n37059_), .A2(new_n37060_), .B(new_n13976_), .ZN(po0786));
  NAND3_X1   g33753(.A1(po0897), .A2(pi0966), .A3(pi1120), .ZN(new_n37062_));
  INV_X1     g33754(.I(pi1120), .ZN(new_n37063_));
  NAND3_X1   g33755(.A1(po0897), .A2(new_n36958_), .A3(new_n37063_), .ZN(new_n37064_));
  AOI21_X1   g33756(.A1(new_n37062_), .A2(new_n37064_), .B(new_n14010_), .ZN(po0787));
  INV_X1     g33757(.I(pi0631), .ZN(new_n37066_));
  NAND3_X1   g33758(.A1(po0954), .A2(pi0962), .A3(pi1113), .ZN(new_n37067_));
  NAND3_X1   g33759(.A1(po0954), .A2(new_n37045_), .A3(new_n36972_), .ZN(new_n37068_));
  AOI21_X1   g33760(.A1(new_n37067_), .A2(new_n37068_), .B(new_n37066_), .ZN(po0788));
  INV_X1     g33761(.I(pi0632), .ZN(new_n37070_));
  NAND3_X1   g33762(.A1(po0954), .A2(pi0962), .A3(pi1115), .ZN(new_n37071_));
  NAND3_X1   g33763(.A1(po0954), .A2(new_n37045_), .A3(new_n36986_), .ZN(new_n37072_));
  AOI21_X1   g33764(.A1(new_n37071_), .A2(new_n37072_), .B(new_n37070_), .ZN(po0789));
  NAND3_X1   g33765(.A1(po0897), .A2(pi0966), .A3(pi1110), .ZN(new_n37074_));
  INV_X1     g33766(.I(pi1110), .ZN(new_n37075_));
  NAND3_X1   g33767(.A1(po0897), .A2(new_n36958_), .A3(new_n37075_), .ZN(new_n37076_));
  AOI21_X1   g33768(.A1(new_n37074_), .A2(new_n37076_), .B(new_n26463_), .ZN(po0790));
  NAND3_X1   g33769(.A1(po0954), .A2(pi0962), .A3(pi1110), .ZN(new_n37078_));
  NAND3_X1   g33770(.A1(po0954), .A2(new_n37045_), .A3(new_n37075_), .ZN(new_n37079_));
  AOI21_X1   g33771(.A1(new_n37078_), .A2(new_n37079_), .B(new_n26624_), .ZN(po0791));
  INV_X1     g33772(.I(pi0635), .ZN(new_n37081_));
  NAND3_X1   g33773(.A1(po0954), .A2(pi0962), .A3(pi1112), .ZN(new_n37082_));
  NAND3_X1   g33774(.A1(po0954), .A2(new_n37045_), .A3(new_n37017_), .ZN(new_n37083_));
  AOI21_X1   g33775(.A1(new_n37082_), .A2(new_n37083_), .B(new_n37081_), .ZN(po0792));
  INV_X1     g33776(.I(pi0636), .ZN(new_n37085_));
  NAND3_X1   g33777(.A1(po0897), .A2(pi0966), .A3(pi1127), .ZN(new_n37086_));
  INV_X1     g33778(.I(pi1127), .ZN(new_n37087_));
  NAND3_X1   g33779(.A1(po0897), .A2(new_n36958_), .A3(new_n37087_), .ZN(new_n37088_));
  AOI21_X1   g33780(.A1(new_n37086_), .A2(new_n37088_), .B(new_n37085_), .ZN(po0793));
  NAND3_X1   g33781(.A1(po0954), .A2(pi0962), .A3(pi1105), .ZN(new_n37090_));
  NAND3_X1   g33782(.A1(po0954), .A2(new_n37045_), .A3(new_n37002_), .ZN(new_n37091_));
  AOI21_X1   g33783(.A1(new_n37090_), .A2(new_n37091_), .B(new_n26983_), .ZN(po0794));
  NAND3_X1   g33784(.A1(po0954), .A2(pi0962), .A3(pi1107), .ZN(new_n37093_));
  NAND3_X1   g33785(.A1(po0954), .A2(new_n37045_), .A3(new_n36959_), .ZN(new_n37094_));
  AOI21_X1   g33786(.A1(new_n37093_), .A2(new_n37094_), .B(new_n28243_), .ZN(po0795));
  NAND3_X1   g33787(.A1(po0954), .A2(pi0962), .A3(pi1109), .ZN(new_n37096_));
  NAND3_X1   g33788(.A1(po0954), .A2(new_n37045_), .A3(new_n37025_), .ZN(new_n37097_));
  AOI21_X1   g33789(.A1(new_n37096_), .A2(new_n37097_), .B(new_n28297_), .ZN(po0796));
  INV_X1     g33790(.I(pi0640), .ZN(new_n37099_));
  NAND3_X1   g33791(.A1(po0897), .A2(pi0966), .A3(pi1128), .ZN(new_n37100_));
  INV_X1     g33792(.I(pi1128), .ZN(new_n37101_));
  NAND3_X1   g33793(.A1(po0897), .A2(new_n36958_), .A3(new_n37101_), .ZN(new_n37102_));
  AOI21_X1   g33794(.A1(new_n37100_), .A2(new_n37102_), .B(new_n37099_), .ZN(po0797));
  NAND3_X1   g33795(.A1(po0954), .A2(pi0962), .A3(pi1121), .ZN(new_n37104_));
  NAND3_X1   g33796(.A1(po0954), .A2(new_n37045_), .A3(new_n37049_), .ZN(new_n37105_));
  AOI21_X1   g33797(.A1(new_n37104_), .A2(new_n37105_), .B(new_n13922_), .ZN(po0798));
  NAND3_X1   g33798(.A1(po0897), .A2(pi0966), .A3(pi1103), .ZN(new_n37107_));
  INV_X1     g33799(.I(pi1103), .ZN(new_n37108_));
  NAND3_X1   g33800(.A1(po0897), .A2(new_n36958_), .A3(new_n37108_), .ZN(new_n37109_));
  AOI21_X1   g33801(.A1(new_n37107_), .A2(new_n37109_), .B(new_n5379_), .ZN(po0799));
  NAND3_X1   g33802(.A1(po0954), .A2(pi0962), .A3(pi1104), .ZN(new_n37111_));
  NAND3_X1   g33803(.A1(po0954), .A2(new_n37045_), .A3(new_n36951_), .ZN(new_n37112_));
  AOI21_X1   g33804(.A1(new_n37111_), .A2(new_n37112_), .B(new_n27295_), .ZN(po0800));
  NAND3_X1   g33805(.A1(po0897), .A2(pi0966), .A3(pi1123), .ZN(new_n37114_));
  INV_X1     g33806(.I(pi1123), .ZN(new_n37115_));
  NAND3_X1   g33807(.A1(po0897), .A2(new_n36958_), .A3(new_n37115_), .ZN(new_n37116_));
  AOI21_X1   g33808(.A1(new_n37114_), .A2(new_n37116_), .B(new_n14204_), .ZN(po0801));
  INV_X1     g33809(.I(pi0645), .ZN(new_n37118_));
  NAND3_X1   g33810(.A1(po0897), .A2(pi0966), .A3(pi1125), .ZN(new_n37119_));
  INV_X1     g33811(.I(pi1125), .ZN(new_n37120_));
  NAND3_X1   g33812(.A1(po0897), .A2(new_n36958_), .A3(new_n37120_), .ZN(new_n37121_));
  AOI21_X1   g33813(.A1(new_n37119_), .A2(new_n37121_), .B(new_n37118_), .ZN(po0802));
  INV_X1     g33814(.I(pi0646), .ZN(new_n37123_));
  NAND3_X1   g33815(.A1(po0954), .A2(pi0962), .A3(pi1114), .ZN(new_n37124_));
  NAND3_X1   g33816(.A1(po0954), .A2(new_n37045_), .A3(new_n36977_), .ZN(new_n37125_));
  AOI21_X1   g33817(.A1(new_n37124_), .A2(new_n37125_), .B(new_n37123_), .ZN(po0803));
  NAND3_X1   g33818(.A1(po0954), .A2(pi0962), .A3(pi1120), .ZN(new_n37127_));
  NAND3_X1   g33819(.A1(po0954), .A2(new_n37045_), .A3(new_n37063_), .ZN(new_n37128_));
  AOI21_X1   g33820(.A1(new_n37127_), .A2(new_n37128_), .B(new_n14005_), .ZN(po0804));
  NAND3_X1   g33821(.A1(po0954), .A2(pi0962), .A3(pi1122), .ZN(new_n37130_));
  NAND3_X1   g33822(.A1(po0954), .A2(new_n37045_), .A3(new_n37012_), .ZN(new_n37131_));
  AOI21_X1   g33823(.A1(new_n37130_), .A2(new_n37131_), .B(new_n13884_), .ZN(po0805));
  INV_X1     g33824(.I(pi0649), .ZN(new_n37133_));
  NAND3_X1   g33825(.A1(po0954), .A2(pi0962), .A3(pi1126), .ZN(new_n37134_));
  INV_X1     g33826(.I(pi1126), .ZN(new_n37135_));
  NAND3_X1   g33827(.A1(po0954), .A2(new_n37045_), .A3(new_n37135_), .ZN(new_n37136_));
  AOI21_X1   g33828(.A1(new_n37134_), .A2(new_n37136_), .B(new_n37133_), .ZN(po0806));
  INV_X1     g33829(.I(pi0650), .ZN(new_n37138_));
  NAND3_X1   g33830(.A1(po0954), .A2(pi0962), .A3(pi1127), .ZN(new_n37139_));
  NAND3_X1   g33831(.A1(po0954), .A2(new_n37045_), .A3(new_n37087_), .ZN(new_n37140_));
  AOI21_X1   g33832(.A1(new_n37139_), .A2(new_n37140_), .B(new_n37138_), .ZN(po0807));
  INV_X1     g33833(.I(pi0651), .ZN(new_n37142_));
  NAND3_X1   g33834(.A1(po0897), .A2(pi0966), .A3(pi1130), .ZN(new_n37143_));
  INV_X1     g33835(.I(pi1130), .ZN(new_n37144_));
  NAND3_X1   g33836(.A1(po0897), .A2(new_n36958_), .A3(new_n37144_), .ZN(new_n37145_));
  AOI21_X1   g33837(.A1(new_n37143_), .A2(new_n37145_), .B(new_n37142_), .ZN(po0808));
  INV_X1     g33838(.I(pi0652), .ZN(new_n37147_));
  NAND3_X1   g33839(.A1(po0897), .A2(pi0966), .A3(pi1131), .ZN(new_n37148_));
  INV_X1     g33840(.I(pi1131), .ZN(new_n37149_));
  NAND3_X1   g33841(.A1(po0897), .A2(new_n36958_), .A3(new_n37149_), .ZN(new_n37150_));
  AOI21_X1   g33842(.A1(new_n37148_), .A2(new_n37150_), .B(new_n37147_), .ZN(po0809));
  INV_X1     g33843(.I(pi0653), .ZN(new_n37152_));
  NAND3_X1   g33844(.A1(po0897), .A2(pi0966), .A3(pi1129), .ZN(new_n37153_));
  INV_X1     g33845(.I(pi1129), .ZN(new_n37154_));
  NAND3_X1   g33846(.A1(po0897), .A2(new_n36958_), .A3(new_n37154_), .ZN(new_n37155_));
  AOI21_X1   g33847(.A1(new_n37153_), .A2(new_n37155_), .B(new_n37152_), .ZN(po0810));
  INV_X1     g33848(.I(pi0654), .ZN(new_n37157_));
  NAND3_X1   g33849(.A1(po0954), .A2(pi0962), .A3(pi1130), .ZN(new_n37158_));
  NAND3_X1   g33850(.A1(po0954), .A2(new_n37045_), .A3(new_n37144_), .ZN(new_n37159_));
  AOI21_X1   g33851(.A1(new_n37158_), .A2(new_n37159_), .B(new_n37157_), .ZN(po0811));
  INV_X1     g33852(.I(pi0655), .ZN(new_n37161_));
  NAND3_X1   g33853(.A1(po0954), .A2(pi0962), .A3(pi1124), .ZN(new_n37162_));
  INV_X1     g33854(.I(pi1124), .ZN(new_n37163_));
  NAND3_X1   g33855(.A1(po0954), .A2(new_n37045_), .A3(new_n37163_), .ZN(new_n37164_));
  AOI21_X1   g33856(.A1(new_n37162_), .A2(new_n37164_), .B(new_n37161_), .ZN(po0812));
  INV_X1     g33857(.I(pi0656), .ZN(new_n37166_));
  NAND3_X1   g33858(.A1(po0897), .A2(pi0966), .A3(pi1126), .ZN(new_n37167_));
  NAND3_X1   g33859(.A1(po0897), .A2(new_n36958_), .A3(new_n37135_), .ZN(new_n37168_));
  AOI21_X1   g33860(.A1(new_n37167_), .A2(new_n37168_), .B(new_n37166_), .ZN(po0813));
  INV_X1     g33861(.I(pi0657), .ZN(new_n37170_));
  NAND3_X1   g33862(.A1(po0954), .A2(pi0962), .A3(pi1131), .ZN(new_n37171_));
  NAND3_X1   g33863(.A1(po0954), .A2(new_n37045_), .A3(new_n37149_), .ZN(new_n37172_));
  AOI21_X1   g33864(.A1(new_n37171_), .A2(new_n37172_), .B(new_n37170_), .ZN(po0814));
  INV_X1     g33865(.I(pi0658), .ZN(new_n37174_));
  NAND3_X1   g33866(.A1(po0897), .A2(pi0966), .A3(pi1124), .ZN(new_n37175_));
  NAND3_X1   g33867(.A1(po0897), .A2(new_n36958_), .A3(new_n37163_), .ZN(new_n37176_));
  AOI21_X1   g33868(.A1(new_n37175_), .A2(new_n37176_), .B(new_n37174_), .ZN(po0815));
  NOR2_X1    g33869(.A1(new_n4786_), .A2(pi0280), .ZN(new_n37178_));
  NAND2_X1   g33870(.A1(new_n37178_), .A2(pi0992), .ZN(new_n37179_));
  NOR3_X1    g33871(.A1(new_n37179_), .A2(pi0269), .A3(pi0281), .ZN(new_n37180_));
  INV_X1     g33872(.I(new_n37180_), .ZN(new_n37181_));
  OR3_X2     g33873(.A1(pi0270), .A2(pi0277), .A3(pi0282), .Z(new_n37182_));
  NOR2_X1    g33874(.A1(new_n37181_), .A2(new_n37182_), .ZN(new_n37183_));
  INV_X1     g33875(.I(new_n37183_), .ZN(new_n37184_));
  NOR3_X1    g33876(.A1(new_n37184_), .A2(pi0264), .A3(pi0265), .ZN(new_n37185_));
  XOR2_X1    g33877(.A1(new_n37185_), .A2(new_n3505_), .Z(po0816));
  NAND3_X1   g33878(.A1(po0954), .A2(pi0962), .A3(pi1118), .ZN(new_n37187_));
  NAND3_X1   g33879(.A1(po0954), .A2(new_n37045_), .A3(new_n36967_), .ZN(new_n37188_));
  AOI21_X1   g33880(.A1(new_n37187_), .A2(new_n37188_), .B(new_n13783_), .ZN(po0817));
  NAND3_X1   g33881(.A1(po0954), .A2(pi0962), .A3(pi1101), .ZN(new_n37190_));
  INV_X1     g33882(.I(pi1101), .ZN(new_n37191_));
  NAND3_X1   g33883(.A1(po0954), .A2(new_n37045_), .A3(new_n37191_), .ZN(new_n37192_));
  AOI21_X1   g33884(.A1(new_n37190_), .A2(new_n37192_), .B(new_n5374_), .ZN(po0818));
  NAND3_X1   g33885(.A1(po0954), .A2(pi0962), .A3(pi1102), .ZN(new_n37194_));
  INV_X1     g33886(.I(pi1102), .ZN(new_n37195_));
  NAND3_X1   g33887(.A1(po0954), .A2(new_n37045_), .A3(new_n37195_), .ZN(new_n37196_));
  AOI21_X1   g33888(.A1(new_n37194_), .A2(new_n37196_), .B(new_n5633_), .ZN(po0819));
  NAND3_X1   g33889(.A1(pi0334), .A2(pi0591), .A3(pi0592), .ZN(new_n37198_));
  NAND3_X1   g33890(.A1(new_n35424_), .A2(new_n6350_), .A3(pi0592), .ZN(new_n37199_));
  XOR2_X1    g33891(.A1(new_n37199_), .A2(new_n37198_), .Z(new_n37200_));
  NOR2_X1    g33892(.A1(new_n7129_), .A2(pi0592), .ZN(new_n37201_));
  NOR2_X1    g33893(.A1(pi0223), .A2(pi0224), .ZN(new_n37202_));
  AOI21_X1   g33894(.A1(pi0588), .A2(new_n37202_), .B(new_n37201_), .ZN(new_n37203_));
  NOR3_X1    g33895(.A1(new_n6933_), .A2(pi0591), .A3(pi0592), .ZN(new_n37204_));
  NAND2_X1   g33896(.A1(new_n37204_), .A2(pi0323), .ZN(new_n37205_));
  NAND3_X1   g33897(.A1(new_n37205_), .A2(pi0464), .A3(new_n9787_), .ZN(new_n37206_));
  OAI21_X1   g33898(.A1(new_n37203_), .A2(new_n37206_), .B(new_n6933_), .ZN(new_n37207_));
  AOI21_X1   g33899(.A1(new_n37207_), .A2(new_n37200_), .B(new_n10169_), .ZN(new_n37208_));
  NOR2_X1    g33900(.A1(new_n4959_), .A2(new_n4785_), .ZN(new_n37209_));
  NAND2_X1   g33901(.A1(new_n26463_), .A2(pi1136), .ZN(new_n37210_));
  XOR2_X1    g33902(.A1(new_n37209_), .A2(new_n37210_), .Z(new_n37211_));
  NOR2_X1    g33903(.A1(pi1137), .A2(pi1138), .ZN(new_n37212_));
  INV_X1     g33904(.I(new_n37212_), .ZN(new_n37213_));
  NOR2_X1    g33905(.A1(new_n37213_), .A2(new_n5132_), .ZN(new_n37214_));
  INV_X1     g33906(.I(new_n37214_), .ZN(new_n37215_));
  NOR2_X1    g33907(.A1(new_n4959_), .A2(pi1136), .ZN(new_n37216_));
  NOR2_X1    g33908(.A1(new_n37215_), .A2(new_n37216_), .ZN(new_n37217_));
  INV_X1     g33909(.I(pi0855), .ZN(new_n37218_));
  OAI22_X1   g33910(.A1(new_n17392_), .A2(new_n4785_), .B1(new_n37218_), .B2(new_n4959_), .ZN(new_n37219_));
  NOR2_X1    g33911(.A1(new_n37217_), .A2(new_n37219_), .ZN(new_n37220_));
  AOI21_X1   g33912(.A1(new_n37212_), .A2(pi1135), .B(new_n4785_), .ZN(new_n37221_));
  NOR2_X1    g33913(.A1(new_n37213_), .A2(pi1134), .ZN(new_n37222_));
  NAND3_X1   g33914(.A1(new_n37222_), .A2(pi0766), .A3(new_n37221_), .ZN(new_n37223_));
  OAI22_X1   g33915(.A1(new_n37220_), .A2(new_n37223_), .B1(new_n35633_), .B2(new_n37211_), .ZN(new_n37224_));
  NOR2_X1    g33916(.A1(new_n8549_), .A2(pi1065), .ZN(new_n37225_));
  INV_X1     g33917(.I(new_n37202_), .ZN(new_n37226_));
  NOR2_X1    g33918(.A1(new_n37226_), .A2(new_n8549_), .ZN(new_n37227_));
  XOR2_X1    g33919(.A1(new_n37227_), .A2(new_n37225_), .Z(new_n37228_));
  NOR2_X1    g33920(.A1(new_n4959_), .A2(pi0634), .ZN(new_n37229_));
  XOR2_X1    g33921(.A1(new_n37209_), .A2(new_n37229_), .Z(new_n37230_));
  AND3_X2    g33922(.A1(new_n7250_), .A2(pi0257), .A3(pi0784), .Z(new_n37231_));
  NAND4_X1   g33923(.A1(new_n37224_), .A2(new_n37228_), .A3(new_n37230_), .A4(new_n37231_), .ZN(new_n37232_));
  XNOR2_X1   g33924(.A1(new_n37232_), .A2(new_n37208_), .ZN(po0820));
  AOI21_X1   g33925(.A1(new_n6933_), .A2(pi0592), .B(pi0588), .ZN(new_n37234_));
  NAND2_X1   g33926(.A1(new_n6773_), .A2(new_n6350_), .ZN(new_n37235_));
  NOR2_X1    g33927(.A1(new_n6933_), .A2(new_n6358_), .ZN(new_n37236_));
  OAI21_X1   g33928(.A1(new_n37234_), .A2(new_n37235_), .B(new_n37236_), .ZN(new_n37237_));
  INV_X1     g33929(.I(new_n37203_), .ZN(new_n37238_));
  NAND3_X1   g33930(.A1(new_n37238_), .A2(pi0429), .A3(pi0591), .ZN(new_n37239_));
  AOI21_X1   g33931(.A1(new_n35460_), .A2(new_n37237_), .B(new_n37239_), .ZN(new_n37240_));
  OAI21_X1   g33932(.A1(new_n37240_), .A2(pi0355), .B(new_n37204_), .ZN(new_n37241_));
  INV_X1     g33933(.I(pi0811), .ZN(new_n37242_));
  NAND2_X1   g33934(.A1(new_n13801_), .A2(pi1135), .ZN(new_n37243_));
  XOR2_X1    g33935(.A1(new_n37209_), .A2(new_n37243_), .Z(new_n37244_));
  NAND2_X1   g33936(.A1(new_n12868_), .A2(pi1136), .ZN(new_n37245_));
  XOR2_X1    g33937(.A1(new_n37209_), .A2(new_n37245_), .Z(new_n37246_));
  OAI22_X1   g33938(.A1(new_n5633_), .A2(new_n37246_), .B1(new_n37244_), .B2(new_n37242_), .ZN(new_n37247_));
  NAND2_X1   g33939(.A1(new_n17866_), .A2(pi1136), .ZN(new_n37248_));
  XOR2_X1    g33940(.A1(new_n37209_), .A2(new_n37248_), .Z(new_n37249_));
  OAI21_X1   g33941(.A1(new_n37249_), .A2(new_n17845_), .B(new_n5132_), .ZN(new_n37250_));
  NOR2_X1    g33942(.A1(pi1135), .A2(pi1136), .ZN(new_n37251_));
  INV_X1     g33943(.I(new_n37251_), .ZN(new_n37252_));
  NOR4_X1    g33944(.A1(new_n37213_), .A2(new_n37252_), .A3(new_n36932_), .A4(pi1134), .ZN(new_n37253_));
  NAND4_X1   g33945(.A1(new_n37247_), .A2(new_n7250_), .A3(new_n37250_), .A4(new_n37253_), .ZN(new_n37254_));
  NOR3_X1    g33946(.A1(new_n37226_), .A2(new_n8549_), .A3(new_n35181_), .ZN(new_n37255_));
  NOR3_X1    g33947(.A1(new_n37202_), .A2(new_n8549_), .A3(pi1084), .ZN(new_n37256_));
  OAI21_X1   g33948(.A1(new_n37255_), .A2(new_n37256_), .B(pi0292), .ZN(new_n37257_));
  AOI21_X1   g33949(.A1(new_n37241_), .A2(new_n37254_), .B(new_n37257_), .ZN(po0821));
  NAND3_X1   g33950(.A1(po0954), .A2(pi0962), .A3(pi1108), .ZN(new_n37259_));
  NAND3_X1   g33951(.A1(po0954), .A2(new_n37045_), .A3(new_n37021_), .ZN(new_n37260_));
  AOI21_X1   g33952(.A1(new_n37259_), .A2(new_n37260_), .B(new_n13124_), .ZN(po0822));
  INV_X1     g33953(.I(pi0441), .ZN(new_n37262_));
  INV_X1     g33954(.I(new_n37236_), .ZN(new_n37263_));
  NOR3_X1    g33955(.A1(new_n37234_), .A2(pi0456), .A3(pi0591), .ZN(new_n37264_));
  OAI21_X1   g33956(.A1(new_n37264_), .A2(new_n37263_), .B(new_n35353_), .ZN(new_n37265_));
  NAND4_X1   g33957(.A1(new_n37238_), .A2(pi0443), .A3(pi0591), .A4(new_n37265_), .ZN(new_n37266_));
  NAND2_X1   g33958(.A1(new_n37266_), .A2(new_n37262_), .ZN(new_n37267_));
  AOI21_X1   g33959(.A1(new_n37267_), .A2(new_n37204_), .B(new_n10169_), .ZN(new_n37268_));
  NOR2_X1    g33960(.A1(new_n4959_), .A2(pi0790), .ZN(new_n37269_));
  XOR2_X1    g33961(.A1(new_n37209_), .A2(new_n37269_), .Z(new_n37270_));
  INV_X1     g33962(.I(new_n37217_), .ZN(new_n37271_));
  AOI22_X1   g33963(.A1(pi0691), .A2(pi1136), .B1(pi0873), .B2(pi1135), .ZN(new_n37272_));
  NAND2_X1   g33964(.A1(new_n37271_), .A2(new_n37272_), .ZN(new_n37273_));
  INV_X1     g33965(.I(new_n37221_), .ZN(new_n37274_));
  INV_X1     g33966(.I(new_n37222_), .ZN(new_n37275_));
  NOR3_X1    g33967(.A1(new_n37275_), .A2(new_n18051_), .A3(new_n37274_), .ZN(new_n37276_));
  AOI22_X1   g33968(.A1(new_n37273_), .A2(new_n37276_), .B1(pi0799), .B2(new_n37270_), .ZN(new_n37277_));
  NAND2_X1   g33969(.A1(new_n34014_), .A2(pi0199), .ZN(new_n37278_));
  XOR2_X1    g33970(.A1(new_n37227_), .A2(new_n37278_), .Z(new_n37279_));
  NAND2_X1   g33971(.A1(new_n28263_), .A2(pi1136), .ZN(new_n37280_));
  XOR2_X1    g33972(.A1(new_n37209_), .A2(new_n37280_), .Z(new_n37281_));
  NAND3_X1   g33973(.A1(new_n7250_), .A2(pi0297), .A3(pi0638), .ZN(new_n37282_));
  NOR4_X1    g33974(.A1(new_n37277_), .A2(new_n37279_), .A3(new_n37281_), .A4(new_n37282_), .ZN(new_n37283_));
  XOR2_X1    g33975(.A1(new_n37283_), .A2(new_n37268_), .Z(po0823));
  NAND2_X1   g33976(.A1(new_n6774_), .A2(new_n6350_), .ZN(new_n37285_));
  OAI21_X1   g33977(.A1(new_n37234_), .A2(new_n37285_), .B(new_n37236_), .ZN(new_n37286_));
  NAND3_X1   g33978(.A1(new_n37238_), .A2(pi0444), .A3(pi0591), .ZN(new_n37287_));
  AOI21_X1   g33979(.A1(new_n35356_), .A2(new_n37286_), .B(new_n37287_), .ZN(new_n37288_));
  OAI21_X1   g33980(.A1(new_n37288_), .A2(pi0458), .B(new_n37204_), .ZN(new_n37289_));
  INV_X1     g33981(.I(pi0809), .ZN(new_n37290_));
  NAND2_X1   g33982(.A1(new_n5379_), .A2(pi1136), .ZN(new_n37291_));
  XOR2_X1    g33983(.A1(new_n37209_), .A2(new_n37291_), .Z(new_n37292_));
  NAND2_X1   g33984(.A1(new_n5632_), .A2(pi1135), .ZN(new_n37293_));
  XOR2_X1    g33985(.A1(new_n37209_), .A2(new_n37293_), .Z(new_n37294_));
  OAI22_X1   g33986(.A1(new_n12777_), .A2(new_n37294_), .B1(new_n37292_), .B2(new_n37290_), .ZN(new_n37295_));
  NAND2_X1   g33987(.A1(new_n17943_), .A2(pi1136), .ZN(new_n37296_));
  XOR2_X1    g33988(.A1(new_n37209_), .A2(new_n37296_), .Z(new_n37297_));
  OAI21_X1   g33989(.A1(new_n37297_), .A2(new_n17912_), .B(new_n5132_), .ZN(new_n37298_));
  NOR4_X1    g33990(.A1(new_n37213_), .A2(new_n37252_), .A3(new_n36931_), .A4(pi1134), .ZN(new_n37299_));
  NAND4_X1   g33991(.A1(new_n37295_), .A2(new_n7250_), .A3(new_n37298_), .A4(new_n37299_), .ZN(new_n37300_));
  NOR3_X1    g33992(.A1(new_n37226_), .A2(new_n8549_), .A3(new_n35187_), .ZN(new_n37301_));
  NOR3_X1    g33993(.A1(new_n37202_), .A2(new_n8549_), .A3(pi1072), .ZN(new_n37302_));
  OAI21_X1   g33994(.A1(new_n37301_), .A2(new_n37302_), .B(pi0294), .ZN(new_n37303_));
  AOI21_X1   g33995(.A1(new_n37289_), .A2(new_n37300_), .B(new_n37303_), .ZN(po0824));
  NOR3_X1    g33996(.A1(new_n37234_), .A2(pi0390), .A3(pi0591), .ZN(new_n37305_));
  OAI21_X1   g33997(.A1(new_n37305_), .A2(new_n37263_), .B(new_n6705_), .ZN(new_n37306_));
  NAND4_X1   g33998(.A1(new_n37238_), .A2(pi0414), .A3(pi0591), .A4(new_n37306_), .ZN(new_n37307_));
  NAND2_X1   g33999(.A1(new_n37307_), .A2(new_n6581_), .ZN(new_n37308_));
  AOI21_X1   g34000(.A1(new_n37308_), .A2(new_n37204_), .B(new_n10169_), .ZN(new_n37309_));
  NOR2_X1    g34001(.A1(new_n4959_), .A2(pi0778), .ZN(new_n37310_));
  XOR2_X1    g34002(.A1(new_n37209_), .A2(new_n37310_), .Z(new_n37311_));
  AOI22_X1   g34003(.A1(pi0696), .A2(pi1136), .B1(pi0837), .B2(pi1135), .ZN(new_n37312_));
  NAND2_X1   g34004(.A1(new_n37271_), .A2(new_n37312_), .ZN(new_n37313_));
  NOR3_X1    g34005(.A1(new_n37275_), .A2(new_n17309_), .A3(new_n37274_), .ZN(new_n37314_));
  AOI22_X1   g34006(.A1(new_n37313_), .A2(new_n37314_), .B1(pi0981), .B2(new_n37311_), .ZN(new_n37315_));
  NAND2_X1   g34007(.A1(new_n35178_), .A2(pi0199), .ZN(new_n37316_));
  XOR2_X1    g34008(.A1(new_n37227_), .A2(new_n37316_), .Z(new_n37317_));
  NAND2_X1   g34009(.A1(new_n5794_), .A2(pi1136), .ZN(new_n37318_));
  XOR2_X1    g34010(.A1(new_n37209_), .A2(new_n37318_), .Z(new_n37319_));
  NAND3_X1   g34011(.A1(new_n7250_), .A2(pi0291), .A3(pi0680), .ZN(new_n37320_));
  NOR4_X1    g34012(.A1(new_n37315_), .A2(new_n37317_), .A3(new_n37319_), .A4(new_n37320_), .ZN(new_n37321_));
  XOR2_X1    g34013(.A1(new_n37321_), .A2(new_n37309_), .Z(po0825));
  INV_X1     g34014(.I(pi0669), .ZN(new_n37323_));
  NAND3_X1   g34015(.A1(po0954), .A2(pi0962), .A3(pi1125), .ZN(new_n37324_));
  NAND3_X1   g34016(.A1(po0954), .A2(new_n37045_), .A3(new_n37120_), .ZN(new_n37325_));
  AOI21_X1   g34017(.A1(new_n37324_), .A2(new_n37325_), .B(new_n37323_), .ZN(po0826));
  NAND3_X1   g34018(.A1(pi0364), .A2(pi0591), .A3(pi0592), .ZN(new_n37327_));
  NOR3_X1    g34019(.A1(new_n6350_), .A2(pi0391), .A3(pi0592), .ZN(new_n37328_));
  XOR2_X1    g34020(.A1(new_n37328_), .A2(new_n37327_), .Z(new_n37329_));
  NAND2_X1   g34021(.A1(new_n37204_), .A2(pi0343), .ZN(new_n37330_));
  AND3_X2    g34022(.A1(new_n37201_), .A2(pi0415), .A3(new_n9787_), .Z(new_n37331_));
  AOI21_X1   g34023(.A1(new_n37331_), .A2(new_n37330_), .B(pi0590), .ZN(new_n37332_));
  OAI21_X1   g34024(.A1(new_n37332_), .A2(new_n37329_), .B(new_n7250_), .ZN(new_n37333_));
  AOI22_X1   g34025(.A1(pi0723), .A2(pi1136), .B1(pi0852), .B2(pi1135), .ZN(new_n37334_));
  NAND2_X1   g34026(.A1(new_n37271_), .A2(new_n37334_), .ZN(new_n37335_));
  NAND3_X1   g34027(.A1(new_n37335_), .A2(pi0745), .A3(new_n37221_), .ZN(new_n37336_));
  NAND2_X1   g34028(.A1(new_n28683_), .A2(pi1135), .ZN(new_n37337_));
  NAND2_X1   g34029(.A1(pi1134), .A2(pi1135), .ZN(new_n37338_));
  XOR2_X1    g34030(.A1(new_n37337_), .A2(new_n37338_), .Z(new_n37339_));
  NOR2_X1    g34031(.A1(new_n37213_), .A2(new_n4785_), .ZN(new_n37340_));
  NAND3_X1   g34032(.A1(new_n37339_), .A2(pi0695), .A3(new_n37340_), .ZN(new_n37341_));
  NOR2_X1    g34033(.A1(new_n8549_), .A2(pi1062), .ZN(new_n37342_));
  XOR2_X1    g34034(.A1(new_n37227_), .A2(new_n37342_), .Z(new_n37343_));
  NOR2_X1    g34035(.A1(new_n10169_), .A2(new_n34002_), .ZN(new_n37344_));
  NAND4_X1   g34036(.A1(new_n37336_), .A2(new_n37341_), .A3(new_n37343_), .A4(new_n37344_), .ZN(new_n37345_));
  XOR2_X1    g34037(.A1(new_n37345_), .A2(new_n37333_), .Z(po0827));
  NAND3_X1   g34038(.A1(pi0333), .A2(pi0591), .A3(pi0592), .ZN(new_n37347_));
  NOR3_X1    g34039(.A1(new_n6358_), .A2(pi0447), .A3(pi0591), .ZN(new_n37348_));
  XOR2_X1    g34040(.A1(new_n37348_), .A2(new_n37347_), .Z(new_n37349_));
  NAND2_X1   g34041(.A1(new_n37204_), .A2(pi0327), .ZN(new_n37350_));
  AND3_X2    g34042(.A1(new_n37201_), .A2(pi0453), .A3(new_n9787_), .Z(new_n37351_));
  AOI21_X1   g34043(.A1(new_n37351_), .A2(new_n37350_), .B(pi0590), .ZN(new_n37352_));
  OAI21_X1   g34044(.A1(new_n37352_), .A2(new_n37349_), .B(new_n7250_), .ZN(new_n37353_));
  AOI22_X1   g34045(.A1(pi0724), .A2(pi1136), .B1(pi0865), .B2(pi1135), .ZN(new_n37354_));
  NAND2_X1   g34046(.A1(new_n37271_), .A2(new_n37354_), .ZN(new_n37355_));
  NAND3_X1   g34047(.A1(new_n37355_), .A2(pi0741), .A3(new_n37221_), .ZN(new_n37356_));
  INV_X1     g34048(.I(pi0261), .ZN(new_n37357_));
  INV_X1     g34049(.I(new_n37340_), .ZN(new_n37358_));
  NOR2_X1    g34050(.A1(new_n4959_), .A2(pi0611), .ZN(new_n37359_));
  XOR2_X1    g34051(.A1(new_n37359_), .A2(new_n37338_), .Z(new_n37360_));
  NOR3_X1    g34052(.A1(new_n37360_), .A2(new_n37123_), .A3(new_n37358_), .ZN(new_n37361_));
  NAND2_X1   g34053(.A1(new_n34023_), .A2(pi0199), .ZN(new_n37362_));
  XOR2_X1    g34054(.A1(new_n37227_), .A2(new_n37362_), .Z(new_n37363_));
  NOR4_X1    g34055(.A1(new_n37361_), .A2(new_n37363_), .A3(new_n37357_), .A4(new_n10169_), .ZN(new_n37364_));
  NAND2_X1   g34056(.A1(new_n37356_), .A2(new_n37364_), .ZN(new_n37365_));
  XOR2_X1    g34057(.A1(new_n37365_), .A2(new_n37353_), .Z(po0828));
  NOR3_X1    g34058(.A1(new_n37234_), .A2(pi0397), .A3(pi0591), .ZN(new_n37367_));
  OAI21_X1   g34059(.A1(new_n37367_), .A2(new_n37263_), .B(new_n6707_), .ZN(new_n37368_));
  NAND4_X1   g34060(.A1(new_n37238_), .A2(pi0422), .A3(pi0591), .A4(new_n37368_), .ZN(new_n37369_));
  NAND2_X1   g34061(.A1(new_n37369_), .A2(new_n6584_), .ZN(new_n37370_));
  AOI21_X1   g34062(.A1(new_n37370_), .A2(new_n37204_), .B(new_n10169_), .ZN(new_n37371_));
  NOR2_X1    g34063(.A1(new_n4959_), .A2(pi0781), .ZN(new_n37372_));
  XOR2_X1    g34064(.A1(new_n37209_), .A2(new_n37372_), .Z(new_n37373_));
  AOI22_X1   g34065(.A1(pi0736), .A2(pi1136), .B1(pi0850), .B2(pi1135), .ZN(new_n37374_));
  NAND2_X1   g34066(.A1(new_n37271_), .A2(new_n37374_), .ZN(new_n37375_));
  NOR3_X1    g34067(.A1(new_n37275_), .A2(new_n16090_), .A3(new_n37274_), .ZN(new_n37376_));
  AOI22_X1   g34068(.A1(new_n37375_), .A2(new_n37376_), .B1(pi0808), .B2(new_n37373_), .ZN(new_n37377_));
  NAND2_X1   g34069(.A1(new_n35175_), .A2(pi0199), .ZN(new_n37378_));
  XOR2_X1    g34070(.A1(new_n37227_), .A2(new_n37378_), .Z(new_n37379_));
  NAND2_X1   g34071(.A1(new_n12841_), .A2(pi1136), .ZN(new_n37380_));
  XOR2_X1    g34072(.A1(new_n37209_), .A2(new_n37380_), .Z(new_n37381_));
  NAND3_X1   g34073(.A1(new_n7250_), .A2(pi0290), .A3(pi0661), .ZN(new_n37382_));
  NOR4_X1    g34074(.A1(new_n37377_), .A2(new_n37379_), .A3(new_n37381_), .A4(new_n37382_), .ZN(new_n37383_));
  XOR2_X1    g34075(.A1(new_n37383_), .A2(new_n37371_), .Z(po0829));
  NOR3_X1    g34076(.A1(new_n37234_), .A2(pi0411), .A3(pi0591), .ZN(new_n37385_));
  OAI21_X1   g34077(.A1(new_n37385_), .A2(new_n37263_), .B(new_n6700_), .ZN(new_n37386_));
  NAND4_X1   g34078(.A1(new_n37238_), .A2(pi0435), .A3(pi0591), .A4(new_n37386_), .ZN(new_n37387_));
  NAND2_X1   g34079(.A1(new_n37387_), .A2(new_n6596_), .ZN(new_n37388_));
  AOI21_X1   g34080(.A1(new_n37388_), .A2(new_n37204_), .B(new_n10169_), .ZN(new_n37389_));
  NOR2_X1    g34081(.A1(new_n4959_), .A2(pi0788), .ZN(new_n37390_));
  XOR2_X1    g34082(.A1(new_n37209_), .A2(new_n37390_), .Z(new_n37391_));
  AOI22_X1   g34083(.A1(pi0706), .A2(pi1136), .B1(pi0866), .B2(pi1135), .ZN(new_n37392_));
  NAND2_X1   g34084(.A1(new_n37271_), .A2(new_n37392_), .ZN(new_n37393_));
  NOR3_X1    g34085(.A1(new_n37275_), .A2(new_n14263_), .A3(new_n37274_), .ZN(new_n37394_));
  AOI22_X1   g34086(.A1(new_n37393_), .A2(new_n37394_), .B1(pi0814), .B2(new_n37391_), .ZN(new_n37395_));
  NAND2_X1   g34087(.A1(new_n33607_), .A2(pi0199), .ZN(new_n37396_));
  XOR2_X1    g34088(.A1(new_n37227_), .A2(new_n37396_), .Z(new_n37397_));
  NAND2_X1   g34089(.A1(new_n26964_), .A2(pi1136), .ZN(new_n37398_));
  XOR2_X1    g34090(.A1(new_n37209_), .A2(new_n37398_), .Z(new_n37399_));
  NAND3_X1   g34091(.A1(new_n7250_), .A2(pi0295), .A3(pi0637), .ZN(new_n37400_));
  NOR4_X1    g34092(.A1(new_n37395_), .A2(new_n37397_), .A3(new_n37399_), .A4(new_n37400_), .ZN(new_n37401_));
  XOR2_X1    g34093(.A1(new_n37401_), .A2(new_n37389_), .Z(po0830));
  NAND3_X1   g34094(.A1(pi0336), .A2(pi0591), .A3(pi0592), .ZN(new_n37403_));
  NOR3_X1    g34095(.A1(new_n6350_), .A2(pi0463), .A3(pi0592), .ZN(new_n37404_));
  XNOR2_X1   g34096(.A1(new_n37404_), .A2(new_n37403_), .ZN(new_n37405_));
  AND2_X2    g34097(.A1(new_n37204_), .A2(pi0362), .Z(new_n37406_));
  NAND3_X1   g34098(.A1(new_n37201_), .A2(pi0437), .A3(new_n9787_), .ZN(new_n37407_));
  OAI21_X1   g34099(.A1(new_n37407_), .A2(new_n37406_), .B(new_n6933_), .ZN(new_n37408_));
  NAND2_X1   g34100(.A1(new_n37408_), .A2(new_n37405_), .ZN(new_n37409_));
  INV_X1     g34101(.I(pi0783), .ZN(new_n37410_));
  NAND2_X1   g34102(.A1(new_n37410_), .A2(pi1135), .ZN(new_n37411_));
  XOR2_X1    g34103(.A1(new_n37209_), .A2(new_n37411_), .Z(new_n37412_));
  NAND2_X1   g34104(.A1(new_n28296_), .A2(pi1136), .ZN(new_n37413_));
  XOR2_X1    g34105(.A1(new_n37209_), .A2(new_n37413_), .Z(new_n37414_));
  OAI22_X1   g34106(.A1(new_n28297_), .A2(new_n37414_), .B1(new_n37412_), .B2(new_n35621_), .ZN(new_n37415_));
  NAND2_X1   g34107(.A1(new_n14833_), .A2(pi1136), .ZN(new_n37416_));
  XOR2_X1    g34108(.A1(new_n37209_), .A2(new_n37416_), .Z(new_n37417_));
  OAI21_X1   g34109(.A1(new_n37417_), .A2(new_n14921_), .B(new_n5132_), .ZN(new_n37418_));
  INV_X1     g34110(.I(pi0859), .ZN(new_n37419_));
  NOR4_X1    g34111(.A1(new_n37213_), .A2(new_n37252_), .A3(new_n37419_), .A4(pi1134), .ZN(new_n37420_));
  NAND4_X1   g34112(.A1(new_n37415_), .A2(new_n7250_), .A3(new_n37418_), .A4(new_n37420_), .ZN(new_n37421_));
  NOR3_X1    g34113(.A1(new_n37226_), .A2(new_n8549_), .A3(new_n33991_), .ZN(new_n37422_));
  NOR3_X1    g34114(.A1(new_n37202_), .A2(new_n8549_), .A3(pi1070), .ZN(new_n37423_));
  OAI21_X1   g34115(.A1(new_n37422_), .A2(new_n37423_), .B(pi0256), .ZN(new_n37424_));
  AOI21_X1   g34116(.A1(new_n37421_), .A2(new_n37409_), .B(new_n37424_), .ZN(po0831));
  INV_X1     g34117(.I(new_n37204_), .ZN(new_n37426_));
  NOR3_X1    g34118(.A1(new_n37234_), .A2(pi0412), .A3(pi0591), .ZN(new_n37427_));
  OAI21_X1   g34119(.A1(new_n37427_), .A2(new_n37263_), .B(new_n6699_), .ZN(new_n37428_));
  NOR3_X1    g34120(.A1(new_n37203_), .A2(new_n7218_), .A3(new_n6350_), .ZN(new_n37429_));
  AOI21_X1   g34121(.A1(new_n37429_), .A2(new_n37428_), .B(pi0455), .ZN(new_n37430_));
  OAI21_X1   g34122(.A1(new_n37430_), .A2(new_n37426_), .B(new_n7250_), .ZN(new_n37431_));
  NAND2_X1   g34123(.A1(new_n18025_), .A2(pi1136), .ZN(new_n37432_));
  XOR2_X1    g34124(.A1(new_n37209_), .A2(new_n37432_), .Z(new_n37433_));
  NOR3_X1    g34125(.A1(new_n37433_), .A2(new_n18000_), .A3(new_n37215_), .ZN(new_n37434_));
  NOR3_X1    g34126(.A1(new_n37275_), .A2(pi1135), .A3(pi1136), .ZN(new_n37438_));
  OAI21_X1   g34127(.A1(new_n37434_), .A2(pi0876), .B(new_n37438_), .ZN(new_n37439_));
  NOR2_X1    g34128(.A1(new_n8549_), .A2(pi1037), .ZN(new_n37440_));
  XOR2_X1    g34129(.A1(new_n37227_), .A2(new_n37440_), .Z(new_n37441_));
  NAND4_X1   g34130(.A1(new_n37441_), .A2(pi0296), .A3(pi0623), .A4(new_n7250_), .ZN(new_n37442_));
  AOI21_X1   g34131(.A1(new_n37274_), .A2(new_n37439_), .B(new_n37442_), .ZN(new_n37443_));
  XNOR2_X1   g34132(.A1(new_n37443_), .A2(new_n37431_), .ZN(po0832));
  INV_X1     g34133(.I(pi0361), .ZN(new_n37445_));
  NOR3_X1    g34134(.A1(new_n37234_), .A2(pi0410), .A3(pi0591), .ZN(new_n37446_));
  OAI21_X1   g34135(.A1(new_n37446_), .A2(new_n37263_), .B(new_n6708_), .ZN(new_n37447_));
  NAND4_X1   g34136(.A1(new_n37238_), .A2(pi0434), .A3(pi0591), .A4(new_n37447_), .ZN(new_n37448_));
  NAND2_X1   g34137(.A1(new_n37448_), .A2(new_n37445_), .ZN(new_n37449_));
  AOI21_X1   g34138(.A1(new_n37449_), .A2(new_n37204_), .B(new_n10169_), .ZN(new_n37450_));
  NOR2_X1    g34139(.A1(new_n4959_), .A2(pi0787), .ZN(new_n37451_));
  XOR2_X1    g34140(.A1(new_n37209_), .A2(new_n37451_), .Z(new_n37452_));
  AOI22_X1   g34141(.A1(pi0729), .A2(pi1136), .B1(pi0881), .B2(pi1135), .ZN(new_n37453_));
  NAND2_X1   g34142(.A1(new_n37271_), .A2(new_n37453_), .ZN(new_n37454_));
  NOR3_X1    g34143(.A1(new_n37275_), .A2(new_n17956_), .A3(new_n37274_), .ZN(new_n37455_));
  AOI22_X1   g34144(.A1(new_n37454_), .A2(new_n37455_), .B1(pi0812), .B2(new_n37452_), .ZN(new_n37456_));
  NAND2_X1   g34145(.A1(new_n35184_), .A2(pi0199), .ZN(new_n37457_));
  XOR2_X1    g34146(.A1(new_n37227_), .A2(new_n37457_), .Z(new_n37458_));
  NAND2_X1   g34147(.A1(new_n27261_), .A2(pi1136), .ZN(new_n37459_));
  XOR2_X1    g34148(.A1(new_n37209_), .A2(new_n37459_), .Z(new_n37460_));
  NAND3_X1   g34149(.A1(new_n7250_), .A2(pi0293), .A3(pi0643), .ZN(new_n37461_));
  NOR4_X1    g34150(.A1(new_n37456_), .A2(new_n37458_), .A3(new_n37460_), .A4(new_n37461_), .ZN(new_n37462_));
  XOR2_X1    g34151(.A1(new_n37462_), .A2(new_n37450_), .Z(po0833));
  NAND3_X1   g34152(.A1(pi0335), .A2(pi0591), .A3(pi0592), .ZN(new_n37464_));
  NOR3_X1    g34153(.A1(new_n6358_), .A2(pi0366), .A3(pi0591), .ZN(new_n37465_));
  XOR2_X1    g34154(.A1(new_n37465_), .A2(new_n37464_), .Z(new_n37466_));
  NAND2_X1   g34155(.A1(new_n37204_), .A2(pi0344), .ZN(new_n37467_));
  INV_X1     g34156(.I(new_n37201_), .ZN(new_n37468_));
  NOR3_X1    g34157(.A1(new_n37468_), .A2(new_n7046_), .A3(pi0588), .ZN(new_n37469_));
  AOI21_X1   g34158(.A1(new_n37469_), .A2(new_n37467_), .B(pi0590), .ZN(new_n37470_));
  OAI21_X1   g34159(.A1(new_n37470_), .A2(new_n37466_), .B(new_n7250_), .ZN(new_n37471_));
  AOI22_X1   g34160(.A1(pi0704), .A2(pi1136), .B1(pi0870), .B2(pi1135), .ZN(new_n37472_));
  NAND2_X1   g34161(.A1(new_n37271_), .A2(new_n37472_), .ZN(new_n37473_));
  NAND3_X1   g34162(.A1(new_n37473_), .A2(pi0742), .A3(new_n37221_), .ZN(new_n37474_));
  INV_X1     g34163(.I(pi0259), .ZN(new_n37475_));
  NOR2_X1    g34164(.A1(new_n4959_), .A2(pi0620), .ZN(new_n37476_));
  XOR2_X1    g34165(.A1(new_n37476_), .A2(new_n37338_), .Z(new_n37477_));
  NOR3_X1    g34166(.A1(new_n37477_), .A2(new_n37081_), .A3(new_n37358_), .ZN(new_n37478_));
  NAND2_X1   g34167(.A1(new_n34009_), .A2(pi0199), .ZN(new_n37479_));
  XOR2_X1    g34168(.A1(new_n37227_), .A2(new_n37479_), .Z(new_n37480_));
  NOR4_X1    g34169(.A1(new_n37478_), .A2(new_n37480_), .A3(new_n37475_), .A4(new_n10169_), .ZN(new_n37481_));
  NAND2_X1   g34170(.A1(new_n37474_), .A2(new_n37481_), .ZN(new_n37482_));
  XOR2_X1    g34171(.A1(new_n37482_), .A2(new_n37471_), .Z(po0834));
  NAND3_X1   g34172(.A1(pi0368), .A2(pi0591), .A3(pi0592), .ZN(new_n37484_));
  NOR3_X1    g34173(.A1(new_n6350_), .A2(pi0393), .A3(pi0592), .ZN(new_n37485_));
  XOR2_X1    g34174(.A1(new_n37485_), .A2(new_n37484_), .Z(new_n37486_));
  NAND2_X1   g34175(.A1(new_n37204_), .A2(pi0346), .ZN(new_n37487_));
  NOR3_X1    g34176(.A1(new_n37468_), .A2(new_n7064_), .A3(pi0588), .ZN(new_n37488_));
  AOI21_X1   g34177(.A1(new_n37488_), .A2(new_n37487_), .B(pi0590), .ZN(new_n37489_));
  OAI21_X1   g34178(.A1(new_n37489_), .A2(new_n37486_), .B(new_n7250_), .ZN(new_n37490_));
  AOI22_X1   g34179(.A1(pi0688), .A2(pi1136), .B1(pi0856), .B2(pi1135), .ZN(new_n37491_));
  NAND2_X1   g34180(.A1(new_n37271_), .A2(new_n37491_), .ZN(new_n37492_));
  NAND3_X1   g34181(.A1(new_n37492_), .A2(pi0760), .A3(new_n37221_), .ZN(new_n37493_));
  NAND2_X1   g34182(.A1(new_n36984_), .A2(pi1135), .ZN(new_n37494_));
  XOR2_X1    g34183(.A1(new_n37494_), .A2(new_n37338_), .Z(new_n37495_));
  NAND3_X1   g34184(.A1(new_n37495_), .A2(pi0632), .A3(new_n37340_), .ZN(new_n37496_));
  NOR2_X1    g34185(.A1(new_n8549_), .A2(pi1067), .ZN(new_n37497_));
  XOR2_X1    g34186(.A1(new_n37227_), .A2(new_n37497_), .Z(new_n37498_));
  AND2_X2    g34187(.A1(new_n7250_), .A2(pi0260), .Z(new_n37499_));
  NAND4_X1   g34188(.A1(new_n37493_), .A2(new_n37496_), .A3(new_n37498_), .A4(new_n37499_), .ZN(new_n37500_));
  XOR2_X1    g34189(.A1(new_n37500_), .A2(new_n37490_), .Z(po0835));
  NAND3_X1   g34190(.A1(pi0389), .A2(pi0591), .A3(pi0592), .ZN(new_n37502_));
  NOR3_X1    g34191(.A1(new_n6350_), .A2(pi0413), .A3(pi0592), .ZN(new_n37503_));
  XOR2_X1    g34192(.A1(new_n37503_), .A2(new_n37502_), .Z(new_n37504_));
  NAND2_X1   g34193(.A1(new_n37204_), .A2(pi0450), .ZN(new_n37505_));
  AND3_X2    g34194(.A1(new_n37201_), .A2(pi0438), .A3(new_n9787_), .Z(new_n37506_));
  AOI21_X1   g34195(.A1(new_n37506_), .A2(new_n37505_), .B(pi0590), .ZN(new_n37507_));
  OAI21_X1   g34196(.A1(new_n37507_), .A2(new_n37504_), .B(new_n7250_), .ZN(new_n37508_));
  NOR2_X1    g34197(.A1(new_n4785_), .A2(pi0621), .ZN(new_n37509_));
  XOR2_X1    g34198(.A1(new_n37209_), .A2(new_n37509_), .Z(new_n37510_));
  AOI22_X1   g34199(.A1(pi0690), .A2(pi1136), .B1(pi0874), .B2(pi1135), .ZN(new_n37511_));
  NAND2_X1   g34200(.A1(new_n37271_), .A2(new_n37511_), .ZN(new_n37512_));
  NOR3_X1    g34201(.A1(new_n37275_), .A2(new_n18095_), .A3(new_n37274_), .ZN(new_n37513_));
  AOI22_X1   g34202(.A1(new_n37512_), .A2(new_n37513_), .B1(pi0810), .B2(new_n37510_), .ZN(new_n37514_));
  NAND2_X1   g34203(.A1(new_n33985_), .A2(pi0199), .ZN(new_n37515_));
  XOR2_X1    g34204(.A1(new_n37227_), .A2(new_n37515_), .Z(new_n37516_));
  NAND2_X1   g34205(.A1(new_n13124_), .A2(pi1135), .ZN(new_n37517_));
  XOR2_X1    g34206(.A1(new_n37209_), .A2(new_n37517_), .Z(new_n37518_));
  NAND3_X1   g34207(.A1(new_n7250_), .A2(pi0255), .A3(pi0791), .ZN(new_n37519_));
  NOR4_X1    g34208(.A1(new_n37514_), .A2(new_n37516_), .A3(new_n37518_), .A4(new_n37519_), .ZN(new_n37520_));
  XNOR2_X1   g34209(.A1(new_n37520_), .A2(new_n37508_), .ZN(po0836));
  NAND3_X1   g34210(.A1(po0954), .A2(pi0962), .A3(pi1100), .ZN(new_n37522_));
  INV_X1     g34211(.I(pi1100), .ZN(new_n37523_));
  NAND3_X1   g34212(.A1(po0954), .A2(new_n37045_), .A3(new_n37523_), .ZN(new_n37524_));
  AOI21_X1   g34213(.A1(new_n37522_), .A2(new_n37524_), .B(new_n5375_), .ZN(po0837));
  NAND3_X1   g34214(.A1(po0954), .A2(pi0962), .A3(pi1103), .ZN(new_n37526_));
  NAND3_X1   g34215(.A1(po0954), .A2(new_n37045_), .A3(new_n37108_), .ZN(new_n37527_));
  AOI21_X1   g34216(.A1(new_n37526_), .A2(new_n37527_), .B(new_n5632_), .ZN(po0838));
  NAND3_X1   g34217(.A1(pi0367), .A2(pi0591), .A3(pi0592), .ZN(new_n37529_));
  NOR3_X1    g34218(.A1(new_n6350_), .A2(pi0392), .A3(pi0592), .ZN(new_n37530_));
  XOR2_X1    g34219(.A1(new_n37530_), .A2(new_n37529_), .Z(new_n37531_));
  NAND2_X1   g34220(.A1(new_n37204_), .A2(pi0345), .ZN(new_n37532_));
  NOR3_X1    g34221(.A1(new_n37468_), .A2(new_n7063_), .A3(pi0588), .ZN(new_n37533_));
  AOI21_X1   g34222(.A1(new_n37533_), .A2(new_n37532_), .B(pi0590), .ZN(new_n37534_));
  OAI21_X1   g34223(.A1(new_n37534_), .A2(new_n37531_), .B(new_n7250_), .ZN(new_n37535_));
  AOI22_X1   g34224(.A1(pi0686), .A2(pi1136), .B1(pi0848), .B2(pi1135), .ZN(new_n37536_));
  NAND2_X1   g34225(.A1(new_n37271_), .A2(new_n37536_), .ZN(new_n37537_));
  NAND3_X1   g34226(.A1(new_n37537_), .A2(pi0757), .A3(new_n37221_), .ZN(new_n37538_));
  NAND2_X1   g34227(.A1(new_n36970_), .A2(pi1135), .ZN(new_n37539_));
  XOR2_X1    g34228(.A1(new_n37539_), .A2(new_n37338_), .Z(new_n37540_));
  NAND3_X1   g34229(.A1(new_n37540_), .A2(pi0631), .A3(new_n37340_), .ZN(new_n37541_));
  NOR2_X1    g34230(.A1(new_n8549_), .A2(pi1039), .ZN(new_n37542_));
  XOR2_X1    g34231(.A1(new_n37227_), .A2(new_n37542_), .Z(new_n37543_));
  AND2_X2    g34232(.A1(new_n7250_), .A2(pi0251), .Z(new_n37544_));
  NAND4_X1   g34233(.A1(new_n37538_), .A2(new_n37541_), .A3(new_n37543_), .A4(new_n37544_), .ZN(new_n37545_));
  XOR2_X1    g34234(.A1(new_n37545_), .A2(new_n37535_), .Z(po0839));
  INV_X1     g34235(.I(pi0684), .ZN(new_n37547_));
  NAND2_X1   g34236(.A1(new_n37041_), .A2(pi0953), .ZN(new_n37548_));
  INV_X1     g34237(.I(new_n37548_), .ZN(po0980));
  NAND3_X1   g34238(.A1(po0980), .A2(pi0962), .A3(pi1130), .ZN(new_n37550_));
  NAND3_X1   g34239(.A1(po0980), .A2(new_n37045_), .A3(new_n37144_), .ZN(new_n37551_));
  AOI21_X1   g34240(.A1(new_n37550_), .A2(new_n37551_), .B(new_n37547_), .ZN(po0841));
  NOR2_X1    g34241(.A1(new_n4785_), .A2(pi0728), .ZN(new_n37553_));
  XOR2_X1    g34242(.A1(new_n37209_), .A2(new_n37553_), .Z(new_n37554_));
  INV_X1     g34243(.I(pi0744), .ZN(new_n37555_));
  NOR2_X1    g34244(.A1(new_n37215_), .A2(new_n37555_), .ZN(new_n37556_));
  AOI21_X1   g34245(.A1(new_n37556_), .A2(new_n37554_), .B(pi0860), .ZN(new_n37557_));
  OAI21_X1   g34246(.A1(new_n37557_), .A2(new_n37252_), .B(new_n7250_), .ZN(new_n37558_));
  NAND3_X1   g34247(.A1(pi0357), .A2(pi0590), .A3(pi0592), .ZN(new_n37559_));
  NAND3_X1   g34248(.A1(new_n35465_), .A2(new_n6933_), .A3(pi0592), .ZN(new_n37560_));
  XOR2_X1    g34249(.A1(new_n37560_), .A2(new_n37559_), .Z(new_n37561_));
  NOR2_X1    g34250(.A1(new_n6935_), .A2(new_n6358_), .ZN(new_n37562_));
  INV_X1     g34251(.I(new_n37562_), .ZN(new_n37563_));
  NAND2_X1   g34252(.A1(pi0406), .A2(pi0588), .ZN(new_n37564_));
  OAI21_X1   g34253(.A1(new_n37563_), .A2(new_n37564_), .B(new_n6350_), .ZN(new_n37565_));
  NOR4_X1    g34254(.A1(new_n8549_), .A2(new_n35404_), .A3(pi0223), .A4(pi0224), .ZN(new_n37566_));
  AOI21_X1   g34255(.A1(new_n37565_), .A2(new_n37561_), .B(new_n37566_), .ZN(new_n37567_));
  NOR3_X1    g34256(.A1(new_n37147_), .A2(new_n4959_), .A3(new_n4785_), .ZN(new_n37568_));
  NOR3_X1    g34257(.A1(new_n4785_), .A2(pi0652), .A3(pi1135), .ZN(new_n37569_));
  OAI21_X1   g34258(.A1(new_n37568_), .A2(new_n37569_), .B(pi0657), .ZN(new_n37570_));
  NOR2_X1    g34259(.A1(new_n37212_), .A2(pi0813), .ZN(new_n37571_));
  NAND2_X1   g34260(.A1(new_n37570_), .A2(new_n37571_), .ZN(new_n37572_));
  AOI21_X1   g34261(.A1(new_n37572_), .A2(new_n37251_), .B(pi1134), .ZN(new_n37573_));
  NAND2_X1   g34262(.A1(new_n7250_), .A2(pi0430), .ZN(new_n37574_));
  NOR2_X1    g34263(.A1(new_n9787_), .A2(pi0590), .ZN(new_n37575_));
  NOR2_X1    g34264(.A1(new_n6350_), .A2(new_n6358_), .ZN(new_n37576_));
  NAND2_X1   g34265(.A1(new_n37576_), .A2(new_n37575_), .ZN(new_n37577_));
  NOR2_X1    g34266(.A1(new_n37358_), .A2(new_n37577_), .ZN(new_n37578_));
  INV_X1     g34267(.I(new_n37578_), .ZN(new_n37579_));
  NOR4_X1    g34268(.A1(new_n37567_), .A2(new_n37573_), .A3(new_n37574_), .A4(new_n37579_), .ZN(new_n37580_));
  XNOR2_X1   g34269(.A1(new_n37580_), .A2(new_n37558_), .ZN(po0842));
  NAND3_X1   g34270(.A1(po0980), .A2(pi0962), .A3(pi1113), .ZN(new_n37582_));
  NAND3_X1   g34271(.A1(po0980), .A2(new_n37045_), .A3(new_n36972_), .ZN(new_n37583_));
  AOI21_X1   g34272(.A1(new_n37582_), .A2(new_n37583_), .B(new_n17440_), .ZN(po0843));
  NAND3_X1   g34273(.A1(po0980), .A2(pi0962), .A3(pi1127), .ZN(new_n37585_));
  NAND3_X1   g34274(.A1(po0980), .A2(new_n37045_), .A3(new_n37087_), .ZN(new_n37586_));
  AOI21_X1   g34275(.A1(new_n37585_), .A2(new_n37586_), .B(new_n15572_), .ZN(po0844));
  NAND3_X1   g34276(.A1(po0980), .A2(pi0962), .A3(pi1115), .ZN(new_n37588_));
  NAND3_X1   g34277(.A1(po0980), .A2(new_n37045_), .A3(new_n36986_), .ZN(new_n37589_));
  AOI21_X1   g34278(.A1(new_n37588_), .A2(new_n37589_), .B(new_n17495_), .ZN(po0845));
  INV_X1     g34279(.I(pi0843), .ZN(new_n37591_));
  OAI22_X1   g34280(.A1(new_n17777_), .A2(new_n4785_), .B1(new_n37591_), .B2(new_n4959_), .ZN(new_n37592_));
  NOR2_X1    g34281(.A1(new_n37217_), .A2(new_n37592_), .ZN(new_n37593_));
  NAND2_X1   g34282(.A1(new_n37221_), .A2(pi0752), .ZN(new_n37594_));
  OAI21_X1   g34283(.A1(new_n37593_), .A2(new_n37594_), .B(new_n7250_), .ZN(new_n37595_));
  NAND3_X1   g34284(.A1(pi0351), .A2(pi0590), .A3(pi0592), .ZN(new_n37596_));
  NAND3_X1   g34285(.A1(new_n35450_), .A2(new_n6933_), .A3(pi0592), .ZN(new_n37597_));
  XOR2_X1    g34286(.A1(new_n37597_), .A2(new_n37596_), .Z(new_n37598_));
  NAND2_X1   g34287(.A1(pi0401), .A2(pi0588), .ZN(new_n37599_));
  OAI21_X1   g34288(.A1(new_n37563_), .A2(new_n37599_), .B(new_n6350_), .ZN(new_n37600_));
  NOR4_X1    g34289(.A1(new_n33987_), .A2(new_n8549_), .A3(new_n35388_), .A4(new_n37226_), .ZN(new_n37601_));
  AOI21_X1   g34290(.A1(new_n37600_), .A2(new_n37598_), .B(new_n37601_), .ZN(new_n37602_));
  NAND2_X1   g34291(.A1(new_n37161_), .A2(pi1136), .ZN(new_n37603_));
  XNOR2_X1   g34292(.A1(new_n37209_), .A2(new_n37603_), .ZN(new_n37604_));
  NOR2_X1    g34293(.A1(new_n37275_), .A2(new_n37174_), .ZN(new_n37605_));
  AOI21_X1   g34294(.A1(new_n37605_), .A2(new_n37604_), .B(pi0798), .ZN(new_n37606_));
  NAND3_X1   g34295(.A1(new_n7250_), .A2(new_n37251_), .A3(pi0426), .ZN(new_n37607_));
  NOR4_X1    g34296(.A1(new_n37602_), .A2(new_n37577_), .A3(new_n37606_), .A4(new_n37607_), .ZN(new_n37608_));
  XNOR2_X1   g34297(.A1(new_n37608_), .A2(new_n37595_), .ZN(po0846));
  NAND3_X1   g34298(.A1(po0980), .A2(pi0962), .A3(pi1108), .ZN(new_n37610_));
  NAND3_X1   g34299(.A1(po0980), .A2(new_n37045_), .A3(new_n37021_), .ZN(new_n37611_));
  AOI21_X1   g34300(.A1(new_n37610_), .A2(new_n37611_), .B(new_n18129_), .ZN(po0847));
  NAND3_X1   g34301(.A1(po0980), .A2(pi0962), .A3(pi1107), .ZN(new_n37613_));
  NAND3_X1   g34302(.A1(po0980), .A2(new_n37045_), .A3(new_n36959_), .ZN(new_n37614_));
  AOI21_X1   g34303(.A1(new_n37613_), .A2(new_n37614_), .B(new_n18082_), .ZN(po0848));
  NAND3_X1   g34304(.A1(pi0726), .A2(pi1135), .A3(pi1136), .ZN(new_n37616_));
  NAND3_X1   g34305(.A1(new_n16962_), .A2(new_n4959_), .A3(pi1136), .ZN(new_n37617_));
  NAND2_X1   g34306(.A1(new_n37617_), .A2(new_n37616_), .ZN(new_n37618_));
  AOI21_X1   g34307(.A1(new_n37618_), .A2(pi0770), .B(pi1134), .ZN(new_n37619_));
  NAND3_X1   g34308(.A1(new_n7250_), .A2(new_n37251_), .A3(pi0844), .ZN(new_n37620_));
  NAND3_X1   g34309(.A1(pi0317), .A2(pi0590), .A3(pi0592), .ZN(new_n37621_));
  NOR3_X1    g34310(.A1(new_n6933_), .A2(pi0352), .A3(pi0592), .ZN(new_n37622_));
  XNOR2_X1   g34311(.A1(new_n37622_), .A2(new_n37621_), .ZN(new_n37623_));
  NAND2_X1   g34312(.A1(pi0402), .A2(pi0588), .ZN(new_n37624_));
  OAI21_X1   g34313(.A1(new_n37563_), .A2(new_n37624_), .B(new_n6350_), .ZN(new_n37625_));
  NOR4_X1    g34314(.A1(new_n33999_), .A2(new_n8549_), .A3(new_n35391_), .A4(new_n37226_), .ZN(new_n37626_));
  AOI21_X1   g34315(.A1(new_n37625_), .A2(new_n37623_), .B(new_n37626_), .ZN(new_n37627_));
  NAND3_X1   g34316(.A1(pi0649), .A2(pi1135), .A3(pi1136), .ZN(new_n37628_));
  NAND3_X1   g34317(.A1(new_n37133_), .A2(new_n4959_), .A3(pi1136), .ZN(new_n37629_));
  AOI21_X1   g34318(.A1(new_n37629_), .A2(new_n37628_), .B(new_n37166_), .ZN(new_n37630_));
  INV_X1     g34319(.I(pi0801), .ZN(new_n37631_));
  NOR2_X1    g34320(.A1(new_n37252_), .A2(new_n37631_), .ZN(new_n37632_));
  OAI21_X1   g34321(.A1(new_n37630_), .A2(pi1134), .B(new_n37632_), .ZN(new_n37633_));
  NOR4_X1    g34322(.A1(new_n37577_), .A2(new_n7231_), .A3(new_n7250_), .A4(new_n37213_), .ZN(new_n37634_));
  NAND2_X1   g34323(.A1(new_n37633_), .A2(new_n37634_), .ZN(new_n37635_));
  OAI22_X1   g34324(.A1(new_n37627_), .A2(new_n37635_), .B1(new_n37619_), .B2(new_n37620_), .ZN(po0849));
  INV_X1     g34325(.I(pi0693), .ZN(new_n37637_));
  NAND3_X1   g34326(.A1(po0954), .A2(pi0962), .A3(pi1129), .ZN(new_n37638_));
  NAND3_X1   g34327(.A1(po0954), .A2(new_n37045_), .A3(new_n37154_), .ZN(new_n37639_));
  AOI21_X1   g34328(.A1(new_n37638_), .A2(new_n37639_), .B(new_n37637_), .ZN(po0850));
  INV_X1     g34329(.I(pi0694), .ZN(new_n37641_));
  NAND3_X1   g34330(.A1(po0980), .A2(pi0962), .A3(pi1128), .ZN(new_n37642_));
  NAND3_X1   g34331(.A1(po0980), .A2(new_n37045_), .A3(new_n37101_), .ZN(new_n37643_));
  AOI21_X1   g34332(.A1(new_n37642_), .A2(new_n37643_), .B(new_n37641_), .ZN(po0851));
  NAND3_X1   g34333(.A1(po0954), .A2(pi0962), .A3(pi1111), .ZN(new_n37645_));
  NAND3_X1   g34334(.A1(po0954), .A2(new_n37045_), .A3(new_n36981_), .ZN(new_n37646_));
  AOI21_X1   g34335(.A1(new_n37645_), .A2(new_n37646_), .B(new_n28682_), .ZN(po0852));
  NAND3_X1   g34336(.A1(po0980), .A2(pi0962), .A3(pi1100), .ZN(new_n37648_));
  NAND3_X1   g34337(.A1(po0980), .A2(new_n37045_), .A3(new_n37523_), .ZN(new_n37649_));
  AOI21_X1   g34338(.A1(new_n37648_), .A2(new_n37649_), .B(new_n17327_), .ZN(po0853));
  INV_X1     g34339(.I(pi0697), .ZN(new_n37651_));
  NAND3_X1   g34340(.A1(po0980), .A2(pi0962), .A3(pi1129), .ZN(new_n37652_));
  NAND3_X1   g34341(.A1(po0980), .A2(new_n37045_), .A3(new_n37154_), .ZN(new_n37653_));
  AOI21_X1   g34342(.A1(new_n37652_), .A2(new_n37653_), .B(new_n37651_), .ZN(po0854));
  NAND3_X1   g34343(.A1(po0980), .A2(pi0962), .A3(pi1116), .ZN(new_n37655_));
  NAND3_X1   g34344(.A1(po0980), .A2(new_n37045_), .A3(new_n36963_), .ZN(new_n37656_));
  AOI21_X1   g34345(.A1(new_n37655_), .A2(new_n37656_), .B(new_n16550_), .ZN(po0855));
  NAND3_X1   g34346(.A1(po0980), .A2(pi0962), .A3(pi1103), .ZN(new_n37658_));
  NAND3_X1   g34347(.A1(po0980), .A2(new_n37045_), .A3(new_n37108_), .ZN(new_n37659_));
  AOI21_X1   g34348(.A1(new_n37658_), .A2(new_n37659_), .B(new_n17943_), .ZN(po0856));
  NAND3_X1   g34349(.A1(po0980), .A2(pi0962), .A3(pi1110), .ZN(new_n37661_));
  NAND3_X1   g34350(.A1(po0980), .A2(new_n37045_), .A3(new_n37075_), .ZN(new_n37662_));
  AOI21_X1   g34351(.A1(new_n37661_), .A2(new_n37662_), .B(new_n17392_), .ZN(po0857));
  NAND3_X1   g34352(.A1(po0980), .A2(pi0962), .A3(pi1123), .ZN(new_n37664_));
  NAND3_X1   g34353(.A1(po0980), .A2(new_n37045_), .A3(new_n37115_), .ZN(new_n37665_));
  AOI21_X1   g34354(.A1(new_n37664_), .A2(new_n37665_), .B(new_n22585_), .ZN(po0858));
  NAND3_X1   g34355(.A1(po0980), .A2(pi0962), .A3(pi1117), .ZN(new_n37667_));
  NAND3_X1   g34356(.A1(po0980), .A2(new_n37045_), .A3(new_n37008_), .ZN(new_n37668_));
  AOI21_X1   g34357(.A1(new_n37667_), .A2(new_n37668_), .B(new_n20724_), .ZN(po0859));
  NAND3_X1   g34358(.A1(po0980), .A2(pi0962), .A3(pi1124), .ZN(new_n37670_));
  NAND3_X1   g34359(.A1(po0980), .A2(new_n37045_), .A3(new_n37163_), .ZN(new_n37671_));
  AOI21_X1   g34360(.A1(new_n37670_), .A2(new_n37671_), .B(new_n17777_), .ZN(po0860));
  NAND3_X1   g34361(.A1(po0980), .A2(pi0962), .A3(pi1112), .ZN(new_n37673_));
  NAND3_X1   g34362(.A1(po0980), .A2(new_n37045_), .A3(new_n37017_), .ZN(new_n37674_));
  AOI21_X1   g34363(.A1(new_n37673_), .A2(new_n37674_), .B(new_n17414_), .ZN(po0861));
  NAND3_X1   g34364(.A1(po0980), .A2(pi0962), .A3(pi1125), .ZN(new_n37676_));
  NAND3_X1   g34365(.A1(po0980), .A2(new_n37045_), .A3(new_n37120_), .ZN(new_n37677_));
  AOI21_X1   g34366(.A1(new_n37676_), .A2(new_n37677_), .B(new_n17880_), .ZN(po0862));
  NAND3_X1   g34367(.A1(po0980), .A2(pi0962), .A3(pi1105), .ZN(new_n37679_));
  NAND3_X1   g34368(.A1(po0980), .A2(new_n37045_), .A3(new_n37002_), .ZN(new_n37680_));
  AOI21_X1   g34369(.A1(new_n37679_), .A2(new_n37680_), .B(new_n14261_), .ZN(po0863));
  INV_X1     g34370(.I(pi0847), .ZN(new_n37682_));
  OAI22_X1   g34371(.A1(new_n20724_), .A2(new_n4785_), .B1(new_n37682_), .B2(new_n4959_), .ZN(new_n37683_));
  NOR2_X1    g34372(.A1(new_n37217_), .A2(new_n37683_), .ZN(new_n37684_));
  NAND2_X1   g34373(.A1(new_n37221_), .A2(pi0753), .ZN(new_n37685_));
  OAI21_X1   g34374(.A1(new_n37684_), .A2(new_n37685_), .B(new_n7250_), .ZN(new_n37686_));
  OAI21_X1   g34375(.A1(pi0223), .A2(pi0224), .B(new_n9787_), .ZN(new_n37692_));
  INV_X1     g34376(.I(pi0347), .ZN(new_n37693_));
  NAND3_X1   g34377(.A1(pi0370), .A2(pi0591), .A3(pi0592), .ZN(new_n37694_));
  NOR3_X1    g34378(.A1(new_n6350_), .A2(pi0395), .A3(pi0592), .ZN(new_n37695_));
  XOR2_X1    g34379(.A1(new_n37695_), .A2(new_n37694_), .Z(new_n37696_));
  NOR2_X1    g34380(.A1(new_n37426_), .A2(new_n6933_), .ZN(new_n37697_));
  INV_X1     g34381(.I(new_n37697_), .ZN(new_n37698_));
  OAI21_X1   g34382(.A1(new_n37696_), .A2(new_n37693_), .B(new_n37698_), .ZN(new_n37699_));
  NOR2_X1    g34383(.A1(new_n4959_), .A2(pi0618), .ZN(new_n37700_));
  XOR2_X1    g34384(.A1(new_n37700_), .A2(new_n37338_), .Z(new_n37701_));
  NOR4_X1    g34385(.A1(new_n37701_), .A2(new_n13823_), .A3(new_n10169_), .A4(new_n37358_), .ZN(new_n37702_));
  NAND3_X1   g34386(.A1(new_n37699_), .A2(new_n37692_), .A3(new_n37702_), .ZN(new_n37703_));
  XOR2_X1    g34387(.A1(new_n37703_), .A2(new_n37686_), .Z(po0864));
  NOR2_X1    g34388(.A1(new_n4959_), .A2(pi0609), .ZN(new_n37705_));
  XOR2_X1    g34389(.A1(new_n37705_), .A2(new_n37338_), .Z(new_n37706_));
  NOR3_X1    g34390(.A1(new_n37706_), .A2(new_n13783_), .A3(new_n37358_), .ZN(new_n37707_));
  NOR2_X1    g34391(.A1(new_n37213_), .A2(new_n37216_), .ZN(new_n37708_));
  OR2_X2     g34392(.A1(pi0857), .A2(pi1136), .Z(new_n37709_));
  AOI21_X1   g34393(.A1(pi1134), .A2(new_n37709_), .B(new_n37708_), .ZN(new_n37710_));
  NAND2_X1   g34394(.A1(pi0709), .A2(pi1135), .ZN(new_n37711_));
  NOR4_X1    g34395(.A1(new_n37707_), .A2(new_n7250_), .A3(new_n37710_), .A4(new_n37711_), .ZN(new_n37712_));
  OAI21_X1   g34396(.A1(new_n37712_), .A2(pi0754), .B(new_n37221_), .ZN(new_n37713_));
  AOI21_X1   g34397(.A1(new_n8555_), .A2(pi0305), .B(new_n8549_), .ZN(new_n37714_));
  OAI21_X1   g34398(.A1(new_n8555_), .A2(new_n35181_), .B(new_n37714_), .ZN(new_n37715_));
  XNOR2_X1   g34399(.A1(new_n37715_), .A2(new_n37227_), .ZN(new_n37716_));
  NAND3_X1   g34400(.A1(new_n37202_), .A2(new_n6350_), .A3(new_n6358_), .ZN(new_n37717_));
  NOR2_X1    g34401(.A1(new_n37575_), .A2(pi0459), .ZN(new_n37718_));
  AOI21_X1   g34402(.A1(new_n37718_), .A2(new_n10169_), .B(new_n37717_), .ZN(new_n37719_));
  AOI21_X1   g34403(.A1(new_n37716_), .A2(pi1058), .B(new_n37719_), .ZN(new_n37720_));
  NAND2_X1   g34404(.A1(new_n37204_), .A2(new_n37202_), .ZN(new_n37721_));
  NAND2_X1   g34405(.A1(pi0321), .A2(pi0588), .ZN(new_n37722_));
  OAI21_X1   g34406(.A1(new_n37721_), .A2(new_n37722_), .B(new_n6933_), .ZN(new_n37723_));
  NAND3_X1   g34407(.A1(new_n37576_), .A2(pi0328), .A3(new_n37202_), .ZN(new_n37724_));
  NOR2_X1    g34408(.A1(new_n6358_), .A2(pi0591), .ZN(new_n37725_));
  NOR2_X1    g34409(.A1(new_n37725_), .A2(pi0442), .ZN(new_n37726_));
  AOI21_X1   g34410(.A1(new_n37724_), .A2(new_n37726_), .B(new_n37226_), .ZN(new_n37727_));
  NAND2_X1   g34411(.A1(new_n37727_), .A2(new_n37723_), .ZN(new_n37728_));
  AOI21_X1   g34412(.A1(new_n37713_), .A2(new_n37720_), .B(new_n37728_), .ZN(po0865));
  NAND3_X1   g34413(.A1(po0980), .A2(pi0962), .A3(pi1118), .ZN(new_n37730_));
  NAND3_X1   g34414(.A1(po0980), .A2(new_n37045_), .A3(new_n36967_), .ZN(new_n37731_));
  AOI21_X1   g34415(.A1(new_n37730_), .A2(new_n37731_), .B(new_n21105_), .ZN(po0866));
  NAND3_X1   g34416(.A1(po0954), .A2(pi0962), .A3(pi1106), .ZN(new_n37733_));
  NAND3_X1   g34417(.A1(po0954), .A2(new_n37045_), .A3(new_n37029_), .ZN(new_n37734_));
  AOI21_X1   g34418(.A1(new_n37733_), .A2(new_n37734_), .B(new_n28176_), .ZN(po0867));
  INV_X1     g34419(.I(pi0858), .ZN(new_n37736_));
  OAI22_X1   g34420(.A1(new_n17148_), .A2(new_n4785_), .B1(new_n37736_), .B2(new_n4959_), .ZN(new_n37737_));
  NOR2_X1    g34421(.A1(new_n37217_), .A2(new_n37737_), .ZN(new_n37738_));
  NAND2_X1   g34422(.A1(new_n37221_), .A2(pi0755), .ZN(new_n37739_));
  OAI21_X1   g34423(.A1(new_n37738_), .A2(new_n37739_), .B(new_n7250_), .ZN(new_n37740_));
  OAI21_X1   g34424(.A1(pi0223), .A2(pi0224), .B(new_n9787_), .ZN(new_n37746_));
  NAND3_X1   g34425(.A1(pi0373), .A2(pi0591), .A3(pi0592), .ZN(new_n37747_));
  NOR3_X1    g34426(.A1(new_n6350_), .A2(pi0398), .A3(pi0592), .ZN(new_n37748_));
  XOR2_X1    g34427(.A1(new_n37748_), .A2(new_n37747_), .Z(new_n37749_));
  OAI21_X1   g34428(.A1(new_n37749_), .A2(new_n6604_), .B(new_n37698_), .ZN(new_n37750_));
  NOR2_X1    g34429(.A1(new_n4959_), .A2(pi0630), .ZN(new_n37751_));
  XOR2_X1    g34430(.A1(new_n37751_), .A2(new_n37338_), .Z(new_n37752_));
  NOR4_X1    g34431(.A1(new_n37752_), .A2(new_n14005_), .A3(new_n10169_), .A4(new_n37358_), .ZN(new_n37753_));
  NAND3_X1   g34432(.A1(new_n37750_), .A2(new_n37746_), .A3(new_n37753_), .ZN(new_n37754_));
  XOR2_X1    g34433(.A1(new_n37754_), .A2(new_n37740_), .Z(po0868));
  NAND3_X1   g34434(.A1(pi0374), .A2(pi0591), .A3(pi0592), .ZN(new_n37756_));
  NAND3_X1   g34435(.A1(new_n6762_), .A2(new_n6358_), .A3(pi0591), .ZN(new_n37757_));
  XOR2_X1    g34436(.A1(new_n37757_), .A2(new_n37756_), .Z(new_n37758_));
  AOI21_X1   g34437(.A1(new_n37758_), .A2(pi0350), .B(new_n37697_), .ZN(new_n37759_));
  INV_X1     g34438(.I(pi0425), .ZN(new_n37760_));
  OAI21_X1   g34439(.A1(new_n37577_), .A2(new_n37760_), .B(new_n37226_), .ZN(new_n37761_));
  NAND2_X1   g34440(.A1(new_n37761_), .A2(pi0588), .ZN(new_n37762_));
  OAI21_X1   g34441(.A1(new_n37759_), .A2(new_n37762_), .B(new_n7250_), .ZN(new_n37763_));
  NAND2_X1   g34442(.A1(new_n37221_), .A2(pi0751), .ZN(new_n37764_));
  INV_X1     g34443(.I(new_n37708_), .ZN(new_n37765_));
  OAI21_X1   g34444(.A1(pi0842), .A2(pi1136), .B(pi1134), .ZN(new_n37766_));
  NAND2_X1   g34445(.A1(new_n37765_), .A2(new_n37766_), .ZN(new_n37767_));
  NAND4_X1   g34446(.A1(new_n37767_), .A2(pi0701), .A3(pi1135), .A4(new_n37764_), .ZN(new_n37768_));
  NOR2_X1    g34447(.A1(new_n4959_), .A2(pi0644), .ZN(new_n37769_));
  XOR2_X1    g34448(.A1(new_n37769_), .A2(new_n37338_), .Z(new_n37770_));
  NOR3_X1    g34449(.A1(new_n37770_), .A2(new_n14200_), .A3(new_n37358_), .ZN(new_n37771_));
  AOI21_X1   g34450(.A1(new_n30650_), .A2(pi1044), .B(new_n37202_), .ZN(new_n37772_));
  NAND2_X1   g34451(.A1(new_n8772_), .A2(pi0298), .ZN(new_n37773_));
  NAND4_X1   g34452(.A1(new_n37773_), .A2(pi0199), .A3(pi1035), .A4(new_n7250_), .ZN(new_n37774_));
  NOR3_X1    g34453(.A1(new_n37771_), .A2(new_n37772_), .A3(new_n37774_), .ZN(new_n37775_));
  NAND2_X1   g34454(.A1(new_n37775_), .A2(new_n37768_), .ZN(new_n37776_));
  XOR2_X1    g34455(.A1(new_n37776_), .A2(new_n37763_), .Z(po0869));
  INV_X1     g34456(.I(pi0854), .ZN(new_n37778_));
  OAI22_X1   g34457(.A1(new_n17604_), .A2(new_n4785_), .B1(new_n37778_), .B2(new_n4959_), .ZN(new_n37779_));
  NOR2_X1    g34458(.A1(new_n37217_), .A2(new_n37779_), .ZN(new_n37780_));
  NAND2_X1   g34459(.A1(new_n37221_), .A2(pi0756), .ZN(new_n37781_));
  OAI21_X1   g34460(.A1(new_n37780_), .A2(new_n37781_), .B(new_n7250_), .ZN(new_n37782_));
  OAI21_X1   g34461(.A1(pi0223), .A2(pi0224), .B(new_n9787_), .ZN(new_n37788_));
  NAND3_X1   g34462(.A1(pi0371), .A2(pi0591), .A3(pi0592), .ZN(new_n37789_));
  NOR3_X1    g34463(.A1(new_n6350_), .A2(pi0396), .A3(pi0592), .ZN(new_n37790_));
  XOR2_X1    g34464(.A1(new_n37790_), .A2(new_n37789_), .Z(new_n37791_));
  OAI21_X1   g34465(.A1(new_n37791_), .A2(new_n6606_), .B(new_n37698_), .ZN(new_n37792_));
  NOR2_X1    g34466(.A1(new_n4959_), .A2(pi0628), .ZN(new_n37793_));
  XOR2_X1    g34467(.A1(new_n37793_), .A2(new_n37338_), .Z(new_n37794_));
  NOR4_X1    g34468(.A1(new_n37794_), .A2(new_n13976_), .A3(new_n10169_), .A4(new_n37358_), .ZN(new_n37795_));
  NAND3_X1   g34469(.A1(new_n37792_), .A2(new_n37788_), .A3(new_n37795_), .ZN(new_n37796_));
  XOR2_X1    g34470(.A1(new_n37796_), .A2(new_n37782_), .Z(po0870));
  NOR2_X1    g34471(.A1(new_n4785_), .A2(pi0697), .ZN(new_n37798_));
  XOR2_X1    g34472(.A1(new_n37209_), .A2(new_n37798_), .Z(new_n37799_));
  INV_X1     g34473(.I(pi0762), .ZN(new_n37800_));
  NOR2_X1    g34474(.A1(new_n37215_), .A2(new_n37800_), .ZN(new_n37801_));
  AOI21_X1   g34475(.A1(new_n37801_), .A2(new_n37799_), .B(pi0867), .ZN(new_n37802_));
  OAI21_X1   g34476(.A1(new_n37802_), .A2(new_n37252_), .B(new_n7250_), .ZN(new_n37803_));
  NAND3_X1   g34477(.A1(pi0439), .A2(pi0590), .A3(pi0592), .ZN(new_n37804_));
  NOR3_X1    g34478(.A1(new_n6933_), .A2(pi0461), .A3(pi0592), .ZN(new_n37805_));
  XOR2_X1    g34479(.A1(new_n37805_), .A2(new_n37804_), .Z(new_n37806_));
  NOR2_X1    g34480(.A1(new_n6820_), .A2(new_n9787_), .ZN(new_n37807_));
  AOI21_X1   g34481(.A1(new_n37562_), .A2(new_n37807_), .B(pi0591), .ZN(new_n37808_));
  NAND4_X1   g34482(.A1(new_n3090_), .A2(new_n3100_), .A3(pi0199), .A4(pi1057), .ZN(new_n37809_));
  OAI21_X1   g34483(.A1(new_n37808_), .A2(new_n37806_), .B(new_n37809_), .ZN(new_n37810_));
  NAND3_X1   g34484(.A1(pi0653), .A2(pi1135), .A3(pi1136), .ZN(new_n37811_));
  NAND3_X1   g34485(.A1(new_n37152_), .A2(new_n4959_), .A3(pi1136), .ZN(new_n37812_));
  AOI21_X1   g34486(.A1(new_n37812_), .A2(new_n37811_), .B(new_n37637_), .ZN(new_n37813_));
  INV_X1     g34487(.I(pi0816), .ZN(new_n37814_));
  NAND2_X1   g34488(.A1(new_n37213_), .A2(new_n37814_), .ZN(new_n37815_));
  OAI21_X1   g34489(.A1(new_n37813_), .A2(new_n37815_), .B(new_n37251_), .ZN(new_n37816_));
  NAND2_X1   g34490(.A1(new_n37816_), .A2(new_n5132_), .ZN(new_n37817_));
  NOR2_X1    g34491(.A1(new_n10169_), .A2(new_n7117_), .ZN(new_n37818_));
  NAND4_X1   g34492(.A1(new_n37810_), .A2(new_n37578_), .A3(new_n37817_), .A4(new_n37818_), .ZN(new_n37819_));
  XOR2_X1    g34493(.A1(new_n37819_), .A2(new_n37803_), .Z(po0871));
  NAND3_X1   g34494(.A1(po0954), .A2(pi0962), .A3(pi1123), .ZN(new_n37821_));
  NAND3_X1   g34495(.A1(po0954), .A2(new_n37045_), .A3(new_n37115_), .ZN(new_n37822_));
  AOI21_X1   g34496(.A1(new_n37821_), .A2(new_n37822_), .B(new_n14200_), .ZN(po0872));
  NOR2_X1    g34497(.A1(new_n4959_), .A2(pi0626), .ZN(new_n37824_));
  XOR2_X1    g34498(.A1(new_n37824_), .A2(new_n37338_), .Z(new_n37825_));
  NOR3_X1    g34499(.A1(new_n37825_), .A2(new_n13922_), .A3(new_n37358_), .ZN(new_n37826_));
  OR2_X2     g34500(.A1(pi0845), .A2(pi1136), .Z(new_n37827_));
  AOI21_X1   g34501(.A1(pi1134), .A2(new_n37827_), .B(new_n37708_), .ZN(new_n37828_));
  NAND2_X1   g34502(.A1(pi0738), .A2(pi1135), .ZN(new_n37829_));
  NOR4_X1    g34503(.A1(new_n37826_), .A2(new_n7250_), .A3(new_n37828_), .A4(new_n37829_), .ZN(new_n37830_));
  OAI21_X1   g34504(.A1(new_n37830_), .A2(pi0761), .B(new_n37221_), .ZN(new_n37831_));
  AOI21_X1   g34505(.A1(new_n8555_), .A2(pi0307), .B(new_n8549_), .ZN(new_n37832_));
  OAI21_X1   g34506(.A1(new_n8555_), .A2(new_n33607_), .B(new_n37832_), .ZN(new_n37833_));
  XNOR2_X1   g34507(.A1(new_n37833_), .A2(new_n37227_), .ZN(new_n37834_));
  NOR2_X1    g34508(.A1(new_n37575_), .A2(pi0454), .ZN(new_n37835_));
  AOI21_X1   g34509(.A1(new_n37835_), .A2(new_n10169_), .B(new_n37717_), .ZN(new_n37836_));
  AOI21_X1   g34510(.A1(new_n37834_), .A2(pi1043), .B(new_n37836_), .ZN(new_n37837_));
  NAND2_X1   g34511(.A1(pi0349), .A2(pi0588), .ZN(new_n37838_));
  OAI21_X1   g34512(.A1(new_n37721_), .A2(new_n37838_), .B(new_n6933_), .ZN(new_n37839_));
  NAND3_X1   g34513(.A1(new_n37576_), .A2(pi0329), .A3(new_n37202_), .ZN(new_n37840_));
  NOR2_X1    g34514(.A1(new_n37725_), .A2(pi0440), .ZN(new_n37841_));
  AOI21_X1   g34515(.A1(new_n37840_), .A2(new_n37841_), .B(new_n37226_), .ZN(new_n37842_));
  NAND2_X1   g34516(.A1(new_n37842_), .A2(new_n37839_), .ZN(new_n37843_));
  AOI21_X1   g34517(.A1(new_n37831_), .A2(new_n37837_), .B(new_n37843_), .ZN(po0873));
  INV_X1     g34518(.I(pi0462), .ZN(new_n37845_));
  NAND3_X1   g34519(.A1(pi0318), .A2(pi0591), .A3(pi0592), .ZN(new_n37846_));
  NOR3_X1    g34520(.A1(new_n6358_), .A2(pi0377), .A3(pi0591), .ZN(new_n37847_));
  XOR2_X1    g34521(.A1(new_n37847_), .A2(new_n37846_), .Z(new_n37848_));
  NOR2_X1    g34522(.A1(new_n37848_), .A2(new_n37845_), .ZN(new_n37849_));
  NAND3_X1   g34523(.A1(new_n37698_), .A2(new_n9787_), .A3(new_n37202_), .ZN(new_n37850_));
  OAI21_X1   g34524(.A1(new_n37850_), .A2(new_n37849_), .B(new_n7250_), .ZN(new_n37851_));
  NOR2_X1    g34525(.A1(new_n4785_), .A2(pi0645), .ZN(new_n37852_));
  XOR2_X1    g34526(.A1(new_n37209_), .A2(new_n37852_), .Z(new_n37853_));
  NOR2_X1    g34527(.A1(new_n37275_), .A2(new_n37323_), .ZN(new_n37854_));
  AOI21_X1   g34528(.A1(new_n37854_), .A2(new_n37853_), .B(pi0800), .ZN(new_n37855_));
  OAI21_X1   g34529(.A1(pi0839), .A2(pi1136), .B(pi1134), .ZN(new_n37856_));
  NAND2_X1   g34530(.A1(new_n37765_), .A2(new_n37856_), .ZN(new_n37857_));
  NAND4_X1   g34531(.A1(new_n37857_), .A2(pi0705), .A3(pi1135), .A4(new_n37251_), .ZN(new_n37858_));
  OAI21_X1   g34532(.A1(new_n37858_), .A2(new_n37855_), .B(new_n17881_), .ZN(new_n37859_));
  NAND2_X1   g34533(.A1(new_n33993_), .A2(pi0199), .ZN(new_n37860_));
  XOR2_X1    g34534(.A1(new_n37860_), .A2(new_n37227_), .Z(new_n37861_));
  NOR2_X1    g34535(.A1(pi0448), .A2(pi0588), .ZN(new_n37862_));
  OAI21_X1   g34536(.A1(new_n37861_), .A2(new_n35289_), .B(new_n37862_), .ZN(new_n37863_));
  NOR4_X1    g34537(.A1(new_n37468_), .A2(new_n10169_), .A3(new_n37226_), .A4(new_n37274_), .ZN(new_n37864_));
  NAND3_X1   g34538(.A1(new_n37863_), .A2(new_n37859_), .A3(new_n37864_), .ZN(new_n37865_));
  XOR2_X1    g34539(.A1(new_n37865_), .A2(new_n37851_), .Z(po0874));
  NOR2_X1    g34540(.A1(new_n4959_), .A2(pi0608), .ZN(new_n37867_));
  XOR2_X1    g34541(.A1(new_n37867_), .A2(new_n37338_), .Z(new_n37868_));
  NOR3_X1    g34542(.A1(new_n37868_), .A2(new_n13613_), .A3(new_n37358_), .ZN(new_n37869_));
  OR2_X2     g34543(.A1(pi0853), .A2(pi1136), .Z(new_n37870_));
  AOI21_X1   g34544(.A1(pi1134), .A2(new_n37870_), .B(new_n37708_), .ZN(new_n37871_));
  NAND2_X1   g34545(.A1(pi0698), .A2(pi1135), .ZN(new_n37872_));
  NOR4_X1    g34546(.A1(new_n37869_), .A2(new_n7250_), .A3(new_n37871_), .A4(new_n37872_), .ZN(new_n37873_));
  OAI21_X1   g34547(.A1(new_n37873_), .A2(pi0767), .B(new_n37221_), .ZN(new_n37874_));
  AOI21_X1   g34548(.A1(new_n8555_), .A2(pi0303), .B(new_n8549_), .ZN(new_n37875_));
  OAI21_X1   g34549(.A1(new_n8555_), .A2(new_n35178_), .B(new_n37875_), .ZN(new_n37876_));
  XNOR2_X1   g34550(.A1(new_n37876_), .A2(new_n37227_), .ZN(new_n37877_));
  NOR2_X1    g34551(.A1(new_n37575_), .A2(pi0419), .ZN(new_n37878_));
  AOI21_X1   g34552(.A1(new_n37878_), .A2(new_n10169_), .B(new_n37717_), .ZN(new_n37879_));
  AOI21_X1   g34553(.A1(new_n37877_), .A2(pi1080), .B(new_n37879_), .ZN(new_n37880_));
  NAND2_X1   g34554(.A1(pi0315), .A2(pi0588), .ZN(new_n37881_));
  OAI21_X1   g34555(.A1(new_n37721_), .A2(new_n37881_), .B(new_n6933_), .ZN(new_n37882_));
  NAND3_X1   g34556(.A1(new_n37576_), .A2(pi0394), .A3(new_n37202_), .ZN(new_n37883_));
  NOR2_X1    g34557(.A1(new_n37725_), .A2(pi0369), .ZN(new_n37884_));
  AOI21_X1   g34558(.A1(new_n37883_), .A2(new_n37884_), .B(new_n37226_), .ZN(new_n37885_));
  NAND2_X1   g34559(.A1(new_n37885_), .A2(new_n37882_), .ZN(new_n37886_));
  AOI21_X1   g34560(.A1(new_n37874_), .A2(new_n37880_), .B(new_n37886_), .ZN(po0875));
  NAND3_X1   g34561(.A1(pi0325), .A2(pi0591), .A3(pi0592), .ZN(new_n37888_));
  NOR3_X1    g34562(.A1(new_n6358_), .A2(pi0378), .A3(pi0591), .ZN(new_n37889_));
  XOR2_X1    g34563(.A1(new_n37889_), .A2(new_n37888_), .Z(new_n37890_));
  NOR2_X1    g34564(.A1(new_n37890_), .A2(new_n6654_), .ZN(new_n37891_));
  OAI21_X1   g34565(.A1(new_n37850_), .A2(new_n37891_), .B(new_n7250_), .ZN(new_n37892_));
  NOR2_X1    g34566(.A1(new_n4785_), .A2(pi0636), .ZN(new_n37893_));
  XOR2_X1    g34567(.A1(new_n37209_), .A2(new_n37893_), .Z(new_n37894_));
  NOR2_X1    g34568(.A1(new_n37275_), .A2(new_n37138_), .ZN(new_n37895_));
  AOI21_X1   g34569(.A1(new_n37895_), .A2(new_n37894_), .B(pi0807), .ZN(new_n37896_));
  OAI21_X1   g34570(.A1(pi0868), .A2(pi1136), .B(pi1134), .ZN(new_n37897_));
  NAND2_X1   g34571(.A1(new_n37765_), .A2(new_n37897_), .ZN(new_n37898_));
  NAND4_X1   g34572(.A1(new_n37898_), .A2(pi0687), .A3(pi1135), .A4(new_n37251_), .ZN(new_n37899_));
  OAI21_X1   g34573(.A1(new_n37899_), .A2(new_n37896_), .B(new_n15573_), .ZN(new_n37900_));
  NAND2_X1   g34574(.A1(new_n34005_), .A2(pi0199), .ZN(new_n37901_));
  XOR2_X1    g34575(.A1(new_n37901_), .A2(new_n37227_), .Z(new_n37902_));
  NOR2_X1    g34576(.A1(pi0451), .A2(pi0588), .ZN(new_n37903_));
  OAI21_X1   g34577(.A1(new_n37902_), .A2(new_n35309_), .B(new_n37903_), .ZN(new_n37904_));
  NAND3_X1   g34578(.A1(new_n37900_), .A2(new_n37904_), .A3(new_n37864_), .ZN(new_n37905_));
  XOR2_X1    g34579(.A1(new_n37905_), .A2(new_n37892_), .Z(po0876));
  NOR2_X1    g34580(.A1(new_n4785_), .A2(pi0684), .ZN(new_n37907_));
  XOR2_X1    g34581(.A1(new_n37209_), .A2(new_n37907_), .Z(new_n37908_));
  INV_X1     g34582(.I(pi0750), .ZN(new_n37909_));
  NOR2_X1    g34583(.A1(new_n37215_), .A2(new_n37909_), .ZN(new_n37910_));
  AOI21_X1   g34584(.A1(new_n37910_), .A2(new_n37908_), .B(pi0880), .ZN(new_n37911_));
  OAI21_X1   g34585(.A1(new_n37911_), .A2(new_n37252_), .B(new_n7250_), .ZN(new_n37912_));
  NAND3_X1   g34586(.A1(pi0356), .A2(pi0590), .A3(pi0592), .ZN(new_n37913_));
  NAND3_X1   g34587(.A1(new_n6678_), .A2(new_n6933_), .A3(pi0592), .ZN(new_n37914_));
  XOR2_X1    g34588(.A1(new_n37914_), .A2(new_n37913_), .Z(new_n37915_));
  NAND2_X1   g34589(.A1(pi0405), .A2(pi0588), .ZN(new_n37916_));
  OAI21_X1   g34590(.A1(new_n37563_), .A2(new_n37916_), .B(new_n6350_), .ZN(new_n37917_));
  NOR4_X1    g34591(.A1(new_n8549_), .A2(new_n35401_), .A3(pi0223), .A4(pi0224), .ZN(new_n37918_));
  AOI21_X1   g34592(.A1(new_n37917_), .A2(new_n37915_), .B(new_n37918_), .ZN(new_n37919_));
  NOR3_X1    g34593(.A1(new_n37142_), .A2(new_n4959_), .A3(new_n4785_), .ZN(new_n37920_));
  NOR3_X1    g34594(.A1(new_n4785_), .A2(pi0651), .A3(pi1135), .ZN(new_n37921_));
  OAI21_X1   g34595(.A1(new_n37920_), .A2(new_n37921_), .B(pi0654), .ZN(new_n37922_));
  NOR2_X1    g34596(.A1(new_n37212_), .A2(pi0794), .ZN(new_n37923_));
  NAND2_X1   g34597(.A1(new_n37922_), .A2(new_n37923_), .ZN(new_n37924_));
  AOI21_X1   g34598(.A1(new_n37924_), .A2(new_n37251_), .B(pi1134), .ZN(new_n37925_));
  NAND2_X1   g34599(.A1(new_n7250_), .A2(pi0445), .ZN(new_n37926_));
  NOR4_X1    g34600(.A1(new_n37919_), .A2(new_n37579_), .A3(new_n37925_), .A4(new_n37926_), .ZN(new_n37927_));
  XNOR2_X1   g34601(.A1(new_n37927_), .A2(new_n37912_), .ZN(po0877));
  INV_X1     g34602(.I(pi0794), .ZN(new_n37929_));
  INV_X1     g34603(.I(pi0721), .ZN(new_n37930_));
  INV_X1     g34604(.I(pi0813), .ZN(new_n37931_));
  NOR2_X1    g34605(.A1(new_n37930_), .A2(new_n37931_), .ZN(new_n37932_));
  INV_X1     g34606(.I(new_n37932_), .ZN(new_n37933_));
  NOR3_X1    g34607(.A1(new_n37933_), .A2(new_n37929_), .A3(new_n37631_), .ZN(new_n37934_));
  XNOR2_X1   g34608(.A1(pi0771), .A2(pi0800), .ZN(new_n37935_));
  INV_X1     g34609(.I(pi0807), .ZN(new_n37936_));
  XOR2_X1    g34610(.A1(pi0765), .A2(pi0798), .Z(new_n37937_));
  NOR2_X1    g34611(.A1(new_n37937_), .A2(new_n37936_), .ZN(new_n37938_));
  INV_X1     g34612(.I(pi0747), .ZN(new_n37939_));
  XNOR2_X1   g34613(.A1(pi0765), .A2(pi0798), .ZN(new_n37940_));
  NOR3_X1    g34614(.A1(new_n37940_), .A2(new_n37939_), .A3(new_n37936_), .ZN(new_n37941_));
  AOI21_X1   g34615(.A1(pi0747), .A2(new_n37938_), .B(new_n37941_), .ZN(new_n37942_));
  INV_X1     g34616(.I(pi0769), .ZN(new_n37943_));
  NAND2_X1   g34617(.A1(new_n37943_), .A2(new_n37929_), .ZN(new_n37944_));
  NAND2_X1   g34618(.A1(pi0769), .A2(pi0794), .ZN(new_n37945_));
  AOI21_X1   g34619(.A1(new_n37944_), .A2(new_n37945_), .B(new_n37942_), .ZN(new_n37946_));
  NAND2_X1   g34620(.A1(new_n37946_), .A2(new_n37935_), .ZN(new_n37947_));
  INV_X1     g34621(.I(pi0773), .ZN(new_n37948_));
  NOR2_X1    g34622(.A1(new_n37948_), .A2(new_n37631_), .ZN(new_n37949_));
  NOR2_X1    g34623(.A1(pi0773), .A2(pi0801), .ZN(new_n37950_));
  NOR2_X1    g34624(.A1(new_n37949_), .A2(new_n37950_), .ZN(new_n37951_));
  NOR2_X1    g34625(.A1(new_n37947_), .A2(new_n37951_), .ZN(new_n37952_));
  INV_X1     g34626(.I(new_n37952_), .ZN(new_n37953_));
  NOR2_X1    g34627(.A1(new_n37953_), .A2(new_n37933_), .ZN(new_n37954_));
  INV_X1     g34628(.I(new_n37954_), .ZN(new_n37955_));
  NOR2_X1    g34629(.A1(new_n37955_), .A2(new_n37814_), .ZN(new_n37956_));
  INV_X1     g34630(.I(new_n37935_), .ZN(new_n37957_));
  INV_X1     g34631(.I(new_n37938_), .ZN(new_n37958_));
  NOR2_X1    g34632(.A1(new_n37958_), .A2(new_n37957_), .ZN(new_n37959_));
  INV_X1     g34633(.I(new_n37959_), .ZN(new_n37960_));
  NOR2_X1    g34634(.A1(new_n37939_), .A2(new_n37948_), .ZN(new_n37961_));
  INV_X1     g34635(.I(pi0775), .ZN(new_n37962_));
  NOR3_X1    g34636(.A1(new_n37930_), .A2(new_n37962_), .A3(pi0769), .ZN(new_n37963_));
  AOI21_X1   g34637(.A1(pi0721), .A2(pi0775), .B(new_n37943_), .ZN(new_n37964_));
  OAI21_X1   g34638(.A1(new_n37964_), .A2(new_n37963_), .B(new_n37961_), .ZN(new_n37965_));
  INV_X1     g34639(.I(pi0731), .ZN(new_n37966_));
  INV_X1     g34640(.I(pi0945), .ZN(new_n37967_));
  NAND2_X1   g34641(.A1(new_n37967_), .A2(pi0988), .ZN(new_n37968_));
  NOR2_X1    g34642(.A1(new_n37968_), .A2(new_n37966_), .ZN(new_n37969_));
  INV_X1     g34643(.I(new_n37969_), .ZN(new_n37970_));
  OAI21_X1   g34644(.A1(new_n37970_), .A2(new_n37965_), .B(new_n37930_), .ZN(new_n37971_));
  NAND3_X1   g34645(.A1(new_n37971_), .A2(pi0775), .A3(pi0795), .ZN(new_n37972_));
  AOI21_X1   g34646(.A1(new_n37972_), .A2(new_n37965_), .B(new_n37960_), .ZN(new_n37973_));
  OAI21_X1   g34647(.A1(new_n37956_), .A2(new_n37934_), .B(new_n37973_), .ZN(new_n37974_));
  NOR2_X1    g34648(.A1(new_n37962_), .A2(new_n37814_), .ZN(new_n37975_));
  INV_X1     g34649(.I(new_n37975_), .ZN(new_n37976_));
  NOR2_X1    g34650(.A1(pi0775), .A2(pi0816), .ZN(new_n37977_));
  INV_X1     g34651(.I(new_n37977_), .ZN(new_n37978_));
  AOI21_X1   g34652(.A1(new_n37976_), .A2(new_n37978_), .B(new_n37955_), .ZN(new_n37979_));
  XNOR2_X1   g34653(.A1(pi0731), .A2(pi0795), .ZN(new_n37980_));
  AOI21_X1   g34654(.A1(new_n37970_), .A2(new_n37930_), .B(new_n37980_), .ZN(new_n37981_));
  NAND2_X1   g34655(.A1(new_n37979_), .A2(new_n37981_), .ZN(new_n37982_));
  OR3_X2     g34656(.A1(new_n37979_), .A2(new_n37930_), .A3(pi0775), .Z(new_n37983_));
  NAND3_X1   g34657(.A1(new_n37983_), .A2(new_n37982_), .A3(new_n37974_), .ZN(po0878));
  NAND3_X1   g34658(.A1(pi0640), .A2(pi1134), .A3(pi1136), .ZN(new_n37985_));
  NAND3_X1   g34659(.A1(new_n37099_), .A2(new_n5132_), .A3(pi1136), .ZN(new_n37986_));
  NAND2_X1   g34660(.A1(new_n37986_), .A2(new_n37985_), .ZN(new_n37987_));
  NAND3_X1   g34661(.A1(new_n37209_), .A2(pi0694), .A3(pi1134), .ZN(new_n37988_));
  NAND3_X1   g34662(.A1(new_n37209_), .A2(new_n37641_), .A3(new_n5132_), .ZN(new_n37989_));
  NAND2_X1   g34663(.A1(new_n37988_), .A2(new_n37989_), .ZN(new_n37990_));
  INV_X1     g34664(.I(pi0732), .ZN(new_n37991_));
  NOR2_X1    g34665(.A1(new_n37991_), .A2(new_n4959_), .ZN(new_n37992_));
  AOI22_X1   g34666(.A1(new_n37990_), .A2(new_n37992_), .B1(pi0776), .B2(new_n37987_), .ZN(new_n37993_));
  INV_X1     g34667(.I(pi0795), .ZN(new_n37994_));
  NOR3_X1    g34668(.A1(new_n37994_), .A2(new_n5132_), .A3(new_n4785_), .ZN(new_n37995_));
  NOR3_X1    g34669(.A1(new_n5132_), .A2(pi0795), .A3(pi1136), .ZN(new_n37996_));
  OAI21_X1   g34670(.A1(new_n37995_), .A2(new_n37996_), .B(pi0851), .ZN(new_n37997_));
  OAI21_X1   g34671(.A1(new_n37993_), .A2(new_n37997_), .B(new_n7250_), .ZN(new_n37998_));
  AOI21_X1   g34672(.A1(new_n3090_), .A2(new_n3100_), .B(pi0588), .ZN(new_n38003_));
  NAND3_X1   g34673(.A1(pi0379), .A2(pi0591), .A3(pi0592), .ZN(new_n38004_));
  NOR3_X1    g34674(.A1(new_n6350_), .A2(pi0403), .A3(pi0592), .ZN(new_n38005_));
  XNOR2_X1   g34675(.A1(new_n38005_), .A2(new_n38004_), .ZN(new_n38006_));
  AOI21_X1   g34676(.A1(new_n38006_), .A2(pi0354), .B(new_n37697_), .ZN(new_n38007_));
  NOR4_X1    g34677(.A1(new_n38007_), .A2(new_n10169_), .A3(new_n37213_), .A4(new_n38003_), .ZN(new_n38008_));
  XNOR2_X1   g34678(.A1(new_n38008_), .A2(new_n37998_), .ZN(po0879));
  NAND3_X1   g34679(.A1(po0980), .A2(pi0962), .A3(pi1111), .ZN(new_n38010_));
  NAND3_X1   g34680(.A1(po0980), .A2(new_n37045_), .A3(new_n36981_), .ZN(new_n38011_));
  AOI21_X1   g34681(.A1(new_n38010_), .A2(new_n38011_), .B(new_n17227_), .ZN(po0880));
  NAND3_X1   g34682(.A1(po0980), .A2(pi0962), .A3(pi1114), .ZN(new_n38013_));
  NAND3_X1   g34683(.A1(po0980), .A2(new_n37045_), .A3(new_n36977_), .ZN(new_n38014_));
  AOI21_X1   g34684(.A1(new_n38013_), .A2(new_n38014_), .B(new_n17474_), .ZN(po0881));
  NAND3_X1   g34685(.A1(po0980), .A2(pi0962), .A3(pi1120), .ZN(new_n38016_));
  NAND3_X1   g34686(.A1(po0980), .A2(new_n37045_), .A3(new_n37063_), .ZN(new_n38017_));
  AOI21_X1   g34687(.A1(new_n38016_), .A2(new_n38017_), .B(new_n17148_), .ZN(po0882));
  NAND3_X1   g34688(.A1(po0980), .A2(pi0962), .A3(pi1126), .ZN(new_n38019_));
  NAND3_X1   g34689(.A1(po0980), .A2(new_n37045_), .A3(new_n37135_), .ZN(new_n38020_));
  AOI21_X1   g34690(.A1(new_n38019_), .A2(new_n38020_), .B(new_n16962_), .ZN(po0883));
  NAND3_X1   g34691(.A1(po0980), .A2(pi0962), .A3(pi1102), .ZN(new_n38022_));
  NAND3_X1   g34692(.A1(po0980), .A2(new_n37045_), .A3(new_n37195_), .ZN(new_n38023_));
  AOI21_X1   g34693(.A1(new_n38022_), .A2(new_n38023_), .B(new_n17866_), .ZN(po0884));
  INV_X1     g34694(.I(pi0728), .ZN(new_n38025_));
  NAND3_X1   g34695(.A1(po0980), .A2(pi0962), .A3(pi1131), .ZN(new_n38026_));
  NAND3_X1   g34696(.A1(po0980), .A2(new_n37045_), .A3(new_n37149_), .ZN(new_n38027_));
  AOI21_X1   g34697(.A1(new_n38026_), .A2(new_n38027_), .B(new_n38025_), .ZN(po0885));
  NAND3_X1   g34698(.A1(po0980), .A2(pi0962), .A3(pi1104), .ZN(new_n38029_));
  NAND3_X1   g34699(.A1(po0980), .A2(new_n37045_), .A3(new_n36951_), .ZN(new_n38030_));
  AOI21_X1   g34700(.A1(new_n38029_), .A2(new_n38030_), .B(new_n17987_), .ZN(po0886));
  NAND3_X1   g34701(.A1(po0980), .A2(pi0962), .A3(pi1106), .ZN(new_n38032_));
  NAND3_X1   g34702(.A1(po0980), .A2(new_n37045_), .A3(new_n37029_), .ZN(new_n38033_));
  AOI21_X1   g34703(.A1(new_n38032_), .A2(new_n38033_), .B(new_n18025_), .ZN(po0887));
  INV_X1     g34704(.I(new_n37961_), .ZN(new_n38035_));
  NOR2_X1    g34705(.A1(pi0721), .A2(pi0813), .ZN(new_n38036_));
  OAI21_X1   g34706(.A1(new_n37932_), .A2(new_n38036_), .B(new_n37952_), .ZN(new_n38037_));
  XOR2_X1    g34707(.A1(new_n38037_), .A2(new_n37994_), .Z(new_n38038_));
  NAND2_X1   g34708(.A1(new_n38038_), .A2(new_n37975_), .ZN(new_n38039_));
  XOR2_X1    g34709(.A1(pi0769), .A2(pi0801), .Z(new_n38040_));
  NAND3_X1   g34710(.A1(new_n38040_), .A2(pi0794), .A3(pi0795), .ZN(new_n38041_));
  XNOR2_X1   g34711(.A1(pi0775), .A2(pi0816), .ZN(new_n38042_));
  XNOR2_X1   g34712(.A1(pi0721), .A2(pi0813), .ZN(new_n38043_));
  NOR2_X1    g34713(.A1(new_n38042_), .A2(new_n38043_), .ZN(new_n38044_));
  INV_X1     g34714(.I(new_n38044_), .ZN(new_n38045_));
  NAND3_X1   g34715(.A1(new_n38045_), .A2(new_n38041_), .A3(new_n38035_), .ZN(new_n38046_));
  NAND2_X1   g34716(.A1(new_n38046_), .A2(new_n37959_), .ZN(new_n38047_));
  INV_X1     g34717(.I(new_n37968_), .ZN(new_n38048_));
  AOI21_X1   g34718(.A1(new_n38046_), .A2(new_n37959_), .B(new_n38048_), .ZN(new_n38049_));
  OAI22_X1   g34719(.A1(new_n38039_), .A2(new_n38049_), .B1(new_n37966_), .B2(new_n38047_), .ZN(new_n38050_));
  NAND2_X1   g34720(.A1(new_n38050_), .A2(new_n37969_), .ZN(new_n38051_));
  AOI21_X1   g34721(.A1(new_n38051_), .A2(new_n38035_), .B(new_n38039_), .ZN(po0888));
  NAND3_X1   g34722(.A1(po0954), .A2(pi0962), .A3(pi1128), .ZN(new_n38053_));
  NAND3_X1   g34723(.A1(po0954), .A2(new_n37045_), .A3(new_n37101_), .ZN(new_n38054_));
  AOI21_X1   g34724(.A1(new_n38053_), .A2(new_n38054_), .B(new_n37991_), .ZN(po0889));
  NOR2_X1    g34725(.A1(new_n4959_), .A2(pi0619), .ZN(new_n38056_));
  XOR2_X1    g34726(.A1(new_n38056_), .A2(new_n37338_), .Z(new_n38057_));
  NOR3_X1    g34727(.A1(new_n38057_), .A2(new_n13884_), .A3(new_n37358_), .ZN(new_n38058_));
  OR2_X2     g34728(.A1(pi0838), .A2(pi1136), .Z(new_n38059_));
  AOI21_X1   g34729(.A1(pi1134), .A2(new_n38059_), .B(new_n37708_), .ZN(new_n38060_));
  NAND2_X1   g34730(.A1(pi0737), .A2(pi1135), .ZN(new_n38061_));
  NOR4_X1    g34731(.A1(new_n38058_), .A2(new_n7250_), .A3(new_n38060_), .A4(new_n38061_), .ZN(new_n38062_));
  OAI21_X1   g34732(.A1(new_n38062_), .A2(pi0777), .B(new_n37221_), .ZN(new_n38063_));
  AOI21_X1   g34733(.A1(new_n8555_), .A2(pi0308), .B(new_n8549_), .ZN(new_n38064_));
  OAI21_X1   g34734(.A1(new_n8555_), .A2(new_n34021_), .B(new_n38064_), .ZN(new_n38065_));
  XNOR2_X1   g34735(.A1(new_n38065_), .A2(new_n37227_), .ZN(new_n38066_));
  NOR2_X1    g34736(.A1(new_n37575_), .A2(pi0424), .ZN(new_n38067_));
  AOI21_X1   g34737(.A1(new_n38067_), .A2(new_n10169_), .B(new_n37717_), .ZN(new_n38068_));
  AOI21_X1   g34738(.A1(new_n38066_), .A2(pi1047), .B(new_n38068_), .ZN(new_n38069_));
  NAND2_X1   g34739(.A1(pi0316), .A2(pi0588), .ZN(new_n38070_));
  OAI21_X1   g34740(.A1(new_n37721_), .A2(new_n38070_), .B(new_n6933_), .ZN(new_n38071_));
  NAND3_X1   g34741(.A1(new_n37576_), .A2(pi0399), .A3(new_n37202_), .ZN(new_n38072_));
  NOR2_X1    g34742(.A1(new_n37725_), .A2(pi0375), .ZN(new_n38073_));
  AOI21_X1   g34743(.A1(new_n38072_), .A2(new_n38073_), .B(new_n37226_), .ZN(new_n38074_));
  NAND2_X1   g34744(.A1(new_n38074_), .A2(new_n38071_), .ZN(new_n38075_));
  AOI21_X1   g34745(.A1(new_n38063_), .A2(new_n38069_), .B(new_n38075_), .ZN(po0890));
  NAND3_X1   g34746(.A1(po0980), .A2(pi0962), .A3(pi1119), .ZN(new_n38077_));
  NAND3_X1   g34747(.A1(po0980), .A2(new_n37045_), .A3(new_n37056_), .ZN(new_n38078_));
  AOI21_X1   g34748(.A1(new_n38077_), .A2(new_n38078_), .B(new_n17604_), .ZN(po0891));
  NAND3_X1   g34749(.A1(po0980), .A2(pi0962), .A3(pi1109), .ZN(new_n38080_));
  NAND3_X1   g34750(.A1(po0980), .A2(new_n37045_), .A3(new_n37025_), .ZN(new_n38081_));
  AOI21_X1   g34751(.A1(new_n38080_), .A2(new_n38081_), .B(new_n14833_), .ZN(po0892));
  NAND3_X1   g34752(.A1(po0980), .A2(pi0962), .A3(pi1101), .ZN(new_n38083_));
  NAND3_X1   g34753(.A1(po0980), .A2(new_n37045_), .A3(new_n37191_), .ZN(new_n38084_));
  AOI21_X1   g34754(.A1(new_n38083_), .A2(new_n38084_), .B(new_n16136_), .ZN(po0893));
  NAND3_X1   g34755(.A1(po0980), .A2(pi0962), .A3(pi1122), .ZN(new_n38086_));
  NAND3_X1   g34756(.A1(po0980), .A2(new_n37045_), .A3(new_n37012_), .ZN(new_n38087_));
  AOI21_X1   g34757(.A1(new_n38086_), .A2(new_n38087_), .B(new_n17730_), .ZN(po0894));
  NAND3_X1   g34758(.A1(po0980), .A2(pi0962), .A3(pi1121), .ZN(new_n38089_));
  NAND3_X1   g34759(.A1(po0980), .A2(new_n37045_), .A3(new_n37049_), .ZN(new_n38090_));
  AOI21_X1   g34760(.A1(new_n38089_), .A2(new_n38090_), .B(new_n13226_), .ZN(po0895));
  NOR3_X1    g34761(.A1(new_n36935_), .A2(pi0952), .A3(pi1061), .ZN(new_n38092_));
  NAND2_X1   g34762(.A1(new_n38092_), .A2(pi0832), .ZN(new_n38093_));
  INV_X1     g34763(.I(new_n38093_), .ZN(po0988));
  NAND3_X1   g34764(.A1(po0988), .A2(pi0966), .A3(pi1108), .ZN(new_n38095_));
  NAND3_X1   g34765(.A1(po0988), .A2(new_n36958_), .A3(new_n37021_), .ZN(new_n38096_));
  AOI21_X1   g34766(.A1(new_n38095_), .A2(new_n38096_), .B(new_n18095_), .ZN(po0896));
  NAND3_X1   g34767(.A1(po0988), .A2(pi0966), .A3(pi1114), .ZN(new_n38098_));
  NAND3_X1   g34768(.A1(po0988), .A2(new_n36958_), .A3(new_n36977_), .ZN(new_n38099_));
  AOI21_X1   g34769(.A1(new_n38098_), .A2(new_n38099_), .B(new_n17475_), .ZN(po0898));
  NAND3_X1   g34770(.A1(po0988), .A2(pi0966), .A3(pi1112), .ZN(new_n38101_));
  NAND3_X1   g34771(.A1(po0988), .A2(new_n36958_), .A3(new_n37017_), .ZN(new_n38102_));
  AOI21_X1   g34772(.A1(new_n38101_), .A2(new_n38102_), .B(new_n17409_), .ZN(po0899));
  NAND3_X1   g34773(.A1(po0988), .A2(pi0966), .A3(pi1109), .ZN(new_n38104_));
  NAND3_X1   g34774(.A1(po0988), .A2(new_n36958_), .A3(new_n37025_), .ZN(new_n38105_));
  AOI21_X1   g34775(.A1(new_n38104_), .A2(new_n38105_), .B(new_n14921_), .ZN(po0900));
  NAND3_X1   g34776(.A1(po0988), .A2(pi0966), .A3(pi1131), .ZN(new_n38107_));
  NAND3_X1   g34777(.A1(po0988), .A2(new_n36958_), .A3(new_n37149_), .ZN(new_n38108_));
  AOI21_X1   g34778(.A1(new_n38107_), .A2(new_n38108_), .B(new_n37555_), .ZN(po0901));
  NAND3_X1   g34779(.A1(po0988), .A2(pi0966), .A3(pi1111), .ZN(new_n38110_));
  NAND3_X1   g34780(.A1(po0988), .A2(new_n36958_), .A3(new_n36981_), .ZN(new_n38111_));
  AOI21_X1   g34781(.A1(new_n38110_), .A2(new_n38111_), .B(new_n18290_), .ZN(po0902));
  NAND3_X1   g34782(.A1(po0988), .A2(pi0966), .A3(pi1104), .ZN(new_n38113_));
  NAND3_X1   g34783(.A1(po0988), .A2(new_n36958_), .A3(new_n36951_), .ZN(new_n38114_));
  AOI21_X1   g34784(.A1(new_n38113_), .A2(new_n38114_), .B(new_n17956_), .ZN(po0903));
  INV_X1     g34785(.I(new_n37980_), .ZN(new_n38116_));
  NOR2_X1    g34786(.A1(new_n38045_), .A2(new_n38116_), .ZN(new_n38117_));
  XOR2_X1    g34787(.A1(new_n38117_), .A2(new_n37929_), .Z(new_n38118_));
  XOR2_X1    g34788(.A1(new_n37938_), .A2(pi0801), .Z(new_n38119_));
  OAI21_X1   g34789(.A1(pi0773), .A2(pi0801), .B(new_n38048_), .ZN(new_n38120_));
  NAND4_X1   g34790(.A1(new_n38119_), .A2(pi0769), .A3(new_n37957_), .A4(new_n38120_), .ZN(new_n38121_));
  OAI21_X1   g34791(.A1(new_n38118_), .A2(new_n38121_), .B(new_n37631_), .ZN(new_n38122_));
  NAND3_X1   g34792(.A1(new_n38122_), .A2(pi0747), .A3(new_n37941_), .ZN(new_n38123_));
  XOR2_X1    g34793(.A1(new_n38123_), .A2(pi0773), .Z(new_n38124_));
  NOR2_X1    g34794(.A1(new_n38124_), .A2(new_n37968_), .ZN(po0904));
  NAND3_X1   g34795(.A1(po0988), .A2(pi0966), .A3(pi1106), .ZN(new_n38126_));
  NAND3_X1   g34796(.A1(po0988), .A2(new_n36958_), .A3(new_n37029_), .ZN(new_n38127_));
  AOI21_X1   g34797(.A1(new_n38126_), .A2(new_n38127_), .B(new_n18000_), .ZN(po0905));
  NAND3_X1   g34798(.A1(po0988), .A2(pi0966), .A3(pi1105), .ZN(new_n38129_));
  NAND3_X1   g34799(.A1(po0988), .A2(new_n36958_), .A3(new_n37002_), .ZN(new_n38130_));
  AOI21_X1   g34800(.A1(new_n38129_), .A2(new_n38130_), .B(new_n14263_), .ZN(po0906));
  NAND3_X1   g34801(.A1(po0988), .A2(pi0966), .A3(pi1130), .ZN(new_n38132_));
  NAND3_X1   g34802(.A1(po0988), .A2(new_n36958_), .A3(new_n37144_), .ZN(new_n38133_));
  AOI21_X1   g34803(.A1(new_n38132_), .A2(new_n38133_), .B(new_n37909_), .ZN(po0907));
  NAND3_X1   g34804(.A1(po0988), .A2(pi0966), .A3(pi1123), .ZN(new_n38135_));
  NAND3_X1   g34805(.A1(po0988), .A2(new_n36958_), .A3(new_n37115_), .ZN(new_n38136_));
  AOI21_X1   g34806(.A1(new_n38135_), .A2(new_n38136_), .B(new_n17192_), .ZN(po0908));
  NAND3_X1   g34807(.A1(po0988), .A2(pi0966), .A3(pi1124), .ZN(new_n38138_));
  NAND3_X1   g34808(.A1(po0988), .A2(new_n36958_), .A3(new_n37163_), .ZN(new_n38139_));
  AOI21_X1   g34809(.A1(new_n38138_), .A2(new_n38139_), .B(new_n17769_), .ZN(po0909));
  NAND3_X1   g34810(.A1(po0988), .A2(pi0966), .A3(pi1117), .ZN(new_n38141_));
  NAND3_X1   g34811(.A1(po0988), .A2(new_n36958_), .A3(new_n37008_), .ZN(new_n38142_));
  AOI21_X1   g34812(.A1(new_n38141_), .A2(new_n38142_), .B(new_n17532_), .ZN(po0910));
  NAND3_X1   g34813(.A1(po0988), .A2(pi0966), .A3(pi1118), .ZN(new_n38144_));
  NAND3_X1   g34814(.A1(po0988), .A2(new_n36958_), .A3(new_n36967_), .ZN(new_n38145_));
  AOI21_X1   g34815(.A1(new_n38144_), .A2(new_n38145_), .B(new_n17569_), .ZN(po0911));
  NAND3_X1   g34816(.A1(po0988), .A2(pi0966), .A3(pi1120), .ZN(new_n38147_));
  NAND3_X1   g34817(.A1(po0988), .A2(new_n36958_), .A3(new_n37063_), .ZN(new_n38148_));
  AOI21_X1   g34818(.A1(new_n38147_), .A2(new_n38148_), .B(new_n17153_), .ZN(po0912));
  NAND3_X1   g34819(.A1(po0988), .A2(pi0966), .A3(pi1119), .ZN(new_n38150_));
  NAND3_X1   g34820(.A1(po0988), .A2(new_n36958_), .A3(new_n37056_), .ZN(new_n38151_));
  AOI21_X1   g34821(.A1(new_n38150_), .A2(new_n38151_), .B(new_n17609_), .ZN(po0913));
  NAND3_X1   g34822(.A1(po0988), .A2(pi0966), .A3(pi1113), .ZN(new_n38153_));
  NAND3_X1   g34823(.A1(po0988), .A2(new_n36958_), .A3(new_n36972_), .ZN(new_n38154_));
  AOI21_X1   g34824(.A1(new_n38153_), .A2(new_n38154_), .B(new_n17446_), .ZN(po0914));
  NAND3_X1   g34825(.A1(po0988), .A2(pi0966), .A3(pi1101), .ZN(new_n38156_));
  NAND3_X1   g34826(.A1(po0988), .A2(new_n36958_), .A3(new_n37191_), .ZN(new_n38157_));
  AOI21_X1   g34827(.A1(new_n38156_), .A2(new_n38157_), .B(new_n16090_), .ZN(po0915));
  NAND3_X1   g34828(.A1(new_n38092_), .A2(pi0966), .A3(new_n36937_), .ZN(new_n38159_));
  AOI21_X1   g34829(.A1(new_n38159_), .A2(new_n17309_), .B(new_n38093_), .ZN(po0916));
  NAND3_X1   g34830(.A1(po0988), .A2(pi0966), .A3(pi1115), .ZN(new_n38161_));
  NAND3_X1   g34831(.A1(po0988), .A2(new_n36958_), .A3(new_n36986_), .ZN(new_n38162_));
  AOI21_X1   g34832(.A1(new_n38161_), .A2(new_n38162_), .B(new_n17500_), .ZN(po0917));
  NAND3_X1   g34833(.A1(po0988), .A2(pi0966), .A3(pi1121), .ZN(new_n38164_));
  NAND3_X1   g34834(.A1(po0988), .A2(new_n36958_), .A3(new_n37049_), .ZN(new_n38165_));
  AOI21_X1   g34835(.A1(new_n38164_), .A2(new_n38165_), .B(new_n13099_), .ZN(po0918));
  NAND3_X1   g34836(.A1(po0988), .A2(pi0966), .A3(pi1129), .ZN(new_n38167_));
  NAND3_X1   g34837(.A1(po0988), .A2(new_n36958_), .A3(new_n37154_), .ZN(new_n38168_));
  AOI21_X1   g34838(.A1(new_n38167_), .A2(new_n38168_), .B(new_n37800_), .ZN(po0919));
  NAND3_X1   g34839(.A1(po0988), .A2(pi0966), .A3(pi1103), .ZN(new_n38170_));
  NAND3_X1   g34840(.A1(po0988), .A2(new_n36958_), .A3(new_n37108_), .ZN(new_n38171_));
  AOI21_X1   g34841(.A1(new_n38170_), .A2(new_n38171_), .B(new_n17912_), .ZN(po0920));
  NAND3_X1   g34842(.A1(po0988), .A2(pi0966), .A3(pi1107), .ZN(new_n38173_));
  NAND3_X1   g34843(.A1(po0988), .A2(new_n36958_), .A3(new_n36959_), .ZN(new_n38174_));
  AOI21_X1   g34844(.A1(new_n38173_), .A2(new_n38174_), .B(new_n18051_), .ZN(po0921));
  NAND2_X1   g34845(.A1(new_n37952_), .A2(new_n38117_), .ZN(new_n38176_));
  INV_X1     g34846(.I(new_n38176_), .ZN(po0978));
  NOR2_X1    g34847(.A1(po0978), .A2(new_n37967_), .ZN(new_n38178_));
  INV_X1     g34848(.I(pi0765), .ZN(new_n38179_));
  XOR2_X1    g34849(.A1(new_n37947_), .A2(new_n37631_), .Z(new_n38180_));
  INV_X1     g34850(.I(pi0771), .ZN(new_n38181_));
  INV_X1     g34851(.I(pi0800), .ZN(new_n38182_));
  NOR2_X1    g34852(.A1(new_n38181_), .A2(new_n38182_), .ZN(new_n38183_));
  OAI22_X1   g34853(.A1(new_n37958_), .A2(new_n37939_), .B1(pi0765), .B2(new_n38183_), .ZN(new_n38184_));
  NOR2_X1    g34854(.A1(new_n37950_), .A2(new_n37945_), .ZN(new_n38185_));
  NAND2_X1   g34855(.A1(new_n38184_), .A2(new_n38185_), .ZN(new_n38186_));
  NAND4_X1   g34856(.A1(new_n38180_), .A2(pi0721), .A3(new_n37978_), .A4(new_n38186_), .ZN(new_n38187_));
  XOR2_X1    g34857(.A1(new_n38187_), .A2(new_n37931_), .Z(new_n38188_));
  INV_X1     g34858(.I(new_n38037_), .ZN(new_n38189_));
  OAI21_X1   g34859(.A1(pi0765), .A2(new_n37978_), .B(new_n38189_), .ZN(new_n38190_));
  NAND2_X1   g34860(.A1(pi0731), .A2(pi0795), .ZN(new_n38191_));
  OAI21_X1   g34861(.A1(new_n37953_), .A2(new_n38036_), .B(pi0795), .ZN(new_n38192_));
  AOI21_X1   g34862(.A1(new_n38190_), .A2(new_n38191_), .B(new_n38192_), .ZN(new_n38193_));
  AOI21_X1   g34863(.A1(new_n38179_), .A2(new_n37994_), .B(new_n37966_), .ZN(new_n38194_));
  AOI22_X1   g34864(.A1(new_n38188_), .A2(new_n38193_), .B1(new_n38039_), .B2(new_n38194_), .ZN(new_n38195_));
  NOR3_X1    g34865(.A1(new_n38195_), .A2(new_n38179_), .A3(new_n37967_), .ZN(new_n38196_));
  XOR2_X1    g34866(.A1(new_n38196_), .A2(new_n38178_), .Z(po0922));
  NAND3_X1   g34867(.A1(po0988), .A2(pi0966), .A3(pi1110), .ZN(new_n38198_));
  NAND3_X1   g34868(.A1(po0988), .A2(new_n36958_), .A3(new_n37075_), .ZN(new_n38199_));
  AOI21_X1   g34869(.A1(new_n38198_), .A2(new_n38199_), .B(new_n17355_), .ZN(po0923));
  NAND3_X1   g34870(.A1(po0988), .A2(pi0966), .A3(pi1116), .ZN(new_n38201_));
  NAND3_X1   g34871(.A1(po0988), .A2(new_n36958_), .A3(new_n36963_), .ZN(new_n38202_));
  AOI21_X1   g34872(.A1(new_n38201_), .A2(new_n38202_), .B(new_n16517_), .ZN(po0924));
  NAND3_X1   g34873(.A1(po0988), .A2(pi0966), .A3(pi1125), .ZN(new_n38204_));
  NAND3_X1   g34874(.A1(po0988), .A2(new_n36958_), .A3(new_n37120_), .ZN(new_n38205_));
  AOI21_X1   g34875(.A1(new_n38204_), .A2(new_n38205_), .B(new_n17881_), .ZN(po0925));
  NAND2_X1   g34876(.A1(new_n38037_), .A2(pi0775), .ZN(new_n38207_));
  XOR2_X1    g34877(.A1(pi0794), .A2(pi0801), .Z(new_n38208_));
  NAND4_X1   g34878(.A1(new_n38044_), .A2(pi0773), .A3(new_n37957_), .A4(new_n38208_), .ZN(new_n38209_));
  NOR2_X1    g34879(.A1(new_n37942_), .A2(new_n38209_), .ZN(new_n38210_));
  NAND2_X1   g34880(.A1(new_n38210_), .A2(new_n37975_), .ZN(new_n38211_));
  XNOR2_X1   g34881(.A1(new_n38207_), .A2(new_n38211_), .ZN(new_n38212_));
  NAND2_X1   g34882(.A1(new_n37969_), .A2(pi0769), .ZN(new_n38213_));
  XOR2_X1    g34883(.A1(new_n38213_), .A2(pi0775), .Z(new_n38214_));
  NOR2_X1    g34884(.A1(new_n37969_), .A2(pi0769), .ZN(new_n38215_));
  NOR4_X1    g34885(.A1(new_n38214_), .A2(new_n38035_), .A3(new_n37980_), .A4(new_n38215_), .ZN(new_n38216_));
  AOI21_X1   g34886(.A1(new_n38216_), .A2(new_n38210_), .B(pi0795), .ZN(new_n38217_));
  NOR2_X1    g34887(.A1(new_n38212_), .A2(new_n38217_), .ZN(po0926));
  NAND3_X1   g34888(.A1(po0988), .A2(pi0966), .A3(pi1126), .ZN(new_n38219_));
  NAND3_X1   g34889(.A1(po0988), .A2(new_n36958_), .A3(new_n37135_), .ZN(new_n38220_));
  AOI21_X1   g34890(.A1(new_n38219_), .A2(new_n38220_), .B(new_n17019_), .ZN(po0927));
  NAND2_X1   g34891(.A1(new_n38116_), .A2(new_n37975_), .ZN(new_n38222_));
  NAND2_X1   g34892(.A1(new_n38187_), .A2(new_n37976_), .ZN(new_n38223_));
  NAND3_X1   g34893(.A1(new_n38223_), .A2(new_n37966_), .A3(new_n37994_), .ZN(new_n38224_));
  AOI21_X1   g34894(.A1(new_n38224_), .A2(new_n38222_), .B(new_n38037_), .ZN(po0963));
  INV_X1     g34895(.I(po0963), .ZN(new_n38226_));
  NOR3_X1    g34896(.A1(po0978), .A2(new_n38181_), .A3(new_n37967_), .ZN(new_n38227_));
  NOR3_X1    g34897(.A1(new_n38227_), .A2(pi0945), .A3(pi0987), .ZN(new_n38228_));
  NOR2_X1    g34898(.A1(new_n38226_), .A2(new_n38228_), .ZN(po0928));
  NAND3_X1   g34899(.A1(po0988), .A2(pi0966), .A3(pi1102), .ZN(new_n38230_));
  NAND3_X1   g34900(.A1(po0988), .A2(new_n36958_), .A3(new_n37195_), .ZN(new_n38231_));
  AOI21_X1   g34901(.A1(new_n38230_), .A2(new_n38231_), .B(new_n17845_), .ZN(po0929));
  NOR4_X1    g34902(.A1(new_n37947_), .A2(new_n37948_), .A3(pi0801), .A4(new_n37968_), .ZN(new_n38233_));
  NAND2_X1   g34903(.A1(po0963), .A2(new_n38233_), .ZN(new_n38234_));
  OAI21_X1   g34904(.A1(new_n37631_), .A2(new_n38117_), .B(new_n37952_), .ZN(new_n38235_));
  NAND3_X1   g34905(.A1(new_n38235_), .A2(pi0773), .A3(new_n37968_), .ZN(new_n38236_));
  XOR2_X1    g34906(.A1(new_n38234_), .A2(new_n38236_), .Z(po0930));
  NAND3_X1   g34907(.A1(po0988), .A2(pi0966), .A3(pi1127), .ZN(new_n38238_));
  NAND3_X1   g34908(.A1(po0988), .A2(new_n36958_), .A3(new_n37087_), .ZN(new_n38239_));
  AOI21_X1   g34909(.A1(new_n38238_), .A2(new_n38239_), .B(new_n15573_), .ZN(po0931));
  NAND4_X1   g34910(.A1(pi0795), .A2(pi0800), .A3(pi0801), .A4(pi0816), .ZN(new_n38241_));
  XOR2_X1    g34911(.A1(new_n37946_), .A2(new_n38241_), .Z(new_n38242_));
  NOR3_X1    g34912(.A1(new_n38035_), .A2(new_n38179_), .A3(new_n38181_), .ZN(new_n38243_));
  NOR3_X1    g34913(.A1(new_n37966_), .A2(new_n37962_), .A3(pi0945), .ZN(new_n38244_));
  NOR2_X1    g34914(.A1(new_n38243_), .A2(new_n38244_), .ZN(new_n38245_));
  OAI21_X1   g34915(.A1(new_n37966_), .A2(pi0945), .B(new_n37962_), .ZN(new_n38246_));
  NAND3_X1   g34916(.A1(new_n38243_), .A2(new_n37932_), .A3(new_n38246_), .ZN(new_n38247_));
  OR4_X2     g34917(.A1(new_n38039_), .A2(new_n38242_), .A3(new_n38245_), .A4(new_n38247_), .Z(new_n38248_));
  AOI21_X1   g34918(.A1(new_n38248_), .A2(new_n37962_), .B(new_n38176_), .ZN(po0932));
  INV_X1     g34919(.I(pi0776), .ZN(new_n38250_));
  NAND3_X1   g34920(.A1(po0988), .A2(pi0966), .A3(pi1128), .ZN(new_n38251_));
  NAND3_X1   g34921(.A1(po0988), .A2(new_n36958_), .A3(new_n37101_), .ZN(new_n38252_));
  AOI21_X1   g34922(.A1(new_n38251_), .A2(new_n38252_), .B(new_n38250_), .ZN(po0933));
  NAND3_X1   g34923(.A1(po0988), .A2(pi0966), .A3(pi1122), .ZN(new_n38254_));
  NAND3_X1   g34924(.A1(po0988), .A2(new_n36958_), .A3(new_n37012_), .ZN(new_n38255_));
  AOI21_X1   g34925(.A1(new_n38254_), .A2(new_n38255_), .B(new_n17735_), .ZN(po0934));
  NOR2_X1    g34926(.A1(pi1046), .A2(pi1083), .ZN(new_n38257_));
  NAND4_X1   g34927(.A1(new_n38257_), .A2(pi0832), .A3(pi0956), .A4(pi1085), .ZN(new_n38258_));
  NOR2_X1    g34928(.A1(new_n38258_), .A2(pi0968), .ZN(new_n38259_));
  NAND2_X1   g34929(.A1(new_n38259_), .A2(pi1100), .ZN(new_n38260_));
  OAI21_X1   g34930(.A1(new_n13748_), .A2(new_n38259_), .B(new_n38260_), .ZN(po0935));
  AOI21_X1   g34931(.A1(new_n36940_), .A2(new_n36994_), .B(new_n7240_), .ZN(po0936));
  AOI21_X1   g34932(.A1(new_n37032_), .A2(new_n36911_), .B(new_n7240_), .ZN(po0937));
  NAND2_X1   g34933(.A1(new_n38259_), .A2(pi1101), .ZN(new_n38264_));
  OAI21_X1   g34934(.A1(new_n13855_), .A2(new_n38259_), .B(new_n38264_), .ZN(po0938));
  OAI22_X1   g34935(.A1(new_n3098_), .A2(new_n5403_), .B1(new_n5405_), .B2(new_n36943_), .ZN(new_n38266_));
  OAI21_X1   g34936(.A1(po1038), .A2(pi0882), .B(new_n38266_), .ZN(po0939));
  NAND2_X1   g34937(.A1(new_n38259_), .A2(pi1109), .ZN(new_n38268_));
  OAI21_X1   g34938(.A1(new_n37410_), .A2(new_n38259_), .B(new_n38268_), .ZN(po0940));
  INV_X1     g34939(.I(pi0784), .ZN(new_n38270_));
  NAND2_X1   g34940(.A1(new_n38259_), .A2(pi1110), .ZN(new_n38271_));
  OAI21_X1   g34941(.A1(new_n38270_), .A2(new_n38259_), .B(new_n38271_), .ZN(po0941));
  NAND2_X1   g34942(.A1(new_n38259_), .A2(pi1102), .ZN(new_n38273_));
  OAI21_X1   g34943(.A1(new_n13801_), .A2(new_n38259_), .B(new_n38273_), .ZN(po0942));
  NAND2_X1   g34944(.A1(new_n8319_), .A2(pi0954), .ZN(new_n38275_));
  OAI21_X1   g34945(.A1(pi0024), .A2(pi0954), .B(new_n38275_), .ZN(po0943));
  NAND2_X1   g34946(.A1(new_n38259_), .A2(pi1104), .ZN(new_n38277_));
  OAI21_X1   g34947(.A1(new_n12776_), .A2(new_n38259_), .B(new_n38277_), .ZN(po0944));
  NAND2_X1   g34948(.A1(new_n38259_), .A2(pi1105), .ZN(new_n38279_));
  OAI21_X1   g34949(.A1(new_n13937_), .A2(new_n38259_), .B(new_n38279_), .ZN(po0945));
  NAND2_X1   g34950(.A1(new_n38259_), .A2(pi1106), .ZN(new_n38281_));
  OAI21_X1   g34951(.A1(new_n13896_), .A2(new_n38259_), .B(new_n38281_), .ZN(po0946));
  NAND2_X1   g34952(.A1(new_n38259_), .A2(pi1107), .ZN(new_n38283_));
  OAI21_X1   g34953(.A1(new_n12775_), .A2(new_n38259_), .B(new_n38283_), .ZN(po0947));
  INV_X1     g34954(.I(pi0791), .ZN(new_n38285_));
  NAND2_X1   g34955(.A1(new_n38259_), .A2(pi1108), .ZN(new_n38286_));
  OAI21_X1   g34956(.A1(new_n38285_), .A2(new_n38259_), .B(new_n38286_), .ZN(po0948));
  NAND2_X1   g34957(.A1(new_n38259_), .A2(pi1103), .ZN(new_n38288_));
  OAI21_X1   g34958(.A1(new_n12777_), .A2(new_n38259_), .B(new_n38288_), .ZN(po0949));
  INV_X1     g34959(.I(pi0968), .ZN(new_n38290_));
  NOR2_X1    g34960(.A1(new_n38258_), .A2(new_n38290_), .ZN(new_n38291_));
  NAND2_X1   g34961(.A1(new_n38291_), .A2(pi1130), .ZN(new_n38292_));
  OAI21_X1   g34962(.A1(new_n37929_), .A2(new_n38291_), .B(new_n38292_), .ZN(po0951));
  NAND2_X1   g34963(.A1(new_n38291_), .A2(pi1128), .ZN(new_n38294_));
  OAI21_X1   g34964(.A1(new_n37994_), .A2(new_n38291_), .B(new_n38294_), .ZN(po0952));
  NAND4_X1   g34965(.A1(new_n37178_), .A2(new_n34586_), .A3(pi0278), .A4(pi0279), .ZN(new_n38296_));
  NOR3_X1    g34966(.A1(new_n38296_), .A2(new_n3669_), .A3(new_n37182_), .ZN(new_n38297_));
  XOR2_X1    g34967(.A1(new_n38297_), .A2(pi0281), .Z(po0953));
  INV_X1     g34968(.I(pi0798), .ZN(new_n38299_));
  NAND2_X1   g34969(.A1(new_n38291_), .A2(pi1124), .ZN(new_n38300_));
  OAI21_X1   g34970(.A1(new_n38299_), .A2(new_n38291_), .B(new_n38300_), .ZN(po0955));
  NAND2_X1   g34971(.A1(new_n38291_), .A2(pi1107), .ZN(new_n38302_));
  OAI21_X1   g34972(.A1(pi0799), .A2(new_n38291_), .B(new_n38302_), .ZN(po0956));
  NAND2_X1   g34973(.A1(new_n38291_), .A2(pi1125), .ZN(new_n38304_));
  OAI21_X1   g34974(.A1(new_n38182_), .A2(new_n38291_), .B(new_n38304_), .ZN(po0957));
  NAND2_X1   g34975(.A1(new_n38291_), .A2(pi1126), .ZN(new_n38306_));
  OAI21_X1   g34976(.A1(new_n37631_), .A2(new_n38291_), .B(new_n38306_), .ZN(po0958));
  NOR4_X1    g34977(.A1(new_n37184_), .A2(pi0264), .A3(pi0265), .A4(pi0274), .ZN(po0959));
  NAND2_X1   g34978(.A1(new_n38291_), .A2(pi1106), .ZN(new_n38309_));
  OAI21_X1   g34979(.A1(pi0803), .A2(new_n38291_), .B(new_n38309_), .ZN(po0960));
  NAND2_X1   g34980(.A1(new_n38291_), .A2(pi1109), .ZN(new_n38311_));
  OAI21_X1   g34981(.A1(new_n35621_), .A2(new_n38291_), .B(new_n38311_), .ZN(po0961));
  NOR2_X1    g34982(.A1(new_n37181_), .A2(pi0282), .ZN(new_n38313_));
  NAND2_X1   g34983(.A1(new_n35070_), .A2(pi0270), .ZN(new_n38314_));
  OAI22_X1   g34984(.A1(new_n38313_), .A2(pi0270), .B1(new_n37181_), .B2(new_n38314_), .ZN(po0962));
  NAND2_X1   g34985(.A1(new_n38291_), .A2(pi1127), .ZN(new_n38316_));
  OAI21_X1   g34986(.A1(new_n37936_), .A2(new_n38291_), .B(new_n38316_), .ZN(po0964));
  INV_X1     g34987(.I(pi0808), .ZN(new_n38318_));
  NAND2_X1   g34988(.A1(new_n38291_), .A2(pi1101), .ZN(new_n38319_));
  OAI21_X1   g34989(.A1(new_n38318_), .A2(new_n38291_), .B(new_n38319_), .ZN(po0965));
  NAND2_X1   g34990(.A1(new_n38291_), .A2(pi1103), .ZN(new_n38321_));
  OAI21_X1   g34991(.A1(pi0809), .A2(new_n38291_), .B(new_n38321_), .ZN(po0966));
  NAND2_X1   g34992(.A1(new_n38291_), .A2(pi1108), .ZN(new_n38323_));
  OAI21_X1   g34993(.A1(new_n35622_), .A2(new_n38291_), .B(new_n38323_), .ZN(po0967));
  NAND2_X1   g34994(.A1(new_n38291_), .A2(pi1102), .ZN(new_n38325_));
  OAI21_X1   g34995(.A1(new_n37242_), .A2(new_n38291_), .B(new_n38325_), .ZN(po0968));
  NAND2_X1   g34996(.A1(new_n38291_), .A2(pi1104), .ZN(new_n38327_));
  OAI21_X1   g34997(.A1(pi0812), .A2(new_n38291_), .B(new_n38327_), .ZN(po0969));
  NAND2_X1   g34998(.A1(new_n38291_), .A2(pi1131), .ZN(new_n38329_));
  OAI21_X1   g34999(.A1(new_n37931_), .A2(new_n38291_), .B(new_n38329_), .ZN(po0970));
  NAND2_X1   g35000(.A1(new_n38291_), .A2(pi1105), .ZN(new_n38331_));
  OAI21_X1   g35001(.A1(pi0814), .A2(new_n38291_), .B(new_n38331_), .ZN(po0971));
  NAND2_X1   g35002(.A1(new_n38291_), .A2(pi1110), .ZN(new_n38333_));
  OAI21_X1   g35003(.A1(new_n35633_), .A2(new_n38291_), .B(new_n38333_), .ZN(po0972));
  NAND2_X1   g35004(.A1(new_n38291_), .A2(pi1129), .ZN(new_n38335_));
  OAI21_X1   g35005(.A1(new_n37814_), .A2(new_n38291_), .B(new_n38335_), .ZN(po0973));
  XOR2_X1    g35006(.A1(new_n37179_), .A2(pi0269), .Z(po0974));
  OAI21_X1   g35007(.A1(new_n11015_), .A2(new_n10169_), .B(new_n10915_), .ZN(po0975));
  NOR2_X1    g35008(.A1(new_n37184_), .A2(pi0264), .ZN(new_n38339_));
  NAND2_X1   g35009(.A1(new_n3669_), .A2(pi0265), .ZN(new_n38340_));
  OAI22_X1   g35010(.A1(new_n38339_), .A2(pi0265), .B1(new_n37184_), .B2(new_n38340_), .ZN(po0976));
  NAND3_X1   g35011(.A1(new_n37180_), .A2(pi0277), .A3(pi0282), .ZN(new_n38342_));
  XOR2_X1    g35012(.A1(new_n38342_), .A2(new_n34630_), .Z(po0977));
  NOR2_X1    g35013(.A1(pi0811), .A2(pi0893), .ZN(po0979));
  INV_X1     g35014(.I(pi0982), .ZN(new_n38345_));
  NAND3_X1   g35015(.A1(new_n2980_), .A2(new_n6940_), .A3(new_n7250_), .ZN(new_n38346_));
  AOI21_X1   g35016(.A1(new_n38346_), .A2(new_n38345_), .B(new_n10461_), .ZN(po0981));
  XOR2_X1    g35017(.A1(pi1125), .A2(pi1128), .Z(new_n38348_));
  XOR2_X1    g35018(.A1(new_n38348_), .A2(new_n37135_), .Z(new_n38349_));
  XOR2_X1    g35019(.A1(new_n38349_), .A2(pi1129), .Z(new_n38350_));
  XNOR2_X1   g35020(.A1(pi1124), .A2(pi1130), .ZN(new_n38351_));
  NAND2_X1   g35021(.A1(new_n38350_), .A2(new_n38351_), .ZN(new_n38352_));
  XNOR2_X1   g35022(.A1(pi1124), .A2(pi1130), .ZN(new_n38353_));
  OR2_X2     g35023(.A1(new_n38350_), .A2(new_n38353_), .Z(new_n38354_));
  NOR2_X1    g35024(.A1(new_n3136_), .A2(new_n34027_), .ZN(new_n38355_));
  NAND4_X1   g35025(.A1(new_n38355_), .A2(pi0825), .A3(pi1127), .A4(pi1131), .ZN(new_n38356_));
  NAND2_X1   g35026(.A1(pi0825), .A2(pi1131), .ZN(new_n38357_));
  NAND3_X1   g35027(.A1(new_n38355_), .A2(new_n37087_), .A3(new_n38357_), .ZN(new_n38358_));
  INV_X1     g35028(.I(new_n38355_), .ZN(new_n38359_));
  NAND3_X1   g35029(.A1(new_n38359_), .A2(pi1127), .A3(pi1131), .ZN(new_n38360_));
  NAND3_X1   g35030(.A1(new_n38360_), .A2(new_n38356_), .A3(new_n38358_), .ZN(new_n38361_));
  AOI21_X1   g35031(.A1(new_n38354_), .A2(new_n38352_), .B(new_n38361_), .ZN(po0982));
  XOR2_X1    g35032(.A1(pi1116), .A2(pi1120), .Z(new_n38363_));
  XOR2_X1    g35033(.A1(new_n38363_), .A2(new_n37008_), .Z(new_n38364_));
  XOR2_X1    g35034(.A1(new_n38364_), .A2(pi1121), .Z(new_n38365_));
  XNOR2_X1   g35035(.A1(pi1118), .A2(pi1119), .ZN(new_n38366_));
  NAND2_X1   g35036(.A1(new_n38365_), .A2(new_n38366_), .ZN(new_n38367_));
  XNOR2_X1   g35037(.A1(pi1118), .A2(pi1119), .ZN(new_n38368_));
  OR2_X2     g35038(.A1(new_n38365_), .A2(new_n38368_), .Z(new_n38369_));
  NAND4_X1   g35039(.A1(new_n38355_), .A2(pi0826), .A3(pi1122), .A4(pi1123), .ZN(new_n38370_));
  NAND2_X1   g35040(.A1(pi0826), .A2(pi1123), .ZN(new_n38371_));
  NAND3_X1   g35041(.A1(new_n38355_), .A2(new_n37012_), .A3(new_n38371_), .ZN(new_n38372_));
  NAND3_X1   g35042(.A1(new_n38359_), .A2(pi1122), .A3(pi1123), .ZN(new_n38373_));
  NAND3_X1   g35043(.A1(new_n38373_), .A2(new_n38370_), .A3(new_n38372_), .ZN(new_n38374_));
  AOI21_X1   g35044(.A1(new_n38369_), .A2(new_n38367_), .B(new_n38374_), .ZN(po0983));
  XOR2_X1    g35045(.A1(pi1101), .A2(pi1104), .Z(new_n38376_));
  XOR2_X1    g35046(.A1(new_n38376_), .A2(new_n37195_), .Z(new_n38377_));
  XOR2_X1    g35047(.A1(new_n38377_), .A2(pi1106), .Z(new_n38378_));
  XNOR2_X1   g35048(.A1(pi1103), .A2(pi1105), .ZN(new_n38379_));
  NAND2_X1   g35049(.A1(new_n38378_), .A2(new_n38379_), .ZN(new_n38380_));
  XNOR2_X1   g35050(.A1(pi1103), .A2(pi1105), .ZN(new_n38381_));
  OR2_X2     g35051(.A1(new_n38378_), .A2(new_n38381_), .Z(new_n38382_));
  NAND4_X1   g35052(.A1(new_n38355_), .A2(pi0827), .A3(pi1100), .A4(pi1107), .ZN(new_n38383_));
  NAND2_X1   g35053(.A1(pi0827), .A2(pi1107), .ZN(new_n38384_));
  NAND3_X1   g35054(.A1(new_n38355_), .A2(new_n37523_), .A3(new_n38384_), .ZN(new_n38385_));
  NAND3_X1   g35055(.A1(new_n38359_), .A2(pi1100), .A3(pi1107), .ZN(new_n38386_));
  NAND3_X1   g35056(.A1(new_n38386_), .A2(new_n38383_), .A3(new_n38385_), .ZN(new_n38387_));
  AOI21_X1   g35057(.A1(new_n38382_), .A2(new_n38380_), .B(new_n38387_), .ZN(po0984));
  XOR2_X1    g35058(.A1(pi1108), .A2(pi1112), .Z(new_n38389_));
  XOR2_X1    g35059(.A1(new_n38389_), .A2(new_n37025_), .Z(new_n38390_));
  XOR2_X1    g35060(.A1(new_n38390_), .A2(pi1113), .Z(new_n38391_));
  XNOR2_X1   g35061(.A1(pi1110), .A2(pi1111), .ZN(new_n38392_));
  NAND2_X1   g35062(.A1(new_n38391_), .A2(new_n38392_), .ZN(new_n38393_));
  XNOR2_X1   g35063(.A1(pi1110), .A2(pi1111), .ZN(new_n38394_));
  OR2_X2     g35064(.A1(new_n38391_), .A2(new_n38394_), .Z(new_n38395_));
  NAND4_X1   g35065(.A1(new_n38355_), .A2(pi0828), .A3(pi1114), .A4(pi1115), .ZN(new_n38396_));
  NAND2_X1   g35066(.A1(pi0828), .A2(pi1115), .ZN(new_n38397_));
  NAND3_X1   g35067(.A1(new_n38355_), .A2(new_n36977_), .A3(new_n38397_), .ZN(new_n38398_));
  NAND3_X1   g35068(.A1(new_n38359_), .A2(pi1114), .A3(pi1115), .ZN(new_n38399_));
  NAND3_X1   g35069(.A1(new_n38399_), .A2(new_n38396_), .A3(new_n38398_), .ZN(new_n38400_));
  AOI21_X1   g35070(.A1(new_n38395_), .A2(new_n38393_), .B(new_n38400_), .ZN(po0985));
  NAND2_X1   g35071(.A1(pi0951), .A2(pi1092), .ZN(new_n38402_));
  AOI21_X1   g35072(.A1(new_n2986_), .A2(new_n38402_), .B(new_n10169_), .ZN(po0986));
  XOR2_X1    g35073(.A1(new_n38296_), .A2(pi0281), .Z(po0987));
  AND4_X2    g35074(.A1(pi0832), .A2(new_n7259_), .A3(pi1091), .A4(pi1162), .Z(po0989));
  NAND3_X1   g35075(.A1(new_n9992_), .A2(pi0833), .A3(pi1091), .ZN(new_n38406_));
  NAND3_X1   g35076(.A1(new_n9992_), .A2(new_n3058_), .A3(new_n2726_), .ZN(new_n38407_));
  NAND2_X1   g35077(.A1(new_n38406_), .A2(new_n38407_), .ZN(po0990));
  INV_X1     g35078(.I(pi0946), .ZN(new_n38409_));
  NOR2_X1    g35079(.A1(new_n2723_), .A2(new_n38409_), .ZN(po0991));
  XOR2_X1    g35080(.A1(new_n37180_), .A2(new_n35070_), .Z(po0992));
  NAND2_X1   g35081(.A1(pi0837), .A2(pi0955), .ZN(new_n38412_));
  OAI21_X1   g35082(.A1(pi0955), .A2(new_n35178_), .B(new_n38412_), .ZN(po0993));
  NAND2_X1   g35083(.A1(pi0838), .A2(pi0955), .ZN(new_n38414_));
  OAI21_X1   g35084(.A1(pi0955), .A2(new_n35282_), .B(new_n38414_), .ZN(po0994));
  NAND2_X1   g35085(.A1(pi0839), .A2(pi0955), .ZN(new_n38416_));
  OAI21_X1   g35086(.A1(pi0955), .A2(new_n35289_), .B(new_n38416_), .ZN(po0995));
  NAND2_X1   g35087(.A1(new_n2723_), .A2(pi0840), .ZN(new_n38418_));
  OAI21_X1   g35088(.A1(new_n6595_), .A2(new_n2723_), .B(new_n38418_), .ZN(po0996));
  INV_X1     g35089(.I(new_n7960_), .ZN(new_n38420_));
  NOR2_X1    g35090(.A1(new_n38420_), .A2(pi0033), .ZN(po0997));
  NAND2_X1   g35091(.A1(pi0842), .A2(pi0955), .ZN(new_n38422_));
  OAI21_X1   g35092(.A1(pi0955), .A2(new_n35385_), .B(new_n38422_), .ZN(po0998));
  NAND2_X1   g35093(.A1(pi0843), .A2(pi0955), .ZN(new_n38424_));
  OAI21_X1   g35094(.A1(pi0955), .A2(new_n35388_), .B(new_n38424_), .ZN(po0999));
  NAND2_X1   g35095(.A1(pi0844), .A2(pi0955), .ZN(new_n38426_));
  OAI21_X1   g35096(.A1(pi0955), .A2(new_n35391_), .B(new_n38426_), .ZN(po1000));
  NAND2_X1   g35097(.A1(pi0845), .A2(pi0955), .ZN(new_n38428_));
  OAI21_X1   g35098(.A1(pi0955), .A2(new_n35319_), .B(new_n38428_), .ZN(po1001));
  NAND2_X1   g35099(.A1(new_n34029_), .A2(pi0846), .ZN(new_n38430_));
  OAI21_X1   g35100(.A1(new_n5132_), .A2(new_n34029_), .B(new_n38430_), .ZN(po1002));
  NAND2_X1   g35101(.A1(pi0847), .A2(pi0955), .ZN(new_n38432_));
  OAI21_X1   g35102(.A1(pi0955), .A2(new_n35377_), .B(new_n38432_), .ZN(po1003));
  NAND2_X1   g35103(.A1(pi0848), .A2(pi0955), .ZN(new_n38434_));
  OAI21_X1   g35104(.A1(pi0955), .A2(new_n33609_), .B(new_n38434_), .ZN(po1004));
  NAND2_X1   g35105(.A1(new_n2723_), .A2(pi0849), .ZN(new_n38436_));
  OAI21_X1   g35106(.A1(new_n6577_), .A2(new_n2723_), .B(new_n38436_), .ZN(po1005));
  NAND2_X1   g35107(.A1(pi0850), .A2(pi0955), .ZN(new_n38438_));
  OAI21_X1   g35108(.A1(pi0955), .A2(new_n35175_), .B(new_n38438_), .ZN(po1006));
  NAND2_X1   g35109(.A1(pi0851), .A2(pi0955), .ZN(new_n38440_));
  OAI21_X1   g35110(.A1(pi0955), .A2(new_n35396_), .B(new_n38440_), .ZN(po1007));
  NAND2_X1   g35111(.A1(pi0852), .A2(pi0955), .ZN(new_n38442_));
  OAI21_X1   g35112(.A1(pi0955), .A2(new_n34003_), .B(new_n38442_), .ZN(po1008));
  NAND2_X1   g35113(.A1(pi0853), .A2(pi0955), .ZN(new_n38444_));
  OAI21_X1   g35114(.A1(pi0955), .A2(new_n35277_), .B(new_n38444_), .ZN(po1009));
  NAND2_X1   g35115(.A1(pi0854), .A2(pi0955), .ZN(new_n38446_));
  OAI21_X1   g35116(.A1(pi0955), .A2(new_n35301_), .B(new_n38446_), .ZN(po1010));
  NAND2_X1   g35117(.A1(pi0855), .A2(pi0955), .ZN(new_n38448_));
  OAI21_X1   g35118(.A1(pi0955), .A2(new_n33997_), .B(new_n38448_), .ZN(po1011));
  NAND2_X1   g35119(.A1(pi0856), .A2(pi0955), .ZN(new_n38450_));
  OAI21_X1   g35120(.A1(pi0955), .A2(new_n34016_), .B(new_n38450_), .ZN(po1012));
  NAND2_X1   g35121(.A1(pi0857), .A2(pi0955), .ZN(new_n38452_));
  OAI21_X1   g35122(.A1(pi0955), .A2(new_n35298_), .B(new_n38452_), .ZN(po1013));
  NAND2_X1   g35123(.A1(pi0858), .A2(pi0955), .ZN(new_n38454_));
  OAI21_X1   g35124(.A1(pi0955), .A2(new_n35380_), .B(new_n38454_), .ZN(po1014));
  NAND2_X1   g35125(.A1(pi0859), .A2(pi0955), .ZN(new_n38456_));
  OAI21_X1   g35126(.A1(pi0955), .A2(new_n33991_), .B(new_n38456_), .ZN(po1015));
  NAND2_X1   g35127(.A1(pi0860), .A2(pi0955), .ZN(new_n38458_));
  OAI21_X1   g35128(.A1(pi0955), .A2(new_n35404_), .B(new_n38458_), .ZN(po1016));
  NAND2_X1   g35129(.A1(pi0228), .A2(pi1093), .ZN(new_n38460_));
  NOR2_X1    g35130(.A1(new_n2984_), .A2(pi0861), .ZN(new_n38461_));
  XOR2_X1    g35131(.A1(new_n38461_), .A2(new_n38460_), .Z(new_n38462_));
  NAND2_X1   g35132(.A1(pi0123), .A2(pi0228), .ZN(new_n38463_));
  NOR2_X1    g35133(.A1(new_n3005_), .A2(pi0861), .ZN(new_n38464_));
  XOR2_X1    g35134(.A1(new_n38464_), .A2(new_n38463_), .Z(new_n38465_));
  AOI21_X1   g35135(.A1(new_n38462_), .A2(new_n38465_), .B(new_n3980_), .ZN(po1017));
  NAND2_X1   g35136(.A1(new_n34029_), .A2(pi0862), .ZN(new_n38467_));
  OAI21_X1   g35137(.A1(new_n4300_), .A2(new_n34029_), .B(new_n38467_), .ZN(po1018));
  NAND2_X1   g35138(.A1(new_n2723_), .A2(pi0863), .ZN(new_n38469_));
  OAI21_X1   g35139(.A1(new_n6356_), .A2(new_n2723_), .B(new_n38469_), .ZN(po1019));
  NAND2_X1   g35140(.A1(new_n2723_), .A2(pi0864), .ZN(new_n38471_));
  OAI21_X1   g35141(.A1(new_n6728_), .A2(new_n2723_), .B(new_n38471_), .ZN(po1020));
  NAND2_X1   g35142(.A1(pi0865), .A2(pi0955), .ZN(new_n38473_));
  OAI21_X1   g35143(.A1(pi0955), .A2(new_n34023_), .B(new_n38473_), .ZN(po1021));
  NAND2_X1   g35144(.A1(pi0866), .A2(pi0955), .ZN(new_n38475_));
  OAI21_X1   g35145(.A1(pi0955), .A2(new_n33607_), .B(new_n38475_), .ZN(po1022));
  NAND2_X1   g35146(.A1(pi0867), .A2(pi0955), .ZN(new_n38477_));
  OAI21_X1   g35147(.A1(pi0955), .A2(new_n35312_), .B(new_n38477_), .ZN(po1023));
  NAND2_X1   g35148(.A1(pi0868), .A2(pi0955), .ZN(new_n38479_));
  OAI21_X1   g35149(.A1(pi0955), .A2(new_n35309_), .B(new_n38479_), .ZN(po1024));
  NOR2_X1    g35150(.A1(new_n2984_), .A2(pi0869), .ZN(new_n38481_));
  XOR2_X1    g35151(.A1(new_n38481_), .A2(new_n38460_), .Z(new_n38482_));
  NOR2_X1    g35152(.A1(new_n3005_), .A2(pi0869), .ZN(new_n38483_));
  XOR2_X1    g35153(.A1(new_n38483_), .A2(new_n38463_), .Z(new_n38484_));
  AOI21_X1   g35154(.A1(new_n38482_), .A2(new_n38484_), .B(new_n4141_), .ZN(po1025));
  NAND2_X1   g35155(.A1(pi0870), .A2(pi0955), .ZN(new_n38486_));
  OAI21_X1   g35156(.A1(pi0955), .A2(new_n34009_), .B(new_n38486_), .ZN(po1026));
  NAND2_X1   g35157(.A1(pi0871), .A2(pi0955), .ZN(new_n38488_));
  OAI21_X1   g35158(.A1(pi0955), .A2(new_n35187_), .B(new_n38488_), .ZN(po1027));
  NAND2_X1   g35159(.A1(pi0872), .A2(pi0955), .ZN(new_n38490_));
  OAI21_X1   g35160(.A1(pi0955), .A2(new_n35181_), .B(new_n38490_), .ZN(po1028));
  NAND2_X1   g35161(.A1(pi0873), .A2(pi0955), .ZN(new_n38492_));
  OAI21_X1   g35162(.A1(pi0955), .A2(new_n34014_), .B(new_n38492_), .ZN(po1029));
  NAND2_X1   g35163(.A1(pi0874), .A2(pi0955), .ZN(new_n38494_));
  OAI21_X1   g35164(.A1(pi0955), .A2(new_n33985_), .B(new_n38494_), .ZN(po1030));
  NAND2_X1   g35165(.A1(new_n4809_), .A2(pi1093), .ZN(new_n38496_));
  XOR2_X1    g35166(.A1(new_n38496_), .A2(new_n38460_), .Z(new_n38497_));
  NAND2_X1   g35167(.A1(new_n4809_), .A2(pi0228), .ZN(new_n38498_));
  XOR2_X1    g35168(.A1(new_n38498_), .A2(new_n38463_), .Z(new_n38499_));
  OAI21_X1   g35169(.A1(new_n38497_), .A2(new_n38499_), .B(pi1136), .ZN(po1031));
  NAND2_X1   g35170(.A1(pi0876), .A2(pi0955), .ZN(new_n38501_));
  OAI21_X1   g35171(.A1(pi0955), .A2(new_n34021_), .B(new_n38501_), .ZN(po1032));
  NOR2_X1    g35172(.A1(new_n2984_), .A2(pi0877), .ZN(new_n38503_));
  XOR2_X1    g35173(.A1(new_n38503_), .A2(new_n38460_), .Z(new_n38504_));
  NOR2_X1    g35174(.A1(new_n3005_), .A2(pi0877), .ZN(new_n38505_));
  XOR2_X1    g35175(.A1(new_n38505_), .A2(new_n38463_), .Z(new_n38506_));
  AOI21_X1   g35176(.A1(new_n38504_), .A2(new_n38506_), .B(new_n4465_), .ZN(po1033));
  NOR2_X1    g35177(.A1(new_n2984_), .A2(pi0878), .ZN(new_n38508_));
  XOR2_X1    g35178(.A1(new_n38508_), .A2(new_n38460_), .Z(new_n38509_));
  NOR2_X1    g35179(.A1(new_n3005_), .A2(pi0878), .ZN(new_n38510_));
  XOR2_X1    g35180(.A1(new_n38510_), .A2(new_n38463_), .Z(new_n38511_));
  AOI21_X1   g35181(.A1(new_n38509_), .A2(new_n38511_), .B(new_n4626_), .ZN(po1034));
  NOR2_X1    g35182(.A1(new_n2984_), .A2(pi0879), .ZN(new_n38513_));
  XOR2_X1    g35183(.A1(new_n38513_), .A2(new_n38460_), .Z(new_n38514_));
  NOR2_X1    g35184(.A1(new_n3005_), .A2(pi0879), .ZN(new_n38515_));
  XOR2_X1    g35185(.A1(new_n38515_), .A2(new_n38463_), .Z(new_n38516_));
  AOI21_X1   g35186(.A1(new_n38514_), .A2(new_n38516_), .B(new_n4959_), .ZN(po1035));
  NAND2_X1   g35187(.A1(pi0880), .A2(pi0955), .ZN(new_n38518_));
  OAI21_X1   g35188(.A1(pi0955), .A2(new_n35401_), .B(new_n38518_), .ZN(po1036));
  NAND2_X1   g35189(.A1(pi0881), .A2(pi0955), .ZN(new_n38520_));
  OAI21_X1   g35190(.A1(pi0955), .A2(new_n35184_), .B(new_n38520_), .ZN(po1037));
  INV_X1     g35191(.I(pi0883), .ZN(po1163));
  NAND2_X1   g35192(.A1(new_n38355_), .A2(po1163), .ZN(new_n38523_));
  OAI21_X1   g35193(.A1(new_n36959_), .A2(new_n38355_), .B(new_n38523_), .ZN(po1039));
  INV_X1     g35194(.I(pi0884), .ZN(po1180));
  NAND2_X1   g35195(.A1(new_n38355_), .A2(po1180), .ZN(new_n38526_));
  OAI21_X1   g35196(.A1(new_n37163_), .A2(new_n38355_), .B(new_n38526_), .ZN(po1040));
  INV_X1     g35197(.I(pi0885), .ZN(po1172));
  NAND2_X1   g35198(.A1(new_n38355_), .A2(po1172), .ZN(new_n38529_));
  OAI21_X1   g35199(.A1(new_n37120_), .A2(new_n38355_), .B(new_n38529_), .ZN(po1041));
  INV_X1     g35200(.I(pi0886), .ZN(po1166));
  NAND2_X1   g35201(.A1(new_n38355_), .A2(po1166), .ZN(new_n38532_));
  OAI21_X1   g35202(.A1(new_n37025_), .A2(new_n38355_), .B(new_n38532_), .ZN(po1042));
  INV_X1     g35203(.I(pi0887), .ZN(po1179));
  NAND2_X1   g35204(.A1(new_n38355_), .A2(po1179), .ZN(new_n38535_));
  OAI21_X1   g35205(.A1(new_n37523_), .A2(new_n38355_), .B(new_n38535_), .ZN(po1043));
  INV_X1     g35206(.I(pi0888), .ZN(po1164));
  NAND2_X1   g35207(.A1(new_n38355_), .A2(po1164), .ZN(new_n38538_));
  OAI21_X1   g35208(.A1(new_n37063_), .A2(new_n38355_), .B(new_n38538_), .ZN(po1044));
  INV_X1     g35209(.I(pi0889), .ZN(po1170));
  NAND2_X1   g35210(.A1(new_n38355_), .A2(po1170), .ZN(new_n38541_));
  OAI21_X1   g35211(.A1(new_n37108_), .A2(new_n38355_), .B(new_n38541_), .ZN(po1045));
  INV_X1     g35212(.I(pi0890), .ZN(po1153));
  NAND2_X1   g35213(.A1(new_n38355_), .A2(po1153), .ZN(new_n38544_));
  OAI21_X1   g35214(.A1(new_n37135_), .A2(new_n38355_), .B(new_n38544_), .ZN(po1046));
  INV_X1     g35215(.I(pi0891), .ZN(po1160));
  NAND2_X1   g35216(.A1(new_n38355_), .A2(po1160), .ZN(new_n38547_));
  OAI21_X1   g35217(.A1(new_n36963_), .A2(new_n38355_), .B(new_n38547_), .ZN(po1047));
  INV_X1     g35218(.I(pi0892), .ZN(po1183));
  NAND2_X1   g35219(.A1(new_n38355_), .A2(po1183), .ZN(new_n38550_));
  OAI21_X1   g35220(.A1(new_n37191_), .A2(new_n38355_), .B(new_n38550_), .ZN(po1048));
  NAND2_X1   g35221(.A1(new_n2539_), .A2(new_n2644_), .ZN(po1049));
  INV_X1     g35222(.I(pi0894), .ZN(po1150));
  NAND2_X1   g35223(.A1(new_n38355_), .A2(po1150), .ZN(new_n38554_));
  OAI21_X1   g35224(.A1(new_n37056_), .A2(new_n38355_), .B(new_n38554_), .ZN(po1050));
  INV_X1     g35225(.I(pi0895), .ZN(po1168));
  NAND2_X1   g35226(.A1(new_n38355_), .A2(po1168), .ZN(new_n38557_));
  OAI21_X1   g35227(.A1(new_n36972_), .A2(new_n38355_), .B(new_n38557_), .ZN(po1051));
  INV_X1     g35228(.I(pi0896), .ZN(po1156));
  NAND2_X1   g35229(.A1(new_n38355_), .A2(po1156), .ZN(new_n38560_));
  OAI21_X1   g35230(.A1(new_n36967_), .A2(new_n38355_), .B(new_n38560_), .ZN(po1052));
  INV_X1     g35231(.I(pi0898), .ZN(po1176));
  NAND2_X1   g35232(.A1(new_n38355_), .A2(po1176), .ZN(new_n38563_));
  OAI21_X1   g35233(.A1(new_n37154_), .A2(new_n38355_), .B(new_n38563_), .ZN(po1054));
  INV_X1     g35234(.I(pi0899), .ZN(po1174));
  NAND2_X1   g35235(.A1(new_n38355_), .A2(po1174), .ZN(new_n38566_));
  OAI21_X1   g35236(.A1(new_n36986_), .A2(new_n38355_), .B(new_n38566_), .ZN(po1055));
  INV_X1     g35237(.I(pi0900), .ZN(po1171));
  NAND2_X1   g35238(.A1(new_n38355_), .A2(po1171), .ZN(new_n38569_));
  OAI21_X1   g35239(.A1(new_n37075_), .A2(new_n38355_), .B(new_n38569_), .ZN(po1056));
  INV_X1     g35240(.I(pi0902), .ZN(po1161));
  NAND2_X1   g35241(.A1(new_n38355_), .A2(po1161), .ZN(new_n38572_));
  OAI21_X1   g35242(.A1(new_n36981_), .A2(new_n38355_), .B(new_n38572_), .ZN(po1058));
  INV_X1     g35243(.I(pi0903), .ZN(po1162));
  NAND2_X1   g35244(.A1(new_n38355_), .A2(po1162), .ZN(new_n38575_));
  OAI21_X1   g35245(.A1(new_n37049_), .A2(new_n38355_), .B(new_n38575_), .ZN(po1059));
  INV_X1     g35246(.I(pi0904), .ZN(po1173));
  NAND2_X1   g35247(.A1(new_n38355_), .A2(po1173), .ZN(new_n38578_));
  OAI21_X1   g35248(.A1(new_n37087_), .A2(new_n38355_), .B(new_n38578_), .ZN(po1060));
  INV_X1     g35249(.I(pi0905), .ZN(po1151));
  NAND2_X1   g35250(.A1(new_n38355_), .A2(po1151), .ZN(new_n38581_));
  OAI21_X1   g35251(.A1(new_n37149_), .A2(new_n38355_), .B(new_n38581_), .ZN(po1061));
  INV_X1     g35252(.I(pi0906), .ZN(po1155));
  NAND2_X1   g35253(.A1(new_n38355_), .A2(po1155), .ZN(new_n38584_));
  OAI21_X1   g35254(.A1(new_n37101_), .A2(new_n38355_), .B(new_n38584_), .ZN(po1062));
  OAI21_X1   g35255(.A1(new_n36942_), .A2(pi0979), .B(pi0782), .ZN(new_n38586_));
  AOI21_X1   g35256(.A1(new_n36993_), .A2(pi0979), .B(new_n38586_), .ZN(new_n38587_));
  INV_X1     g35257(.I(pi0782), .ZN(new_n38588_));
  NOR3_X1    g35258(.A1(new_n36910_), .A2(new_n38588_), .A3(new_n5405_), .ZN(new_n38589_));
  NOR3_X1    g35259(.A1(new_n38588_), .A2(pi0598), .A3(pi0979), .ZN(new_n38590_));
  OAI21_X1   g35260(.A1(new_n38589_), .A2(new_n38590_), .B(pi0624), .ZN(new_n38591_));
  NOR2_X1    g35261(.A1(new_n38591_), .A2(new_n38588_), .ZN(new_n38592_));
  XNOR2_X1   g35262(.A1(new_n38592_), .A2(new_n38587_), .ZN(new_n38593_));
  NOR2_X1    g35263(.A1(new_n38593_), .A2(new_n5741_), .ZN(po1063));
  INV_X1     g35264(.I(pi0908), .ZN(po1159));
  NAND2_X1   g35265(.A1(new_n38355_), .A2(po1159), .ZN(new_n38596_));
  OAI21_X1   g35266(.A1(new_n37012_), .A2(new_n38355_), .B(new_n38596_), .ZN(po1064));
  INV_X1     g35267(.I(pi0909), .ZN(po1157));
  NAND2_X1   g35268(.A1(new_n38355_), .A2(po1157), .ZN(new_n38599_));
  OAI21_X1   g35269(.A1(new_n37002_), .A2(new_n38355_), .B(new_n38599_), .ZN(po1065));
  INV_X1     g35270(.I(pi0910), .ZN(po1181));
  NAND2_X1   g35271(.A1(new_n38355_), .A2(po1181), .ZN(new_n38602_));
  OAI21_X1   g35272(.A1(new_n37008_), .A2(new_n38355_), .B(new_n38602_), .ZN(po1066));
  INV_X1     g35273(.I(pi0911), .ZN(po1158));
  NAND2_X1   g35274(.A1(new_n38355_), .A2(po1158), .ZN(new_n38605_));
  OAI21_X1   g35275(.A1(new_n37144_), .A2(new_n38355_), .B(new_n38605_), .ZN(po1067));
  INV_X1     g35276(.I(pi0912), .ZN(po1167));
  NAND2_X1   g35277(.A1(new_n38355_), .A2(po1167), .ZN(new_n38608_));
  OAI21_X1   g35278(.A1(new_n36977_), .A2(new_n38355_), .B(new_n38608_), .ZN(po1068));
  INV_X1     g35279(.I(pi0913), .ZN(po1149));
  NAND2_X1   g35280(.A1(new_n38355_), .A2(po1149), .ZN(new_n38611_));
  OAI21_X1   g35281(.A1(new_n37029_), .A2(new_n38355_), .B(new_n38611_), .ZN(po1069));
  NAND2_X1   g35282(.A1(pi0266), .A2(pi0992), .ZN(new_n38613_));
  XOR2_X1    g35283(.A1(new_n38613_), .A2(pi0280), .Z(po1070));
  INV_X1     g35284(.I(pi0915), .ZN(po1146));
  NAND2_X1   g35285(.A1(new_n38355_), .A2(po1146), .ZN(new_n38616_));
  OAI21_X1   g35286(.A1(new_n37021_), .A2(new_n38355_), .B(new_n38616_), .ZN(po1071));
  INV_X1     g35287(.I(pi0916), .ZN(po1169));
  NAND2_X1   g35288(.A1(new_n38355_), .A2(po1169), .ZN(new_n38619_));
  OAI21_X1   g35289(.A1(new_n37115_), .A2(new_n38355_), .B(new_n38619_), .ZN(po1072));
  INV_X1     g35290(.I(pi0917), .ZN(po1177));
  NAND2_X1   g35291(.A1(new_n38355_), .A2(po1177), .ZN(new_n38622_));
  OAI21_X1   g35292(.A1(new_n37017_), .A2(new_n38355_), .B(new_n38622_), .ZN(po1073));
  INV_X1     g35293(.I(pi0918), .ZN(po1175));
  NAND2_X1   g35294(.A1(new_n38355_), .A2(po1175), .ZN(new_n38625_));
  OAI21_X1   g35295(.A1(new_n36951_), .A2(new_n38355_), .B(new_n38625_), .ZN(po1074));
  INV_X1     g35296(.I(pi0919), .ZN(po1165));
  NAND2_X1   g35297(.A1(new_n38355_), .A2(po1165), .ZN(new_n38628_));
  OAI21_X1   g35298(.A1(new_n37195_), .A2(new_n38355_), .B(new_n38628_), .ZN(po1075));
  NAND2_X1   g35299(.A1(pi1093), .A2(pi1139), .ZN(new_n38630_));
  OAI21_X1   g35300(.A1(new_n4302_), .A2(pi1093), .B(new_n38630_), .ZN(po1076));
  NAND2_X1   g35301(.A1(pi1093), .A2(pi1140), .ZN(new_n38632_));
  OAI21_X1   g35302(.A1(new_n4143_), .A2(pi1093), .B(new_n38632_), .ZN(po1077));
  NAND2_X1   g35303(.A1(pi1093), .A2(pi1152), .ZN(new_n38634_));
  OAI21_X1   g35304(.A1(new_n35770_), .A2(pi1093), .B(new_n38634_), .ZN(po1078));
  NAND2_X1   g35305(.A1(new_n2984_), .A2(pi0923), .ZN(new_n38636_));
  OAI21_X1   g35306(.A1(new_n2984_), .A2(new_n13817_), .B(new_n38636_), .ZN(po1079));
  AND4_X2    g35307(.A1(pi0300), .A2(pi0301), .A3(pi0311), .A4(pi0312), .Z(po1080));
  NAND2_X1   g35308(.A1(new_n2984_), .A2(pi0925), .ZN(new_n38639_));
  OAI21_X1   g35309(.A1(new_n2984_), .A2(new_n13778_), .B(new_n38639_), .ZN(po1081));
  NAND2_X1   g35310(.A1(new_n2984_), .A2(pi0926), .ZN(new_n38641_));
  OAI21_X1   g35311(.A1(new_n2984_), .A2(new_n14006_), .B(new_n38641_), .ZN(po1082));
  NAND2_X1   g35312(.A1(pi1093), .A2(pi1145), .ZN(new_n38643_));
  OAI21_X1   g35313(.A1(new_n3506_), .A2(pi1093), .B(new_n38643_), .ZN(po1083));
  NAND2_X1   g35314(.A1(pi1093), .A2(pi1136), .ZN(new_n38645_));
  OAI21_X1   g35315(.A1(new_n4792_), .A2(pi1093), .B(new_n38645_), .ZN(po1084));
  NAND2_X1   g35316(.A1(pi1093), .A2(pi1144), .ZN(new_n38647_));
  OAI21_X1   g35317(.A1(new_n3061_), .A2(pi1093), .B(new_n38647_), .ZN(po1085));
  NAND2_X1   g35318(.A1(pi1093), .A2(pi1134), .ZN(new_n38649_));
  OAI21_X1   g35319(.A1(new_n5150_), .A2(pi1093), .B(new_n38649_), .ZN(po1086));
  NAND2_X1   g35320(.A1(pi1093), .A2(pi1150), .ZN(new_n38651_));
  OAI21_X1   g35321(.A1(new_n35777_), .A2(pi1093), .B(new_n38651_), .ZN(po1087));
  NAND2_X1   g35322(.A1(pi1093), .A2(pi1142), .ZN(new_n38653_));
  OAI21_X1   g35323(.A1(new_n3816_), .A2(pi1093), .B(new_n38653_), .ZN(po1088));
  NAND2_X1   g35324(.A1(pi1093), .A2(pi1137), .ZN(new_n38655_));
  OAI21_X1   g35325(.A1(new_n4628_), .A2(pi1093), .B(new_n38655_), .ZN(po1089));
  NAND2_X1   g35326(.A1(new_n2984_), .A2(pi0934), .ZN(new_n38657_));
  OAI21_X1   g35327(.A1(new_n2984_), .A2(new_n31940_), .B(new_n38657_), .ZN(po1090));
  NAND2_X1   g35328(.A1(pi1093), .A2(pi1141), .ZN(new_n38659_));
  OAI21_X1   g35329(.A1(new_n3982_), .A2(pi1093), .B(new_n38659_), .ZN(po1091));
  NAND2_X1   g35330(.A1(pi1093), .A2(pi1149), .ZN(new_n38661_));
  OAI21_X1   g35331(.A1(new_n35784_), .A2(pi1093), .B(new_n38661_), .ZN(po1092));
  NAND2_X1   g35332(.A1(new_n2984_), .A2(pi0937), .ZN(new_n38663_));
  OAI21_X1   g35333(.A1(new_n2984_), .A2(new_n31953_), .B(new_n38663_), .ZN(po1093));
  NAND2_X1   g35334(.A1(pi1093), .A2(pi1135), .ZN(new_n38665_));
  OAI21_X1   g35335(.A1(new_n4961_), .A2(pi1093), .B(new_n38665_), .ZN(po1094));
  NAND2_X1   g35336(.A1(pi1093), .A2(pi1146), .ZN(new_n38667_));
  OAI21_X1   g35337(.A1(new_n3342_), .A2(pi1093), .B(new_n38667_), .ZN(po1095));
  NAND2_X1   g35338(.A1(pi1093), .A2(pi1138), .ZN(new_n38669_));
  OAI21_X1   g35339(.A1(new_n4467_), .A2(pi1093), .B(new_n38669_), .ZN(po1096));
  NAND2_X1   g35340(.A1(new_n2984_), .A2(pi0941), .ZN(new_n38671_));
  OAI21_X1   g35341(.A1(new_n2984_), .A2(new_n13614_), .B(new_n38671_), .ZN(po1097));
  NAND2_X1   g35342(.A1(new_n2984_), .A2(pi0942), .ZN(new_n38673_));
  OAI21_X1   g35343(.A1(new_n2984_), .A2(new_n13969_), .B(new_n38673_), .ZN(po1098));
  NAND2_X1   g35344(.A1(pi1093), .A2(pi1151), .ZN(new_n38675_));
  OAI21_X1   g35345(.A1(new_n35683_), .A2(pi1093), .B(new_n38675_), .ZN(po1099));
  NAND2_X1   g35346(.A1(pi1093), .A2(pi1143), .ZN(new_n38677_));
  OAI21_X1   g35347(.A1(new_n3652_), .A2(pi1093), .B(new_n38677_), .ZN(po1100));
  NOR2_X1    g35348(.A1(new_n2723_), .A2(new_n30557_), .ZN(po1102));
  OAI21_X1   g35349(.A1(pi0782), .A2(new_n5800_), .B(new_n38591_), .ZN(po1103));
  XOR2_X1    g35350(.A1(pi0266), .A2(pi0992), .Z(po1104));
  NAND2_X1   g35351(.A1(pi0949), .A2(pi0954), .ZN(new_n38682_));
  OAI21_X1   g35352(.A1(pi0313), .A2(pi0954), .B(new_n38682_), .ZN(po1105));
  NOR3_X1    g35353(.A1(new_n6940_), .A2(new_n2721_), .A3(new_n2979_), .ZN(po1107));
  OAI21_X1   g35354(.A1(new_n2727_), .A2(new_n2979_), .B(new_n6349_), .ZN(po1112));
  NOR2_X1    g35355(.A1(new_n6045_), .A2(pi0782), .ZN(po1115));
  NOR2_X1    g35356(.A1(new_n5394_), .A2(pi0230), .ZN(po1116));
  NOR2_X1    g35357(.A1(new_n6100_), .A2(pi0782), .ZN(po1118));
  NOR2_X1    g35358(.A1(new_n5395_), .A2(pi0230), .ZN(po1122));
  NOR2_X1    g35359(.A1(new_n5387_), .A2(pi0230), .ZN(po1124));
  NOR2_X1    g35360(.A1(new_n5446_), .A2(pi0782), .ZN(po1125));
  NOR2_X1    g35361(.A1(new_n5388_), .A2(pi0230), .ZN(po1126));
  NOR2_X1    g35362(.A1(new_n5447_), .A2(pi0782), .ZN(po1127));
  NOR2_X1    g35363(.A1(new_n5389_), .A2(pi0230), .ZN(po1128));
  NOR2_X1    g35364(.A1(new_n5448_), .A2(pi0782), .ZN(po1129));
  NOR2_X1    g35365(.A1(new_n5390_), .A2(pi0230), .ZN(po1131));
  NOR2_X1    g35366(.A1(new_n5449_), .A2(pi0782), .ZN(po1132));
  NAND2_X1   g35367(.A1(new_n36910_), .A2(pi0615), .ZN(po1133));
  NOR2_X1    g35368(.A1(new_n5683_), .A2(new_n2979_), .ZN(po1135));
  NAND2_X1   g35369(.A1(new_n36942_), .A2(new_n37034_), .ZN(po1137));
  INV_X1     g35370(.I(pi0825), .ZN(po1147));
  INV_X1     g35371(.I(pi0826), .ZN(po1148));
  INV_X1     g35372(.I(pi0827), .ZN(po1178));
  INV_X1     g35373(.I(pi0828), .ZN(po1182));
  assign     po0166 = 1'b1;
  BUF_X16    g35374(.I(pi0668), .Z(po0000));
  BUF_X16    g35375(.I(pi0672), .Z(po0001));
  BUF_X16    g35376(.I(pi0664), .Z(po0002));
  BUF_X16    g35377(.I(pi0667), .Z(po0003));
  BUF_X16    g35378(.I(pi0676), .Z(po0004));
  BUF_X16    g35379(.I(pi0673), .Z(po0005));
  BUF_X16    g35380(.I(pi0675), .Z(po0006));
  BUF_X16    g35381(.I(pi0666), .Z(po0007));
  BUF_X16    g35382(.I(pi0679), .Z(po0008));
  BUF_X16    g35383(.I(pi0674), .Z(po0009));
  BUF_X16    g35384(.I(pi0663), .Z(po0010));
  BUF_X16    g35385(.I(pi0670), .Z(po0011));
  BUF_X16    g35386(.I(pi0677), .Z(po0012));
  BUF_X16    g35387(.I(pi0682), .Z(po0013));
  BUF_X16    g35388(.I(pi0671), .Z(po0014));
  BUF_X16    g35389(.I(pi0678), .Z(po0015));
  BUF_X16    g35390(.I(pi0718), .Z(po0016));
  BUF_X16    g35391(.I(pi0707), .Z(po0017));
  BUF_X16    g35392(.I(pi0708), .Z(po0018));
  BUF_X16    g35393(.I(pi0713), .Z(po0019));
  BUF_X16    g35394(.I(pi0711), .Z(po0020));
  BUF_X16    g35395(.I(pi0716), .Z(po0021));
  BUF_X16    g35396(.I(pi0733), .Z(po0022));
  BUF_X16    g35397(.I(pi0712), .Z(po0023));
  BUF_X16    g35398(.I(pi0689), .Z(po0024));
  BUF_X16    g35399(.I(pi0717), .Z(po0025));
  BUF_X16    g35400(.I(pi0692), .Z(po0026));
  BUF_X16    g35401(.I(pi0719), .Z(po0027));
  BUF_X16    g35402(.I(pi0722), .Z(po0028));
  BUF_X16    g35403(.I(pi0714), .Z(po0029));
  BUF_X16    g35404(.I(pi0720), .Z(po0030));
  BUF_X16    g35405(.I(pi0685), .Z(po0031));
  BUF_X16    g35406(.I(pi0837), .Z(po0032));
  BUF_X16    g35407(.I(pi0850), .Z(po0033));
  BUF_X16    g35408(.I(pi0872), .Z(po0034));
  BUF_X16    g35409(.I(pi0871), .Z(po0035));
  BUF_X16    g35410(.I(pi0881), .Z(po0036));
  BUF_X16    g35411(.I(pi0866), .Z(po0037));
  BUF_X16    g35412(.I(pi0876), .Z(po0038));
  BUF_X16    g35413(.I(pi0873), .Z(po0039));
  BUF_X16    g35414(.I(pi0874), .Z(po0040));
  BUF_X16    g35415(.I(pi0859), .Z(po0041));
  BUF_X16    g35416(.I(pi0855), .Z(po0042));
  BUF_X16    g35417(.I(pi0852), .Z(po0043));
  BUF_X16    g35418(.I(pi0870), .Z(po0044));
  BUF_X16    g35419(.I(pi0848), .Z(po0045));
  BUF_X16    g35420(.I(pi0865), .Z(po0046));
  BUF_X16    g35421(.I(pi0856), .Z(po0047));
  BUF_X16    g35422(.I(pi0853), .Z(po0048));
  BUF_X16    g35423(.I(pi0847), .Z(po0049));
  BUF_X16    g35424(.I(pi0857), .Z(po0050));
  BUF_X16    g35425(.I(pi0854), .Z(po0051));
  BUF_X16    g35426(.I(pi0858), .Z(po0052));
  BUF_X16    g35427(.I(pi0845), .Z(po0053));
  BUF_X16    g35428(.I(pi0838), .Z(po0054));
  BUF_X16    g35429(.I(pi0842), .Z(po0055));
  BUF_X16    g35430(.I(pi0843), .Z(po0056));
  BUF_X16    g35431(.I(pi0839), .Z(po0057));
  BUF_X16    g35432(.I(pi0844), .Z(po0058));
  BUF_X16    g35433(.I(pi0868), .Z(po0059));
  BUF_X16    g35434(.I(pi0851), .Z(po0060));
  BUF_X16    g35435(.I(pi0867), .Z(po0061));
  BUF_X16    g35436(.I(pi0880), .Z(po0062));
  BUF_X16    g35437(.I(pi0860), .Z(po0063));
  BUF_X16    g35438(.I(pi1030), .Z(po0064));
  BUF_X16    g35439(.I(pi1034), .Z(po0065));
  BUF_X16    g35440(.I(pi1015), .Z(po0066));
  BUF_X16    g35441(.I(pi1020), .Z(po0067));
  BUF_X16    g35442(.I(pi1025), .Z(po0068));
  BUF_X16    g35443(.I(pi1005), .Z(po0069));
  BUF_X16    g35444(.I(pi0996), .Z(po0070));
  BUF_X16    g35445(.I(pi1012), .Z(po0071));
  BUF_X16    g35446(.I(pi0993), .Z(po0072));
  BUF_X16    g35447(.I(pi1016), .Z(po0073));
  BUF_X16    g35448(.I(pi1021), .Z(po0074));
  BUF_X16    g35449(.I(pi1010), .Z(po0075));
  BUF_X16    g35450(.I(pi1027), .Z(po0076));
  BUF_X16    g35451(.I(pi1018), .Z(po0077));
  BUF_X16    g35452(.I(pi1017), .Z(po0078));
  BUF_X16    g35453(.I(pi1024), .Z(po0079));
  BUF_X16    g35454(.I(pi1009), .Z(po0080));
  BUF_X16    g35455(.I(pi1032), .Z(po0081));
  BUF_X16    g35456(.I(pi1003), .Z(po0082));
  BUF_X16    g35457(.I(pi0997), .Z(po0083));
  BUF_X16    g35458(.I(pi1013), .Z(po0084));
  BUF_X16    g35459(.I(pi1011), .Z(po0085));
  BUF_X16    g35460(.I(pi1008), .Z(po0086));
  BUF_X16    g35461(.I(pi1019), .Z(po0087));
  BUF_X16    g35462(.I(pi1031), .Z(po0088));
  BUF_X16    g35463(.I(pi1022), .Z(po0089));
  BUF_X16    g35464(.I(pi1000), .Z(po0090));
  BUF_X16    g35465(.I(pi1023), .Z(po0091));
  BUF_X16    g35466(.I(pi1002), .Z(po0092));
  BUF_X16    g35467(.I(pi1026), .Z(po0093));
  BUF_X16    g35468(.I(pi1006), .Z(po0094));
  BUF_X16    g35469(.I(pi0998), .Z(po0095));
  BUF_X16    g35470(.I(pi0031), .Z(po0096));
  BUF_X16    g35471(.I(pi0080), .Z(po0097));
  BUF_X16    g35472(.I(pi0893), .Z(po0098));
  BUF_X16    g35473(.I(pi0467), .Z(po0099));
  BUF_X16    g35474(.I(pi0078), .Z(po0100));
  BUF_X16    g35475(.I(pi0112), .Z(po0101));
  BUF_X16    g35476(.I(pi0013), .Z(po0102));
  BUF_X16    g35477(.I(pi0025), .Z(po0103));
  BUF_X16    g35478(.I(pi0226), .Z(po0104));
  BUF_X16    g35479(.I(pi0127), .Z(po0105));
  BUF_X16    g35480(.I(pi0822), .Z(po0106));
  BUF_X16    g35481(.I(pi0808), .Z(po0107));
  BUF_X16    g35482(.I(pi0227), .Z(po0108));
  BUF_X16    g35483(.I(pi0477), .Z(po0109));
  BUF_X16    g35484(.I(pi0834), .Z(po0110));
  BUF_X16    g35485(.I(pi0229), .Z(po0111));
  BUF_X16    g35486(.I(pi0012), .Z(po0112));
  BUF_X16    g35487(.I(pi0011), .Z(po0113));
  BUF_X16    g35488(.I(pi0010), .Z(po0114));
  BUF_X16    g35489(.I(pi0009), .Z(po0115));
  BUF_X16    g35490(.I(pi0008), .Z(po0116));
  BUF_X16    g35491(.I(pi0007), .Z(po0117));
  BUF_X16    g35492(.I(pi0006), .Z(po0118));
  BUF_X16    g35493(.I(pi0005), .Z(po0119));
  BUF_X16    g35494(.I(pi0004), .Z(po0120));
  BUF_X16    g35495(.I(pi0003), .Z(po0121));
  BUF_X16    g35496(.I(pi0000), .Z(po0122));
  BUF_X16    g35497(.I(pi0002), .Z(po0123));
  BUF_X16    g35498(.I(pi0001), .Z(po0124));
  BUF_X16    g35499(.I(pi0310), .Z(po0125));
  BUF_X16    g35500(.I(pi0302), .Z(po0126));
  BUF_X16    g35501(.I(pi0475), .Z(po0127));
  BUF_X16    g35502(.I(pi0474), .Z(po0128));
  BUF_X16    g35503(.I(pi0466), .Z(po0129));
  BUF_X16    g35504(.I(pi0473), .Z(po0130));
  BUF_X16    g35505(.I(pi0471), .Z(po0131));
  BUF_X16    g35506(.I(pi0472), .Z(po0132));
  BUF_X16    g35507(.I(pi0470), .Z(po0133));
  BUF_X16    g35508(.I(pi0469), .Z(po0134));
  BUF_X16    g35509(.I(pi0465), .Z(po0135));
  BUF_X16    g35510(.I(pi1028), .Z(po0136));
  BUF_X16    g35511(.I(pi1033), .Z(po0137));
  BUF_X16    g35512(.I(pi0995), .Z(po0138));
  BUF_X16    g35513(.I(pi0994), .Z(po0139));
  BUF_X16    g35514(.I(pi0028), .Z(po0140));
  BUF_X16    g35515(.I(pi0027), .Z(po0141));
  BUF_X16    g35516(.I(pi0026), .Z(po0142));
  BUF_X16    g35517(.I(pi0029), .Z(po0143));
  BUF_X16    g35518(.I(pi0015), .Z(po0144));
  BUF_X16    g35519(.I(pi0014), .Z(po0145));
  BUF_X16    g35520(.I(pi0021), .Z(po0146));
  BUF_X16    g35521(.I(pi0020), .Z(po0147));
  BUF_X16    g35522(.I(pi0019), .Z(po0148));
  BUF_X16    g35523(.I(pi0018), .Z(po0149));
  BUF_X16    g35524(.I(pi0017), .Z(po0150));
  BUF_X16    g35525(.I(pi0016), .Z(po0151));
  BUF_X16    g35526(.I(pi1096), .Z(po0152));
  BUF_X16    g35527(.I(pi0228), .Z(po0168));
  BUF_X16    g35528(.I(pi0022), .Z(po0169));
  BUF_X16    g35529(.I(pi1089), .Z(po0179));
  BUF_X16    g35530(.I(pi0023), .Z(po0180));
  OAI22_X1   g35531(.A1(new_n5543_), .A2(new_n5545_), .B1(new_n5371_), .B2(new_n5548_), .ZN(po0181));
  BUF_X16    g35532(.I(pi0037), .Z(po0188));
  BUF_X16    g35533(.I(pi0117), .Z(po0263));
  BUF_X16    g35534(.I(pi0131), .Z(po0285));
  BUF_X16    g35535(.I(pi0232), .Z(po0386));
  BUF_X16    g35536(.I(pi0236), .Z(po0388));
  BUF_X16    g35537(.I(pi0583), .Z(po0636));
  BUF_X16    g35538(.I(pi0067), .Z(po1053));
  BUF_X16    g35539(.I(pi1134), .Z(po1108));
  BUF_X16    g35540(.I(pi0964), .Z(po1109));
  BUF_X16    g35541(.I(pi0965), .Z(po1111));
  BUF_X16    g35542(.I(pi0991), .Z(po1113));
  BUF_X16    g35543(.I(pi0985), .Z(po1114));
  BUF_X16    g35544(.I(pi1014), .Z(po1117));
  BUF_X16    g35545(.I(pi1029), .Z(po1119));
  BUF_X16    g35546(.I(pi1004), .Z(po1120));
  BUF_X16    g35547(.I(pi1007), .Z(po1121));
  BUF_X16    g35548(.I(pi1135), .Z(po1123));
  BUF_X16    g35549(.I(pi1064), .Z(po1134));
  BUF_X16    g35550(.I(pi0299), .Z(po1136));
  BUF_X16    g35551(.I(pi1075), .Z(po1138));
  BUF_X16    g35552(.I(pi1052), .Z(po1139));
  BUF_X16    g35553(.I(pi0771), .Z(po1140));
  BUF_X16    g35554(.I(pi0765), .Z(po1141));
  BUF_X16    g35555(.I(pi0605), .Z(po1142));
  BUF_X16    g35556(.I(pi0601), .Z(po1143));
  BUF_X16    g35557(.I(pi0278), .Z(po1144));
  BUF_X16    g35558(.I(pi0279), .Z(po1145));
  BUF_X16    g35559(.I(pi1095), .Z(po1152));
  BUF_X16    g35560(.I(pi1094), .Z(po1154));
  BUF_X16    g35561(.I(pi1187), .Z(po1184));
  BUF_X16    g35562(.I(pi1172), .Z(po1185));
  BUF_X16    g35563(.I(pi1170), .Z(po1186));
  BUF_X16    g35564(.I(pi1138), .Z(po1187));
  BUF_X16    g35565(.I(pi1177), .Z(po1188));
  BUF_X16    g35566(.I(pi1178), .Z(po1189));
  BUF_X16    g35567(.I(pi0863), .Z(po1190));
  BUF_X16    g35568(.I(pi1203), .Z(po1191));
  BUF_X16    g35569(.I(pi1185), .Z(po1192));
  BUF_X16    g35570(.I(pi1171), .Z(po1193));
  BUF_X16    g35571(.I(pi1192), .Z(po1194));
  BUF_X16    g35572(.I(pi1137), .Z(po1195));
  BUF_X16    g35573(.I(pi1186), .Z(po1196));
  BUF_X16    g35574(.I(pi1165), .Z(po1197));
  BUF_X16    g35575(.I(pi1164), .Z(po1198));
  BUF_X16    g35576(.I(pi1098), .Z(po1199));
  BUF_X16    g35577(.I(pi1183), .Z(po1200));
  BUF_X16    g35578(.I(pi0230), .Z(po1201));
  BUF_X16    g35579(.I(pi1169), .Z(po1202));
  BUF_X16    g35580(.I(pi1136), .Z(po1203));
  BUF_X16    g35581(.I(pi1181), .Z(po1204));
  BUF_X16    g35582(.I(pi0849), .Z(po1205));
  BUF_X16    g35583(.I(pi1193), .Z(po1206));
  BUF_X16    g35584(.I(pi1182), .Z(po1207));
  BUF_X16    g35585(.I(pi1168), .Z(po1208));
  BUF_X16    g35586(.I(pi1175), .Z(po1209));
  BUF_X16    g35587(.I(pi1191), .Z(po1210));
  BUF_X16    g35588(.I(pi1099), .Z(po1211));
  BUF_X16    g35589(.I(pi1174), .Z(po1212));
  BUF_X16    g35590(.I(pi1179), .Z(po1213));
  BUF_X16    g35591(.I(pi1202), .Z(po1214));
  BUF_X16    g35592(.I(pi1176), .Z(po1215));
  BUF_X16    g35593(.I(pi1173), .Z(po1216));
  BUF_X16    g35594(.I(pi1201), .Z(po1217));
  BUF_X16    g35595(.I(pi1167), .Z(po1218));
  BUF_X16    g35596(.I(pi0840), .Z(po1219));
  BUF_X16    g35597(.I(pi1189), .Z(po1220));
  BUF_X16    g35598(.I(pi1195), .Z(po1221));
  BUF_X16    g35599(.I(pi0864), .Z(po1222));
  BUF_X16    g35600(.I(pi1190), .Z(po1223));
  BUF_X16    g35601(.I(pi1188), .Z(po1224));
  BUF_X16    g35602(.I(pi1180), .Z(po1225));
  BUF_X16    g35603(.I(pi1194), .Z(po1226));
  BUF_X16    g35604(.I(pi1097), .Z(po1227));
  BUF_X16    g35605(.I(pi1166), .Z(po1228));
  BUF_X16    g35606(.I(pi1200), .Z(po1229));
  BUF_X16    g35607(.I(pi1184), .Z(po1230));
endmodule


