// Benchmark "i2c" written by ABC on Thu Sep 14 22:41:19 2023

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n453_, new_n454_, new_n455_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n479_, new_n480_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n489_, new_n490_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n499_, new_n500_, new_n501_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n525_, new_n526_, new_n527_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n534_, new_n535_, new_n537_, new_n538_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n559_,
    new_n560_, new_n561_, new_n563_, new_n564_, new_n565_, new_n567_,
    new_n568_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n616_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n900_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n955_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n987_, new_n989_, new_n990_, new_n992_,
    new_n994_, new_n995_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1007_, new_n1008_,
    new_n1009_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1031_,
    new_n1032_, new_n1033_, new_n1035_, new_n1036_, new_n1037_, new_n1039_,
    new_n1040_, new_n1041_, new_n1043_, new_n1044_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1064_, new_n1065_, new_n1066_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1073_, new_n1074_,
    new_n1075_, new_n1077_, new_n1078_, new_n1079_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1086_, new_n1087_, new_n1089_, new_n1090_,
    new_n1092_, new_n1093_, new_n1095_, new_n1096_, new_n1098_, new_n1099_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1113_, new_n1115_,
    new_n1117_, new_n1118_, new_n1120_, new_n1121_, new_n1123_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1189_, new_n1190_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1231_, new_n1232_, new_n1234_, new_n1235_, new_n1236_, new_n1238_,
    new_n1240_, new_n1241_, new_n1242_, new_n1244_, new_n1245_, new_n1247_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1256_, new_n1262_,
    new_n1264_;
  INV_X1     g000(.I(pi054), .ZN(new_n291_));
  NOR2_X1    g001(.A1(pi005), .A2(pi022), .ZN(new_n292_));
  NAND2_X1   g002(.A1(new_n292_), .A2(pi056), .ZN(new_n293_));
  INV_X1     g003(.I(pi014), .ZN(new_n294_));
  NOR2_X1    g004(.A1(new_n294_), .A2(pi013), .ZN(new_n295_));
  NOR3_X1    g005(.A1(pi007), .A2(pi008), .A3(pi021), .ZN(new_n296_));
  NAND2_X1   g006(.A1(pi007), .A2(pi013), .ZN(new_n297_));
  NAND3_X1   g007(.A1(new_n296_), .A2(pi014), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1   g008(.A1(pi008), .A2(pi021), .ZN(new_n299_));
  NAND2_X1   g009(.A1(pi013), .A2(pi021), .ZN(new_n300_));
  NAND2_X1   g010(.A1(pi007), .A2(pi008), .ZN(new_n301_));
  XOR2_X1    g011(.A1(new_n300_), .A2(new_n301_), .Z(new_n302_));
  NOR4_X1    g012(.A1(new_n302_), .A2(new_n295_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n303_));
  INV_X1     g013(.I(new_n295_), .ZN(new_n304_));
  INV_X1     g014(.I(new_n298_), .ZN(new_n305_));
  AOI21_X1   g015(.A1(pi013), .A2(pi021), .B(new_n301_), .ZN(new_n306_));
  AOI21_X1   g016(.A1(pi007), .A2(pi008), .B(new_n300_), .ZN(new_n307_));
  NOR3_X1    g017(.A1(new_n307_), .A2(new_n299_), .A3(new_n306_), .ZN(new_n308_));
  AOI21_X1   g018(.A1(new_n308_), .A2(new_n305_), .B(new_n304_), .ZN(new_n309_));
  INV_X1     g019(.I(pi010), .ZN(new_n310_));
  INV_X1     g020(.I(pi006), .ZN(new_n311_));
  INV_X1     g021(.I(pi013), .ZN(new_n312_));
  NOR4_X1    g022(.A1(new_n311_), .A2(new_n312_), .A3(new_n294_), .A4(pi017), .ZN(new_n313_));
  INV_X1     g023(.I(pi012), .ZN(new_n314_));
  NOR4_X1    g024(.A1(new_n310_), .A2(new_n314_), .A3(pi005), .A4(pi022), .ZN(new_n315_));
  INV_X1     g025(.I(pi004), .ZN(new_n316_));
  INV_X1     g026(.I(pi016), .ZN(new_n317_));
  INV_X1     g027(.I(pi018), .ZN(new_n318_));
  INV_X1     g028(.I(pi019), .ZN(new_n319_));
  NOR4_X1    g029(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .A4(new_n319_), .ZN(new_n320_));
  NAND4_X1   g030(.A1(new_n320_), .A2(new_n313_), .A3(new_n315_), .A4(new_n296_), .ZN(new_n321_));
  NOR2_X1    g031(.A1(pi009), .A2(pi011), .ZN(new_n322_));
  XNOR2_X1   g032(.A1(new_n322_), .A2(pi056), .ZN(new_n323_));
  AOI21_X1   g033(.A1(new_n321_), .A2(new_n310_), .B(new_n323_), .ZN(new_n324_));
  OAI21_X1   g034(.A1(new_n309_), .A2(new_n303_), .B(new_n324_), .ZN(new_n325_));
  AOI21_X1   g035(.A1(new_n325_), .A2(new_n293_), .B(new_n291_), .ZN(new_n326_));
  NAND4_X1   g036(.A1(new_n292_), .A2(new_n322_), .A3(pi006), .A4(pi007), .ZN(new_n327_));
  NOR3_X1    g037(.A1(pi008), .A2(pi017), .A3(pi021), .ZN(new_n328_));
  NOR2_X1    g038(.A1(new_n314_), .A2(pi013), .ZN(new_n329_));
  NAND4_X1   g039(.A1(new_n320_), .A2(new_n294_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  NOR2_X1    g040(.A1(new_n291_), .A2(pi000), .ZN(new_n331_));
  OAI21_X1   g041(.A1(new_n330_), .A2(new_n327_), .B(new_n331_), .ZN(new_n332_));
  NOR2_X1    g042(.A1(pi003), .A2(pi129), .ZN(new_n333_));
  OAI21_X1   g043(.A1(new_n326_), .A2(new_n332_), .B(new_n333_), .ZN(po015));
  INV_X1     g044(.I(pi001), .ZN(new_n335_));
  NOR2_X1    g045(.A1(new_n312_), .A2(pi007), .ZN(new_n336_));
  NOR3_X1    g046(.A1(pi005), .A2(pi006), .A3(pi012), .ZN(new_n337_));
  NAND2_X1   g047(.A1(pi005), .A2(pi007), .ZN(new_n338_));
  NAND3_X1   g048(.A1(new_n337_), .A2(pi013), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1    g049(.A1(pi006), .A2(pi012), .Z(new_n340_));
  NAND2_X1   g050(.A1(pi007), .A2(pi012), .ZN(new_n341_));
  NAND3_X1   g051(.A1(new_n341_), .A2(pi005), .A3(pi006), .ZN(new_n342_));
  NAND2_X1   g052(.A1(pi005), .A2(pi006), .ZN(new_n343_));
  NAND3_X1   g053(.A1(new_n343_), .A2(pi007), .A3(pi012), .ZN(new_n344_));
  NAND3_X1   g054(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1   g055(.A1(new_n345_), .A2(new_n339_), .B(new_n336_), .ZN(new_n346_));
  INV_X1     g056(.I(new_n336_), .ZN(new_n347_));
  XNOR2_X1   g057(.A1(pi006), .A2(pi012), .ZN(new_n348_));
  AOI21_X1   g058(.A1(pi007), .A2(pi012), .B(new_n343_), .ZN(new_n349_));
  AOI21_X1   g059(.A1(pi005), .A2(pi006), .B(new_n341_), .ZN(new_n350_));
  NOR4_X1    g060(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .A4(new_n339_), .ZN(new_n351_));
  NOR4_X1    g061(.A1(new_n291_), .A2(pi010), .A3(pi014), .A4(pi022), .ZN(new_n352_));
  INV_X1     g062(.I(pi017), .ZN(new_n353_));
  INV_X1     g063(.I(pi021), .ZN(new_n354_));
  NAND2_X1   g064(.A1(pi008), .A2(pi011), .ZN(new_n355_));
  NOR3_X1    g065(.A1(new_n355_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n356_));
  NAND3_X1   g066(.A1(new_n320_), .A2(new_n356_), .A3(new_n352_), .ZN(new_n357_));
  AOI21_X1   g067(.A1(new_n351_), .A2(new_n347_), .B(new_n357_), .ZN(new_n358_));
  NAND4_X1   g068(.A1(new_n320_), .A2(new_n356_), .A3(new_n352_), .A4(pi009), .ZN(new_n359_));
  AOI21_X1   g069(.A1(new_n358_), .A2(new_n346_), .B(new_n359_), .ZN(new_n360_));
  INV_X1     g070(.I(new_n339_), .ZN(new_n361_));
  NOR3_X1    g071(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n362_));
  AOI21_X1   g072(.A1(new_n362_), .A2(new_n361_), .B(new_n347_), .ZN(new_n363_));
  NOR3_X1    g073(.A1(new_n345_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n364_));
  NOR4_X1    g074(.A1(new_n363_), .A2(pi009), .A3(new_n364_), .A4(new_n357_), .ZN(new_n365_));
  INV_X1     g075(.I(new_n333_), .ZN(new_n366_));
  NOR2_X1    g076(.A1(pi007), .A2(pi013), .ZN(new_n367_));
  NAND2_X1   g077(.A1(new_n337_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1    g078(.A1(new_n368_), .A2(new_n366_), .ZN(new_n369_));
  OAI21_X1   g079(.A1(new_n360_), .A2(new_n365_), .B(new_n369_), .ZN(new_n370_));
  NAND4_X1   g080(.A1(pi005), .A2(pi006), .A3(pi007), .A4(pi013), .ZN(new_n371_));
  NOR2_X1    g081(.A1(pi008), .A2(pi021), .ZN(new_n372_));
  NOR2_X1    g082(.A1(pi011), .A2(pi012), .ZN(new_n373_));
  INV_X1     g083(.I(new_n373_), .ZN(new_n374_));
  NOR3_X1    g084(.A1(new_n374_), .A2(pi010), .A3(pi022), .ZN(new_n375_));
  NAND4_X1   g085(.A1(new_n375_), .A2(pi014), .A3(new_n320_), .A4(new_n372_), .ZN(new_n376_));
  NOR2_X1    g086(.A1(new_n291_), .A2(pi017), .ZN(new_n377_));
  OAI21_X1   g087(.A1(new_n376_), .A2(new_n371_), .B(new_n377_), .ZN(new_n378_));
  AOI21_X1   g088(.A1(new_n370_), .A2(new_n335_), .B(new_n378_), .ZN(po016));
  INV_X1     g089(.I(pi002), .ZN(new_n380_));
  NOR3_X1    g090(.A1(pi015), .A2(pi020), .A3(pi049), .ZN(new_n381_));
  NOR2_X1    g091(.A1(pi047), .A2(pi048), .ZN(new_n382_));
  INV_X1     g092(.I(pi024), .ZN(new_n383_));
  INV_X1     g093(.I(pi045), .ZN(new_n384_));
  NOR2_X1    g094(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1   g095(.A1(new_n385_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n386_));
  NAND2_X1   g096(.A1(new_n386_), .A2(pi082), .ZN(new_n387_));
  INV_X1     g097(.I(pi043), .ZN(new_n388_));
  NAND4_X1   g098(.A1(pi038), .A2(pi040), .A3(pi042), .A4(pi044), .ZN(new_n389_));
  NAND3_X1   g099(.A1(pi041), .A2(pi046), .A3(pi050), .ZN(new_n390_));
  NOR2_X1    g100(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1   g101(.A1(new_n391_), .A2(new_n388_), .ZN(new_n392_));
  NAND2_X1   g102(.A1(pi122), .A2(pi127), .ZN(new_n393_));
  INV_X1     g103(.I(new_n393_), .ZN(new_n394_));
  NAND2_X1   g104(.A1(new_n394_), .A2(pi082), .ZN(new_n395_));
  NOR2_X1    g105(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  XOR2_X1    g106(.A1(new_n396_), .A2(new_n387_), .Z(new_n397_));
  INV_X1     g107(.I(pi082), .ZN(new_n398_));
  INV_X1     g108(.I(pi129), .ZN(new_n399_));
  NOR3_X1    g109(.A1(new_n398_), .A2(new_n399_), .A3(pi048), .ZN(new_n400_));
  NOR2_X1    g110(.A1(pi002), .A2(pi045), .ZN(new_n401_));
  INV_X1     g111(.I(new_n401_), .ZN(new_n402_));
  NOR3_X1    g112(.A1(new_n402_), .A2(pi043), .A3(pi047), .ZN(new_n403_));
  INV_X1     g113(.I(pi065), .ZN(new_n404_));
  NAND4_X1   g114(.A1(pi038), .A2(pi041), .A3(pi046), .A4(pi050), .ZN(new_n405_));
  AOI21_X1   g115(.A1(new_n404_), .A2(new_n393_), .B(new_n405_), .ZN(new_n406_));
  INV_X1     g116(.I(pi044), .ZN(new_n407_));
  NOR2_X1    g117(.A1(pi040), .A2(pi042), .ZN(new_n408_));
  NAND2_X1   g118(.A1(new_n408_), .A2(new_n407_), .ZN(new_n409_));
  INV_X1     g119(.I(pi015), .ZN(new_n410_));
  INV_X1     g120(.I(pi020), .ZN(new_n411_));
  INV_X1     g121(.I(pi049), .ZN(new_n412_));
  NOR4_X1    g122(.A1(new_n410_), .A2(new_n411_), .A3(new_n383_), .A4(new_n412_), .ZN(new_n413_));
  INV_X1     g123(.I(new_n413_), .ZN(new_n414_));
  NOR2_X1    g124(.A1(new_n414_), .A2(new_n409_), .ZN(new_n415_));
  NAND4_X1   g125(.A1(new_n415_), .A2(new_n400_), .A3(new_n403_), .A4(new_n406_), .ZN(new_n416_));
  AOI21_X1   g126(.A1(new_n380_), .A2(new_n416_), .B(new_n397_), .ZN(po017));
  INV_X1     g127(.I(new_n320_), .ZN(new_n418_));
  NAND4_X1   g128(.A1(new_n373_), .A2(pi008), .A3(pi017), .A4(pi021), .ZN(new_n419_));
  NOR4_X1    g129(.A1(pi009), .A2(pi010), .A3(pi014), .A4(pi022), .ZN(new_n420_));
  INV_X1     g130(.I(new_n420_), .ZN(new_n421_));
  NOR3_X1    g131(.A1(new_n418_), .A2(new_n419_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1     g132(.I(pi113), .ZN(new_n423_));
  INV_X1     g133(.I(pi123), .ZN(new_n424_));
  NAND3_X1   g134(.A1(new_n423_), .A2(new_n424_), .A3(pi000), .ZN(new_n425_));
  NOR2_X1    g135(.A1(pi061), .A2(pi118), .ZN(new_n426_));
  AOI21_X1   g136(.A1(new_n425_), .A2(new_n426_), .B(new_n371_), .ZN(new_n427_));
  AOI21_X1   g137(.A1(new_n422_), .A2(new_n427_), .B(pi129), .ZN(po018));
  INV_X1     g138(.I(new_n368_), .ZN(new_n429_));
  INV_X1     g139(.I(new_n356_), .ZN(new_n430_));
  NOR3_X1    g140(.A1(new_n418_), .A2(new_n430_), .A3(new_n291_), .ZN(new_n431_));
  INV_X1     g141(.I(pi009), .ZN(new_n432_));
  INV_X1     g142(.I(pi022), .ZN(new_n433_));
  NOR2_X1    g143(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NOR3_X1    g144(.A1(new_n366_), .A2(new_n310_), .A3(new_n294_), .ZN(new_n435_));
  NAND4_X1   g145(.A1(new_n431_), .A2(new_n429_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  AOI21_X1   g146(.A1(new_n436_), .A2(new_n316_), .B(new_n291_), .ZN(po019));
  INV_X1     g147(.I(pi005), .ZN(new_n438_));
  NAND2_X1   g148(.A1(new_n420_), .A2(new_n312_), .ZN(new_n439_));
  NAND2_X1   g149(.A1(new_n317_), .A2(pi054), .ZN(new_n440_));
  NOR4_X1    g150(.A1(new_n430_), .A2(pi059), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  NAND4_X1   g151(.A1(pi005), .A2(pi006), .A3(pi007), .A4(pi012), .ZN(new_n442_));
  INV_X1     g152(.I(new_n442_), .ZN(new_n443_));
  NOR2_X1    g153(.A1(pi004), .A2(pi019), .ZN(new_n444_));
  NAND2_X1   g154(.A1(new_n444_), .A2(new_n318_), .ZN(new_n445_));
  INV_X1     g155(.I(new_n445_), .ZN(new_n446_));
  INV_X1     g156(.I(pi025), .ZN(new_n447_));
  INV_X1     g157(.I(pi028), .ZN(new_n448_));
  INV_X1     g158(.I(pi029), .ZN(new_n449_));
  NOR4_X1    g159(.A1(new_n366_), .A2(new_n447_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND4_X1   g160(.A1(new_n441_), .A2(new_n443_), .A3(new_n446_), .A4(new_n450_), .ZN(new_n451_));
  AOI21_X1   g161(.A1(new_n451_), .A2(new_n438_), .B(new_n291_), .ZN(po020));
  NOR3_X1    g162(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n453_));
  NOR2_X1    g163(.A1(new_n366_), .A2(new_n447_), .ZN(new_n454_));
  NAND4_X1   g164(.A1(new_n441_), .A2(new_n443_), .A3(new_n453_), .A4(new_n454_), .ZN(new_n455_));
  AOI21_X1   g165(.A1(new_n455_), .A2(new_n311_), .B(new_n291_), .ZN(po021));
  INV_X1     g166(.I(pi007), .ZN(new_n457_));
  INV_X1     g167(.I(new_n439_), .ZN(new_n458_));
  NAND2_X1   g168(.A1(new_n318_), .A2(new_n354_), .ZN(new_n459_));
  NAND2_X1   g169(.A1(pi005), .A2(pi017), .ZN(new_n460_));
  NOR4_X1    g170(.A1(new_n366_), .A2(new_n459_), .A3(new_n301_), .A4(new_n460_), .ZN(new_n461_));
  NAND3_X1   g171(.A1(new_n444_), .A2(new_n317_), .A3(pi054), .ZN(new_n462_));
  NOR3_X1    g172(.A1(new_n462_), .A2(pi006), .A3(new_n374_), .ZN(new_n463_));
  NAND3_X1   g173(.A1(new_n458_), .A2(new_n463_), .A3(new_n461_), .ZN(new_n464_));
  AOI21_X1   g174(.A1(new_n464_), .A2(new_n457_), .B(new_n291_), .ZN(po022));
  INV_X1     g175(.I(pi008), .ZN(new_n466_));
  INV_X1     g176(.I(new_n462_), .ZN(new_n467_));
  NOR2_X1    g177(.A1(new_n421_), .A2(new_n368_), .ZN(new_n468_));
  NAND3_X1   g178(.A1(new_n333_), .A2(new_n353_), .A3(new_n318_), .ZN(new_n469_));
  NOR4_X1    g179(.A1(new_n469_), .A2(pi008), .A3(pi011), .A4(new_n354_), .ZN(new_n470_));
  NAND3_X1   g180(.A1(new_n470_), .A2(new_n468_), .A3(new_n467_), .ZN(new_n471_));
  AOI21_X1   g181(.A1(new_n471_), .A2(new_n466_), .B(new_n291_), .ZN(po023));
  NAND4_X1   g182(.A1(pi009), .A2(pi011), .A3(pi013), .A4(pi014), .ZN(new_n473_));
  NOR4_X1    g183(.A1(new_n366_), .A2(new_n473_), .A3(pi010), .A4(pi022), .ZN(new_n474_));
  NAND4_X1   g184(.A1(pi008), .A2(pi017), .A3(pi018), .A4(pi021), .ZN(new_n475_));
  NOR2_X1    g185(.A1(new_n462_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1   g186(.A1(new_n474_), .A2(new_n476_), .A3(new_n443_), .ZN(new_n477_));
  AOI21_X1   g187(.A1(new_n477_), .A2(new_n432_), .B(new_n291_), .ZN(po024));
  INV_X1     g188(.I(new_n475_), .ZN(new_n479_));
  NOR4_X1    g189(.A1(new_n374_), .A2(pi005), .A3(pi006), .A4(pi007), .ZN(new_n480_));
  NOR2_X1    g190(.A1(new_n310_), .A2(new_n291_), .ZN(po025));
  INV_X1     g191(.I(pi011), .ZN(new_n484_));
  NAND3_X1   g192(.A1(pi010), .A2(pi011), .A3(pi022), .ZN(new_n485_));
  NOR4_X1    g193(.A1(new_n366_), .A2(pi009), .A3(pi014), .A4(new_n485_), .ZN(new_n486_));
  NAND3_X1   g194(.A1(new_n476_), .A2(new_n486_), .A3(new_n429_), .ZN(new_n487_));
  AOI21_X1   g195(.A1(new_n487_), .A2(new_n484_), .B(new_n291_), .ZN(po026));
  NOR4_X1    g196(.A1(new_n366_), .A2(new_n374_), .A3(new_n371_), .A4(new_n318_), .ZN(new_n489_));
  NAND4_X1   g197(.A1(new_n489_), .A2(new_n328_), .A3(new_n467_), .A4(new_n420_), .ZN(new_n490_));
  AOI21_X1   g198(.A1(new_n490_), .A2(new_n314_), .B(new_n291_), .ZN(po027));
  NAND3_X1   g199(.A1(new_n447_), .A2(new_n448_), .A3(pi029), .ZN(new_n492_));
  NOR3_X1    g200(.A1(new_n421_), .A2(new_n445_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1     g201(.I(new_n367_), .ZN(new_n494_));
  NAND2_X1   g202(.A1(new_n333_), .A2(pi059), .ZN(new_n495_));
  NOR3_X1    g203(.A1(new_n495_), .A2(new_n494_), .A3(new_n440_), .ZN(new_n496_));
  NAND4_X1   g204(.A1(new_n493_), .A2(new_n496_), .A3(new_n337_), .A4(new_n356_), .ZN(new_n497_));
  AOI21_X1   g205(.A1(new_n497_), .A2(new_n312_), .B(new_n291_), .ZN(po028));
  NAND2_X1   g206(.A1(new_n333_), .A2(new_n444_), .ZN(new_n499_));
  NOR4_X1    g207(.A1(new_n499_), .A2(new_n432_), .A3(new_n312_), .A4(new_n317_), .ZN(new_n500_));
  NAND4_X1   g208(.A1(new_n500_), .A2(new_n352_), .A3(new_n480_), .A4(new_n479_), .ZN(new_n501_));
  AOI21_X1   g209(.A1(new_n501_), .A2(new_n294_), .B(new_n291_), .ZN(po029));
  NOR3_X1    g210(.A1(pi038), .A2(pi046), .A3(pi050), .ZN(new_n503_));
  NAND3_X1   g211(.A1(new_n503_), .A2(new_n408_), .A3(new_n407_), .ZN(new_n504_));
  NOR2_X1    g212(.A1(pi024), .A2(pi049), .ZN(new_n505_));
  INV_X1     g213(.I(new_n382_), .ZN(new_n506_));
  NOR3_X1    g214(.A1(new_n506_), .A2(new_n410_), .A3(new_n384_), .ZN(new_n507_));
  INV_X1     g215(.I(pi070), .ZN(new_n508_));
  NAND2_X1   g216(.A1(new_n393_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1     g217(.I(pi041), .ZN(new_n510_));
  NOR3_X1    g218(.A1(new_n510_), .A2(new_n388_), .A3(new_n398_), .ZN(new_n511_));
  NAND4_X1   g219(.A1(new_n507_), .A2(new_n505_), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  NOR2_X1    g220(.A1(new_n394_), .A2(pi015), .ZN(new_n513_));
  OAI21_X1   g221(.A1(new_n512_), .A2(new_n504_), .B(new_n513_), .ZN(new_n514_));
  NOR2_X1    g222(.A1(new_n398_), .A2(new_n399_), .ZN(new_n515_));
  AOI21_X1   g223(.A1(new_n514_), .A2(new_n515_), .B(pi082), .ZN(new_n516_));
  NOR3_X1    g224(.A1(pi043), .A2(pi047), .A3(pi048), .ZN(new_n517_));
  INV_X1     g225(.I(new_n517_), .ZN(new_n518_));
  NAND2_X1   g226(.A1(new_n505_), .A2(new_n384_), .ZN(new_n519_));
  OAI21_X1   g227(.A1(pi024), .A2(pi049), .B(new_n410_), .ZN(new_n520_));
  NAND4_X1   g228(.A1(new_n507_), .A2(new_n520_), .A3(pi002), .A4(pi020), .ZN(new_n521_));
  OAI22_X1   g229(.A1(new_n521_), .A2(new_n392_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n522_));
  NAND2_X1   g230(.A1(new_n522_), .A2(new_n391_), .ZN(new_n523_));
  NOR2_X1    g231(.A1(new_n516_), .A2(new_n523_), .ZN(po030));
  NOR3_X1    g232(.A1(new_n311_), .A2(pi005), .A3(pi012), .ZN(new_n525_));
  NOR2_X1    g233(.A1(new_n366_), .A2(new_n494_), .ZN(new_n526_));
  NAND4_X1   g234(.A1(new_n431_), .A2(new_n420_), .A3(new_n525_), .A4(new_n526_), .ZN(new_n527_));
  AOI21_X1   g235(.A1(new_n527_), .A2(new_n317_), .B(new_n291_), .ZN(po031));
  NAND4_X1   g236(.A1(pi006), .A2(pi007), .A3(pi012), .A4(pi016), .ZN(new_n529_));
  NOR4_X1    g237(.A1(new_n529_), .A2(new_n447_), .A3(new_n291_), .A4(new_n460_), .ZN(new_n530_));
  NOR4_X1    g238(.A1(new_n495_), .A2(pi008), .A3(new_n484_), .A4(pi021), .ZN(new_n531_));
  NAND4_X1   g239(.A1(new_n531_), .A2(new_n458_), .A3(new_n453_), .A4(new_n530_), .ZN(new_n532_));
  AOI21_X1   g240(.A1(new_n532_), .A2(new_n353_), .B(new_n291_), .ZN(po032));
  NOR3_X1    g241(.A1(new_n366_), .A2(new_n317_), .A3(new_n291_), .ZN(new_n534_));
  NAND4_X1   g242(.A1(new_n468_), .A2(new_n356_), .A3(new_n446_), .A4(new_n534_), .ZN(new_n535_));
  AOI21_X1   g243(.A1(new_n535_), .A2(new_n318_), .B(new_n291_), .ZN(po033));
  NOR4_X1    g244(.A1(new_n462_), .A2(new_n353_), .A3(new_n366_), .A4(new_n318_), .ZN(new_n537_));
  NAND4_X1   g245(.A1(new_n537_), .A2(new_n468_), .A3(pi011), .A4(new_n372_), .ZN(new_n538_));
  AOI21_X1   g246(.A1(new_n538_), .A2(new_n319_), .B(new_n291_), .ZN(po034));
  NAND4_X1   g247(.A1(pi041), .A2(pi043), .A3(pi046), .A4(pi047), .ZN(new_n540_));
  INV_X1     g248(.I(new_n540_), .ZN(new_n541_));
  NAND3_X1   g249(.A1(new_n541_), .A2(pi048), .A3(new_n385_), .ZN(new_n542_));
  NOR2_X1    g250(.A1(pi038), .A2(pi050), .ZN(new_n543_));
  NAND2_X1   g251(.A1(new_n408_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1   g252(.A1(new_n381_), .A2(pi044), .ZN(new_n545_));
  NOR3_X1    g253(.A1(new_n542_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1     g254(.I(pi040), .ZN(new_n547_));
  NAND2_X1   g255(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1    g256(.A1(pi042), .A2(pi044), .ZN(new_n549_));
  INV_X1     g257(.I(new_n549_), .ZN(new_n550_));
  NAND2_X1   g258(.A1(new_n410_), .A2(new_n412_), .ZN(new_n551_));
  NOR4_X1    g259(.A1(new_n542_), .A2(new_n548_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  AOI22_X1   g260(.A1(new_n552_), .A2(new_n546_), .B1(pi002), .B2(pi020), .ZN(new_n553_));
  OAI21_X1   g261(.A1(new_n394_), .A2(pi071), .B(pi082), .ZN(new_n554_));
  NOR4_X1    g262(.A1(new_n542_), .A2(new_n544_), .A3(new_n545_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1   g263(.A1(new_n393_), .A2(new_n411_), .ZN(new_n556_));
  OAI21_X1   g264(.A1(new_n555_), .A2(new_n556_), .B(new_n515_), .ZN(new_n557_));
  AOI21_X1   g265(.A1(new_n398_), .A2(new_n557_), .B(new_n553_), .ZN(po035));
  NOR2_X1    g266(.A1(new_n319_), .A2(pi021), .ZN(new_n559_));
  NOR4_X1    g267(.A1(new_n469_), .A2(new_n316_), .A3(new_n317_), .A4(new_n355_), .ZN(new_n560_));
  NAND4_X1   g268(.A1(new_n560_), .A2(new_n468_), .A3(pi054), .A4(new_n559_), .ZN(new_n561_));
  AOI21_X1   g269(.A1(new_n561_), .A2(new_n354_), .B(new_n291_), .ZN(po036));
  NOR4_X1    g270(.A1(new_n475_), .A2(new_n432_), .A3(new_n310_), .A4(new_n433_), .ZN(new_n563_));
  NOR4_X1    g271(.A1(new_n366_), .A2(new_n312_), .A3(new_n294_), .A4(new_n338_), .ZN(new_n564_));
  NAND3_X1   g272(.A1(new_n463_), .A2(new_n564_), .A3(new_n563_), .ZN(new_n565_));
  AOI21_X1   g273(.A1(new_n565_), .A2(new_n433_), .B(new_n291_), .ZN(po037));
  NOR2_X1    g274(.A1(pi061), .A2(pi129), .ZN(new_n567_));
  NAND2_X1   g275(.A1(pi023), .A2(pi055), .ZN(new_n568_));
  NOR2_X1    g276(.A1(new_n567_), .A2(new_n568_), .ZN(po038));
  INV_X1     g277(.I(new_n381_), .ZN(new_n570_));
  NAND3_X1   g278(.A1(new_n392_), .A2(new_n398_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1   g279(.A1(new_n571_), .A2(new_n382_), .A3(new_n401_), .ZN(new_n572_));
  NAND3_X1   g280(.A1(new_n572_), .A2(pi063), .A3(new_n393_), .ZN(new_n573_));
  NAND2_X1   g281(.A1(new_n510_), .A2(new_n388_), .ZN(new_n574_));
  NOR2_X1    g282(.A1(new_n574_), .A2(pi046), .ZN(new_n575_));
  NAND3_X1   g283(.A1(new_n575_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n576_));
  NAND3_X1   g284(.A1(new_n576_), .A2(new_n399_), .A3(new_n548_), .ZN(new_n577_));
  NAND4_X1   g285(.A1(new_n577_), .A2(pi024), .A3(pi082), .A4(new_n549_), .ZN(new_n578_));
  INV_X1     g286(.I(new_n504_), .ZN(new_n579_));
  NOR2_X1    g287(.A1(new_n574_), .A2(pi047), .ZN(new_n580_));
  INV_X1     g288(.I(pi048), .ZN(new_n581_));
  NOR2_X1    g289(.A1(new_n384_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1   g290(.A1(new_n579_), .A2(pi082), .A3(new_n580_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1   g291(.A1(new_n393_), .A2(pi082), .ZN(new_n584_));
  INV_X1     g292(.I(new_n584_), .ZN(new_n585_));
  NAND4_X1   g293(.A1(pi002), .A2(pi015), .A3(pi020), .A4(pi049), .ZN(new_n586_));
  NAND4_X1   g294(.A1(new_n583_), .A2(pi024), .A3(new_n585_), .A4(new_n586_), .ZN(new_n587_));
  AOI21_X1   g295(.A1(new_n573_), .A2(new_n578_), .B(new_n587_), .ZN(po039));
  INV_X1     g296(.I(pi085), .ZN(new_n589_));
  INV_X1     g297(.I(pi100), .ZN(new_n590_));
  INV_X1     g298(.I(pi096), .ZN(new_n591_));
  INV_X1     g299(.I(pi116), .ZN(new_n592_));
  INV_X1     g300(.I(pi110), .ZN(new_n593_));
  NAND4_X1   g301(.A1(new_n591_), .A2(new_n592_), .A3(pi025), .A4(pi085), .ZN(new_n595_));
  OAI21_X1   g302(.A1(new_n589_), .A2(new_n590_), .B(new_n595_), .ZN(new_n596_));
  INV_X1     g303(.I(pi026), .ZN(new_n597_));
  NOR3_X1    g304(.A1(pi039), .A2(pi051), .A3(pi052), .ZN(new_n598_));
  INV_X1     g305(.I(new_n598_), .ZN(new_n599_));
  NOR3_X1    g306(.A1(new_n599_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n600_));
  INV_X1     g307(.I(pi097), .ZN(new_n601_));
  NOR2_X1    g308(.A1(pi095), .A2(pi100), .ZN(new_n602_));
  AOI21_X1   g309(.A1(new_n602_), .A2(new_n593_), .B(new_n601_), .ZN(new_n603_));
  INV_X1     g310(.I(new_n603_), .ZN(new_n604_));
  NOR2_X1    g311(.A1(new_n604_), .A2(new_n589_), .ZN(new_n605_));
  OAI21_X1   g312(.A1(pi025), .A2(new_n600_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1    g313(.A1(new_n447_), .A2(pi116), .ZN(new_n607_));
  NAND2_X1   g314(.A1(new_n607_), .A2(pi027), .ZN(new_n608_));
  OAI21_X1   g315(.A1(new_n606_), .A2(new_n608_), .B(new_n597_), .ZN(new_n609_));
  NAND2_X1   g316(.A1(new_n609_), .A2(new_n596_), .ZN(new_n610_));
  NAND2_X1   g317(.A1(new_n607_), .A2(new_n597_), .ZN(new_n611_));
  INV_X1     g318(.I(new_n611_), .ZN(new_n612_));
  NAND4_X1   g319(.A1(new_n612_), .A2(pi027), .A3(pi053), .A4(pi085), .ZN(new_n613_));
  INV_X1     g320(.I(pi027), .ZN(new_n614_));
  NAND2_X1   g321(.A1(pi027), .A2(pi116), .ZN(new_n616_));
  OAI21_X1   g322(.A1(pi025), .A2(new_n598_), .B(new_n603_), .ZN(new_n618_));
  INV_X1     g323(.I(pi058), .ZN(new_n619_));
  NOR2_X1    g324(.A1(new_n619_), .A2(pi053), .ZN(new_n620_));
  NOR2_X1    g325(.A1(new_n614_), .A2(new_n589_), .ZN(new_n621_));
  NAND3_X1   g326(.A1(new_n621_), .A2(new_n620_), .A3(new_n333_), .ZN(new_n622_));
  OAI21_X1   g327(.A1(new_n622_), .A2(new_n611_), .B(new_n619_), .ZN(new_n623_));
  NOR2_X1    g328(.A1(pi026), .A2(pi085), .ZN(new_n624_));
  NAND3_X1   g329(.A1(new_n623_), .A2(new_n618_), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1   g330(.A1(new_n610_), .A2(new_n613_), .B(new_n625_), .ZN(po040));
  NOR2_X1    g331(.A1(new_n589_), .A2(new_n592_), .ZN(new_n627_));
  AOI21_X1   g332(.A1(new_n592_), .A2(pi085), .B(pi110), .ZN(new_n628_));
  NOR2_X1    g333(.A1(new_n597_), .A2(new_n592_), .ZN(new_n629_));
  NOR3_X1    g334(.A1(new_n629_), .A2(pi096), .A3(new_n590_), .ZN(new_n630_));
  AOI21_X1   g335(.A1(new_n630_), .A2(new_n628_), .B(new_n627_), .ZN(new_n631_));
  INV_X1     g336(.I(new_n624_), .ZN(new_n632_));
  NOR2_X1    g337(.A1(new_n599_), .A2(new_n592_), .ZN(new_n633_));
  NOR3_X1    g338(.A1(pi027), .A2(pi053), .A3(pi058), .ZN(new_n634_));
  OR2_X2     g339(.A1(new_n634_), .A2(new_n333_), .Z(new_n635_));
  NAND4_X1   g340(.A1(new_n633_), .A2(new_n635_), .A3(pi026), .A4(new_n632_), .ZN(new_n636_));
  NOR2_X1    g341(.A1(new_n636_), .A2(new_n631_), .ZN(po041));
  NAND2_X1   g342(.A1(new_n628_), .A2(pi027), .ZN(new_n638_));
  INV_X1     g343(.I(pi095), .ZN(new_n639_));
  NOR2_X1    g344(.A1(new_n639_), .A2(pi096), .ZN(new_n640_));
  NAND3_X1   g345(.A1(new_n627_), .A2(new_n640_), .A3(new_n616_), .ZN(new_n641_));
  NOR2_X1    g346(.A1(new_n366_), .A2(pi026), .ZN(new_n642_));
  NAND2_X1   g347(.A1(new_n614_), .A2(new_n589_), .ZN(new_n643_));
  NOR2_X1    g348(.A1(pi053), .A2(pi058), .ZN(new_n644_));
  NAND4_X1   g349(.A1(new_n633_), .A2(new_n642_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  AOI22_X1   g350(.A1(new_n645_), .A2(new_n590_), .B1(new_n638_), .B2(new_n641_), .ZN(po042));
  INV_X1     g351(.I(pi039), .ZN(new_n647_));
  INV_X1     g352(.I(pi052), .ZN(new_n648_));
  NOR2_X1    g353(.A1(pi026), .A2(pi051), .ZN(new_n649_));
  AOI21_X1   g354(.A1(new_n649_), .A2(new_n648_), .B(new_n647_), .ZN(new_n650_));
  NOR2_X1    g355(.A1(new_n650_), .A2(new_n614_), .ZN(new_n651_));
  NOR3_X1    g356(.A1(pi026), .A2(pi100), .A3(pi110), .ZN(new_n652_));
  AOI22_X1   g357(.A1(new_n629_), .A2(new_n652_), .B1(new_n640_), .B2(new_n598_), .ZN(new_n653_));
  OR3_X2     g358(.A1(new_n653_), .A2(new_n651_), .A3(new_n616_), .Z(new_n654_));
  OAI21_X1   g359(.A1(new_n653_), .A2(new_n616_), .B(new_n651_), .ZN(new_n655_));
  AOI21_X1   g360(.A1(new_n654_), .A2(new_n655_), .B(new_n589_), .ZN(new_n656_));
  AOI21_X1   g361(.A1(new_n603_), .A2(new_n650_), .B(new_n598_), .ZN(new_n657_));
  AOI21_X1   g362(.A1(new_n657_), .A2(pi027), .B(pi026), .ZN(new_n658_));
  NOR2_X1    g363(.A1(new_n658_), .A2(new_n592_), .ZN(new_n659_));
  OAI21_X1   g364(.A1(new_n656_), .A2(pi028), .B(new_n659_), .ZN(new_n660_));
  NOR3_X1    g365(.A1(new_n448_), .A2(pi027), .A3(pi116), .ZN(new_n661_));
  NAND4_X1   g366(.A1(new_n661_), .A2(pi026), .A3(pi053), .A4(pi085), .ZN(new_n662_));
  INV_X1     g367(.I(new_n661_), .ZN(new_n663_));
  NAND4_X1   g368(.A1(new_n620_), .A2(pi026), .A3(pi085), .A4(new_n333_), .ZN(new_n664_));
  OAI21_X1   g369(.A1(new_n664_), .A2(new_n663_), .B(new_n619_), .ZN(new_n665_));
  NOR2_X1    g370(.A1(pi026), .A2(pi027), .ZN(new_n666_));
  NAND4_X1   g371(.A1(new_n666_), .A2(pi028), .A3(pi085), .A4(pi116), .ZN(new_n667_));
  NAND4_X1   g372(.A1(new_n666_), .A2(new_n448_), .A3(new_n592_), .A4(pi085), .ZN(new_n668_));
  AOI21_X1   g373(.A1(new_n667_), .A2(new_n668_), .B(new_n590_), .ZN(new_n669_));
  NAND2_X1   g374(.A1(new_n665_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1   g375(.A1(new_n660_), .A2(new_n662_), .B(new_n670_), .ZN(po043));
  NAND4_X1   g376(.A1(new_n644_), .A2(pi026), .A3(pi027), .A4(pi085), .ZN(new_n672_));
  OR3_X2     g377(.A1(new_n672_), .A2(new_n449_), .A3(pi116), .Z(new_n673_));
  NOR2_X1    g378(.A1(pi029), .A2(pi116), .ZN(new_n674_));
  AOI21_X1   g379(.A1(new_n601_), .A2(pi116), .B(new_n674_), .ZN(new_n675_));
  NAND4_X1   g380(.A1(pi029), .A2(pi096), .A3(pi097), .A4(pi110), .ZN(new_n676_));
  NAND3_X1   g381(.A1(pi029), .A2(pi097), .A3(pi110), .ZN(new_n677_));
  NAND3_X1   g382(.A1(new_n677_), .A2(new_n591_), .A3(pi097), .ZN(new_n678_));
  AOI21_X1   g383(.A1(new_n678_), .A2(new_n676_), .B(new_n593_), .ZN(new_n679_));
  AOI21_X1   g384(.A1(new_n602_), .A2(pi029), .B(new_n619_), .ZN(new_n680_));
  INV_X1     g385(.I(new_n680_), .ZN(new_n681_));
  INV_X1     g386(.I(pi053), .ZN(new_n682_));
  NOR2_X1    g387(.A1(new_n682_), .A2(new_n619_), .ZN(new_n683_));
  OAI21_X1   g388(.A1(new_n679_), .A2(new_n681_), .B(new_n683_), .ZN(new_n684_));
  NAND2_X1   g389(.A1(new_n678_), .A2(new_n676_), .ZN(new_n685_));
  NAND2_X1   g390(.A1(new_n685_), .A2(pi110), .ZN(new_n686_));
  INV_X1     g391(.I(new_n683_), .ZN(new_n687_));
  NAND3_X1   g392(.A1(new_n686_), .A2(new_n680_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1   g393(.A1(new_n688_), .A2(new_n684_), .B(new_n675_), .ZN(new_n689_));
  INV_X1     g394(.I(new_n644_), .ZN(new_n690_));
  NOR3_X1    g395(.A1(new_n690_), .A2(new_n449_), .A3(new_n616_), .ZN(new_n691_));
  NAND4_X1   g396(.A1(new_n627_), .A2(pi026), .A3(pi029), .A4(new_n634_), .ZN(new_n692_));
  NOR2_X1    g397(.A1(new_n619_), .A2(new_n592_), .ZN(new_n693_));
  NAND3_X1   g398(.A1(new_n693_), .A2(pi029), .A3(pi053), .ZN(new_n694_));
  AOI21_X1   g399(.A1(new_n692_), .A2(new_n589_), .B(new_n694_), .ZN(new_n695_));
  OAI21_X1   g400(.A1(new_n689_), .A2(new_n691_), .B(new_n695_), .ZN(new_n696_));
  AOI21_X1   g401(.A1(new_n696_), .A2(new_n673_), .B(new_n366_), .ZN(po044));
  INV_X1     g402(.I(pi088), .ZN(new_n698_));
  INV_X1     g403(.I(pi109), .ZN(new_n699_));
  NOR2_X1    g404(.A1(new_n699_), .A2(pi060), .ZN(new_n700_));
  OAI21_X1   g405(.A1(pi030), .A2(pi109), .B(pi106), .ZN(new_n701_));
  NOR2_X1    g406(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1   g407(.A1(pi106), .A2(pi129), .ZN(new_n703_));
  XOR2_X1    g408(.A1(new_n702_), .A2(new_n703_), .Z(new_n704_));
  NOR2_X1    g409(.A1(new_n704_), .A2(new_n698_), .ZN(po045));
  INV_X1     g410(.I(pi089), .ZN(new_n706_));
  INV_X1     g411(.I(pi030), .ZN(new_n707_));
  OAI21_X1   g412(.A1(pi031), .A2(pi109), .B(pi106), .ZN(new_n708_));
  AOI21_X1   g413(.A1(new_n707_), .A2(pi109), .B(new_n708_), .ZN(new_n709_));
  XOR2_X1    g414(.A1(new_n709_), .A2(new_n703_), .Z(new_n710_));
  NOR2_X1    g415(.A1(new_n710_), .A2(new_n706_), .ZN(po046));
  INV_X1     g416(.I(pi099), .ZN(new_n712_));
  NOR2_X1    g417(.A1(new_n699_), .A2(pi031), .ZN(new_n713_));
  OAI21_X1   g418(.A1(pi032), .A2(pi109), .B(pi106), .ZN(new_n714_));
  NOR2_X1    g419(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XOR2_X1    g420(.A1(new_n715_), .A2(new_n703_), .Z(new_n716_));
  NOR2_X1    g421(.A1(new_n716_), .A2(new_n712_), .ZN(po047));
  INV_X1     g422(.I(pi090), .ZN(new_n718_));
  INV_X1     g423(.I(pi032), .ZN(new_n719_));
  OAI21_X1   g424(.A1(pi033), .A2(pi109), .B(pi106), .ZN(new_n720_));
  AOI21_X1   g425(.A1(new_n719_), .A2(pi109), .B(new_n720_), .ZN(new_n721_));
  XOR2_X1    g426(.A1(new_n721_), .A2(new_n703_), .Z(new_n722_));
  NOR2_X1    g427(.A1(new_n722_), .A2(new_n718_), .ZN(po048));
  INV_X1     g428(.I(pi091), .ZN(new_n724_));
  INV_X1     g429(.I(pi033), .ZN(new_n725_));
  OAI21_X1   g430(.A1(pi034), .A2(pi109), .B(pi106), .ZN(new_n726_));
  AOI21_X1   g431(.A1(new_n725_), .A2(pi109), .B(new_n726_), .ZN(new_n727_));
  XOR2_X1    g432(.A1(new_n727_), .A2(new_n703_), .Z(new_n728_));
  NOR2_X1    g433(.A1(new_n728_), .A2(new_n724_), .ZN(po049));
  INV_X1     g434(.I(pi092), .ZN(new_n730_));
  INV_X1     g435(.I(pi034), .ZN(new_n731_));
  OAI21_X1   g436(.A1(pi035), .A2(pi109), .B(pi106), .ZN(new_n732_));
  AOI21_X1   g437(.A1(new_n731_), .A2(pi109), .B(new_n732_), .ZN(new_n733_));
  XOR2_X1    g438(.A1(new_n733_), .A2(new_n703_), .Z(new_n734_));
  NOR2_X1    g439(.A1(new_n734_), .A2(new_n730_), .ZN(po050));
  INV_X1     g440(.I(pi098), .ZN(new_n736_));
  INV_X1     g441(.I(pi035), .ZN(new_n737_));
  OAI21_X1   g442(.A1(pi036), .A2(pi109), .B(pi106), .ZN(new_n738_));
  AOI21_X1   g443(.A1(new_n737_), .A2(pi109), .B(new_n738_), .ZN(new_n739_));
  XOR2_X1    g444(.A1(new_n739_), .A2(new_n703_), .Z(new_n740_));
  NOR2_X1    g445(.A1(new_n740_), .A2(new_n736_), .ZN(po051));
  INV_X1     g446(.I(pi093), .ZN(new_n742_));
  INV_X1     g447(.I(pi036), .ZN(new_n743_));
  OAI21_X1   g448(.A1(pi037), .A2(pi109), .B(pi106), .ZN(new_n744_));
  AOI21_X1   g449(.A1(new_n743_), .A2(pi109), .B(new_n744_), .ZN(new_n745_));
  XOR2_X1    g450(.A1(new_n745_), .A2(new_n703_), .Z(new_n746_));
  NOR2_X1    g451(.A1(new_n746_), .A2(new_n742_), .ZN(po052));
  INV_X1     g452(.I(new_n390_), .ZN(new_n748_));
  NAND2_X1   g453(.A1(new_n748_), .A2(new_n517_), .ZN(new_n749_));
  NAND2_X1   g454(.A1(new_n749_), .A2(new_n395_), .ZN(new_n750_));
  INV_X1     g455(.I(pi038), .ZN(new_n751_));
  NAND2_X1   g456(.A1(new_n413_), .A2(new_n401_), .ZN(new_n752_));
  NOR2_X1    g457(.A1(new_n752_), .A2(new_n751_), .ZN(new_n753_));
  AOI21_X1   g458(.A1(new_n753_), .A2(new_n750_), .B(pi082), .ZN(new_n754_));
  INV_X1     g459(.I(pi074), .ZN(new_n755_));
  NAND2_X1   g460(.A1(new_n393_), .A2(new_n755_), .ZN(new_n756_));
  NOR2_X1    g461(.A1(new_n409_), .A2(new_n540_), .ZN(new_n757_));
  NAND4_X1   g462(.A1(pi002), .A2(pi024), .A3(pi045), .A4(pi048), .ZN(new_n758_));
  NOR2_X1    g463(.A1(new_n570_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1     g464(.I(new_n408_), .ZN(new_n760_));
  NAND3_X1   g465(.A1(new_n515_), .A2(pi038), .A3(pi050), .ZN(new_n761_));
  NOR2_X1    g466(.A1(new_n398_), .A2(pi044), .ZN(new_n762_));
  INV_X1     g467(.I(new_n762_), .ZN(new_n763_));
  NOR3_X1    g468(.A1(new_n761_), .A2(new_n760_), .A3(new_n763_), .ZN(new_n764_));
  NAND4_X1   g469(.A1(new_n764_), .A2(new_n756_), .A3(new_n757_), .A4(new_n759_), .ZN(new_n765_));
  NOR2_X1    g470(.A1(new_n754_), .A2(new_n765_), .ZN(po053));
  INV_X1     g471(.I(pi051), .ZN(new_n767_));
  NOR4_X1    g472(.A1(new_n647_), .A2(new_n767_), .A3(new_n648_), .A4(new_n699_), .ZN(po054));
  NOR2_X1    g473(.A1(new_n752_), .A2(new_n518_), .ZN(new_n770_));
  AOI21_X1   g474(.A1(pi082), .A2(new_n394_), .B(new_n770_), .ZN(new_n771_));
  NOR2_X1    g475(.A1(new_n771_), .A2(new_n405_), .ZN(new_n772_));
  INV_X1     g476(.I(new_n543_), .ZN(new_n773_));
  OAI21_X1   g477(.A1(pi073), .A2(new_n394_), .B(new_n541_), .ZN(new_n774_));
  NOR4_X1    g478(.A1(new_n774_), .A2(new_n398_), .A3(new_n773_), .A4(new_n550_), .ZN(new_n775_));
  NOR2_X1    g479(.A1(pi082), .A2(pi129), .ZN(new_n776_));
  NAND2_X1   g480(.A1(new_n550_), .A2(new_n776_), .ZN(new_n777_));
  AOI22_X1   g481(.A1(new_n775_), .A2(new_n759_), .B1(pi040), .B2(new_n777_), .ZN(new_n778_));
  NOR2_X1    g482(.A1(new_n549_), .A2(new_n398_), .ZN(new_n779_));
  NOR4_X1    g483(.A1(new_n772_), .A2(new_n778_), .A3(new_n547_), .A4(new_n779_), .ZN(po055));
  NOR4_X1    g484(.A1(new_n770_), .A2(new_n398_), .A3(new_n394_), .A4(new_n579_), .ZN(new_n781_));
  NOR2_X1    g485(.A1(new_n781_), .A2(pi041), .ZN(new_n782_));
  INV_X1     g486(.I(pi046), .ZN(new_n783_));
  NAND3_X1   g487(.A1(pi047), .A2(pi050), .A3(pi082), .ZN(new_n784_));
  INV_X1     g488(.I(new_n389_), .ZN(new_n785_));
  OAI21_X1   g489(.A1(pi076), .A2(new_n394_), .B(new_n785_), .ZN(new_n786_));
  NOR4_X1    g490(.A1(new_n786_), .A2(new_n388_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n787_));
  AOI21_X1   g491(.A1(new_n787_), .A2(new_n759_), .B(pi129), .ZN(new_n788_));
  INV_X1     g492(.I(pi050), .ZN(new_n789_));
  NOR4_X1    g493(.A1(new_n751_), .A2(new_n547_), .A3(new_n783_), .A4(new_n789_), .ZN(new_n790_));
  NAND4_X1   g494(.A1(new_n790_), .A2(pi041), .A3(pi082), .A4(new_n549_), .ZN(new_n791_));
  NOR3_X1    g495(.A1(new_n782_), .A2(new_n788_), .A3(new_n791_), .ZN(po056));
  NAND2_X1   g496(.A1(pi044), .A2(pi082), .ZN(new_n793_));
  NOR2_X1    g497(.A1(new_n394_), .A2(pi072), .ZN(new_n794_));
  NOR4_X1    g498(.A1(new_n794_), .A2(new_n540_), .A3(new_n548_), .A4(new_n793_), .ZN(new_n795_));
  NAND2_X1   g499(.A1(new_n762_), .A2(pi042), .ZN(new_n796_));
  AOI22_X1   g500(.A1(new_n795_), .A2(new_n759_), .B1(new_n399_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1   g501(.A1(new_n759_), .A2(new_n580_), .A3(new_n790_), .ZN(new_n798_));
  NAND4_X1   g502(.A1(new_n798_), .A2(pi042), .A3(new_n585_), .A4(new_n793_), .ZN(new_n799_));
  NOR2_X1    g503(.A1(new_n797_), .A2(new_n799_), .ZN(po057));
  NAND3_X1   g504(.A1(new_n762_), .A2(pi043), .A3(new_n408_), .ZN(new_n801_));
  OAI21_X1   g505(.A1(new_n801_), .A2(new_n405_), .B(new_n399_), .ZN(new_n802_));
  NAND2_X1   g506(.A1(new_n391_), .A2(pi082), .ZN(new_n803_));
  NOR3_X1    g507(.A1(new_n414_), .A2(new_n506_), .A3(new_n402_), .ZN(new_n804_));
  NOR3_X1    g508(.A1(new_n804_), .A2(new_n388_), .A3(new_n584_), .ZN(new_n805_));
  NAND3_X1   g509(.A1(new_n805_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n806_));
  NOR2_X1    g510(.A1(new_n394_), .A2(pi077), .ZN(new_n807_));
  OR3_X2     g511(.A1(new_n759_), .A2(pi082), .A3(new_n391_), .Z(new_n808_));
  NAND2_X1   g512(.A1(new_n808_), .A2(pi047), .ZN(new_n809_));
  AOI21_X1   g513(.A1(new_n806_), .A2(new_n807_), .B(new_n809_), .ZN(po058));
  NAND3_X1   g514(.A1(new_n544_), .A2(new_n398_), .A3(new_n540_), .ZN(new_n811_));
  NAND3_X1   g515(.A1(new_n811_), .A2(new_n759_), .A3(new_n394_), .ZN(new_n812_));
  AOI21_X1   g516(.A1(new_n407_), .A2(new_n394_), .B(new_n812_), .ZN(new_n813_));
  AND3_X2    g517(.A1(new_n812_), .A2(new_n407_), .A3(new_n394_), .Z(new_n814_));
  OAI21_X1   g518(.A1(new_n814_), .A2(new_n813_), .B(pi067), .ZN(new_n815_));
  AOI21_X1   g519(.A1(new_n815_), .A2(new_n399_), .B(new_n793_), .ZN(po059));
  NAND2_X1   g520(.A1(new_n395_), .A2(new_n586_), .ZN(new_n817_));
  AOI21_X1   g521(.A1(new_n817_), .A2(new_n385_), .B(pi082), .ZN(new_n818_));
  INV_X1     g522(.I(new_n749_), .ZN(new_n819_));
  NOR2_X1    g523(.A1(new_n409_), .A2(new_n773_), .ZN(new_n820_));
  NOR4_X1    g524(.A1(new_n380_), .A2(new_n384_), .A3(new_n398_), .A4(new_n399_), .ZN(new_n821_));
  NOR2_X1    g525(.A1(new_n763_), .A2(new_n506_), .ZN(new_n822_));
  NAND4_X1   g526(.A1(new_n819_), .A2(new_n820_), .A3(new_n822_), .A4(new_n821_), .ZN(new_n823_));
  INV_X1     g527(.I(pi068), .ZN(new_n824_));
  NAND2_X1   g528(.A1(new_n393_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1    g529(.A1(new_n760_), .A2(pi038), .ZN(new_n826_));
  NAND4_X1   g530(.A1(new_n575_), .A2(new_n826_), .A3(new_n413_), .A4(new_n825_), .ZN(new_n827_));
  NOR4_X1    g531(.A1(new_n823_), .A2(new_n818_), .A3(new_n392_), .A4(new_n827_), .ZN(po060));
  NAND2_X1   g532(.A1(new_n759_), .A2(new_n580_), .ZN(new_n829_));
  NOR2_X1    g533(.A1(new_n389_), .A2(pi050), .ZN(new_n830_));
  INV_X1     g534(.I(new_n830_), .ZN(new_n831_));
  OAI21_X1   g535(.A1(new_n829_), .A2(new_n831_), .B(pi082), .ZN(new_n832_));
  NAND3_X1   g536(.A1(new_n832_), .A2(pi075), .A3(new_n393_), .ZN(new_n833_));
  NAND2_X1   g537(.A1(new_n831_), .A2(new_n776_), .ZN(new_n834_));
  NAND2_X1   g538(.A1(new_n834_), .A2(pi046), .ZN(new_n835_));
  NAND2_X1   g539(.A1(new_n820_), .A2(pi082), .ZN(new_n836_));
  NAND4_X1   g540(.A1(new_n829_), .A2(new_n836_), .A3(pi046), .A4(new_n585_), .ZN(new_n837_));
  AOI21_X1   g541(.A1(new_n833_), .A2(new_n835_), .B(new_n837_), .ZN(po061));
  INV_X1     g542(.I(new_n759_), .ZN(new_n839_));
  INV_X1     g543(.I(new_n392_), .ZN(new_n840_));
  NAND2_X1   g544(.A1(new_n840_), .A2(pi082), .ZN(new_n841_));
  NOR2_X1    g545(.A1(new_n763_), .A2(new_n574_), .ZN(new_n842_));
  NAND4_X1   g546(.A1(new_n842_), .A2(pi047), .A3(new_n408_), .A4(new_n503_), .ZN(new_n843_));
  NAND2_X1   g547(.A1(new_n843_), .A2(new_n399_), .ZN(new_n844_));
  INV_X1     g548(.I(pi047), .ZN(new_n845_));
  NOR2_X1    g549(.A1(new_n584_), .A2(new_n845_), .ZN(new_n846_));
  NAND4_X1   g550(.A1(new_n844_), .A2(new_n839_), .A3(new_n841_), .A4(new_n846_), .ZN(new_n847_));
  NOR2_X1    g551(.A1(new_n394_), .A2(pi064), .ZN(new_n848_));
  OAI21_X1   g552(.A1(new_n839_), .A2(new_n392_), .B(pi082), .ZN(new_n849_));
  AOI21_X1   g553(.A1(new_n847_), .A2(new_n848_), .B(new_n849_), .ZN(po062));
  NOR3_X1    g554(.A1(new_n570_), .A2(pi024), .A3(pi045), .ZN(new_n851_));
  INV_X1     g555(.I(pi062), .ZN(new_n852_));
  NAND2_X1   g556(.A1(new_n393_), .A2(new_n852_), .ZN(new_n853_));
  NOR3_X1    g557(.A1(new_n380_), .A2(new_n845_), .A3(new_n398_), .ZN(new_n854_));
  AND3_X2    g558(.A1(new_n851_), .A2(new_n853_), .A3(new_n854_), .Z(new_n855_));
  NOR3_X1    g559(.A1(new_n388_), .A2(new_n845_), .A3(new_n581_), .ZN(new_n856_));
  NAND4_X1   g560(.A1(new_n826_), .A2(new_n748_), .A3(new_n762_), .A4(new_n856_), .ZN(new_n857_));
  AOI22_X1   g561(.A1(new_n855_), .A2(new_n840_), .B1(new_n399_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1   g562(.A1(new_n820_), .A2(pi082), .A3(new_n541_), .ZN(new_n859_));
  NAND4_X1   g563(.A1(new_n859_), .A2(pi048), .A3(new_n585_), .A4(new_n752_), .ZN(new_n860_));
  NOR2_X1    g564(.A1(new_n858_), .A2(new_n860_), .ZN(po063));
  NOR2_X1    g565(.A1(new_n394_), .A2(pi069), .ZN(new_n862_));
  NAND2_X1   g566(.A1(new_n505_), .A2(pi082), .ZN(new_n863_));
  NOR4_X1    g567(.A1(new_n576_), .A2(new_n831_), .A3(new_n862_), .A4(new_n863_), .ZN(new_n864_));
  NAND2_X1   g568(.A1(new_n393_), .A2(new_n412_), .ZN(new_n865_));
  OAI21_X1   g569(.A1(new_n864_), .A2(new_n865_), .B(new_n515_), .ZN(new_n866_));
  NOR2_X1    g570(.A1(pi024), .A2(pi042), .ZN(new_n867_));
  NAND4_X1   g571(.A1(new_n575_), .A2(new_n384_), .A3(new_n382_), .A4(new_n867_), .ZN(new_n868_));
  AOI21_X1   g572(.A1(new_n543_), .A2(new_n547_), .B(pi049), .ZN(new_n869_));
  AOI21_X1   g573(.A1(new_n868_), .A2(new_n869_), .B(new_n407_), .ZN(new_n870_));
  NOR2_X1    g574(.A1(pi002), .A2(pi015), .ZN(new_n871_));
  NAND4_X1   g575(.A1(new_n871_), .A2(new_n411_), .A3(pi045), .A4(pi048), .ZN(new_n872_));
  OAI22_X1   g576(.A1(new_n872_), .A2(new_n540_), .B1(pi024), .B2(pi049), .ZN(new_n873_));
  OAI21_X1   g577(.A1(new_n870_), .A2(new_n873_), .B(new_n830_), .ZN(new_n874_));
  AOI21_X1   g578(.A1(new_n398_), .A2(new_n866_), .B(new_n874_), .ZN(po064));
  NAND2_X1   g579(.A1(new_n540_), .A2(new_n398_), .ZN(new_n876_));
  OAI21_X1   g580(.A1(new_n759_), .A2(new_n876_), .B(new_n785_), .ZN(new_n877_));
  NAND3_X1   g581(.A1(new_n877_), .A2(pi066), .A3(new_n393_), .ZN(new_n878_));
  NAND2_X1   g582(.A1(new_n789_), .A2(new_n399_), .ZN(new_n879_));
  OAI21_X1   g583(.A1(new_n826_), .A2(new_n879_), .B(new_n762_), .ZN(new_n880_));
  NAND4_X1   g584(.A1(new_n851_), .A2(pi002), .A3(new_n382_), .A4(new_n575_), .ZN(new_n881_));
  NOR4_X1    g585(.A1(new_n785_), .A2(new_n789_), .A3(new_n398_), .A4(new_n394_), .ZN(new_n882_));
  NAND2_X1   g586(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1   g587(.A1(new_n878_), .A2(new_n880_), .B(new_n883_), .ZN(po065));
  INV_X1     g588(.I(pi106), .ZN(new_n885_));
  NAND2_X1   g589(.A1(new_n399_), .A2(pi109), .ZN(new_n886_));
  AOI21_X1   g590(.A1(new_n699_), .A2(pi129), .B(pi051), .ZN(new_n887_));
  AOI21_X1   g591(.A1(new_n887_), .A2(new_n886_), .B(new_n885_), .ZN(po066));
  NAND2_X1   g592(.A1(pi052), .A2(pi106), .ZN(new_n889_));
  XOR2_X1    g593(.A1(new_n889_), .A2(new_n699_), .Z(new_n890_));
  AOI21_X1   g594(.A1(new_n890_), .A2(pi051), .B(pi129), .ZN(po067));
  NOR3_X1    g595(.A1(new_n619_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n892_));
  NAND2_X1   g596(.A1(new_n682_), .A2(new_n601_), .ZN(new_n893_));
  NAND4_X1   g597(.A1(new_n892_), .A2(new_n693_), .A3(new_n893_), .A4(new_n602_), .ZN(new_n894_));
  NOR2_X1    g598(.A1(pi053), .A2(pi116), .ZN(new_n895_));
  NAND3_X1   g599(.A1(new_n642_), .A2(pi058), .A3(new_n621_), .ZN(new_n896_));
  AOI21_X1   g600(.A1(new_n894_), .A2(new_n895_), .B(new_n896_), .ZN(po068));
  AOI21_X1   g601(.A1(new_n804_), .A2(new_n840_), .B(new_n398_), .ZN(new_n898_));
  OAI21_X1   g602(.A1(new_n898_), .A2(new_n394_), .B(new_n399_), .ZN(po069));
  INV_X1     g603(.I(pi114), .ZN(new_n900_));
  NAND2_X1   g604(.A1(new_n424_), .A2(new_n399_), .ZN(po129));
  NOR3_X1    g605(.A1(po129), .A2(new_n900_), .A3(pi122), .ZN(po070));
  NAND2_X1   g606(.A1(new_n597_), .A2(pi037), .ZN(new_n903_));
  NAND2_X1   g607(.A1(new_n597_), .A2(new_n619_), .ZN(new_n904_));
  NAND2_X1   g608(.A1(new_n597_), .A2(pi094), .ZN(new_n905_));
  INV_X1     g609(.I(pi094), .ZN(new_n906_));
  NAND2_X1   g610(.A1(new_n906_), .A2(pi026), .ZN(new_n907_));
  AOI22_X1   g611(.A1(pi116), .A2(new_n904_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n908_));
  NOR3_X1    g612(.A1(new_n592_), .A2(pi037), .A3(pi058), .ZN(new_n909_));
  NOR2_X1    g613(.A1(pi037), .A2(pi058), .ZN(new_n910_));
  NOR4_X1    g614(.A1(new_n910_), .A2(new_n597_), .A3(new_n619_), .A4(new_n592_), .ZN(new_n911_));
  NOR3_X1    g615(.A1(new_n908_), .A2(new_n911_), .A3(new_n909_), .ZN(new_n912_));
  NAND2_X1   g616(.A1(new_n682_), .A2(pi085), .ZN(new_n913_));
  OAI21_X1   g617(.A1(new_n912_), .A2(new_n913_), .B(new_n903_), .ZN(new_n914_));
  OAI21_X1   g618(.A1(new_n690_), .A2(new_n903_), .B(pi027), .ZN(new_n916_));
  AOI21_X1   g619(.A1(new_n914_), .A2(pi058), .B(new_n916_), .ZN(po071));
  NAND2_X1   g620(.A1(new_n624_), .A2(new_n682_), .ZN(new_n918_));
  INV_X1     g621(.I(new_n918_), .ZN(new_n919_));
  INV_X1     g622(.I(pi057), .ZN(new_n920_));
  AOI21_X1   g623(.A1(pi058), .A2(pi085), .B(pi053), .ZN(new_n921_));
  NOR2_X1    g624(.A1(pi058), .A2(pi085), .ZN(new_n922_));
  NOR4_X1    g625(.A1(new_n921_), .A2(new_n597_), .A3(new_n922_), .A4(new_n920_), .ZN(new_n923_));
  OAI21_X1   g626(.A1(new_n919_), .A2(new_n923_), .B(pi116), .ZN(new_n924_));
  NOR2_X1    g627(.A1(new_n919_), .A2(pi060), .ZN(new_n925_));
  NOR4_X1    g628(.A1(new_n918_), .A2(new_n366_), .A3(new_n920_), .A4(pi058), .ZN(new_n926_));
  OAI21_X1   g629(.A1(new_n926_), .A2(pi027), .B(new_n693_), .ZN(new_n927_));
  AOI21_X1   g630(.A1(new_n924_), .A2(new_n925_), .B(new_n927_), .ZN(po072));
  NOR3_X1    g631(.A1(new_n597_), .A2(new_n619_), .A3(pi116), .ZN(new_n929_));
  NOR2_X1    g632(.A1(new_n597_), .A2(new_n614_), .ZN(new_n930_));
  NAND4_X1   g633(.A1(new_n930_), .A2(new_n619_), .A3(pi116), .A4(new_n598_), .ZN(new_n931_));
  OR2_X2     g634(.A1(new_n931_), .A2(new_n929_), .Z(new_n932_));
  NAND2_X1   g635(.A1(new_n931_), .A2(new_n929_), .ZN(new_n933_));
  NAND3_X1   g636(.A1(new_n333_), .A2(pi053), .A3(pi085), .ZN(new_n934_));
  AOI21_X1   g637(.A1(new_n932_), .A2(new_n933_), .B(new_n934_), .ZN(po073));
  NOR2_X1    g638(.A1(new_n604_), .A2(new_n682_), .ZN(new_n936_));
  NOR2_X1    g639(.A1(new_n687_), .A2(new_n603_), .ZN(new_n937_));
  NOR2_X1    g640(.A1(new_n604_), .A2(new_n683_), .ZN(new_n938_));
  OAI21_X1   g641(.A1(new_n938_), .A2(new_n937_), .B(pi116), .ZN(new_n939_));
  NOR2_X1    g642(.A1(new_n939_), .A2(new_n936_), .ZN(new_n940_));
  INV_X1     g643(.I(new_n936_), .ZN(new_n941_));
  XOR2_X1    g644(.A1(new_n603_), .A2(new_n683_), .Z(new_n942_));
  AOI21_X1   g645(.A1(new_n942_), .A2(pi116), .B(new_n941_), .ZN(new_n943_));
  NOR4_X1    g646(.A1(new_n604_), .A2(new_n589_), .A3(new_n591_), .A4(new_n690_), .ZN(new_n944_));
  OAI22_X1   g647(.A1(new_n943_), .A2(new_n940_), .B1(pi059), .B2(new_n944_), .ZN(new_n945_));
  NAND4_X1   g648(.A1(new_n621_), .A2(pi059), .A3(new_n592_), .A4(new_n644_), .ZN(new_n946_));
  INV_X1     g649(.I(pi059), .ZN(new_n947_));
  NOR4_X1    g650(.A1(new_n672_), .A2(new_n947_), .A3(pi116), .A4(new_n366_), .ZN(new_n948_));
  NOR4_X1    g651(.A1(new_n690_), .A2(new_n947_), .A3(new_n589_), .A4(pi116), .ZN(new_n949_));
  OAI21_X1   g652(.A1(new_n948_), .A2(pi026), .B(new_n949_), .ZN(new_n950_));
  AOI21_X1   g653(.A1(new_n945_), .A2(new_n946_), .B(new_n950_), .ZN(po074));
  NAND3_X1   g654(.A1(new_n424_), .A2(pi117), .A3(pi122), .ZN(new_n952_));
  NAND3_X1   g655(.A1(pi060), .A2(pi117), .A3(pi122), .ZN(new_n953_));
  XOR2_X1    g656(.A1(new_n952_), .A2(new_n953_), .Z(po075));
  INV_X1     g657(.I(pi122), .ZN(new_n955_));
  NOR4_X1    g658(.A1(new_n900_), .A2(new_n955_), .A3(new_n424_), .A4(new_n399_), .ZN(po076));
  NAND3_X1   g659(.A1(pi131), .A2(pi132), .A3(pi133), .ZN(new_n957_));
  INV_X1     g660(.I(new_n957_), .ZN(new_n958_));
  NAND4_X1   g661(.A1(new_n958_), .A2(pi136), .A3(pi137), .A4(pi138), .ZN(new_n959_));
  INV_X1     g662(.I(pi137), .ZN(new_n960_));
  INV_X1     g663(.I(pi138), .ZN(new_n961_));
  NAND2_X1   g664(.A1(new_n958_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1    g665(.A1(new_n962_), .A2(new_n960_), .ZN(new_n963_));
  INV_X1     g666(.I(pi136), .ZN(new_n964_));
  NOR2_X1    g667(.A1(new_n399_), .A2(new_n964_), .ZN(new_n965_));
  NAND3_X1   g668(.A1(new_n963_), .A2(pi140), .A3(new_n965_), .ZN(new_n966_));
  AOI21_X1   g669(.A1(new_n966_), .A2(new_n852_), .B(new_n959_), .ZN(po077));
  INV_X1     g670(.I(pi063), .ZN(new_n968_));
  NAND3_X1   g671(.A1(new_n963_), .A2(pi142), .A3(new_n965_), .ZN(new_n969_));
  AOI21_X1   g672(.A1(new_n969_), .A2(new_n968_), .B(new_n959_), .ZN(po078));
  INV_X1     g673(.I(pi064), .ZN(new_n971_));
  NAND3_X1   g674(.A1(new_n963_), .A2(pi139), .A3(new_n965_), .ZN(new_n972_));
  AOI21_X1   g675(.A1(new_n972_), .A2(new_n971_), .B(new_n959_), .ZN(po079));
  NAND3_X1   g676(.A1(new_n963_), .A2(pi146), .A3(new_n965_), .ZN(new_n974_));
  AOI21_X1   g677(.A1(new_n974_), .A2(new_n404_), .B(new_n959_), .ZN(po080));
  INV_X1     g678(.I(pi066), .ZN(new_n976_));
  NOR3_X1    g679(.A1(new_n962_), .A2(pi136), .A3(pi137), .ZN(new_n977_));
  NAND3_X1   g680(.A1(new_n977_), .A2(pi129), .A3(pi143), .ZN(new_n978_));
  INV_X1     g681(.I(pi143), .ZN(new_n979_));
  NAND3_X1   g682(.A1(new_n977_), .A2(new_n399_), .A3(new_n979_), .ZN(new_n980_));
  AOI21_X1   g683(.A1(new_n978_), .A2(new_n980_), .B(new_n976_), .ZN(po081));
  INV_X1     g684(.I(pi067), .ZN(new_n982_));
  NAND3_X1   g685(.A1(new_n977_), .A2(pi129), .A3(pi139), .ZN(new_n983_));
  INV_X1     g686(.I(pi139), .ZN(new_n984_));
  NAND3_X1   g687(.A1(new_n977_), .A2(new_n399_), .A3(new_n984_), .ZN(new_n985_));
  AOI21_X1   g688(.A1(new_n983_), .A2(new_n985_), .B(new_n982_), .ZN(po082));
  NAND3_X1   g689(.A1(new_n963_), .A2(pi141), .A3(new_n965_), .ZN(new_n987_));
  AOI21_X1   g690(.A1(new_n987_), .A2(new_n824_), .B(new_n959_), .ZN(po083));
  INV_X1     g691(.I(pi069), .ZN(new_n989_));
  NAND3_X1   g692(.A1(new_n963_), .A2(pi143), .A3(new_n965_), .ZN(new_n990_));
  AOI21_X1   g693(.A1(new_n990_), .A2(new_n989_), .B(new_n959_), .ZN(po084));
  NAND3_X1   g694(.A1(new_n963_), .A2(pi144), .A3(new_n965_), .ZN(new_n992_));
  AOI21_X1   g695(.A1(new_n992_), .A2(new_n508_), .B(new_n959_), .ZN(po085));
  INV_X1     g696(.I(pi071), .ZN(new_n994_));
  NAND3_X1   g697(.A1(new_n963_), .A2(pi145), .A3(new_n965_), .ZN(new_n995_));
  AOI21_X1   g698(.A1(new_n995_), .A2(new_n994_), .B(new_n959_), .ZN(po086));
  INV_X1     g699(.I(pi072), .ZN(new_n997_));
  NAND3_X1   g700(.A1(new_n977_), .A2(pi129), .A3(pi140), .ZN(new_n998_));
  INV_X1     g701(.I(pi140), .ZN(new_n999_));
  NAND3_X1   g702(.A1(new_n977_), .A2(new_n399_), .A3(new_n999_), .ZN(new_n1000_));
  AOI21_X1   g703(.A1(new_n998_), .A2(new_n1000_), .B(new_n997_), .ZN(po087));
  INV_X1     g704(.I(pi073), .ZN(new_n1002_));
  NAND3_X1   g705(.A1(new_n977_), .A2(pi129), .A3(pi141), .ZN(new_n1003_));
  INV_X1     g706(.I(pi141), .ZN(new_n1004_));
  NAND3_X1   g707(.A1(new_n977_), .A2(new_n399_), .A3(new_n1004_), .ZN(new_n1005_));
  AOI21_X1   g708(.A1(new_n1003_), .A2(new_n1005_), .B(new_n1002_), .ZN(po088));
  NAND3_X1   g709(.A1(new_n977_), .A2(pi129), .A3(pi142), .ZN(new_n1007_));
  INV_X1     g710(.I(pi142), .ZN(new_n1008_));
  NAND3_X1   g711(.A1(new_n977_), .A2(new_n399_), .A3(new_n1008_), .ZN(new_n1009_));
  AOI21_X1   g712(.A1(new_n1007_), .A2(new_n1009_), .B(new_n755_), .ZN(po089));
  INV_X1     g713(.I(pi075), .ZN(new_n1011_));
  NAND3_X1   g714(.A1(new_n977_), .A2(pi129), .A3(pi144), .ZN(new_n1012_));
  INV_X1     g715(.I(pi144), .ZN(new_n1013_));
  NAND3_X1   g716(.A1(new_n977_), .A2(new_n399_), .A3(new_n1013_), .ZN(new_n1014_));
  AOI21_X1   g717(.A1(new_n1012_), .A2(new_n1014_), .B(new_n1011_), .ZN(po090));
  INV_X1     g718(.I(pi076), .ZN(new_n1016_));
  NAND3_X1   g719(.A1(new_n977_), .A2(pi129), .A3(pi145), .ZN(new_n1017_));
  INV_X1     g720(.I(pi145), .ZN(new_n1018_));
  NAND3_X1   g721(.A1(new_n977_), .A2(new_n399_), .A3(new_n1018_), .ZN(new_n1019_));
  AOI21_X1   g722(.A1(new_n1017_), .A2(new_n1019_), .B(new_n1016_), .ZN(po091));
  INV_X1     g723(.I(pi077), .ZN(new_n1021_));
  NAND3_X1   g724(.A1(new_n977_), .A2(pi129), .A3(pi146), .ZN(new_n1022_));
  INV_X1     g725(.I(pi146), .ZN(new_n1023_));
  NAND3_X1   g726(.A1(new_n977_), .A2(new_n399_), .A3(new_n1023_), .ZN(new_n1024_));
  AOI21_X1   g727(.A1(new_n1022_), .A2(new_n1024_), .B(new_n1021_), .ZN(po092));
  INV_X1     g728(.I(pi078), .ZN(new_n1026_));
  NOR3_X1    g729(.A1(new_n962_), .A2(pi136), .A3(new_n960_), .ZN(new_n1027_));
  NAND3_X1   g730(.A1(new_n1027_), .A2(pi129), .A3(pi142), .ZN(new_n1028_));
  NAND3_X1   g731(.A1(new_n1027_), .A2(new_n399_), .A3(new_n1008_), .ZN(new_n1029_));
  AOI21_X1   g732(.A1(new_n1028_), .A2(new_n1029_), .B(new_n1026_), .ZN(po093));
  INV_X1     g733(.I(pi079), .ZN(new_n1031_));
  NAND3_X1   g734(.A1(new_n1027_), .A2(pi129), .A3(pi143), .ZN(new_n1032_));
  NAND3_X1   g735(.A1(new_n1027_), .A2(new_n399_), .A3(new_n979_), .ZN(new_n1033_));
  AOI21_X1   g736(.A1(new_n1032_), .A2(new_n1033_), .B(new_n1031_), .ZN(po094));
  INV_X1     g737(.I(pi080), .ZN(new_n1035_));
  NAND3_X1   g738(.A1(new_n1027_), .A2(pi129), .A3(pi144), .ZN(new_n1036_));
  NAND3_X1   g739(.A1(new_n1027_), .A2(new_n399_), .A3(new_n1013_), .ZN(new_n1037_));
  AOI21_X1   g740(.A1(new_n1036_), .A2(new_n1037_), .B(new_n1035_), .ZN(po095));
  INV_X1     g741(.I(pi081), .ZN(new_n1039_));
  NAND3_X1   g742(.A1(new_n1027_), .A2(pi129), .A3(pi145), .ZN(new_n1040_));
  NAND3_X1   g743(.A1(new_n1027_), .A2(new_n399_), .A3(new_n1018_), .ZN(new_n1041_));
  AOI21_X1   g744(.A1(new_n1040_), .A2(new_n1041_), .B(new_n1039_), .ZN(po096));
  NAND3_X1   g745(.A1(new_n1027_), .A2(pi129), .A3(pi146), .ZN(new_n1043_));
  NAND3_X1   g746(.A1(new_n1027_), .A2(new_n399_), .A3(new_n1023_), .ZN(new_n1044_));
  AOI21_X1   g747(.A1(new_n1043_), .A2(new_n1044_), .B(new_n398_), .ZN(po097));
  NAND2_X1   g748(.A1(new_n852_), .A2(pi136), .ZN(new_n1046_));
  NAND2_X1   g749(.A1(pi136), .A2(pi138), .ZN(new_n1047_));
  XOR2_X1    g750(.A1(new_n1046_), .A2(new_n1047_), .Z(new_n1048_));
  AOI21_X1   g751(.A1(new_n1048_), .A2(pi089), .B(new_n960_), .ZN(new_n1049_));
  INV_X1     g752(.I(new_n1049_), .ZN(new_n1050_));
  NAND2_X1   g753(.A1(new_n961_), .A2(pi136), .ZN(new_n1051_));
  NAND2_X1   g754(.A1(pi115), .A2(pi138), .ZN(new_n1052_));
  OAI21_X1   g755(.A1(pi087), .A2(pi138), .B(new_n1052_), .ZN(new_n1053_));
  NAND3_X1   g756(.A1(new_n1053_), .A2(pi031), .A3(pi136), .ZN(new_n1054_));
  XOR2_X1    g757(.A1(new_n1054_), .A2(new_n1051_), .Z(new_n1055_));
  NOR2_X1    g758(.A1(new_n961_), .A2(pi072), .ZN(new_n1056_));
  XOR2_X1    g759(.A1(new_n1056_), .A2(new_n1047_), .Z(new_n1057_));
  NAND2_X1   g760(.A1(pi119), .A2(pi137), .ZN(new_n1058_));
  NOR2_X1    g761(.A1(new_n1057_), .A2(new_n1058_), .ZN(new_n1059_));
  NAND3_X1   g762(.A1(new_n1055_), .A2(new_n1050_), .A3(new_n1059_), .ZN(new_n1060_));
  NAND2_X1   g763(.A1(new_n1055_), .A2(new_n1059_), .ZN(new_n1061_));
  NAND2_X1   g764(.A1(new_n1061_), .A2(new_n1049_), .ZN(new_n1062_));
  NAND2_X1   g765(.A1(new_n1062_), .A2(new_n1060_), .ZN(po098));
  INV_X1     g766(.I(pi084), .ZN(new_n1064_));
  NAND3_X1   g767(.A1(new_n1027_), .A2(pi129), .A3(pi141), .ZN(new_n1065_));
  NAND3_X1   g768(.A1(new_n1027_), .A2(new_n399_), .A3(new_n1004_), .ZN(new_n1066_));
  AOI21_X1   g769(.A1(new_n1065_), .A2(new_n1066_), .B(new_n1064_), .ZN(po099));
  NAND2_X1   g770(.A1(new_n602_), .A2(pi097), .ZN(new_n1068_));
  AOI21_X1   g771(.A1(new_n589_), .A2(new_n593_), .B(new_n1068_), .ZN(new_n1069_));
  NAND2_X1   g772(.A1(pi096), .A2(pi116), .ZN(new_n1070_));
  NAND3_X1   g773(.A1(new_n642_), .A2(new_n634_), .A3(new_n1070_), .ZN(new_n1071_));
  AOI21_X1   g774(.A1(pi085), .A2(new_n1069_), .B(new_n1071_), .ZN(po100));
  INV_X1     g775(.I(pi086), .ZN(new_n1073_));
  NAND3_X1   g776(.A1(new_n1027_), .A2(pi129), .A3(pi139), .ZN(new_n1074_));
  NAND3_X1   g777(.A1(new_n1027_), .A2(new_n399_), .A3(new_n984_), .ZN(new_n1075_));
  AOI21_X1   g778(.A1(new_n1074_), .A2(new_n1075_), .B(new_n1073_), .ZN(po101));
  INV_X1     g779(.I(pi087), .ZN(new_n1077_));
  NAND3_X1   g780(.A1(new_n1027_), .A2(pi129), .A3(pi140), .ZN(new_n1078_));
  NAND3_X1   g781(.A1(new_n1027_), .A2(new_n399_), .A3(new_n999_), .ZN(new_n1079_));
  AOI21_X1   g782(.A1(new_n1078_), .A2(new_n1079_), .B(new_n1077_), .ZN(po102));
  NAND2_X1   g783(.A1(pi136), .A2(pi137), .ZN(new_n1081_));
  NOR2_X1    g784(.A1(new_n962_), .A2(new_n1081_), .ZN(new_n1082_));
  NAND3_X1   g785(.A1(new_n1082_), .A2(pi129), .A3(pi139), .ZN(new_n1083_));
  NAND3_X1   g786(.A1(new_n1082_), .A2(new_n399_), .A3(new_n984_), .ZN(new_n1084_));
  AOI21_X1   g787(.A1(new_n1083_), .A2(new_n1084_), .B(new_n698_), .ZN(po103));
  NAND3_X1   g788(.A1(new_n1082_), .A2(pi129), .A3(pi140), .ZN(new_n1086_));
  NAND3_X1   g789(.A1(new_n1082_), .A2(new_n399_), .A3(new_n999_), .ZN(new_n1087_));
  AOI21_X1   g790(.A1(new_n1086_), .A2(new_n1087_), .B(new_n706_), .ZN(po104));
  NAND3_X1   g791(.A1(new_n1082_), .A2(pi129), .A3(pi142), .ZN(new_n1089_));
  NAND3_X1   g792(.A1(new_n1082_), .A2(new_n399_), .A3(new_n1008_), .ZN(new_n1090_));
  AOI21_X1   g793(.A1(new_n1089_), .A2(new_n1090_), .B(new_n718_), .ZN(po105));
  NAND3_X1   g794(.A1(new_n1082_), .A2(pi129), .A3(pi143), .ZN(new_n1092_));
  NAND3_X1   g795(.A1(new_n1082_), .A2(new_n399_), .A3(new_n979_), .ZN(new_n1093_));
  AOI21_X1   g796(.A1(new_n1092_), .A2(new_n1093_), .B(new_n724_), .ZN(po106));
  NAND3_X1   g797(.A1(new_n1082_), .A2(pi129), .A3(pi144), .ZN(new_n1095_));
  NAND3_X1   g798(.A1(new_n1082_), .A2(new_n399_), .A3(new_n1013_), .ZN(new_n1096_));
  AOI21_X1   g799(.A1(new_n1095_), .A2(new_n1096_), .B(new_n730_), .ZN(po107));
  NAND3_X1   g800(.A1(new_n1082_), .A2(pi129), .A3(pi146), .ZN(new_n1098_));
  NAND3_X1   g801(.A1(new_n1082_), .A2(new_n399_), .A3(new_n1023_), .ZN(new_n1099_));
  AOI21_X1   g802(.A1(new_n1098_), .A2(new_n1099_), .B(new_n742_), .ZN(po108));
  NOR3_X1    g803(.A1(new_n398_), .A2(pi136), .A3(pi137), .ZN(new_n1101_));
  NAND3_X1   g804(.A1(new_n958_), .A2(new_n1101_), .A3(pi138), .ZN(new_n1102_));
  INV_X1     g805(.I(new_n1102_), .ZN(new_n1103_));
  NAND3_X1   g806(.A1(new_n1103_), .A2(pi129), .A3(pi142), .ZN(new_n1104_));
  NAND3_X1   g807(.A1(new_n1103_), .A2(new_n399_), .A3(new_n1008_), .ZN(new_n1105_));
  AOI21_X1   g808(.A1(new_n1104_), .A2(new_n1105_), .B(new_n906_), .ZN(po109));
  NOR2_X1    g809(.A1(new_n957_), .A2(pi003), .ZN(new_n1107_));
  NAND2_X1   g810(.A1(new_n1101_), .A2(pi138), .ZN(new_n1108_));
  NOR3_X1    g811(.A1(new_n1108_), .A2(new_n593_), .A3(new_n957_), .ZN(new_n1109_));
  XOR2_X1    g812(.A1(new_n1109_), .A2(new_n1107_), .Z(new_n1110_));
  OAI21_X1   g813(.A1(new_n1102_), .A2(new_n639_), .B(new_n399_), .ZN(new_n1111_));
  AOI21_X1   g814(.A1(new_n1110_), .A2(pi143), .B(new_n1111_), .ZN(po110));
  OAI21_X1   g815(.A1(new_n1102_), .A2(new_n591_), .B(new_n399_), .ZN(new_n1113_));
  AOI21_X1   g816(.A1(new_n1110_), .A2(pi146), .B(new_n1113_), .ZN(po111));
  OAI21_X1   g817(.A1(new_n1102_), .A2(new_n601_), .B(new_n399_), .ZN(new_n1115_));
  AOI21_X1   g818(.A1(new_n1110_), .A2(pi145), .B(new_n1115_), .ZN(po112));
  NAND3_X1   g819(.A1(new_n1082_), .A2(pi129), .A3(pi145), .ZN(new_n1117_));
  NAND3_X1   g820(.A1(new_n1082_), .A2(new_n399_), .A3(new_n1018_), .ZN(new_n1118_));
  AOI21_X1   g821(.A1(new_n1117_), .A2(new_n1118_), .B(new_n736_), .ZN(po113));
  NAND3_X1   g822(.A1(new_n1082_), .A2(pi129), .A3(pi141), .ZN(new_n1120_));
  NAND3_X1   g823(.A1(new_n1082_), .A2(new_n399_), .A3(new_n1004_), .ZN(new_n1121_));
  AOI21_X1   g824(.A1(new_n1120_), .A2(new_n1121_), .B(new_n712_), .ZN(po114));
  OAI21_X1   g825(.A1(new_n1102_), .A2(new_n590_), .B(new_n399_), .ZN(new_n1123_));
  AOI21_X1   g826(.A1(new_n1110_), .A2(pi144), .B(new_n1123_), .ZN(po115));
  NAND2_X1   g827(.A1(new_n1021_), .A2(pi138), .ZN(new_n1125_));
  XOR2_X1    g828(.A1(new_n1125_), .A2(new_n1047_), .Z(new_n1126_));
  AOI21_X1   g829(.A1(new_n1126_), .A2(pi124), .B(new_n960_), .ZN(new_n1127_));
  INV_X1     g830(.I(pi037), .ZN(new_n1128_));
  NOR2_X1    g831(.A1(pi082), .A2(pi138), .ZN(new_n1129_));
  AOI21_X1   g832(.A1(new_n591_), .A2(pi138), .B(new_n1129_), .ZN(new_n1130_));
  NOR4_X1    g833(.A1(new_n1130_), .A2(new_n1128_), .A3(new_n964_), .A4(new_n961_), .ZN(new_n1131_));
  NOR3_X1    g834(.A1(new_n1130_), .A2(new_n1128_), .A3(new_n964_), .ZN(new_n1132_));
  NOR2_X1    g835(.A1(new_n1132_), .A2(new_n1051_), .ZN(new_n1133_));
  NOR2_X1    g836(.A1(new_n1133_), .A2(new_n1131_), .ZN(new_n1134_));
  NOR2_X1    g837(.A1(new_n964_), .A2(pi065), .ZN(new_n1135_));
  XOR2_X1    g838(.A1(new_n1135_), .A2(new_n1047_), .Z(new_n1136_));
  NAND2_X1   g839(.A1(pi093), .A2(pi137), .ZN(new_n1137_));
  OR2_X2     g840(.A1(new_n1136_), .A2(new_n1137_), .Z(new_n1138_));
  OR3_X2     g841(.A1(new_n1138_), .A2(new_n1127_), .A3(new_n1134_), .Z(new_n1139_));
  OAI21_X1   g842(.A1(new_n1138_), .A2(new_n1134_), .B(new_n1127_), .ZN(new_n1140_));
  NAND2_X1   g843(.A1(new_n1139_), .A2(new_n1140_), .ZN(po116));
  NAND2_X1   g844(.A1(new_n731_), .A2(pi137), .ZN(new_n1142_));
  XOR2_X1    g845(.A1(new_n1142_), .A2(new_n1081_), .Z(new_n1143_));
  AOI21_X1   g846(.A1(new_n1143_), .A2(pi079), .B(new_n961_), .ZN(new_n1144_));
  NAND3_X1   g847(.A1(pi091), .A2(pi136), .A3(pi137), .ZN(new_n1145_));
  NAND3_X1   g848(.A1(new_n639_), .A2(new_n964_), .A3(pi137), .ZN(new_n1146_));
  XOR2_X1    g849(.A1(new_n1146_), .A2(new_n1145_), .Z(new_n1147_));
  NAND2_X1   g850(.A1(new_n976_), .A2(pi136), .ZN(new_n1148_));
  XOR2_X1    g851(.A1(new_n1148_), .A2(new_n1081_), .Z(new_n1149_));
  NAND4_X1   g852(.A1(new_n1147_), .A2(pi069), .A3(new_n1149_), .A4(pi138), .ZN(new_n1150_));
  XNOR2_X1   g853(.A1(new_n1150_), .A2(new_n1144_), .ZN(po117));
  NAND2_X1   g854(.A1(new_n725_), .A2(pi137), .ZN(new_n1152_));
  XOR2_X1    g855(.A1(new_n1152_), .A2(new_n1081_), .Z(new_n1153_));
  AOI21_X1   g856(.A1(new_n1153_), .A2(pi078), .B(new_n961_), .ZN(new_n1154_));
  NAND3_X1   g857(.A1(pi090), .A2(pi136), .A3(pi137), .ZN(new_n1155_));
  NAND3_X1   g858(.A1(new_n906_), .A2(new_n964_), .A3(pi137), .ZN(new_n1156_));
  XOR2_X1    g859(.A1(new_n1156_), .A2(new_n1155_), .Z(new_n1157_));
  NAND2_X1   g860(.A1(new_n968_), .A2(pi136), .ZN(new_n1158_));
  XOR2_X1    g861(.A1(new_n1158_), .A2(new_n1081_), .Z(new_n1159_));
  NAND4_X1   g862(.A1(new_n1157_), .A2(pi074), .A3(new_n1159_), .A4(pi138), .ZN(new_n1160_));
  XNOR2_X1   g863(.A1(new_n1160_), .A2(new_n1154_), .ZN(po118));
  NAND2_X1   g864(.A1(new_n824_), .A2(pi136), .ZN(new_n1162_));
  XOR2_X1    g865(.A1(new_n1162_), .A2(new_n1081_), .Z(new_n1163_));
  AOI21_X1   g866(.A1(new_n1163_), .A2(pi073), .B(new_n961_), .ZN(new_n1164_));
  NAND3_X1   g867(.A1(pi099), .A2(pi136), .A3(pi137), .ZN(new_n1165_));
  INV_X1     g868(.I(pi112), .ZN(new_n1166_));
  NAND3_X1   g869(.A1(new_n1166_), .A2(new_n964_), .A3(pi137), .ZN(new_n1167_));
  XOR2_X1    g870(.A1(new_n1167_), .A2(new_n1165_), .Z(new_n1168_));
  NAND2_X1   g871(.A1(new_n719_), .A2(pi137), .ZN(new_n1169_));
  XOR2_X1    g872(.A1(new_n1169_), .A2(new_n1081_), .Z(new_n1170_));
  NAND4_X1   g873(.A1(new_n1168_), .A2(pi084), .A3(new_n1170_), .A4(pi138), .ZN(new_n1171_));
  XNOR2_X1   g874(.A1(new_n1171_), .A2(new_n1164_), .ZN(po119));
  NAND2_X1   g875(.A1(new_n508_), .A2(pi136), .ZN(new_n1173_));
  XOR2_X1    g876(.A1(new_n1173_), .A2(new_n1047_), .Z(new_n1174_));
  AOI21_X1   g877(.A1(new_n1174_), .A2(pi092), .B(new_n960_), .ZN(new_n1175_));
  NOR2_X1    g878(.A1(pi080), .A2(pi138), .ZN(new_n1176_));
  AOI21_X1   g879(.A1(new_n590_), .A2(pi138), .B(new_n1176_), .ZN(new_n1177_));
  NOR4_X1    g880(.A1(new_n1177_), .A2(new_n737_), .A3(new_n964_), .A4(new_n961_), .ZN(new_n1178_));
  NOR3_X1    g881(.A1(new_n1177_), .A2(new_n737_), .A3(new_n964_), .ZN(new_n1179_));
  NOR2_X1    g882(.A1(new_n1179_), .A2(new_n1051_), .ZN(new_n1180_));
  NOR2_X1    g883(.A1(new_n1180_), .A2(new_n1178_), .ZN(new_n1181_));
  NOR2_X1    g884(.A1(new_n961_), .A2(pi075), .ZN(new_n1182_));
  XOR2_X1    g885(.A1(new_n1182_), .A2(new_n1047_), .Z(new_n1183_));
  NAND2_X1   g886(.A1(pi125), .A2(pi137), .ZN(new_n1184_));
  OR2_X2     g887(.A1(new_n1183_), .A2(new_n1184_), .Z(new_n1185_));
  OR3_X2     g888(.A1(new_n1185_), .A2(new_n1175_), .A3(new_n1181_), .Z(new_n1186_));
  OAI21_X1   g889(.A1(new_n1185_), .A2(new_n1181_), .B(new_n1175_), .ZN(new_n1187_));
  NAND2_X1   g890(.A1(new_n1186_), .A2(new_n1187_), .ZN(po120));
  INV_X1     g891(.I(new_n627_), .ZN(new_n1189_));
  NAND3_X1   g892(.A1(new_n1069_), .A2(new_n644_), .A3(new_n930_), .ZN(new_n1190_));
  AOI21_X1   g893(.A1(new_n1190_), .A2(new_n1189_), .B(new_n366_), .ZN(po121));
  NAND2_X1   g894(.A1(new_n994_), .A2(pi136), .ZN(new_n1192_));
  XOR2_X1    g895(.A1(new_n1192_), .A2(new_n1047_), .Z(new_n1193_));
  AOI21_X1   g896(.A1(new_n1193_), .A2(pi098), .B(new_n960_), .ZN(new_n1194_));
  NOR2_X1    g897(.A1(pi081), .A2(pi138), .ZN(new_n1195_));
  AOI21_X1   g898(.A1(new_n601_), .A2(pi138), .B(new_n1195_), .ZN(new_n1196_));
  NOR4_X1    g899(.A1(new_n1196_), .A2(new_n743_), .A3(new_n964_), .A4(new_n961_), .ZN(new_n1197_));
  NOR3_X1    g900(.A1(new_n1196_), .A2(new_n743_), .A3(new_n964_), .ZN(new_n1198_));
  NOR2_X1    g901(.A1(new_n1198_), .A2(new_n1051_), .ZN(new_n1199_));
  NOR2_X1    g902(.A1(new_n1199_), .A2(new_n1197_), .ZN(new_n1200_));
  NOR2_X1    g903(.A1(new_n961_), .A2(pi023), .ZN(new_n1201_));
  XOR2_X1    g904(.A1(new_n1201_), .A2(new_n1047_), .Z(new_n1202_));
  NAND2_X1   g905(.A1(pi076), .A2(pi137), .ZN(new_n1203_));
  OR2_X2     g906(.A1(new_n1202_), .A2(new_n1203_), .Z(new_n1204_));
  OR3_X2     g907(.A1(new_n1204_), .A2(new_n1194_), .A3(new_n1200_), .Z(new_n1205_));
  OAI21_X1   g908(.A1(new_n1204_), .A2(new_n1200_), .B(new_n1194_), .ZN(new_n1206_));
  NAND2_X1   g909(.A1(new_n1205_), .A2(new_n1206_), .ZN(po122));
  NAND2_X1   g910(.A1(new_n971_), .A2(pi136), .ZN(new_n1208_));
  XOR2_X1    g911(.A1(new_n1208_), .A2(new_n1047_), .Z(new_n1209_));
  AOI21_X1   g912(.A1(new_n1209_), .A2(pi088), .B(new_n960_), .ZN(new_n1210_));
  INV_X1     g913(.I(pi111), .ZN(new_n1211_));
  NOR2_X1    g914(.A1(pi086), .A2(pi138), .ZN(new_n1212_));
  AOI21_X1   g915(.A1(new_n1211_), .A2(pi138), .B(new_n1212_), .ZN(new_n1213_));
  NOR4_X1    g916(.A1(new_n1213_), .A2(new_n707_), .A3(new_n964_), .A4(new_n961_), .ZN(new_n1214_));
  NOR3_X1    g917(.A1(new_n1213_), .A2(new_n707_), .A3(new_n964_), .ZN(new_n1215_));
  NOR2_X1    g918(.A1(new_n1215_), .A2(new_n1051_), .ZN(new_n1216_));
  NOR2_X1    g919(.A1(new_n1216_), .A2(new_n1214_), .ZN(new_n1217_));
  NOR2_X1    g920(.A1(new_n961_), .A2(pi067), .ZN(new_n1218_));
  XOR2_X1    g921(.A1(new_n1218_), .A2(new_n1047_), .Z(new_n1219_));
  NAND2_X1   g922(.A1(pi120), .A2(pi137), .ZN(new_n1220_));
  OR2_X2     g923(.A1(new_n1219_), .A2(new_n1220_), .Z(new_n1221_));
  OR3_X2     g924(.A1(new_n1221_), .A2(new_n1210_), .A3(new_n1217_), .Z(new_n1222_));
  OAI21_X1   g925(.A1(new_n1221_), .A2(new_n1217_), .B(new_n1210_), .ZN(new_n1223_));
  NAND2_X1   g926(.A1(new_n1222_), .A2(new_n1223_), .ZN(po123));
  INV_X1     g927(.I(new_n666_), .ZN(new_n1225_));
  NOR2_X1    g928(.A1(new_n366_), .A2(new_n592_), .ZN(new_n1226_));
  NAND2_X1   g929(.A1(new_n1226_), .A2(new_n614_), .ZN(new_n1227_));
  INV_X1     g930(.I(new_n1226_), .ZN(new_n1228_));
  NAND2_X1   g931(.A1(new_n1228_), .A2(pi027), .ZN(new_n1229_));
  AOI22_X1   g932(.A1(new_n1229_), .A2(new_n1227_), .B1(new_n598_), .B2(new_n1225_), .ZN(po124));
  NAND2_X1   g933(.A1(new_n1226_), .A2(new_n619_), .ZN(new_n1231_));
  NAND2_X1   g934(.A1(new_n1228_), .A2(pi058), .ZN(new_n1232_));
  AOI22_X1   g935(.A1(new_n1232_), .A2(new_n1231_), .B1(pi097), .B2(new_n690_), .ZN(po125));
  NOR2_X1    g936(.A1(new_n957_), .A2(pi129), .ZN(new_n1234_));
  NOR4_X1    g937(.A1(new_n398_), .A2(new_n961_), .A3(pi136), .A4(pi137), .ZN(new_n1235_));
  NAND3_X1   g938(.A1(new_n1234_), .A2(new_n1235_), .A3(pi139), .ZN(new_n1236_));
  AOI21_X1   g939(.A1(new_n1236_), .A2(new_n1211_), .B(new_n1108_), .ZN(po126));
  NAND3_X1   g940(.A1(new_n1234_), .A2(new_n1235_), .A3(pi141), .ZN(new_n1238_));
  AOI21_X1   g941(.A1(new_n1238_), .A2(new_n1166_), .B(new_n1108_), .ZN(po127));
  NOR2_X1    g942(.A1(new_n291_), .A2(pi022), .ZN(new_n1240_));
  NAND3_X1   g943(.A1(pi011), .A2(pi054), .A3(pi113), .ZN(new_n1241_));
  OAI21_X1   g944(.A1(new_n1240_), .A2(new_n1241_), .B(new_n333_), .ZN(new_n1242_));
  AOI21_X1   g945(.A1(new_n1240_), .A2(new_n1241_), .B(new_n1242_), .ZN(po128));
  INV_X1     g946(.I(pi115), .ZN(new_n1244_));
  NAND3_X1   g947(.A1(new_n1234_), .A2(new_n1235_), .A3(pi140), .ZN(new_n1245_));
  AOI21_X1   g948(.A1(new_n1245_), .A2(new_n1244_), .B(new_n1108_), .ZN(po130));
  NOR4_X1    g949(.A1(new_n316_), .A2(new_n457_), .A3(new_n432_), .A4(new_n314_), .ZN(new_n1247_));
  NOR3_X1    g950(.A1(new_n1247_), .A2(new_n291_), .A3(new_n366_), .ZN(po131));
  NAND2_X1   g951(.A1(new_n399_), .A2(pi122), .ZN(po132));
  INV_X1     g952(.I(pi118), .ZN(new_n1250_));
  NOR3_X1    g953(.A1(new_n492_), .A2(new_n291_), .A3(new_n1250_), .ZN(new_n1251_));
  NOR3_X1    g954(.A1(new_n1251_), .A2(new_n291_), .A3(pi059), .ZN(new_n1252_));
  NOR4_X1    g955(.A1(new_n492_), .A2(new_n291_), .A3(new_n947_), .A4(new_n1250_), .ZN(new_n1253_));
  NOR3_X1    g956(.A1(new_n1252_), .A2(pi129), .A3(new_n1253_), .ZN(po133));
  NOR2_X1    g957(.A1(new_n602_), .A2(pi129), .ZN(po134));
  NOR3_X1    g958(.A1(pi003), .A2(pi110), .A3(pi120), .ZN(new_n1256_));
  NOR3_X1    g959(.A1(new_n1256_), .A2(pi111), .A3(pi129), .ZN(po135));
  AND3_X2    g960(.A1(new_n399_), .A2(pi081), .A3(pi120), .Z(po136));
  OR2_X2     g961(.A1(pi129), .A2(pi134), .Z(po137));
  OR2_X2     g962(.A1(pi129), .A2(pi135), .Z(po138));
  NOR2_X1    g963(.A1(new_n920_), .A2(pi129), .ZN(po139));
  AOI21_X1   g964(.A1(pi003), .A2(pi129), .B(pi125), .ZN(new_n1262_));
  NOR2_X1    g965(.A1(new_n1262_), .A2(new_n591_), .ZN(po140));
  INV_X1     g966(.I(pi126), .ZN(new_n1264_));
  AND3_X2    g967(.A1(new_n1264_), .A2(pi132), .A3(pi133), .Z(po141));
  assign     po012 = 1'b1;
  BUF_X16    g968(.I(pi108), .Z(po000));
  BUF_X16    g969(.I(pi083), .Z(po001));
  BUF_X16    g970(.I(pi104), .Z(po002));
  BUF_X16    g971(.I(pi103), .Z(po003));
  BUF_X16    g972(.I(pi102), .Z(po004));
  BUF_X16    g973(.I(pi105), .Z(po005));
  BUF_X16    g974(.I(pi107), .Z(po006));
  BUF_X16    g975(.I(pi101), .Z(po007));
  BUF_X16    g976(.I(pi126), .Z(po008));
  BUF_X16    g977(.I(pi121), .Z(po009));
  BUF_X16    g978(.I(pi001), .Z(po010));
  BUF_X16    g979(.I(pi000), .Z(po011));
  BUF_X16    g980(.I(pi130), .Z(po013));
  BUF_X16    g981(.I(pi128), .Z(po014));
endmodule


