// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:30 2022

module misex3  ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n,
    r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n;
  output r2, s2, t2, u2, n2, o2, p2, q2, h2, i2, j2, k2, m2, l2;
  wire new_n29_, new_n30_, new_n31_, new_n32_, new_n33_, new_n34_, new_n35_,
    new_n36_, new_n37_, new_n38_, new_n39_, new_n40_, new_n41_, new_n42_,
    new_n43_, new_n44_, new_n45_, new_n46_, new_n47_, new_n48_, new_n49_,
    new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_;
  assign new_n29_ = ~j & l;
  assign new_n30_ = ~k & ~new_n29_;
  assign new_n31_ = ~c & f;
  assign new_n32_ = ~c & ~new_n31_;
  assign new_n33_ = a & ~new_n32_;
  assign new_n34_ = f & ~new_n33_;
  assign new_n35_ = ~d & ~new_n34_;
  assign new_n36_ = a & ~new_n35_;
  assign new_n37_ = ~n & ~new_n36_;
  assign new_n38_ = m & new_n37_;
  assign new_n39_ = h & new_n38_;
  assign new_n40_ = ~f & ~h;
  assign new_n41_ = c & new_n40_;
  assign new_n42_ = ~m & n;
  assign new_n43_ = i & new_n42_;
  assign new_n44_ = new_n41_ & new_n43_;
  assign new_n45_ = ~new_n39_ & ~new_n44_;
  assign new_n46_ = e & ~new_n45_;
  assign new_n47_ = f & ~h;
  assign new_n48_ = new_n43_ & new_n47_;
  assign new_n49_ = a & ~e;
  assign new_n50_ = m & ~n;
  assign new_n51_ = h & new_n50_;
  assign new_n52_ = new_n49_ & new_n51_;
  assign new_n53_ = ~new_n48_ & ~new_n52_;
  assign new_n54_ = ~c & ~new_n53_;
  assign new_n55_ = ~e & new_n51_;
  assign new_n56_ = a & new_n55_;
  assign new_n57_ = ~new_n54_ & ~new_n56_;
  assign new_n58_ = d & ~new_n57_;
  assign new_n59_ = ~e & new_n47_;
  assign new_n60_ = new_n43_ & new_n59_;
  assign new_n61_ = ~new_n58_ & ~new_n60_;
  assign new_n62_ = ~new_n46_ & new_n61_;
  assign new_n63_ = ~g & ~new_n62_;
  assign new_n64_ = ~c & g;
  assign new_n65_ = e & ~new_n64_;
  assign new_n66_ = d & ~new_n65_;
  assign new_n67_ = e & g;
  assign new_n68_ = ~d & new_n67_;
  assign new_n69_ = ~new_n66_ & ~new_n68_;
  assign new_n70_ = f & ~new_n69_;
  assign new_n71_ = e & ~f;
  assign new_n72_ = ~e & g;
  assign new_n73_ = ~new_n71_ & ~new_n72_;
  assign new_n74_ = ~d & ~new_n73_;
  assign new_n75_ = ~f & g;
  assign new_n76_ = e & new_n75_;
  assign new_n77_ = ~new_n74_ & ~new_n76_;
  assign new_n78_ = c & ~new_n77_;
  assign new_n79_ = ~new_n70_ & ~new_n78_;
  assign new_n80_ = n & ~new_n79_;
  assign new_n81_ = ~m & new_n80_;
  assign new_n82_ = i & new_n81_;
  assign new_n83_ = ~h & new_n82_;
  assign new_n84_ = ~new_n63_ & ~new_n83_;
  assign new_n85_ = b & ~new_n84_;
  assign new_n86_ = d & e;
  assign new_n87_ = f & ~new_n86_;
  assign new_n88_ = d & new_n71_;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = ~n & ~new_n89_;
  assign new_n91_ = ~m & new_n90_;
  assign new_n92_ = i & new_n91_;
  assign new_n93_ = ~h & new_n92_;
  assign new_n94_ = c & new_n93_;
  assign new_n95_ = ~new_n85_ & ~new_n94_;
  assign new_n96_ = ~new_n30_ & ~new_n95_;
  assign new_n97_ = d & ~e;
  assign new_n98_ = e & f;
  assign new_n99_ = ~d & new_n98_;
  assign new_n100_ = ~new_n97_ & ~new_n99_;
  assign new_n101_ = ~c & ~new_n100_;
  assign new_n102_ = ~d & e;
  assign new_n103_ = c & new_n102_;
  assign new_n104_ = ~new_n97_ & ~new_n103_;
  assign new_n105_ = ~new_n101_ & new_n104_;
  assign new_n106_ = a & ~new_n105_;
  assign new_n107_ = ~d & ~f;
  assign new_n108_ = a & ~new_n107_;
  assign new_n109_ = e & ~new_n108_;
  assign new_n110_ = ~new_n106_ & ~new_n109_;
  assign new_n111_ = ~i & l;
  assign new_n112_ = j & ~l;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = h & ~new_n113_;
  assign new_n115_ = k & ~l;
  assign new_n116_ = ~i & ~new_n115_;
  assign new_n117_ = ~k & l;
  assign new_n118_ = ~new_n116_ & ~new_n117_;
  assign new_n119_ = j & ~new_n118_;
  assign new_n120_ = j & l;
  assign new_n121_ = i & ~new_n120_;
  assign new_n122_ = ~j & ~l;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = k & ~new_n123_;
  assign new_n125_ = i & l;
  assign new_n126_ = ~h & new_n125_;
  assign new_n127_ = ~new_n124_ & ~new_n126_;
  assign new_n128_ = ~new_n119_ & new_n127_;
  assign new_n129_ = ~new_n114_ & new_n128_;
  assign new_n130_ = g & ~new_n129_;
  assign new_n131_ = h & new_n115_;
  assign new_n132_ = ~new_n130_ & ~new_n131_;
  assign new_n133_ = ~new_n110_ & ~new_n132_;
  assign new_n134_ = ~n & new_n133_;
  assign new_n135_ = m & new_n134_;
  assign new_n136_ = d & f;
  assign new_n137_ = ~c & new_n136_;
  assign new_n138_ = c & new_n71_;
  assign new_n139_ = ~new_n137_ & ~new_n138_;
  assign new_n140_ = i & new_n120_;
  assign new_n141_ = k & ~new_n140_;
  assign new_n142_ = j & ~k;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = ~new_n139_ & ~new_n143_;
  assign new_n145_ = c & ~new_n73_;
  assign new_n146_ = f & g;
  assign new_n147_ = e & new_n146_;
  assign new_n148_ = ~new_n145_ & ~new_n147_;
  assign new_n149_ = ~d & ~new_n148_;
  assign new_n150_ = ~d & g;
  assign new_n151_ = f & ~new_n150_;
  assign new_n152_ = ~e & new_n151_;
  assign new_n153_ = ~new_n149_ & ~new_n152_;
  assign new_n154_ = ~new_n143_ & ~new_n153_;
  assign new_n155_ = ~new_n144_ & ~new_n154_;
  assign new_n156_ = n & ~new_n155_;
  assign new_n157_ = ~m & new_n156_;
  assign new_n158_ = h & new_n157_;
  assign new_n159_ = ~new_n135_ & ~new_n158_;
  assign new_n160_ = b & ~new_n159_;
  assign new_n161_ = ~new_n89_ & ~new_n143_;
  assign new_n162_ = ~n & new_n161_;
  assign new_n163_ = ~m & new_n162_;
  assign new_n164_ = h & new_n163_;
  assign new_n165_ = c & new_n164_;
  assign new_n166_ = ~new_n160_ & ~new_n165_;
  assign r2 = new_n96_ | ~new_n166_;
  assign new_n168_ = ~e & new_n146_;
  assign new_n169_ = ~new_n71_ & ~new_n168_;
  assign new_n170_ = ~d & ~new_n169_;
  assign new_n171_ = ~e & f;
  assign new_n172_ = d & new_n171_;
  assign new_n173_ = ~new_n71_ & ~new_n172_;
  assign new_n174_ = ~new_n170_ & new_n173_;
  assign new_n175_ = b & ~new_n174_;
  assign new_n176_ = ~e & ~g;
  assign new_n177_ = b & ~new_n176_;
  assign new_n178_ = f & ~new_n177_;
  assign new_n179_ = ~new_n175_ & ~new_n178_;
  assign new_n180_ = n & ~new_n179_;
  assign new_n181_ = ~new_n71_ & ~new_n171_;
  assign new_n182_ = ~n & ~new_n181_;
  assign new_n183_ = d & new_n182_;
  assign new_n184_ = ~new_n180_ & ~new_n183_;
  assign new_n185_ = ~m & ~new_n184_;
  assign new_n186_ = i & new_n185_;
  assign new_n187_ = ~h & new_n186_;
  assign new_n188_ = ~new_n86_ & ~new_n171_;
  assign new_n189_ = ~n & ~new_n188_;
  assign new_n190_ = m & new_n189_;
  assign new_n191_ = h & new_n190_;
  assign new_n192_ = ~g & new_n191_;
  assign new_n193_ = ~b & new_n192_;
  assign new_n194_ = a & new_n193_;
  assign new_n195_ = ~new_n187_ & ~new_n194_;
  assign new_n196_ = c & ~new_n195_;
  assign new_n197_ = ~b & c;
  assign new_n198_ = ~e & ~new_n197_;
  assign new_n199_ = ~new_n31_ & ~new_n198_;
  assign new_n200_ = a & ~new_n199_;
  assign new_n201_ = b & e;
  assign new_n202_ = ~a & new_n201_;
  assign new_n203_ = ~new_n200_ & ~new_n202_;
  assign new_n204_ = m & ~new_n203_;
  assign new_n205_ = h & new_n204_;
  assign new_n206_ = ~g & new_n205_;
  assign new_n207_ = i & ~m;
  assign new_n208_ = ~h & new_n207_;
  assign new_n209_ = new_n31_ & new_n208_;
  assign new_n210_ = ~new_n206_ & ~new_n209_;
  assign new_n211_ = ~n & ~new_n210_;
  assign new_n212_ = d & new_n211_;
  assign new_n213_ = ~new_n196_ & ~new_n212_;
  assign new_n214_ = ~new_n30_ & ~new_n213_;
  assign new_n215_ = g & ~new_n113_;
  assign new_n216_ = ~new_n115_ & ~new_n215_;
  assign new_n217_ = c & e;
  assign new_n218_ = ~b & new_n217_;
  assign new_n219_ = b & ~e;
  assign new_n220_ = ~new_n218_ & ~new_n219_;
  assign new_n221_ = ~c & ~new_n71_;
  assign new_n222_ = new_n220_ & ~new_n221_;
  assign new_n223_ = d & ~new_n222_;
  assign new_n224_ = new_n171_ & new_n197_;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = a & ~new_n225_;
  assign new_n227_ = ~a & b;
  assign new_n228_ = new_n86_ & new_n227_;
  assign new_n229_ = ~new_n226_ & ~new_n228_;
  assign new_n230_ = ~new_n216_ & ~new_n229_;
  assign new_n231_ = m & new_n230_;
  assign new_n232_ = c & ~new_n181_;
  assign new_n233_ = ~new_n31_ & ~new_n232_;
  assign new_n234_ = ~new_n143_ & ~new_n233_;
  assign new_n235_ = ~m & new_n234_;
  assign new_n236_ = d & new_n235_;
  assign new_n237_ = ~new_n231_ & ~new_n236_;
  assign new_n238_ = ~n & ~new_n237_;
  assign new_n239_ = ~new_n143_ & ~new_n179_;
  assign new_n240_ = n & new_n239_;
  assign new_n241_ = ~m & new_n240_;
  assign new_n242_ = c & new_n241_;
  assign new_n243_ = ~new_n238_ & ~new_n242_;
  assign new_n244_ = h & ~new_n243_;
  assign new_n245_ = ~new_n128_ & ~new_n229_;
  assign new_n246_ = ~n & new_n245_;
  assign new_n247_ = m & new_n246_;
  assign new_n248_ = g & new_n247_;
  assign new_n249_ = ~new_n244_ & ~new_n248_;
  assign s2 = new_n214_ | ~new_n249_;
  assign new_n251_ = ~a & ~new_n97_;
  assign new_n252_ = ~c & ~d;
  assign new_n253_ = a & new_n252_;
  assign new_n254_ = ~new_n251_ & ~new_n253_;
  assign new_n255_ = b & ~new_n254_;
  assign new_n256_ = d & ~new_n201_;
  assign new_n257_ = ~new_n103_ & ~new_n256_;
  assign new_n258_ = a & ~new_n257_;
  assign new_n259_ = ~new_n255_ & ~new_n258_;
  assign new_n260_ = m & ~new_n259_;
  assign new_n261_ = h & new_n260_;
  assign new_n262_ = ~g & new_n261_;
  assign new_n263_ = ~c & d;
  assign new_n264_ = c & ~d;
  assign new_n265_ = ~new_n263_ & ~new_n264_;
  assign new_n266_ = ~m & ~new_n265_;
  assign new_n267_ = i & new_n266_;
  assign new_n268_ = ~h & new_n267_;
  assign new_n269_ = e & new_n268_;
  assign new_n270_ = ~new_n262_ & ~new_n269_;
  assign new_n271_ = ~n & ~new_n270_;
  assign new_n272_ = b & new_n263_;
  assign new_n273_ = ~new_n197_ & ~new_n272_;
  assign new_n274_ = n & ~new_n273_;
  assign new_n275_ = ~m & new_n274_;
  assign new_n276_ = i & new_n275_;
  assign new_n277_ = ~h & new_n276_;
  assign new_n278_ = e & new_n277_;
  assign new_n279_ = ~new_n271_ & ~new_n278_;
  assign new_n280_ = f & ~new_n279_;
  assign new_n281_ = ~f & ~new_n263_;
  assign new_n282_ = ~new_n150_ & ~new_n281_;
  assign new_n283_ = e & ~new_n282_;
  assign new_n284_ = new_n75_ & new_n263_;
  assign new_n285_ = ~new_n283_ & ~new_n284_;
  assign new_n286_ = n & ~new_n285_;
  assign new_n287_ = b & new_n286_;
  assign new_n288_ = ~f & ~n;
  assign new_n289_ = new_n217_ & new_n288_;
  assign new_n290_ = ~new_n287_ & ~new_n289_;
  assign new_n291_ = ~m & ~new_n290_;
  assign new_n292_ = i & new_n291_;
  assign new_n293_ = ~h & new_n292_;
  assign new_n294_ = ~new_n280_ & ~new_n293_;
  assign new_n295_ = ~new_n30_ & ~new_n294_;
  assign new_n296_ = ~new_n143_ & ~new_n265_;
  assign new_n297_ = ~m & new_n296_;
  assign new_n298_ = a & new_n264_;
  assign new_n299_ = ~new_n227_ & ~new_n298_;
  assign new_n300_ = ~new_n216_ & ~new_n299_;
  assign new_n301_ = m & new_n300_;
  assign new_n302_ = ~new_n297_ & ~new_n301_;
  assign new_n303_ = e & ~new_n302_;
  assign new_n304_ = a & ~c;
  assign new_n305_ = a & ~new_n304_;
  assign new_n306_ = ~d & ~new_n305_;
  assign new_n307_ = b & new_n306_;
  assign new_n308_ = a & new_n256_;
  assign new_n309_ = ~new_n307_ & ~new_n308_;
  assign new_n310_ = ~new_n216_ & ~new_n309_;
  assign new_n311_ = m & new_n310_;
  assign new_n312_ = ~new_n303_ & ~new_n311_;
  assign new_n313_ = ~n & ~new_n312_;
  assign new_n314_ = ~new_n143_ & ~new_n273_;
  assign new_n315_ = n & new_n314_;
  assign new_n316_ = ~m & new_n315_;
  assign new_n317_ = e & new_n316_;
  assign new_n318_ = ~new_n313_ & ~new_n317_;
  assign new_n319_ = h & ~new_n318_;
  assign new_n320_ = ~new_n128_ & ~new_n259_;
  assign new_n321_ = ~n & new_n320_;
  assign new_n322_ = m & new_n321_;
  assign new_n323_ = g & new_n322_;
  assign new_n324_ = ~new_n319_ & ~new_n323_;
  assign new_n325_ = f & ~new_n324_;
  assign new_n326_ = ~new_n143_ & ~new_n290_;
  assign new_n327_ = ~m & new_n326_;
  assign new_n328_ = h & new_n327_;
  assign new_n329_ = ~new_n325_ & ~new_n328_;
  assign t2 = new_n295_ | ~new_n329_;
  assign new_n331_ = a & ~g;
  assign new_n332_ = h & m;
  assign new_n333_ = new_n331_ & new_n332_;
  assign new_n334_ = ~h & ~m;
  assign new_n335_ = g & new_n334_;
  assign new_n336_ = ~new_n333_ & ~new_n335_;
  assign new_n337_ = ~n & ~new_n336_;
  assign new_n338_ = d & new_n337_;
  assign new_n339_ = ~c & new_n338_;
  assign new_n340_ = c & g;
  assign new_n341_ = ~b & new_n340_;
  assign new_n342_ = ~h & new_n42_;
  assign new_n343_ = new_n341_ & new_n342_;
  assign new_n344_ = ~new_n339_ & ~new_n343_;
  assign new_n345_ = ~new_n30_ & ~new_n344_;
  assign new_n346_ = h & ~l;
  assign new_n347_ = ~new_n117_ & ~new_n346_;
  assign new_n348_ = j & ~new_n347_;
  assign new_n349_ = k & ~new_n120_;
  assign new_n350_ = ~h & l;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign new_n352_ = ~new_n348_ & new_n351_;
  assign new_n353_ = ~n & ~new_n352_;
  assign new_n354_ = m & new_n353_;
  assign new_n355_ = g & new_n354_;
  assign new_n356_ = d & new_n355_;
  assign new_n357_ = ~c & new_n356_;
  assign new_n358_ = a & new_n357_;
  assign new_n359_ = ~new_n345_ & ~new_n358_;
  assign new_n360_ = i & ~new_n359_;
  assign new_n361_ = c & n;
  assign new_n362_ = ~b & new_n361_;
  assign new_n363_ = d & ~n;
  assign new_n364_ = ~c & new_n363_;
  assign new_n365_ = ~new_n362_ & ~new_n364_;
  assign new_n366_ = ~new_n143_ & ~new_n365_;
  assign new_n367_ = ~m & new_n366_;
  assign new_n368_ = h & new_n367_;
  assign new_n369_ = g & new_n368_;
  assign new_n370_ = ~new_n360_ & ~new_n369_;
  assign new_n371_ = ~new_n71_ & ~new_n370_;
  assign new_n372_ = d & ~f;
  assign new_n373_ = ~new_n31_ & ~new_n372_;
  assign new_n374_ = a & ~new_n373_;
  assign new_n375_ = ~d & f;
  assign new_n376_ = ~e & ~new_n375_;
  assign new_n377_ = ~a & ~new_n376_;
  assign new_n378_ = ~new_n71_ & ~new_n377_;
  assign new_n379_ = ~new_n374_ & new_n378_;
  assign new_n380_ = b & ~new_n379_;
  assign new_n381_ = c & ~new_n136_;
  assign new_n382_ = ~new_n107_ & ~new_n381_;
  assign new_n383_ = e & ~new_n382_;
  assign new_n384_ = ~new_n97_ & ~new_n197_;
  assign new_n385_ = f & ~new_n384_;
  assign new_n386_ = ~new_n383_ & ~new_n385_;
  assign new_n387_ = a & ~new_n386_;
  assign new_n388_ = ~new_n380_ & ~new_n387_;
  assign new_n389_ = m & ~new_n388_;
  assign new_n390_ = h & new_n389_;
  assign new_n391_ = ~g & new_n390_;
  assign new_n392_ = f & ~new_n375_;
  assign new_n393_ = e & ~new_n392_;
  assign new_n394_ = ~new_n171_ & ~new_n393_;
  assign new_n395_ = ~m & ~new_n394_;
  assign new_n396_ = ~h & new_n395_;
  assign new_n397_ = g & new_n396_;
  assign new_n398_ = c & new_n397_;
  assign new_n399_ = ~new_n391_ & ~new_n398_;
  assign new_n400_ = ~n & ~new_n399_;
  assign new_n401_ = c & f;
  assign new_n402_ = e & ~new_n401_;
  assign new_n403_ = ~new_n136_ & ~new_n264_;
  assign new_n404_ = ~e & ~new_n403_;
  assign new_n405_ = ~new_n402_ & ~new_n404_;
  assign new_n406_ = n & ~new_n405_;
  assign new_n407_ = ~m & new_n406_;
  assign new_n408_ = ~h & new_n407_;
  assign new_n409_ = g & new_n408_;
  assign new_n410_ = b & new_n409_;
  assign new_n411_ = ~new_n400_ & ~new_n410_;
  assign new_n412_ = ~new_n30_ & ~new_n411_;
  assign new_n413_ = ~new_n352_ & ~new_n388_;
  assign new_n414_ = ~n & new_n413_;
  assign new_n415_ = m & new_n414_;
  assign new_n416_ = g & new_n415_;
  assign new_n417_ = ~new_n412_ & ~new_n416_;
  assign new_n418_ = i & ~new_n417_;
  assign new_n419_ = b & new_n406_;
  assign new_n420_ = ~n & ~new_n394_;
  assign new_n421_ = c & new_n420_;
  assign new_n422_ = ~new_n419_ & ~new_n421_;
  assign new_n423_ = ~new_n143_ & ~new_n422_;
  assign new_n424_ = ~m & new_n423_;
  assign new_n425_ = h & new_n424_;
  assign new_n426_ = g & new_n425_;
  assign new_n427_ = ~new_n418_ & ~new_n426_;
  assign u2 = new_n371_ | ~new_n427_;
  assign new_n429_ = i & j;
  assign new_n430_ = ~m & ~new_n429_;
  assign new_n431_ = h & new_n430_;
  assign new_n432_ = h & j;
  assign new_n433_ = i & ~new_n432_;
  assign new_n434_ = ~i & new_n120_;
  assign new_n435_ = ~new_n122_ & ~new_n434_;
  assign new_n436_ = ~new_n433_ & new_n435_;
  assign new_n437_ = m & ~new_n436_;
  assign new_n438_ = a & new_n437_;
  assign new_n439_ = ~new_n431_ & ~new_n438_;
  assign new_n440_ = ~e & ~new_n439_;
  assign new_n441_ = f & new_n437_;
  assign new_n442_ = a & new_n441_;
  assign new_n443_ = ~new_n440_ & ~new_n442_;
  assign new_n444_ = ~c & ~new_n443_;
  assign new_n445_ = b & ~f;
  assign new_n446_ = ~new_n171_ & ~new_n445_;
  assign new_n447_ = ~new_n436_ & ~new_n446_;
  assign new_n448_ = m & new_n447_;
  assign new_n449_ = a & new_n448_;
  assign new_n450_ = ~new_n444_ & ~new_n449_;
  assign new_n451_ = d & ~new_n450_;
  assign new_n452_ = a & new_n31_;
  assign new_n453_ = ~new_n71_ & ~new_n452_;
  assign new_n454_ = ~new_n377_ & new_n453_;
  assign new_n455_ = b & ~new_n454_;
  assign new_n456_ = ~b & new_n401_;
  assign new_n457_ = ~new_n383_ & ~new_n456_;
  assign new_n458_ = a & ~new_n457_;
  assign new_n459_ = ~new_n455_ & ~new_n458_;
  assign new_n460_ = ~new_n436_ & ~new_n459_;
  assign new_n461_ = m & new_n460_;
  assign new_n462_ = ~new_n451_ & ~new_n461_;
  assign new_n463_ = k & ~new_n462_;
  assign new_n464_ = ~new_n29_ & ~new_n142_;
  assign new_n465_ = ~i & ~new_n464_;
  assign new_n466_ = ~new_n142_ & ~new_n465_;
  assign new_n467_ = ~new_n171_ & ~new_n221_;
  assign new_n468_ = d & ~new_n467_;
  assign new_n469_ = new_n457_ & ~new_n468_;
  assign new_n470_ = a & ~new_n469_;
  assign new_n471_ = ~new_n380_ & ~new_n470_;
  assign new_n472_ = ~new_n466_ & ~new_n471_;
  assign new_n473_ = m & new_n472_;
  assign new_n474_ = ~c & new_n97_;
  assign new_n475_ = ~k & ~m;
  assign new_n476_ = new_n429_ & new_n475_;
  assign new_n477_ = new_n474_ & new_n476_;
  assign new_n478_ = ~new_n473_ & ~new_n477_;
  assign new_n479_ = h & ~new_n478_;
  assign new_n480_ = ~new_n463_ & ~new_n479_;
  assign new_n481_ = ~n & ~new_n480_;
  assign new_n482_ = k & ~new_n429_;
  assign new_n483_ = i & new_n142_;
  assign new_n484_ = ~new_n482_ & ~new_n483_;
  assign new_n485_ = b & ~d;
  assign new_n486_ = ~b & ~e;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = c & ~new_n487_;
  assign new_n489_ = e & ~new_n136_;
  assign new_n490_ = ~new_n263_ & ~new_n489_;
  assign new_n491_ = b & ~new_n490_;
  assign new_n492_ = ~new_n488_ & ~new_n491_;
  assign new_n493_ = ~new_n484_ & ~new_n492_;
  assign new_n494_ = n & new_n493_;
  assign new_n495_ = ~m & new_n494_;
  assign new_n496_ = h & new_n495_;
  assign new_n497_ = ~new_n481_ & ~new_n496_;
  assign new_n498_ = g & ~new_n497_;
  assign new_n499_ = ~f & n;
  assign new_n500_ = new_n201_ & new_n499_;
  assign new_n501_ = f & ~n;
  assign new_n502_ = c & new_n501_;
  assign new_n503_ = ~new_n500_ & ~new_n502_;
  assign new_n504_ = ~d & ~new_n503_;
  assign new_n505_ = ~g & n;
  assign new_n506_ = b & new_n505_;
  assign new_n507_ = ~new_n288_ & ~new_n506_;
  assign new_n508_ = e & ~new_n507_;
  assign new_n509_ = ~b & n;
  assign new_n510_ = ~e & ~n;
  assign new_n511_ = ~new_n509_ & ~new_n510_;
  assign new_n512_ = g & new_n511_;
  assign new_n513_ = f & ~new_n512_;
  assign new_n514_ = ~new_n508_ & ~new_n513_;
  assign new_n515_ = c & ~new_n514_;
  assign new_n516_ = d & ~new_n67_;
  assign new_n517_ = ~new_n176_ & ~new_n516_;
  assign new_n518_ = n & ~new_n517_;
  assign new_n519_ = b & new_n518_;
  assign new_n520_ = ~new_n364_ & ~new_n519_;
  assign new_n521_ = f & ~new_n520_;
  assign new_n522_ = ~new_n515_ & ~new_n521_;
  assign new_n523_ = ~new_n504_ & new_n522_;
  assign new_n524_ = ~new_n484_ & ~new_n523_;
  assign new_n525_ = ~m & new_n524_;
  assign new_n526_ = h & new_n525_;
  assign n2 = new_n498_ | new_n526_;
  assign new_n528_ = m & ~new_n471_;
  assign new_n529_ = ~e & ~m;
  assign new_n530_ = new_n263_ & new_n529_;
  assign new_n531_ = ~new_n528_ & ~new_n530_;
  assign new_n532_ = ~n & ~new_n531_;
  assign new_n533_ = n & ~new_n492_;
  assign new_n534_ = ~m & new_n533_;
  assign new_n535_ = ~new_n532_ & ~new_n534_;
  assign new_n536_ = g & ~new_n535_;
  assign new_n537_ = ~m & ~new_n523_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = k & ~new_n538_;
  assign new_n540_ = ~j & new_n539_;
  assign new_n541_ = ~f & ~new_n72_;
  assign new_n542_ = ~new_n365_ & ~new_n541_;
  assign new_n543_ = d & n;
  assign new_n544_ = b & new_n543_;
  assign new_n545_ = c & ~n;
  assign new_n546_ = ~new_n544_ & ~new_n545_;
  assign new_n547_ = ~new_n67_ & ~new_n546_;
  assign new_n548_ = ~d & ~n;
  assign new_n549_ = ~new_n505_ & ~new_n548_;
  assign new_n550_ = c & ~new_n549_;
  assign new_n551_ = new_n219_ & new_n505_;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~new_n547_ & new_n552_;
  assign new_n554_ = f & ~new_n553_;
  assign new_n555_ = e & ~g;
  assign new_n556_ = ~new_n150_ & ~new_n555_;
  assign new_n557_ = c & ~new_n556_;
  assign new_n558_ = f & ~g;
  assign new_n559_ = ~d & ~new_n558_;
  assign new_n560_ = ~new_n75_ & ~new_n559_;
  assign new_n561_ = e & ~new_n560_;
  assign new_n562_ = d & g;
  assign new_n563_ = ~c & new_n562_;
  assign new_n564_ = ~new_n561_ & ~new_n563_;
  assign new_n565_ = ~new_n557_ & new_n564_;
  assign new_n566_ = n & ~new_n565_;
  assign new_n567_ = b & new_n566_;
  assign new_n568_ = ~new_n289_ & ~new_n567_;
  assign new_n569_ = ~new_n554_ & new_n568_;
  assign new_n570_ = ~new_n542_ & new_n569_;
  assign new_n571_ = ~m & ~new_n570_;
  assign new_n572_ = ~k & new_n571_;
  assign new_n573_ = j & new_n572_;
  assign new_n574_ = ~new_n540_ & ~new_n573_;
  assign new_n575_ = h & ~new_n574_;
  assign new_n576_ = k & new_n571_;
  assign new_n577_ = ~h & new_n576_;
  assign new_n578_ = ~new_n575_ & ~new_n577_;
  assign new_n579_ = i & ~new_n578_;
  assign new_n580_ = k & l;
  assign new_n581_ = ~j & new_n580_;
  assign new_n582_ = ~new_n142_ & ~new_n581_;
  assign new_n583_ = ~i & ~new_n582_;
  assign new_n584_ = ~new_n142_ & ~new_n583_;
  assign new_n585_ = g & ~new_n584_;
  assign new_n586_ = g & ~new_n122_;
  assign new_n587_ = k & ~new_n586_;
  assign new_n588_ = ~new_n585_ & ~new_n587_;
  assign new_n589_ = ~new_n471_ & ~new_n588_;
  assign new_n590_ = ~n & new_n589_;
  assign new_n591_ = m & new_n590_;
  assign new_n592_ = h & new_n591_;
  assign o2 = new_n579_ | new_n592_;
  assign new_n594_ = i & k;
  assign new_n595_ = ~h & new_n594_;
  assign new_n596_ = h & ~k;
  assign new_n597_ = ~new_n595_ & ~new_n596_;
  assign new_n598_ = ~new_n538_ & ~new_n597_;
  assign new_n599_ = ~new_n115_ & ~new_n471_;
  assign new_n600_ = m & new_n599_;
  assign new_n601_ = k & ~m;
  assign new_n602_ = h & new_n601_;
  assign new_n603_ = new_n474_ & new_n602_;
  assign new_n604_ = ~new_n600_ & ~new_n603_;
  assign new_n605_ = ~n & ~new_n604_;
  assign new_n606_ = k & new_n534_;
  assign new_n607_ = h & new_n606_;
  assign new_n608_ = ~new_n605_ & ~new_n607_;
  assign new_n609_ = g & ~new_n608_;
  assign new_n610_ = k & new_n537_;
  assign new_n611_ = h & new_n610_;
  assign new_n612_ = ~new_n609_ & ~new_n611_;
  assign new_n613_ = ~i & ~new_n612_;
  assign new_n614_ = ~n & ~new_n471_;
  assign new_n615_ = m & new_n614_;
  assign new_n616_ = k & new_n615_;
  assign new_n617_ = h & new_n616_;
  assign new_n618_ = ~g & new_n617_;
  assign new_n619_ = ~new_n613_ & ~new_n618_;
  assign new_n620_ = ~new_n598_ & new_n619_;
  assign new_n621_ = j & ~new_n620_;
  assign new_n622_ = l & new_n615_;
  assign new_n623_ = ~k & new_n622_;
  assign new_n624_ = i & new_n623_;
  assign new_n625_ = ~h & new_n624_;
  assign new_n626_ = g & new_n625_;
  assign p2 = new_n621_ | new_n626_;
  assign new_n628_ = h & new_n528_;
  assign new_n629_ = new_n208_ & new_n401_;
  assign new_n630_ = ~new_n628_ & ~new_n629_;
  assign new_n631_ = ~g & ~new_n630_;
  assign new_n632_ = d & ~new_n541_;
  assign new_n633_ = ~c & new_n632_;
  assign new_n634_ = ~new_n71_ & ~new_n87_;
  assign new_n635_ = c & ~new_n634_;
  assign new_n636_ = ~new_n633_ & ~new_n635_;
  assign new_n637_ = ~m & ~new_n636_;
  assign new_n638_ = i & new_n637_;
  assign new_n639_ = ~h & new_n638_;
  assign new_n640_ = ~new_n631_ & ~new_n639_;
  assign new_n641_ = ~new_n142_ & ~new_n640_;
  assign new_n642_ = ~j & new_n528_;
  assign new_n643_ = j & new_n601_;
  assign new_n644_ = new_n474_ & new_n643_;
  assign new_n645_ = ~new_n642_ & ~new_n644_;
  assign new_n646_ = g & ~new_n645_;
  assign new_n647_ = d & new_n67_;
  assign new_n648_ = f & ~new_n647_;
  assign new_n649_ = ~new_n71_ & ~new_n648_;
  assign new_n650_ = c & ~new_n649_;
  assign new_n651_ = ~new_n137_ & ~new_n650_;
  assign new_n652_ = ~m & ~new_n651_;
  assign new_n653_ = k & new_n652_;
  assign new_n654_ = j & new_n653_;
  assign new_n655_ = ~new_n646_ & ~new_n654_;
  assign new_n656_ = ~i & ~new_n655_;
  assign new_n657_ = ~j & k;
  assign new_n658_ = ~new_n142_ & ~new_n657_;
  assign new_n659_ = ~new_n633_ & ~new_n650_;
  assign new_n660_ = ~new_n658_ & ~new_n659_;
  assign new_n661_ = ~m & new_n660_;
  assign new_n662_ = ~new_n656_ & ~new_n661_;
  assign new_n663_ = h & ~new_n662_;
  assign new_n664_ = h & k;
  assign new_n665_ = j & ~new_n664_;
  assign new_n666_ = i & new_n657_;
  assign new_n667_ = ~new_n665_ & ~new_n666_;
  assign new_n668_ = ~new_n471_ & ~new_n667_;
  assign new_n669_ = m & new_n668_;
  assign new_n670_ = g & new_n669_;
  assign new_n671_ = ~new_n663_ & ~new_n670_;
  assign new_n672_ = ~new_n641_ & new_n671_;
  assign new_n673_ = ~n & ~new_n672_;
  assign new_n674_ = i & ~new_n142_;
  assign new_n675_ = ~h & new_n674_;
  assign new_n676_ = ~i & k;
  assign new_n677_ = k & ~new_n676_;
  assign new_n678_ = j & ~new_n677_;
  assign new_n679_ = ~new_n657_ & ~new_n678_;
  assign new_n680_ = h & ~new_n679_;
  assign new_n681_ = ~new_n675_ & ~new_n680_;
  assign new_n682_ = b & ~new_n556_;
  assign new_n683_ = ~b & ~new_n541_;
  assign new_n684_ = ~new_n558_ & ~new_n683_;
  assign new_n685_ = ~new_n682_ & new_n684_;
  assign new_n686_ = c & ~new_n685_;
  assign new_n687_ = f & ~new_n517_;
  assign new_n688_ = ~new_n563_ & ~new_n687_;
  assign new_n689_ = ~new_n561_ & new_n688_;
  assign new_n690_ = b & ~new_n689_;
  assign new_n691_ = ~new_n686_ & ~new_n690_;
  assign new_n692_ = ~new_n681_ & ~new_n691_;
  assign new_n693_ = n & new_n692_;
  assign new_n694_ = ~m & new_n693_;
  assign new_n695_ = ~new_n673_ & ~new_n694_;
  assign q2 = l & ~new_n695_;
  assign new_n697_ = ~h & ~i;
  assign new_n698_ = j & k;
  assign new_n699_ = new_n697_ & new_n698_;
  assign new_n700_ = h & i;
  assign new_n701_ = ~j & ~k;
  assign new_n702_ = new_n700_ & new_n701_;
  assign new_n703_ = ~new_n699_ & ~new_n702_;
  assign new_n704_ = ~m & ~new_n703_;
  assign new_n705_ = f & new_n704_;
  assign new_n706_ = ~c & new_n705_;
  assign new_n707_ = ~h & ~j;
  assign new_n708_ = ~i & ~new_n707_;
  assign new_n709_ = ~h & i;
  assign new_n710_ = ~new_n142_ & ~new_n709_;
  assign new_n711_ = ~new_n708_ & new_n710_;
  assign new_n712_ = m & ~new_n711_;
  assign new_n713_ = c & new_n712_;
  assign new_n714_ = a & new_n713_;
  assign new_n715_ = ~new_n706_ & ~new_n714_;
  assign new_n716_ = ~d & ~new_n715_;
  assign new_n717_ = a & ~f;
  assign new_n718_ = ~new_n227_ & ~new_n717_;
  assign new_n719_ = ~new_n711_ & ~new_n718_;
  assign new_n720_ = m & new_n719_;
  assign new_n721_ = c & new_n720_;
  assign new_n722_ = ~new_n716_ & ~new_n721_;
  assign new_n723_ = e & ~new_n722_;
  assign new_n724_ = ~a & new_n375_;
  assign new_n725_ = a & new_n372_;
  assign new_n726_ = ~new_n724_ & ~new_n725_;
  assign new_n727_ = b & ~new_n726_;
  assign new_n728_ = b & ~new_n97_;
  assign new_n729_ = f & ~new_n728_;
  assign new_n730_ = a & new_n729_;
  assign new_n731_ = ~new_n727_ & ~new_n730_;
  assign new_n732_ = ~new_n711_ & ~new_n731_;
  assign new_n733_ = m & new_n732_;
  assign new_n734_ = c & new_n733_;
  assign new_n735_ = ~new_n723_ & ~new_n734_;
  assign new_n736_ = l & ~new_n735_;
  assign new_n737_ = ~i & ~k;
  assign new_n738_ = ~new_n346_ & ~new_n737_;
  assign new_n739_ = j & ~new_n738_;
  assign new_n740_ = ~new_n124_ & ~new_n739_;
  assign new_n741_ = ~new_n377_ & ~new_n725_;
  assign new_n742_ = b & ~new_n741_;
  assign new_n743_ = ~new_n489_ & ~new_n729_;
  assign new_n744_ = a & ~new_n743_;
  assign new_n745_ = ~new_n742_ & ~new_n744_;
  assign new_n746_ = ~new_n740_ & ~new_n745_;
  assign new_n747_ = m & new_n746_;
  assign new_n748_ = c & new_n747_;
  assign new_n749_ = ~new_n736_ & ~new_n748_;
  assign new_n750_ = g & ~new_n749_;
  assign new_n751_ = ~new_n30_ & ~new_n745_;
  assign new_n752_ = m & new_n751_;
  assign new_n753_ = c & new_n752_;
  assign new_n754_ = ~f & i;
  assign new_n755_ = new_n252_ & new_n754_;
  assign new_n756_ = l & ~m;
  assign new_n757_ = new_n698_ & new_n756_;
  assign new_n758_ = new_n755_ & new_n757_;
  assign new_n759_ = ~new_n753_ & ~new_n758_;
  assign new_n760_ = h & ~new_n759_;
  assign new_n761_ = new_n40_ & new_n252_;
  assign new_n762_ = ~l & ~m;
  assign new_n763_ = new_n737_ & new_n762_;
  assign new_n764_ = new_n761_ & new_n763_;
  assign new_n765_ = ~new_n760_ & ~new_n764_;
  assign new_n766_ = ~g & ~new_n765_;
  assign new_n767_ = m & ~new_n745_;
  assign new_n768_ = ~l & new_n767_;
  assign new_n769_ = k & new_n768_;
  assign new_n770_ = h & new_n769_;
  assign new_n771_ = c & new_n770_;
  assign new_n772_ = ~new_n766_ & ~new_n771_;
  assign new_n773_ = ~new_n750_ & new_n772_;
  assign h2 = ~n & ~new_n773_;
  assign new_n775_ = b & n;
  assign new_n776_ = n & ~new_n775_;
  assign new_n777_ = l & ~new_n703_;
  assign new_n778_ = ~f & new_n777_;
  assign new_n779_ = ~e & new_n778_;
  assign new_n780_ = e & new_n47_;
  assign new_n781_ = ~i & j;
  assign new_n782_ = ~k & ~l;
  assign new_n783_ = new_n781_ & new_n782_;
  assign new_n784_ = new_n780_ & new_n783_;
  assign new_n785_ = ~new_n779_ & ~new_n784_;
  assign new_n786_ = ~new_n776_ & ~new_n785_;
  assign new_n787_ = i & ~new_n30_;
  assign new_n788_ = ~h & new_n787_;
  assign new_n789_ = h & ~new_n143_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = ~e & ~new_n790_;
  assign new_n792_ = e & new_n40_;
  assign new_n793_ = new_n580_ & new_n781_;
  assign new_n794_ = new_n792_ & new_n793_;
  assign new_n795_ = ~new_n791_ & ~new_n794_;
  assign new_n796_ = n & ~new_n795_;
  assign new_n797_ = ~b & new_n796_;
  assign new_n798_ = ~new_n786_ & ~new_n797_;
  assign new_n799_ = c & ~new_n798_;
  assign new_n800_ = c & ~new_n71_;
  assign new_n801_ = ~new_n790_ & ~new_n800_;
  assign new_n802_ = n & new_n801_;
  assign new_n803_ = b & new_n802_;
  assign new_n804_ = ~c & e;
  assign new_n805_ = new_n40_ & new_n804_;
  assign new_n806_ = l & ~n;
  assign new_n807_ = k & new_n806_;
  assign new_n808_ = new_n781_ & new_n807_;
  assign new_n809_ = new_n805_ & new_n808_;
  assign new_n810_ = ~new_n803_ & ~new_n809_;
  assign new_n811_ = ~new_n799_ & new_n810_;
  assign new_n812_ = ~m & ~new_n811_;
  assign new_n813_ = ~new_n98_ & ~new_n219_;
  assign new_n814_ = ~c & ~new_n813_;
  assign new_n815_ = ~new_n219_ & ~new_n814_;
  assign new_n816_ = ~new_n129_ & ~new_n815_;
  assign new_n817_ = ~n & new_n816_;
  assign new_n818_ = m & new_n817_;
  assign new_n819_ = a & new_n818_;
  assign new_n820_ = ~new_n812_ & ~new_n819_;
  assign new_n821_ = d & ~new_n820_;
  assign new_n822_ = b & d;
  assign new_n823_ = c & ~new_n822_;
  assign new_n824_ = ~new_n107_ & ~new_n823_;
  assign new_n825_ = e & ~new_n824_;
  assign new_n826_ = b & ~c;
  assign new_n827_ = new_n375_ & new_n826_;
  assign new_n828_ = ~new_n825_ & ~new_n827_;
  assign new_n829_ = ~new_n129_ & ~new_n828_;
  assign new_n830_ = m & new_n829_;
  assign new_n831_ = a & new_n830_;
  assign new_n832_ = f & h;
  assign new_n833_ = e & new_n832_;
  assign new_n834_ = new_n252_ & new_n833_;
  assign new_n835_ = i & ~j;
  assign new_n836_ = ~k & new_n756_;
  assign new_n837_ = new_n835_ & new_n836_;
  assign new_n838_ = new_n834_ & new_n837_;
  assign new_n839_ = ~new_n831_ & ~new_n838_;
  assign new_n840_ = ~n & ~new_n839_;
  assign new_n841_ = ~new_n821_ & ~new_n840_;
  assign new_n842_ = g & ~new_n841_;
  assign new_n843_ = ~b & f;
  assign new_n844_ = b & new_n555_;
  assign new_n845_ = ~new_n843_ & ~new_n844_;
  assign new_n846_ = c & ~new_n845_;
  assign new_n847_ = f & ~new_n67_;
  assign new_n848_ = b & new_n847_;
  assign new_n849_ = ~new_n846_ & ~new_n848_;
  assign new_n850_ = n & ~new_n849_;
  assign new_n851_ = ~m & new_n850_;
  assign new_n852_ = i & new_n851_;
  assign new_n853_ = ~h & new_n852_;
  assign new_n854_ = ~n & ~new_n815_;
  assign new_n855_ = m & new_n854_;
  assign new_n856_ = h & new_n855_;
  assign new_n857_ = ~g & new_n856_;
  assign new_n858_ = a & new_n857_;
  assign new_n859_ = ~new_n853_ & ~new_n858_;
  assign new_n860_ = ~new_n30_ & ~new_n859_;
  assign new_n861_ = a & new_n855_;
  assign new_n862_ = ~new_n851_ & ~new_n861_;
  assign new_n863_ = ~l & ~new_n862_;
  assign new_n864_ = ~new_n429_ & ~new_n849_;
  assign new_n865_ = n & new_n864_;
  assign new_n866_ = ~m & new_n865_;
  assign new_n867_ = ~new_n863_ & ~new_n866_;
  assign new_n868_ = k & ~new_n867_;
  assign new_n869_ = ~k & new_n851_;
  assign new_n870_ = j & new_n869_;
  assign new_n871_ = ~new_n868_ & ~new_n870_;
  assign new_n872_ = h & ~new_n871_;
  assign new_n873_ = ~new_n860_ & ~new_n872_;
  assign new_n874_ = d & ~new_n873_;
  assign new_n875_ = ~new_n30_ & ~new_n828_;
  assign new_n876_ = m & new_n875_;
  assign new_n877_ = a & new_n876_;
  assign new_n878_ = ~e & ~f;
  assign new_n879_ = new_n252_ & new_n878_;
  assign new_n880_ = k & new_n756_;
  assign new_n881_ = new_n429_ & new_n880_;
  assign new_n882_ = new_n879_ & new_n881_;
  assign new_n883_ = ~new_n877_ & ~new_n882_;
  assign new_n884_ = h & ~new_n883_;
  assign new_n885_ = ~k & new_n762_;
  assign new_n886_ = new_n697_ & new_n885_;
  assign new_n887_ = new_n879_ & new_n886_;
  assign new_n888_ = ~new_n884_ & ~new_n887_;
  assign new_n889_ = ~g & ~new_n888_;
  assign new_n890_ = m & ~new_n828_;
  assign new_n891_ = ~l & new_n890_;
  assign new_n892_ = k & new_n891_;
  assign new_n893_ = h & new_n892_;
  assign new_n894_ = a & new_n893_;
  assign new_n895_ = ~new_n889_ & ~new_n894_;
  assign new_n896_ = ~n & ~new_n895_;
  assign new_n897_ = ~new_n874_ & ~new_n896_;
  assign i2 = new_n842_ | ~new_n897_;
  assign new_n899_ = ~g & j;
  assign new_n900_ = g & ~j;
  assign new_n901_ = ~new_n899_ & ~new_n900_;
  assign new_n902_ = ~n & ~new_n901_;
  assign new_n903_ = m & new_n902_;
  assign new_n904_ = f & new_n903_;
  assign new_n905_ = ~a & new_n904_;
  assign new_n906_ = ~j & new_n42_;
  assign new_n907_ = new_n75_ & new_n906_;
  assign new_n908_ = ~new_n905_ & ~new_n907_;
  assign new_n909_ = ~k & ~new_n908_;
  assign new_n910_ = i & new_n909_;
  assign new_n911_ = h & new_n910_;
  assign new_n912_ = new_n75_ & new_n697_;
  assign new_n913_ = new_n42_ & new_n698_;
  assign new_n914_ = new_n912_ & new_n913_;
  assign new_n915_ = ~new_n911_ & ~new_n914_;
  assign new_n916_ = b & ~new_n915_;
  assign new_n917_ = ~n & ~new_n703_;
  assign new_n918_ = ~m & new_n917_;
  assign new_n919_ = g & new_n918_;
  assign new_n920_ = ~f & new_n919_;
  assign new_n921_ = ~new_n916_ & ~new_n920_;
  assign new_n922_ = ~e & ~new_n921_;
  assign new_n923_ = ~h & j;
  assign new_n924_ = h & ~j;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = n & ~new_n925_;
  assign new_n927_ = ~m & new_n926_;
  assign new_n928_ = ~k & new_n927_;
  assign new_n929_ = i & new_n928_;
  assign new_n930_ = g & new_n929_;
  assign new_n931_ = ~f & new_n930_;
  assign new_n932_ = e & new_n931_;
  assign new_n933_ = ~b & new_n932_;
  assign new_n934_ = ~new_n922_ & ~new_n933_;
  assign new_n935_ = c & ~new_n934_;
  assign new_n936_ = ~n & ~new_n925_;
  assign new_n937_ = ~m & new_n936_;
  assign new_n938_ = ~k & new_n937_;
  assign new_n939_ = i & new_n938_;
  assign new_n940_ = g & new_n939_;
  assign new_n941_ = ~f & new_n940_;
  assign new_n942_ = e & new_n941_;
  assign new_n943_ = ~c & new_n942_;
  assign new_n944_ = ~new_n935_ & ~new_n943_;
  assign new_n945_ = d & ~new_n944_;
  assign new_n946_ = ~g & new_n700_;
  assign new_n947_ = new_n878_ & new_n946_;
  assign new_n948_ = g & new_n697_;
  assign new_n949_ = new_n98_ & new_n948_;
  assign new_n950_ = ~new_n947_ & ~new_n949_;
  assign new_n951_ = ~n & ~new_n950_;
  assign new_n952_ = ~m & new_n951_;
  assign new_n953_ = k & new_n952_;
  assign new_n954_ = j & new_n953_;
  assign new_n955_ = ~d & new_n954_;
  assign new_n956_ = ~c & new_n955_;
  assign new_n957_ = ~new_n945_ & ~new_n956_;
  assign new_n958_ = l & ~new_n957_;
  assign new_n959_ = ~g & ~h;
  assign new_n960_ = ~f & new_n959_;
  assign new_n961_ = new_n252_ & new_n960_;
  assign new_n962_ = ~i & new_n701_;
  assign new_n963_ = ~m & ~n;
  assign new_n964_ = ~l & new_n963_;
  assign new_n965_ = new_n962_ & new_n964_;
  assign new_n966_ = new_n961_ & new_n965_;
  assign j2 = new_n958_ | new_n966_;
  assign new_n968_ = new_n98_ & new_n698_;
  assign new_n969_ = new_n701_ & new_n878_;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = ~new_n776_ & ~new_n970_;
  assign new_n972_ = ~b & new_n71_;
  assign new_n973_ = ~k & n;
  assign new_n974_ = ~j & new_n973_;
  assign new_n975_ = new_n972_ & new_n974_;
  assign new_n976_ = ~new_n971_ & ~new_n975_;
  assign new_n977_ = i & ~new_n976_;
  assign new_n978_ = h & new_n977_;
  assign new_n979_ = ~b & e;
  assign new_n980_ = new_n40_ & new_n979_;
  assign new_n981_ = k & n;
  assign new_n982_ = new_n781_ & new_n981_;
  assign new_n983_ = new_n980_ & new_n982_;
  assign new_n984_ = ~new_n978_ & ~new_n983_;
  assign new_n985_ = c & ~new_n984_;
  assign new_n986_ = ~f & new_n917_;
  assign new_n987_ = e & new_n986_;
  assign new_n988_ = ~c & new_n987_;
  assign new_n989_ = ~new_n985_ & ~new_n988_;
  assign new_n990_ = ~m & ~new_n989_;
  assign new_n991_ = a & e;
  assign new_n992_ = new_n698_ & new_n991_;
  assign new_n993_ = ~a & ~e;
  assign new_n994_ = new_n701_ & new_n993_;
  assign new_n995_ = ~new_n992_ & ~new_n994_;
  assign new_n996_ = ~n & ~new_n995_;
  assign new_n997_ = m & new_n996_;
  assign new_n998_ = i & new_n997_;
  assign new_n999_ = h & new_n998_;
  assign new_n1000_ = f & new_n999_;
  assign new_n1001_ = c & new_n1000_;
  assign new_n1002_ = b & new_n1001_;
  assign new_n1003_ = ~new_n990_ & ~new_n1002_;
  assign new_n1004_ = d & ~new_n1003_;
  assign new_n1005_ = new_n252_ & new_n780_;
  assign new_n1006_ = k & new_n963_;
  assign new_n1007_ = new_n781_ & new_n1006_;
  assign new_n1008_ = new_n1005_ & new_n1007_;
  assign new_n1009_ = ~new_n1004_ & ~new_n1008_;
  assign new_n1010_ = g & ~new_n1009_;
  assign new_n1011_ = ~f & ~g;
  assign new_n1012_ = e & new_n1011_;
  assign new_n1013_ = new_n252_ & new_n1012_;
  assign new_n1014_ = h & new_n429_;
  assign new_n1015_ = new_n1006_ & new_n1014_;
  assign new_n1016_ = new_n1013_ & new_n1015_;
  assign new_n1017_ = ~new_n1010_ & ~new_n1016_;
  assign new_n1018_ = l & ~new_n1017_;
  assign new_n1019_ = ~e & new_n1011_;
  assign new_n1020_ = new_n252_ & new_n1019_;
  assign new_n1021_ = ~h & new_n737_;
  assign new_n1022_ = new_n964_ & new_n1021_;
  assign new_n1023_ = new_n1020_ & new_n1022_;
  assign k2 = new_n1018_ | new_n1023_;
  assign new_n1025_ = ~k & ~new_n901_;
  assign new_n1026_ = ~e & new_n1025_;
  assign new_n1027_ = ~a & new_n1026_;
  assign new_n1028_ = g & new_n698_;
  assign new_n1029_ = new_n991_ & new_n1028_;
  assign new_n1030_ = ~new_n1027_ & ~new_n1029_;
  assign new_n1031_ = ~n & ~new_n1030_;
  assign new_n1032_ = m & new_n1031_;
  assign new_n1033_ = g & j;
  assign new_n1034_ = e & new_n1033_;
  assign new_n1035_ = k & new_n42_;
  assign new_n1036_ = new_n1034_ & new_n1035_;
  assign new_n1037_ = ~new_n1032_ & ~new_n1036_;
  assign new_n1038_ = f & ~new_n1037_;
  assign new_n1039_ = ~e & new_n75_;
  assign new_n1040_ = new_n42_ & new_n701_;
  assign new_n1041_ = new_n1039_ & new_n1040_;
  assign new_n1042_ = ~new_n1038_ & ~new_n1041_;
  assign new_n1043_ = b & ~new_n1042_;
  assign new_n1044_ = ~b & ~f;
  assign new_n1045_ = new_n974_ & new_n1044_;
  assign new_n1046_ = f & j;
  assign new_n1047_ = k & ~n;
  assign new_n1048_ = new_n1046_ & new_n1047_;
  assign new_n1049_ = ~new_n1045_ & ~new_n1048_;
  assign new_n1050_ = e & ~new_n1049_;
  assign new_n1051_ = ~k & ~n;
  assign new_n1052_ = ~j & new_n1051_;
  assign new_n1053_ = new_n878_ & new_n1052_;
  assign new_n1054_ = ~new_n1050_ & ~new_n1053_;
  assign new_n1055_ = ~m & ~new_n1054_;
  assign new_n1056_ = g & new_n1055_;
  assign new_n1057_ = ~new_n1043_ & ~new_n1056_;
  assign new_n1058_ = i & ~new_n1057_;
  assign new_n1059_ = n & ~new_n509_;
  assign new_n1060_ = ~m & ~new_n1059_;
  assign new_n1061_ = ~k & new_n1060_;
  assign new_n1062_ = ~j & new_n1061_;
  assign new_n1063_ = ~i & new_n1062_;
  assign new_n1064_ = ~g & new_n1063_;
  assign new_n1065_ = ~f & new_n1064_;
  assign new_n1066_ = ~e & new_n1065_;
  assign new_n1067_ = ~new_n1058_ & ~new_n1066_;
  assign new_n1068_ = h & ~new_n1067_;
  assign new_n1069_ = i & ~k;
  assign new_n1070_ = ~new_n676_ & ~new_n1069_;
  assign new_n1071_ = e & ~new_n1070_;
  assign new_n1072_ = ~b & new_n1071_;
  assign new_n1073_ = new_n219_ & new_n676_;
  assign new_n1074_ = ~new_n1072_ & ~new_n1073_;
  assign new_n1075_ = n & ~new_n1074_;
  assign new_n1076_ = ~e & ~i;
  assign new_n1077_ = new_n1047_ & new_n1076_;
  assign new_n1078_ = ~new_n1075_ & ~new_n1077_;
  assign new_n1079_ = ~m & ~new_n1078_;
  assign new_n1080_ = j & new_n1079_;
  assign new_n1081_ = ~h & new_n1080_;
  assign new_n1082_ = g & new_n1081_;
  assign new_n1083_ = ~f & new_n1082_;
  assign new_n1084_ = ~new_n1068_ & ~new_n1083_;
  assign new_n1085_ = c & ~new_n1084_;
  assign new_n1086_ = j & ~new_n1070_;
  assign new_n1087_ = ~h & new_n1086_;
  assign new_n1088_ = ~new_n702_ & ~new_n1087_;
  assign new_n1089_ = ~n & ~new_n1088_;
  assign new_n1090_ = ~m & new_n1089_;
  assign new_n1091_ = g & new_n1090_;
  assign new_n1092_ = ~f & new_n1091_;
  assign new_n1093_ = e & new_n1092_;
  assign new_n1094_ = ~c & new_n1093_;
  assign new_n1095_ = ~new_n1085_ & ~new_n1094_;
  assign new_n1096_ = d & ~new_n1095_;
  assign new_n1097_ = g & ~new_n703_;
  assign new_n1098_ = f & new_n1097_;
  assign new_n1099_ = e & new_n1098_;
  assign new_n1100_ = ~g & h;
  assign new_n1101_ = ~f & new_n1100_;
  assign new_n1102_ = i & new_n698_;
  assign new_n1103_ = new_n1101_ & new_n1102_;
  assign new_n1104_ = ~new_n1099_ & ~new_n1103_;
  assign new_n1105_ = ~m & ~new_n1104_;
  assign new_n1106_ = ~c & new_n1105_;
  assign new_n1107_ = c & new_n878_;
  assign new_n1108_ = new_n227_ & new_n1107_;
  assign new_n1109_ = k & m;
  assign new_n1110_ = ~j & new_n1109_;
  assign new_n1111_ = new_n948_ & new_n1110_;
  assign new_n1112_ = new_n1108_ & new_n1111_;
  assign new_n1113_ = ~new_n1106_ & ~new_n1112_;
  assign new_n1114_ = ~n & ~new_n1113_;
  assign new_n1115_ = ~d & new_n1114_;
  assign new_n1116_ = ~new_n1096_ & ~new_n1115_;
  assign new_n1117_ = l & ~new_n1116_;
  assign new_n1118_ = j & ~new_n776_;
  assign new_n1119_ = g & new_n1118_;
  assign new_n1120_ = f & new_n1119_;
  assign new_n1121_ = e & new_n1120_;
  assign new_n1122_ = d & new_n1121_;
  assign new_n1123_ = c & new_n1122_;
  assign new_n1124_ = ~g & ~n;
  assign new_n1125_ = ~f & new_n1124_;
  assign new_n1126_ = new_n252_ & new_n1125_;
  assign new_n1127_ = ~new_n1123_ & ~new_n1126_;
  assign new_n1128_ = ~m & ~new_n1127_;
  assign new_n1129_ = ~l & new_n1128_;
  assign new_n1130_ = ~k & new_n1129_;
  assign new_n1131_ = ~i & new_n1130_;
  assign new_n1132_ = ~h & new_n1131_;
  assign m2 = new_n1117_ | new_n1132_;
  assign new_n1134_ = ~new_n88_ & ~new_n375_;
  assign new_n1135_ = ~c & ~new_n1134_;
  assign new_n1136_ = ~e & new_n281_;
  assign new_n1137_ = j & new_n580_;
  assign new_n1138_ = ~new_n701_ & ~new_n1137_;
  assign new_n1139_ = i & ~new_n1138_;
  assign new_n1140_ = h & new_n1139_;
  assign new_n1141_ = g & new_n1140_;
  assign new_n1142_ = h & ~new_n142_;
  assign new_n1143_ = ~g & ~new_n1142_;
  assign new_n1144_ = new_n29_ & new_n697_;
  assign new_n1145_ = a & ~new_n1144_;
  assign new_n1146_ = ~new_n1143_ & new_n1145_;
  assign new_n1147_ = ~new_n1141_ & new_n1146_;
  assign new_n1148_ = ~new_n1136_ & new_n1147_;
  assign new_n1149_ = ~new_n1135_ & new_n1148_;
  assign new_n1150_ = ~b & ~new_n1149_;
  assign new_n1151_ = g & ~k;
  assign new_n1152_ = d & new_n1151_;
  assign new_n1153_ = f & ~new_n1152_;
  assign new_n1154_ = ~a & ~new_n1153_;
  assign new_n1155_ = g & h;
  assign new_n1156_ = f & new_n1155_;
  assign new_n1157_ = i & new_n580_;
  assign new_n1158_ = new_n1156_ & new_n1157_;
  assign new_n1159_ = ~new_n107_ & ~new_n1158_;
  assign new_n1160_ = ~new_n1154_ & new_n1159_;
  assign new_n1161_ = j & ~new_n1160_;
  assign new_n1162_ = a & d;
  assign new_n1163_ = ~g & ~new_n142_;
  assign new_n1164_ = c & ~h;
  assign new_n1165_ = ~i & new_n580_;
  assign new_n1166_ = new_n1164_ & new_n1165_;
  assign new_n1167_ = ~new_n1163_ & new_n1166_;
  assign new_n1168_ = ~new_n1162_ & ~new_n1167_;
  assign new_n1169_ = ~a & d;
  assign new_n1170_ = a & ~d;
  assign new_n1171_ = ~new_n1169_ & ~new_n1170_;
  assign new_n1172_ = ~new_n1168_ & new_n1171_;
  assign new_n1173_ = ~f & ~new_n1172_;
  assign new_n1174_ = ~f & k;
  assign new_n1175_ = d & ~new_n700_;
  assign new_n1176_ = ~a & new_n1175_;
  assign new_n1177_ = a & b;
  assign new_n1178_ = new_n264_ & new_n1177_;
  assign new_n1179_ = ~new_n1176_ & ~new_n1178_;
  assign new_n1180_ = ~new_n1174_ & ~new_n1179_;
  assign new_n1181_ = ~new_n1169_ & ~new_n1178_;
  assign new_n1182_ = l & ~new_n1163_;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1184_ = f & k;
  assign new_n1185_ = c & ~new_n1184_;
  assign new_n1186_ = d & ~new_n1185_;
  assign new_n1187_ = ~a & new_n1186_;
  assign new_n1188_ = ~new_n1183_ & ~new_n1187_;
  assign new_n1189_ = ~new_n1180_ & new_n1188_;
  assign new_n1190_ = ~new_n1173_ & new_n1189_;
  assign new_n1191_ = ~new_n1161_ & new_n1190_;
  assign new_n1192_ = ~e & ~new_n1191_;
  assign new_n1193_ = ~new_n401_ & ~new_n1138_;
  assign new_n1194_ = new_n580_ & new_n1046_;
  assign new_n1195_ = ~new_n701_ & ~new_n1194_;
  assign new_n1196_ = ~d & ~new_n1195_;
  assign new_n1197_ = ~k & ~new_n993_;
  assign new_n1198_ = ~j & new_n1197_;
  assign new_n1199_ = ~a & f;
  assign new_n1200_ = new_n1137_ & new_n1199_;
  assign new_n1201_ = ~new_n1198_ & ~new_n1200_;
  assign new_n1202_ = ~new_n1196_ & new_n1201_;
  assign new_n1203_ = ~new_n1193_ & new_n1202_;
  assign new_n1204_ = h & ~new_n1203_;
  assign new_n1205_ = g & new_n1204_;
  assign new_n1206_ = ~new_n782_ & ~new_n1011_;
  assign new_n1207_ = ~h & ~new_n1206_;
  assign new_n1208_ = ~new_n1205_ & ~new_n1207_;
  assign new_n1209_ = i & ~new_n1208_;
  assign new_n1210_ = b & c;
  assign new_n1211_ = a & new_n1210_;
  assign new_n1212_ = d & new_n98_;
  assign new_n1213_ = new_n1211_ & new_n1212_;
  assign new_n1214_ = h & ~new_n1213_;
  assign new_n1215_ = ~new_n142_ & ~new_n1214_;
  assign new_n1216_ = ~new_n40_ & ~new_n142_;
  assign new_n1217_ = ~new_n993_ & ~new_n1216_;
  assign new_n1218_ = ~c & ~new_n1142_;
  assign new_n1219_ = ~f & j;
  assign new_n1220_ = l & ~new_n1219_;
  assign new_n1221_ = ~new_n664_ & ~new_n1220_;
  assign new_n1222_ = d & i;
  assign new_n1223_ = j & ~new_n1222_;
  assign new_n1224_ = h & ~new_n1223_;
  assign new_n1225_ = ~k & ~new_n1224_;
  assign new_n1226_ = ~f & ~new_n372_;
  assign new_n1227_ = ~h & ~new_n1226_;
  assign new_n1228_ = ~new_n1225_ & ~new_n1227_;
  assign new_n1229_ = ~new_n1221_ & new_n1228_;
  assign new_n1230_ = ~new_n1218_ & new_n1229_;
  assign new_n1231_ = ~new_n1217_ & new_n1230_;
  assign new_n1232_ = ~new_n1215_ & new_n1231_;
  assign new_n1233_ = ~g & ~new_n1232_;
  assign new_n1234_ = f & ~j;
  assign new_n1235_ = new_n86_ & new_n1234_;
  assign new_n1236_ = new_n1211_ & new_n1235_;
  assign new_n1237_ = new_n112_ & new_n697_;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = k & ~new_n1238_;
  assign new_n1240_ = ~new_n701_ & ~new_n1213_;
  assign new_n1241_ = ~l & ~new_n1240_;
  assign new_n1242_ = ~new_n1144_ & ~new_n1213_;
  assign new_n1243_ = ~k & ~new_n1242_;
  assign new_n1244_ = f & ~new_n700_;
  assign new_n1245_ = e & new_n1244_;
  assign new_n1246_ = d & new_n1245_;
  assign new_n1247_ = c & new_n1246_;
  assign new_n1248_ = b & new_n1247_;
  assign new_n1249_ = ~i & new_n29_;
  assign new_n1250_ = new_n40_ & new_n1249_;
  assign new_n1251_ = ~new_n1248_ & ~new_n1250_;
  assign new_n1252_ = a & ~new_n1251_;
  assign new_n1253_ = ~d & ~e;
  assign new_n1254_ = ~f & ~new_n1253_;
  assign new_n1255_ = c & ~f;
  assign new_n1256_ = ~new_n1254_ & new_n1255_;
  assign new_n1257_ = l & ~new_n1256_;
  assign new_n1258_ = ~j & new_n1257_;
  assign new_n1259_ = ~i & new_n1258_;
  assign new_n1260_ = ~h & new_n1259_;
  assign new_n1261_ = ~new_n1252_ & ~new_n1260_;
  assign new_n1262_ = ~new_n1243_ & new_n1261_;
  assign new_n1263_ = ~new_n1241_ & new_n1262_;
  assign new_n1264_ = ~new_n1239_ & new_n1263_;
  assign new_n1265_ = ~new_n1233_ & new_n1264_;
  assign new_n1266_ = ~new_n1209_ & new_n1265_;
  assign new_n1267_ = ~new_n1192_ & new_n1266_;
  assign new_n1268_ = ~new_n1150_ & new_n1267_;
  assign new_n1269_ = m & ~new_n1268_;
  assign new_n1270_ = g & ~i;
  assign new_n1271_ = f & new_n1270_;
  assign new_n1272_ = new_n217_ & new_n1271_;
  assign new_n1273_ = new_n140_ & new_n1100_;
  assign new_n1274_ = ~new_n1272_ & ~new_n1273_;
  assign new_n1275_ = k & ~new_n1274_;
  assign new_n1276_ = new_n217_ & new_n1033_;
  assign new_n1277_ = ~new_n924_ & ~new_n1276_;
  assign new_n1278_ = i & ~new_n1277_;
  assign new_n1279_ = f & new_n1278_;
  assign new_n1280_ = ~h & ~new_n29_;
  assign new_n1281_ = ~new_n924_ & ~new_n1280_;
  assign new_n1282_ = ~g & ~new_n1281_;
  assign new_n1283_ = ~c & new_n1282_;
  assign new_n1284_ = ~new_n1279_ & ~new_n1283_;
  assign new_n1285_ = ~k & ~new_n1284_;
  assign new_n1286_ = f & ~new_n697_;
  assign new_n1287_ = ~g & ~new_n1286_;
  assign new_n1288_ = f & new_n697_;
  assign new_n1289_ = ~new_n1287_ & ~new_n1288_;
  assign new_n1290_ = ~c & ~new_n1289_;
  assign new_n1291_ = h & l;
  assign new_n1292_ = i & ~new_n1291_;
  assign new_n1293_ = ~h & ~l;
  assign new_n1294_ = ~i & ~new_n1293_;
  assign new_n1295_ = ~new_n1292_ & ~new_n1294_;
  assign new_n1296_ = j & new_n1295_;
  assign new_n1297_ = g & ~new_n1296_;
  assign new_n1298_ = f & new_n1297_;
  assign new_n1299_ = e & new_n1298_;
  assign new_n1300_ = c & new_n1299_;
  assign new_n1301_ = ~new_n1290_ & ~new_n1300_;
  assign new_n1302_ = ~new_n1285_ & new_n1301_;
  assign new_n1303_ = ~new_n1275_ & new_n1302_;
  assign new_n1304_ = d & ~new_n1303_;
  assign new_n1305_ = ~i & ~new_n782_;
  assign new_n1306_ = h & new_n698_;
  assign new_n1307_ = i & ~new_n1306_;
  assign new_n1308_ = ~new_n1305_ & ~new_n1307_;
  assign new_n1309_ = ~g & ~new_n1308_;
  assign new_n1310_ = ~c & new_n1309_;
  assign new_n1311_ = g & new_n700_;
  assign new_n1312_ = new_n1137_ & new_n1311_;
  assign new_n1313_ = ~new_n1310_ & ~new_n1312_;
  assign new_n1314_ = ~new_n136_ & ~new_n1313_;
  assign new_n1315_ = ~g & new_n697_;
  assign new_n1316_ = new_n832_ & new_n1102_;
  assign new_n1317_ = ~new_n1315_ & ~new_n1316_;
  assign new_n1318_ = l & ~new_n1317_;
  assign new_n1319_ = h & ~i;
  assign new_n1320_ = i & ~l;
  assign new_n1321_ = ~new_n1319_ & ~new_n1320_;
  assign new_n1322_ = ~new_n632_ & ~new_n1321_;
  assign new_n1323_ = d & ~new_n71_;
  assign new_n1324_ = ~new_n698_ & ~new_n1323_;
  assign new_n1325_ = ~d & ~new_n98_;
  assign new_n1326_ = e & new_n580_;
  assign new_n1327_ = ~h & ~new_n1326_;
  assign new_n1328_ = ~new_n1325_ & ~new_n1327_;
  assign new_n1329_ = ~new_n1324_ & new_n1328_;
  assign new_n1330_ = ~i & ~new_n1329_;
  assign new_n1331_ = ~new_n432_ & ~new_n594_;
  assign new_n1332_ = ~new_n97_ & ~new_n1331_;
  assign new_n1333_ = e & ~l;
  assign new_n1334_ = ~new_n1332_ & ~new_n1333_;
  assign new_n1335_ = ~f & ~new_n1334_;
  assign new_n1336_ = l & ~new_n429_;
  assign new_n1337_ = ~d & ~new_n1336_;
  assign new_n1338_ = h & ~new_n924_;
  assign new_n1339_ = ~l & ~new_n1338_;
  assign new_n1340_ = ~k & new_n1339_;
  assign new_n1341_ = ~new_n1337_ & ~new_n1340_;
  assign new_n1342_ = ~new_n1335_ & new_n1341_;
  assign new_n1343_ = ~new_n1330_ & new_n1342_;
  assign new_n1344_ = g & ~new_n1343_;
  assign new_n1345_ = ~new_n596_ & ~new_n1323_;
  assign new_n1346_ = ~e & new_n596_;
  assign new_n1347_ = ~new_n1325_ & ~new_n1346_;
  assign new_n1348_ = ~new_n1345_ & new_n1347_;
  assign new_n1349_ = ~j & ~new_n1348_;
  assign new_n1350_ = f & ~new_n924_;
  assign new_n1351_ = ~d & new_n1350_;
  assign new_n1352_ = ~new_n1349_ & ~new_n1351_;
  assign new_n1353_ = i & ~new_n1352_;
  assign new_n1354_ = ~e & ~new_n429_;
  assign new_n1355_ = g & ~new_n1354_;
  assign new_n1356_ = f & ~new_n1355_;
  assign new_n1357_ = ~d & new_n1356_;
  assign new_n1358_ = new_n701_ & new_n1319_;
  assign new_n1359_ = ~new_n1357_ & ~new_n1358_;
  assign new_n1360_ = ~new_n1353_ & new_n1359_;
  assign new_n1361_ = ~new_n1344_ & new_n1360_;
  assign new_n1362_ = ~new_n1322_ & new_n1361_;
  assign new_n1363_ = ~new_n1318_ & new_n1362_;
  assign new_n1364_ = ~c & ~new_n1363_;
  assign new_n1365_ = i & ~new_n835_;
  assign new_n1366_ = ~d & ~new_n1365_;
  assign new_n1367_ = h & ~new_n835_;
  assign new_n1368_ = ~i & ~new_n698_;
  assign new_n1369_ = ~new_n594_ & ~new_n1368_;
  assign new_n1370_ = ~new_n1367_ & new_n1369_;
  assign new_n1371_ = g & ~new_n1370_;
  assign new_n1372_ = g & ~new_n835_;
  assign new_n1373_ = ~h & ~new_n1372_;
  assign new_n1374_ = j & ~new_n1270_;
  assign new_n1375_ = ~i & ~new_n676_;
  assign new_n1376_ = ~g & ~new_n1375_;
  assign new_n1377_ = l & ~new_n666_;
  assign new_n1378_ = ~new_n1376_ & new_n1377_;
  assign new_n1379_ = ~new_n1374_ & new_n1378_;
  assign new_n1380_ = ~new_n1373_ & new_n1379_;
  assign new_n1381_ = ~new_n1371_ & new_n1380_;
  assign new_n1382_ = ~new_n1366_ & new_n1381_;
  assign new_n1383_ = ~e & ~new_n1382_;
  assign new_n1384_ = h & new_n701_;
  assign new_n1385_ = h & ~new_n1384_;
  assign new_n1386_ = e & ~new_n1385_;
  assign new_n1387_ = ~new_n1293_ & ~new_n1386_;
  assign new_n1388_ = ~i & ~new_n1387_;
  assign new_n1389_ = new_n429_ & new_n580_;
  assign new_n1390_ = ~j & new_n782_;
  assign new_n1391_ = ~new_n1389_ & ~new_n1390_;
  assign new_n1392_ = h & ~new_n1391_;
  assign new_n1393_ = ~k & ~new_n1336_;
  assign new_n1394_ = ~h & new_n1393_;
  assign new_n1395_ = ~new_n1392_ & ~new_n1394_;
  assign new_n1396_ = ~new_n1388_ & new_n1395_;
  assign new_n1397_ = ~new_n1383_ & new_n1396_;
  assign new_n1398_ = ~f & ~new_n1397_;
  assign new_n1399_ = f & l;
  assign new_n1400_ = d & ~new_n1399_;
  assign new_n1401_ = ~new_n1385_ & ~new_n1400_;
  assign new_n1402_ = g & ~new_n1184_;
  assign new_n1403_ = ~h & ~new_n1402_;
  assign new_n1404_ = ~new_n1401_ & ~new_n1403_;
  assign new_n1405_ = ~i & ~new_n1404_;
  assign new_n1406_ = e & ~new_n1270_;
  assign new_n1407_ = f & i;
  assign new_n1408_ = ~g & ~l;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1410_ = ~new_n1406_ & new_n1409_;
  assign new_n1411_ = ~j & ~new_n1410_;
  assign new_n1412_ = h & new_n1411_;
  assign new_n1413_ = ~g & new_n1280_;
  assign new_n1414_ = ~new_n1412_ & ~new_n1413_;
  assign new_n1415_ = ~k & ~new_n1414_;
  assign new_n1416_ = new_n946_ & new_n1137_;
  assign new_n1417_ = ~new_n1415_ & ~new_n1416_;
  assign new_n1418_ = ~new_n1405_ & new_n1417_;
  assign new_n1419_ = ~new_n1398_ & new_n1418_;
  assign new_n1420_ = c & ~new_n1419_;
  assign new_n1421_ = g & new_n923_;
  assign new_n1422_ = ~f & new_n924_;
  assign new_n1423_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1424_ = ~d & ~new_n1423_;
  assign new_n1425_ = ~g & ~new_n925_;
  assign new_n1426_ = j & ~new_n541_;
  assign new_n1427_ = l & ~new_n1426_;
  assign new_n1428_ = ~h & ~new_n1427_;
  assign new_n1429_ = h & new_n122_;
  assign new_n1430_ = ~new_n1428_ & ~new_n1429_;
  assign new_n1431_ = ~new_n1425_ & new_n1430_;
  assign new_n1432_ = ~new_n1424_ & new_n1431_;
  assign new_n1433_ = ~k & ~new_n1432_;
  assign new_n1434_ = ~new_n72_ & ~new_n558_;
  assign new_n1435_ = l & ~new_n1434_;
  assign new_n1436_ = k & new_n1435_;
  assign new_n1437_ = j & new_n1436_;
  assign new_n1438_ = h & new_n1437_;
  assign new_n1439_ = ~new_n1433_ & ~new_n1438_;
  assign new_n1440_ = i & ~new_n1439_;
  assign new_n1441_ = i & ~new_n1390_;
  assign new_n1442_ = ~e & ~new_n1441_;
  assign new_n1443_ = ~g & ~new_n787_;
  assign new_n1444_ = ~new_n1442_ & ~new_n1443_;
  assign new_n1445_ = f & ~new_n1444_;
  assign new_n1446_ = d & k;
  assign new_n1447_ = ~f & ~new_n1446_;
  assign new_n1448_ = j & ~new_n1447_;
  assign new_n1449_ = g & ~new_n1448_;
  assign new_n1450_ = ~g & k;
  assign new_n1451_ = ~new_n1449_ & ~new_n1450_;
  assign new_n1452_ = ~i & ~new_n1451_;
  assign new_n1453_ = ~new_n1445_ & ~new_n1452_;
  assign new_n1454_ = ~h & ~new_n1453_;
  assign new_n1455_ = ~new_n847_ & ~new_n1270_;
  assign new_n1456_ = ~k & ~new_n1455_;
  assign new_n1457_ = ~j & new_n1456_;
  assign new_n1458_ = h & new_n1457_;
  assign new_n1459_ = ~new_n1454_ & ~new_n1458_;
  assign new_n1460_ = ~new_n1440_ & new_n1459_;
  assign new_n1461_ = ~new_n1420_ & new_n1460_;
  assign new_n1462_ = ~new_n1364_ & new_n1461_;
  assign new_n1463_ = ~new_n1314_ & new_n1462_;
  assign new_n1464_ = ~new_n1304_ & new_n1463_;
  assign new_n1465_ = ~m & ~new_n1464_;
  assign new_n1466_ = ~new_n1269_ & ~new_n1465_;
  assign new_n1467_ = ~n & ~new_n1466_;
  assign new_n1468_ = new_n647_ & new_n1210_;
  assign new_n1469_ = h & ~new_n1468_;
  assign new_n1470_ = ~new_n782_ & ~new_n1469_;
  assign new_n1471_ = ~h & ~new_n201_;
  assign new_n1472_ = c & d;
  assign new_n1473_ = b & new_n1472_;
  assign new_n1474_ = e & new_n1155_;
  assign new_n1475_ = new_n1473_ & new_n1474_;
  assign new_n1476_ = ~new_n1471_ & ~new_n1475_;
  assign new_n1477_ = ~new_n1470_ & new_n1476_;
  assign new_n1478_ = f & ~new_n1477_;
  assign new_n1479_ = ~b & k;
  assign new_n1480_ = e & ~new_n1479_;
  assign new_n1481_ = l & ~new_n1480_;
  assign new_n1482_ = ~f & ~new_n1481_;
  assign new_n1483_ = b & k;
  assign new_n1484_ = g & ~new_n1483_;
  assign new_n1485_ = l & ~new_n1484_;
  assign new_n1486_ = ~e & ~new_n1485_;
  assign new_n1487_ = new_n1033_ & new_n1472_;
  assign new_n1488_ = ~new_n1486_ & new_n1487_;
  assign new_n1489_ = ~new_n1482_ & new_n1488_;
  assign new_n1490_ = ~h & ~new_n1489_;
  assign new_n1491_ = d & new_n72_;
  assign new_n1492_ = new_n1210_ & new_n1491_;
  assign new_n1493_ = ~new_n979_ & ~new_n1492_;
  assign new_n1494_ = ~h & new_n698_;
  assign new_n1495_ = ~new_n1493_ & ~new_n1494_;
  assign new_n1496_ = ~f & new_n1495_;
  assign new_n1497_ = ~k & ~new_n176_;
  assign new_n1498_ = ~j & new_n1497_;
  assign new_n1499_ = h & new_n1498_;
  assign new_n1500_ = ~new_n1496_ & ~new_n1499_;
  assign new_n1501_ = ~new_n1490_ & new_n1500_;
  assign new_n1502_ = ~new_n1478_ & new_n1501_;
  assign new_n1503_ = ~i & ~new_n1502_;
  assign new_n1504_ = c & new_n86_;
  assign new_n1505_ = new_n146_ & ~new_n843_;
  assign new_n1506_ = new_n1504_ & new_n1505_;
  assign new_n1507_ = new_n700_ & new_n1137_;
  assign new_n1508_ = ~h & new_n782_;
  assign new_n1509_ = ~new_n1507_ & ~new_n1508_;
  assign new_n1510_ = ~new_n1506_ & ~new_n1509_;
  assign new_n1511_ = new_n97_ & new_n1210_;
  assign new_n1512_ = ~new_n979_ & ~new_n1511_;
  assign new_n1513_ = k & ~new_n1512_;
  assign new_n1514_ = ~f & new_n1513_;
  assign new_n1515_ = ~new_n1508_ & ~new_n1514_;
  assign new_n1516_ = ~new_n781_ & ~new_n1515_;
  assign new_n1517_ = f & new_n142_;
  assign new_n1518_ = ~new_n1011_ & ~new_n1517_;
  assign new_n1519_ = ~h & ~new_n1518_;
  assign new_n1520_ = d & ~i;
  assign new_n1521_ = ~j & new_n117_;
  assign new_n1522_ = new_n1520_ & new_n1521_;
  assign new_n1523_ = ~g & ~new_n1522_;
  assign new_n1524_ = ~f & new_n1523_;
  assign new_n1525_ = ~new_n1519_ & ~new_n1524_;
  assign new_n1526_ = ~new_n201_ & ~new_n1525_;
  assign new_n1527_ = e & new_n558_;
  assign new_n1528_ = ~new_n72_ & ~new_n1527_;
  assign new_n1529_ = ~d & ~new_n1528_;
  assign new_n1530_ = ~g & ~new_n102_;
  assign new_n1531_ = ~f & new_n1530_;
  assign new_n1532_ = ~k & ~new_n925_;
  assign new_n1533_ = b & ~new_n1532_;
  assign new_n1534_ = ~new_n1531_ & new_n1533_;
  assign new_n1535_ = ~new_n1529_ & new_n1534_;
  assign new_n1536_ = ~c & ~new_n1535_;
  assign new_n1537_ = ~b & new_n72_;
  assign new_n1538_ = d & ~new_n1537_;
  assign new_n1539_ = ~new_n925_ & ~new_n1538_;
  assign new_n1540_ = b & ~new_n72_;
  assign new_n1541_ = ~b & i;
  assign new_n1542_ = l & ~new_n1541_;
  assign new_n1543_ = ~e & ~new_n1542_;
  assign new_n1544_ = ~g & ~new_n1076_;
  assign new_n1545_ = f & ~i;
  assign new_n1546_ = ~l & ~new_n1545_;
  assign new_n1547_ = ~f & ~new_n1546_;
  assign new_n1548_ = ~new_n1544_ & new_n1547_;
  assign new_n1549_ = ~new_n1543_ & new_n1548_;
  assign new_n1550_ = ~new_n1540_ & new_n1549_;
  assign new_n1551_ = ~j & ~new_n1550_;
  assign new_n1552_ = h & new_n1551_;
  assign new_n1553_ = g & i;
  assign new_n1554_ = f & new_n1553_;
  assign new_n1555_ = new_n1472_ & new_n1554_;
  assign new_n1556_ = ~f & new_n923_;
  assign new_n1557_ = ~new_n1555_ & ~new_n1556_;
  assign new_n1558_ = e & ~new_n1557_;
  assign new_n1559_ = new_n40_ & new_n429_;
  assign new_n1560_ = ~new_n1558_ & ~new_n1559_;
  assign new_n1561_ = b & ~new_n1560_;
  assign new_n1562_ = i & ~new_n71_;
  assign new_n1563_ = g & ~new_n1562_;
  assign new_n1564_ = j & ~new_n1563_;
  assign new_n1565_ = ~h & new_n1564_;
  assign new_n1566_ = ~new_n1561_ & ~new_n1565_;
  assign new_n1567_ = ~new_n1552_ & new_n1566_;
  assign new_n1568_ = ~new_n1539_ & new_n1567_;
  assign new_n1569_ = ~k & ~new_n1568_;
  assign new_n1570_ = ~new_n219_ & ~new_n979_;
  assign new_n1571_ = ~g & ~new_n1570_;
  assign new_n1572_ = l & ~new_n707_;
  assign new_n1573_ = ~new_n432_ & new_n1572_;
  assign new_n1574_ = ~new_n1512_ & ~new_n1573_;
  assign new_n1575_ = ~b & new_n102_;
  assign new_n1576_ = ~e & new_n429_;
  assign new_n1577_ = new_n1473_ & new_n1576_;
  assign new_n1578_ = ~new_n1575_ & ~new_n1577_;
  assign new_n1579_ = ~new_n1574_ & new_n1578_;
  assign new_n1580_ = ~new_n1571_ & new_n1579_;
  assign new_n1581_ = ~f & ~new_n1580_;
  assign new_n1582_ = j & ~new_n1292_;
  assign new_n1583_ = g & ~new_n1582_;
  assign new_n1584_ = f & new_n1583_;
  assign new_n1585_ = e & new_n1584_;
  assign new_n1586_ = d & new_n1585_;
  assign new_n1587_ = c & new_n1586_;
  assign new_n1588_ = b & new_n1587_;
  assign new_n1589_ = ~new_n1581_ & ~new_n1588_;
  assign new_n1590_ = ~new_n1569_ & new_n1589_;
  assign new_n1591_ = ~new_n1536_ & new_n1590_;
  assign new_n1592_ = ~new_n1526_ & new_n1591_;
  assign new_n1593_ = ~new_n1516_ & new_n1592_;
  assign new_n1594_ = ~new_n1510_ & new_n1593_;
  assign new_n1595_ = ~new_n1503_ & new_n1594_;
  assign new_n1596_ = n & ~new_n1595_;
  assign new_n1597_ = ~m & new_n1596_;
  assign l2 = new_n1467_ | new_n1597_;
endmodule


