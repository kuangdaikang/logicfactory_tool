// Benchmark "i5" written by ABC on Fri Feb 25 15:13:09 2022

module i5 ( 
    \V4(0) , \V2(1) , \V4(1) , \V2(0) , \V28(1) , \V16(2) , \V28(2) ,
    \V16(3) , \V28(3) , \V28(5) , \V16(6) , \V28(6) , \V16(7) , \V28(7) ,
    \V28(9) , \V16(10) , \V28(10) , \V16(11) , \V28(11) , \V28(13) ,
    \V16(14) , \V28(14) , \V16(15) , \V28(15) , \V16(1) , \V16(5) ,
    \V16(9) , \V16(13) , \V52(1) , \V40(2) , \V52(2) , \V40(3) , \V52(3) ,
    \V52(5) , \V40(6) , \V52(6) , \V40(7) , \V52(7) , \V52(9) , \V40(10) ,
    \V52(10) , \V40(11) , \V52(11) , \V52(13) , \V40(14) , \V52(14) ,
    \V40(15) , \V52(15) , \V40(1) , \V40(5) , \V40(9) , \V40(13) ,
    \V76(1) , \V64(2) , \V76(2) , \V64(3) , \V76(3) , \V76(5) , \V64(6) ,
    \V76(6) , \V64(7) , \V76(7) , \V76(9) , \V64(10) , \V76(10) ,
    \V64(11) , \V76(11) , \V76(13) , \V64(14) , \V76(14) , \V64(15) ,
    \V76(15) , \V64(1) , \V64(5) , \V64(9) , \V64(13) , \V100(1) ,
    \V88(2) , \V100(2) , \V88(3) , \V100(3) , \V100(5) , \V88(6) ,
    \V100(6) , \V88(7) , \V100(7) , \V100(9) , \V88(10) , \V100(10) ,
    \V88(11) , \V100(11) , \V100(13) , \V88(14) , \V100(14) , \V88(15) ,
    \V133(0) , \V100(15) , \V88(1) , \V88(5) , \V88(9) , \V88(13) ,
    \V106(1) , \V103(2) , \V106(2) , \V103(3) , \V106(3) , \V112(1) ,
    \V109(2) , \V112(2) , \V109(3) , \V112(3) , \V118(1) , \V115(2) ,
    \V118(2) , \V115(3) , \V118(3) , \V124(1) , \V121(2) , \V124(2) ,
    \V121(3) , \V124(3) , \V103(1) , \V109(1) , \V115(1) , \V121(1) ,
    \V132(0) , \V128(1) , \V132(1) , \V128(2) , \V132(2) , \V128(3) ,
    \V132(3) , \V128(0) ,
    \V135(0) , \V135(1) , \V151(1) , \V151(2) , \V151(3) , \V151(5) ,
    \V151(6) , \V151(7) , \V151(9) , \V151(10) , \V151(11) , \V151(13) ,
    \V151(14) , \V151(15) , \V167(1) , \V167(2) , \V167(3) , \V167(5) ,
    \V167(6) , \V167(7) , \V167(9) , \V167(10) , \V167(11) , \V167(13) ,
    \V167(14) , \V167(15) , \V183(1) , \V183(2) , \V183(3) , \V183(5) ,
    \V183(6) , \V183(7) , \V183(9) , \V183(10) , \V183(11) , \V183(13) ,
    \V183(14) , \V183(15) , \V199(1) , \V199(2) , \V199(3) , \V199(5) ,
    \V199(6) , \V199(7) , \V199(9) , \V199(10) , \V199(11) , \V199(13) ,
    \V199(14) , \V199(15) , \V151(4) , \V151(8) , \V151(12) , \V167(4) ,
    \V167(8) , \V167(12) , \V183(4) , \V183(8) , \V183(12) , \V199(4) ,
    \V199(8) , \V199(12) , \V151(0) , \V167(0) , \V183(0) , \V199(0)   );
  input  \V4(0) , \V2(1) , \V4(1) , \V2(0) , \V28(1) , \V16(2) ,
    \V28(2) , \V16(3) , \V28(3) , \V28(5) , \V16(6) , \V28(6) , \V16(7) ,
    \V28(7) , \V28(9) , \V16(10) , \V28(10) , \V16(11) , \V28(11) ,
    \V28(13) , \V16(14) , \V28(14) , \V16(15) , \V28(15) , \V16(1) ,
    \V16(5) , \V16(9) , \V16(13) , \V52(1) , \V40(2) , \V52(2) , \V40(3) ,
    \V52(3) , \V52(5) , \V40(6) , \V52(6) , \V40(7) , \V52(7) , \V52(9) ,
    \V40(10) , \V52(10) , \V40(11) , \V52(11) , \V52(13) , \V40(14) ,
    \V52(14) , \V40(15) , \V52(15) , \V40(1) , \V40(5) , \V40(9) ,
    \V40(13) , \V76(1) , \V64(2) , \V76(2) , \V64(3) , \V76(3) , \V76(5) ,
    \V64(6) , \V76(6) , \V64(7) , \V76(7) , \V76(9) , \V64(10) , \V76(10) ,
    \V64(11) , \V76(11) , \V76(13) , \V64(14) , \V76(14) , \V64(15) ,
    \V76(15) , \V64(1) , \V64(5) , \V64(9) , \V64(13) , \V100(1) ,
    \V88(2) , \V100(2) , \V88(3) , \V100(3) , \V100(5) , \V88(6) ,
    \V100(6) , \V88(7) , \V100(7) , \V100(9) , \V88(10) , \V100(10) ,
    \V88(11) , \V100(11) , \V100(13) , \V88(14) , \V100(14) , \V88(15) ,
    \V133(0) , \V100(15) , \V88(1) , \V88(5) , \V88(9) , \V88(13) ,
    \V106(1) , \V103(2) , \V106(2) , \V103(3) , \V106(3) , \V112(1) ,
    \V109(2) , \V112(2) , \V109(3) , \V112(3) , \V118(1) , \V115(2) ,
    \V118(2) , \V115(3) , \V118(3) , \V124(1) , \V121(2) , \V124(2) ,
    \V121(3) , \V124(3) , \V103(1) , \V109(1) , \V115(1) , \V121(1) ,
    \V132(0) , \V128(1) , \V132(1) , \V128(2) , \V132(2) , \V128(3) ,
    \V132(3) , \V128(0) ;
  output \V135(0) , \V135(1) , \V151(1) , \V151(2) , \V151(3) , \V151(5) ,
    \V151(6) , \V151(7) , \V151(9) , \V151(10) , \V151(11) , \V151(13) ,
    \V151(14) , \V151(15) , \V167(1) , \V167(2) , \V167(3) , \V167(5) ,
    \V167(6) , \V167(7) , \V167(9) , \V167(10) , \V167(11) , \V167(13) ,
    \V167(14) , \V167(15) , \V183(1) , \V183(2) , \V183(3) , \V183(5) ,
    \V183(6) , \V183(7) , \V183(9) , \V183(10) , \V183(11) , \V183(13) ,
    \V183(14) , \V183(15) , \V199(1) , \V199(2) , \V199(3) , \V199(5) ,
    \V199(6) , \V199(7) , \V199(9) , \V199(10) , \V199(11) , \V199(13) ,
    \V199(14) , \V199(15) , \V151(4) , \V151(8) , \V151(12) , \V167(4) ,
    \V167(8) , \V167(12) , \V183(4) , \V183(8) , \V183(12) , \V199(4) ,
    \V199(8) , \V199(12) , \V151(0) , \V167(0) , \V183(0) , \V199(0) ;
  wire new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_,
    new_n212_, new_n214_, new_n215_, new_n216_, new_n217_, new_n219_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n246_, new_n247_,
    new_n249_, new_n251_, new_n252_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n263_,
    new_n264_, new_n266_, new_n268_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n279_,
    new_n280_, new_n282_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n293_, new_n294_,
    new_n296_, new_n298_, new_n299_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n319_, new_n320_, new_n322_, new_n324_, new_n325_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n336_, new_n337_, new_n339_, new_n341_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n352_, new_n353_, new_n355_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n366_, new_n367_, new_n369_, new_n371_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n391_, new_n392_, new_n394_,
    new_n396_, new_n397_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n408_, new_n409_,
    new_n411_, new_n413_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n424_, new_n425_,
    new_n427_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n438_, new_n439_, new_n441_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n461_, new_n462_,
    new_n464_, new_n466_, new_n467_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n478_,
    new_n479_, new_n481_, new_n483_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n494_,
    new_n495_, new_n497_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n508_, new_n509_,
    new_n511_;
  assign new_n200_ = \V133(0)  & \V132(2) ;
  assign new_n201_ = \V132(0)  & new_n200_;
  assign new_n202_ = \V132(1)  & new_n201_;
  assign new_n203_ = \V132(3)  & new_n202_;
  assign new_n204_ = \V132(1)  & \V128(2) ;
  assign new_n205_ = \V132(0)  & new_n204_;
  assign new_n206_ = \V132(0)  & \V128(1) ;
  assign new_n207_ = \V132(0)  & \V132(2) ;
  assign new_n208_ = \V128(3)  & new_n207_;
  assign new_n209_ = \V132(1)  & new_n208_;
  assign new_n210_ = ~new_n203_ & ~new_n205_;
  assign new_n211_ = ~\V128(0)  & new_n210_;
  assign new_n212_ = ~new_n206_ & ~new_n209_;
  assign \V151(0)  = ~new_n211_ | ~new_n212_;
  assign new_n214_ = \V4(0)  & \V151(0) ;
  assign new_n215_ = \V4(1)  & new_n214_;
  assign new_n216_ = \V4(0)  & \V2(1) ;
  assign new_n217_ = ~\V2(0)  & ~new_n215_;
  assign \V135(0)  = new_n216_ | ~new_n217_;
  assign new_n219_ = \V4(1)  & \V151(0) ;
  assign \V135(1)  = \V2(1)  | new_n219_;
  assign new_n221_ = \V132(1)  & new_n200_;
  assign new_n222_ = \V132(3)  & new_n221_;
  assign new_n223_ = \V132(2)  & \V128(3) ;
  assign new_n224_ = \V132(1)  & new_n223_;
  assign new_n225_ = ~new_n204_ & ~new_n222_;
  assign new_n226_ = ~\V128(1)  & ~new_n224_;
  assign \V167(0)  = ~new_n225_ | ~new_n226_;
  assign new_n228_ = \V106(2)  & \V167(0) ;
  assign new_n229_ = \V106(1)  & new_n228_;
  assign new_n230_ = \V106(3)  & new_n229_;
  assign new_n231_ = \V106(1)  & \V103(2) ;
  assign new_n232_ = \V106(2)  & \V103(3) ;
  assign new_n233_ = \V106(1)  & new_n232_;
  assign new_n234_ = ~new_n230_ & ~new_n231_;
  assign new_n235_ = ~\V103(1)  & ~new_n233_;
  assign \V151(4)  = ~new_n234_ | ~new_n235_;
  assign new_n237_ = \V28(2)  & \V151(4) ;
  assign new_n238_ = \V28(1)  & new_n237_;
  assign new_n239_ = \V28(3)  & new_n238_;
  assign new_n240_ = \V28(1)  & \V16(2) ;
  assign new_n241_ = \V28(2)  & \V16(3) ;
  assign new_n242_ = \V28(1)  & new_n241_;
  assign new_n243_ = ~new_n239_ & ~new_n240_;
  assign new_n244_ = ~\V16(1)  & ~new_n242_;
  assign \V151(1)  = ~new_n243_ | ~new_n244_;
  assign new_n246_ = \V28(3)  & new_n237_;
  assign new_n247_ = ~\V16(2)  & ~new_n246_;
  assign \V151(2)  = new_n241_ | ~new_n247_;
  assign new_n249_ = \V28(3)  & \V151(4) ;
  assign \V151(3)  = \V16(3)  | new_n249_;
  assign new_n251_ = \V106(3)  & new_n228_;
  assign new_n252_ = ~\V103(2)  & ~new_n251_;
  assign \V151(8)  = new_n232_ | ~new_n252_;
  assign new_n254_ = \V28(6)  & \V151(8) ;
  assign new_n255_ = \V28(5)  & new_n254_;
  assign new_n256_ = \V28(7)  & new_n255_;
  assign new_n257_ = \V28(5)  & \V16(6) ;
  assign new_n258_ = \V28(6)  & \V16(7) ;
  assign new_n259_ = \V28(5)  & new_n258_;
  assign new_n260_ = ~new_n256_ & ~new_n257_;
  assign new_n261_ = ~\V16(5)  & ~new_n259_;
  assign \V151(5)  = ~new_n260_ | ~new_n261_;
  assign new_n263_ = \V28(7)  & new_n254_;
  assign new_n264_ = ~\V16(6)  & ~new_n263_;
  assign \V151(6)  = new_n258_ | ~new_n264_;
  assign new_n266_ = \V28(7)  & \V151(8) ;
  assign \V151(7)  = \V16(7)  | new_n266_;
  assign new_n268_ = \V106(3)  & \V167(0) ;
  assign \V151(12)  = \V103(3)  | new_n268_;
  assign new_n270_ = \V28(10)  & \V151(12) ;
  assign new_n271_ = \V28(9)  & new_n270_;
  assign new_n272_ = \V28(11)  & new_n271_;
  assign new_n273_ = \V28(9)  & \V16(10) ;
  assign new_n274_ = \V28(10)  & \V16(11) ;
  assign new_n275_ = \V28(9)  & new_n274_;
  assign new_n276_ = ~new_n272_ & ~new_n273_;
  assign new_n277_ = ~\V16(9)  & ~new_n275_;
  assign \V151(9)  = ~new_n276_ | ~new_n277_;
  assign new_n279_ = \V28(11)  & new_n270_;
  assign new_n280_ = ~\V16(10)  & ~new_n279_;
  assign \V151(10)  = new_n274_ | ~new_n280_;
  assign new_n282_ = \V28(11)  & \V151(12) ;
  assign \V151(11)  = \V16(11)  | new_n282_;
  assign new_n284_ = \V28(14)  & \V167(0) ;
  assign new_n285_ = \V28(13)  & new_n284_;
  assign new_n286_ = \V28(15)  & new_n285_;
  assign new_n287_ = \V28(13)  & \V16(14) ;
  assign new_n288_ = \V28(14)  & \V16(15) ;
  assign new_n289_ = \V28(13)  & new_n288_;
  assign new_n290_ = ~new_n286_ & ~new_n287_;
  assign new_n291_ = ~\V16(13)  & ~new_n289_;
  assign \V151(13)  = ~new_n290_ | ~new_n291_;
  assign new_n293_ = \V28(15)  & new_n284_;
  assign new_n294_ = ~\V16(14)  & ~new_n293_;
  assign \V151(14)  = new_n288_ | ~new_n294_;
  assign new_n296_ = \V28(15)  & \V167(0) ;
  assign \V151(15)  = \V16(15)  | new_n296_;
  assign new_n298_ = \V132(3)  & new_n200_;
  assign new_n299_ = ~\V128(2)  & ~new_n298_;
  assign \V183(0)  = new_n223_ | ~new_n299_;
  assign new_n301_ = \V112(2)  & \V183(0) ;
  assign new_n302_ = \V112(1)  & new_n301_;
  assign new_n303_ = \V112(3)  & new_n302_;
  assign new_n304_ = \V112(1)  & \V109(2) ;
  assign new_n305_ = \V112(2)  & \V109(3) ;
  assign new_n306_ = \V112(1)  & new_n305_;
  assign new_n307_ = ~new_n303_ & ~new_n304_;
  assign new_n308_ = ~\V109(1)  & ~new_n306_;
  assign \V167(4)  = ~new_n307_ | ~new_n308_;
  assign new_n310_ = \V52(2)  & \V167(4) ;
  assign new_n311_ = \V52(1)  & new_n310_;
  assign new_n312_ = \V52(3)  & new_n311_;
  assign new_n313_ = \V52(1)  & \V40(2) ;
  assign new_n314_ = \V52(2)  & \V40(3) ;
  assign new_n315_ = \V52(1)  & new_n314_;
  assign new_n316_ = ~new_n312_ & ~new_n313_;
  assign new_n317_ = ~\V40(1)  & ~new_n315_;
  assign \V167(1)  = ~new_n316_ | ~new_n317_;
  assign new_n319_ = \V52(3)  & new_n310_;
  assign new_n320_ = ~\V40(2)  & ~new_n319_;
  assign \V167(2)  = new_n314_ | ~new_n320_;
  assign new_n322_ = \V52(3)  & \V167(4) ;
  assign \V167(3)  = \V40(3)  | new_n322_;
  assign new_n324_ = \V112(3)  & new_n301_;
  assign new_n325_ = ~\V109(2)  & ~new_n324_;
  assign \V167(8)  = new_n305_ | ~new_n325_;
  assign new_n327_ = \V52(6)  & \V167(8) ;
  assign new_n328_ = \V52(5)  & new_n327_;
  assign new_n329_ = \V52(7)  & new_n328_;
  assign new_n330_ = \V52(5)  & \V40(6) ;
  assign new_n331_ = \V52(6)  & \V40(7) ;
  assign new_n332_ = \V52(5)  & new_n331_;
  assign new_n333_ = ~new_n329_ & ~new_n330_;
  assign new_n334_ = ~\V40(5)  & ~new_n332_;
  assign \V167(5)  = ~new_n333_ | ~new_n334_;
  assign new_n336_ = \V52(7)  & new_n327_;
  assign new_n337_ = ~\V40(6)  & ~new_n336_;
  assign \V167(6)  = new_n331_ | ~new_n337_;
  assign new_n339_ = \V52(7)  & \V167(8) ;
  assign \V167(7)  = \V40(7)  | new_n339_;
  assign new_n341_ = \V112(3)  & \V183(0) ;
  assign \V167(12)  = \V109(3)  | new_n341_;
  assign new_n343_ = \V52(10)  & \V167(12) ;
  assign new_n344_ = \V52(9)  & new_n343_;
  assign new_n345_ = \V52(11)  & new_n344_;
  assign new_n346_ = \V52(9)  & \V40(10) ;
  assign new_n347_ = \V52(10)  & \V40(11) ;
  assign new_n348_ = \V52(9)  & new_n347_;
  assign new_n349_ = ~new_n345_ & ~new_n346_;
  assign new_n350_ = ~\V40(9)  & ~new_n348_;
  assign \V167(9)  = ~new_n349_ | ~new_n350_;
  assign new_n352_ = \V52(11)  & new_n343_;
  assign new_n353_ = ~\V40(10)  & ~new_n352_;
  assign \V167(10)  = new_n347_ | ~new_n353_;
  assign new_n355_ = \V52(11)  & \V167(12) ;
  assign \V167(11)  = \V40(11)  | new_n355_;
  assign new_n357_ = \V52(14)  & \V183(0) ;
  assign new_n358_ = \V52(13)  & new_n357_;
  assign new_n359_ = \V52(15)  & new_n358_;
  assign new_n360_ = \V52(13)  & \V40(14) ;
  assign new_n361_ = \V52(14)  & \V40(15) ;
  assign new_n362_ = \V52(13)  & new_n361_;
  assign new_n363_ = ~new_n359_ & ~new_n360_;
  assign new_n364_ = ~\V40(13)  & ~new_n362_;
  assign \V167(13)  = ~new_n363_ | ~new_n364_;
  assign new_n366_ = \V52(15)  & new_n357_;
  assign new_n367_ = ~\V40(14)  & ~new_n366_;
  assign \V167(14)  = new_n361_ | ~new_n367_;
  assign new_n369_ = \V52(15)  & \V183(0) ;
  assign \V167(15)  = \V40(15)  | new_n369_;
  assign new_n371_ = \V133(0)  & \V132(3) ;
  assign \V199(0)  = \V128(3)  | new_n371_;
  assign new_n373_ = \V118(2)  & \V199(0) ;
  assign new_n374_ = \V118(1)  & new_n373_;
  assign new_n375_ = \V118(3)  & new_n374_;
  assign new_n376_ = \V118(1)  & \V115(2) ;
  assign new_n377_ = \V118(2)  & \V115(3) ;
  assign new_n378_ = \V118(1)  & new_n377_;
  assign new_n379_ = ~new_n375_ & ~new_n376_;
  assign new_n380_ = ~\V115(1)  & ~new_n378_;
  assign \V183(4)  = ~new_n379_ | ~new_n380_;
  assign new_n382_ = \V76(2)  & \V183(4) ;
  assign new_n383_ = \V76(1)  & new_n382_;
  assign new_n384_ = \V76(3)  & new_n383_;
  assign new_n385_ = \V76(1)  & \V64(2) ;
  assign new_n386_ = \V76(2)  & \V64(3) ;
  assign new_n387_ = \V76(1)  & new_n386_;
  assign new_n388_ = ~new_n384_ & ~new_n385_;
  assign new_n389_ = ~\V64(1)  & ~new_n387_;
  assign \V183(1)  = ~new_n388_ | ~new_n389_;
  assign new_n391_ = \V76(3)  & new_n382_;
  assign new_n392_ = ~\V64(2)  & ~new_n391_;
  assign \V183(2)  = new_n386_ | ~new_n392_;
  assign new_n394_ = \V76(3)  & \V183(4) ;
  assign \V183(3)  = \V64(3)  | new_n394_;
  assign new_n396_ = \V118(3)  & new_n373_;
  assign new_n397_ = ~\V115(2)  & ~new_n396_;
  assign \V183(8)  = new_n377_ | ~new_n397_;
  assign new_n399_ = \V76(6)  & \V183(8) ;
  assign new_n400_ = \V76(5)  & new_n399_;
  assign new_n401_ = \V76(7)  & new_n400_;
  assign new_n402_ = \V76(5)  & \V64(6) ;
  assign new_n403_ = \V76(6)  & \V64(7) ;
  assign new_n404_ = \V76(5)  & new_n403_;
  assign new_n405_ = ~new_n401_ & ~new_n402_;
  assign new_n406_ = ~\V64(5)  & ~new_n404_;
  assign \V183(5)  = ~new_n405_ | ~new_n406_;
  assign new_n408_ = \V76(7)  & new_n399_;
  assign new_n409_ = ~\V64(6)  & ~new_n408_;
  assign \V183(6)  = new_n403_ | ~new_n409_;
  assign new_n411_ = \V76(7)  & \V183(8) ;
  assign \V183(7)  = \V64(7)  | new_n411_;
  assign new_n413_ = \V118(3)  & \V199(0) ;
  assign \V183(12)  = \V115(3)  | new_n413_;
  assign new_n415_ = \V76(10)  & \V183(12) ;
  assign new_n416_ = \V76(9)  & new_n415_;
  assign new_n417_ = \V76(11)  & new_n416_;
  assign new_n418_ = \V76(9)  & \V64(10) ;
  assign new_n419_ = \V76(10)  & \V64(11) ;
  assign new_n420_ = \V76(9)  & new_n419_;
  assign new_n421_ = ~new_n417_ & ~new_n418_;
  assign new_n422_ = ~\V64(9)  & ~new_n420_;
  assign \V183(9)  = ~new_n421_ | ~new_n422_;
  assign new_n424_ = \V76(11)  & new_n415_;
  assign new_n425_ = ~\V64(10)  & ~new_n424_;
  assign \V183(10)  = new_n419_ | ~new_n425_;
  assign new_n427_ = \V76(11)  & \V183(12) ;
  assign \V183(11)  = \V64(11)  | new_n427_;
  assign new_n429_ = \V76(14)  & \V199(0) ;
  assign new_n430_ = \V76(13)  & new_n429_;
  assign new_n431_ = \V76(15)  & new_n430_;
  assign new_n432_ = \V76(13)  & \V64(14) ;
  assign new_n433_ = \V76(14)  & \V64(15) ;
  assign new_n434_ = \V76(13)  & new_n433_;
  assign new_n435_ = ~new_n431_ & ~new_n432_;
  assign new_n436_ = ~\V64(13)  & ~new_n434_;
  assign \V183(13)  = ~new_n435_ | ~new_n436_;
  assign new_n438_ = \V76(15)  & new_n429_;
  assign new_n439_ = ~\V64(14)  & ~new_n438_;
  assign \V183(14)  = new_n433_ | ~new_n439_;
  assign new_n441_ = \V76(15)  & \V199(0) ;
  assign \V183(15)  = \V64(15)  | new_n441_;
  assign new_n443_ = \V133(0)  & \V124(2) ;
  assign new_n444_ = \V124(1)  & new_n443_;
  assign new_n445_ = \V124(3)  & new_n444_;
  assign new_n446_ = \V124(1)  & \V121(2) ;
  assign new_n447_ = \V124(2)  & \V121(3) ;
  assign new_n448_ = \V124(1)  & new_n447_;
  assign new_n449_ = ~new_n445_ & ~new_n446_;
  assign new_n450_ = ~\V121(1)  & ~new_n448_;
  assign \V199(4)  = ~new_n449_ | ~new_n450_;
  assign new_n452_ = \V100(2)  & \V199(4) ;
  assign new_n453_ = \V100(1)  & new_n452_;
  assign new_n454_ = \V100(3)  & new_n453_;
  assign new_n455_ = \V100(1)  & \V88(2) ;
  assign new_n456_ = \V100(2)  & \V88(3) ;
  assign new_n457_ = \V100(1)  & new_n456_;
  assign new_n458_ = ~new_n454_ & ~new_n455_;
  assign new_n459_ = ~\V88(1)  & ~new_n457_;
  assign \V199(1)  = ~new_n458_ | ~new_n459_;
  assign new_n461_ = \V100(3)  & new_n452_;
  assign new_n462_ = ~\V88(2)  & ~new_n461_;
  assign \V199(2)  = new_n456_ | ~new_n462_;
  assign new_n464_ = \V100(3)  & \V199(4) ;
  assign \V199(3)  = \V88(3)  | new_n464_;
  assign new_n466_ = \V124(3)  & new_n443_;
  assign new_n467_ = ~\V121(2)  & ~new_n466_;
  assign \V199(8)  = new_n447_ | ~new_n467_;
  assign new_n469_ = \V100(6)  & \V199(8) ;
  assign new_n470_ = \V100(5)  & new_n469_;
  assign new_n471_ = \V100(7)  & new_n470_;
  assign new_n472_ = \V100(5)  & \V88(6) ;
  assign new_n473_ = \V100(6)  & \V88(7) ;
  assign new_n474_ = \V100(5)  & new_n473_;
  assign new_n475_ = ~new_n471_ & ~new_n472_;
  assign new_n476_ = ~\V88(5)  & ~new_n474_;
  assign \V199(5)  = ~new_n475_ | ~new_n476_;
  assign new_n478_ = \V100(7)  & new_n469_;
  assign new_n479_ = ~\V88(6)  & ~new_n478_;
  assign \V199(6)  = new_n473_ | ~new_n479_;
  assign new_n481_ = \V100(7)  & \V199(8) ;
  assign \V199(7)  = \V88(7)  | new_n481_;
  assign new_n483_ = \V133(0)  & \V124(3) ;
  assign \V199(12)  = \V121(3)  | new_n483_;
  assign new_n485_ = \V100(10)  & \V199(12) ;
  assign new_n486_ = \V100(9)  & new_n485_;
  assign new_n487_ = \V100(11)  & new_n486_;
  assign new_n488_ = \V100(9)  & \V88(10) ;
  assign new_n489_ = \V100(10)  & \V88(11) ;
  assign new_n490_ = \V100(9)  & new_n489_;
  assign new_n491_ = ~new_n487_ & ~new_n488_;
  assign new_n492_ = ~\V88(9)  & ~new_n490_;
  assign \V199(9)  = ~new_n491_ | ~new_n492_;
  assign new_n494_ = \V100(11)  & new_n485_;
  assign new_n495_ = ~\V88(10)  & ~new_n494_;
  assign \V199(10)  = new_n489_ | ~new_n495_;
  assign new_n497_ = \V100(11)  & \V199(12) ;
  assign \V199(11)  = \V88(11)  | new_n497_;
  assign new_n499_ = \V100(14)  & \V133(0) ;
  assign new_n500_ = \V100(13)  & new_n499_;
  assign new_n501_ = \V100(15)  & new_n500_;
  assign new_n502_ = \V100(13)  & \V88(14) ;
  assign new_n503_ = \V100(14)  & \V88(15) ;
  assign new_n504_ = \V100(13)  & new_n503_;
  assign new_n505_ = ~new_n501_ & ~new_n502_;
  assign new_n506_ = ~\V88(13)  & ~new_n504_;
  assign \V199(13)  = ~new_n505_ | ~new_n506_;
  assign new_n508_ = \V100(15)  & new_n499_;
  assign new_n509_ = ~\V88(14)  & ~new_n508_;
  assign \V199(14)  = new_n503_ | ~new_n509_;
  assign new_n511_ = \V133(0)  & \V100(15) ;
  assign \V199(15)  = \V88(15)  | new_n511_;
endmodule


