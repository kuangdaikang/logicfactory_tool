// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:57 2022

module t2  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16,
    \v17.0 , \v17.1 , \v17.2 , \v17.3 , \v17.4 , \v17.5 , \v17.6 , \v17.7 ,
    \v17.8 , \v17.9 , \v17.10 , \v17.11 , \v17.12 , \v17.13 , \v17.14 ,
    \v17.15   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16;
  output \v17.0 , \v17.1 , \v17.2 , \v17.3 , \v17.4 , \v17.5 , \v17.6 ,
    \v17.7 , \v17.8 , \v17.9 , \v17.10 , \v17.11 , \v17.12 , \v17.13 ,
    \v17.14 , \v17.15 ;
  wire new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n60_, new_n61_, new_n62_,
    new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_,
    new_n194_, new_n196_, new_n197_, new_n198_, new_n199_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n237_, new_n239_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_;
  assign new_n34_ = ~v2 & ~v6;
  assign new_n35_ = ~v6 & ~new_n34_;
  assign new_n36_ = ~v11 & ~new_n35_;
  assign new_n37_ = ~v4 & new_n36_;
  assign new_n38_ = v3 & new_n37_;
  assign new_n39_ = v1 & new_n38_;
  assign new_n40_ = ~v11 & ~new_n39_;
  assign new_n41_ = ~v16 & ~new_n40_;
  assign new_n42_ = v11 & v16;
  assign new_n43_ = ~new_n41_ & ~new_n42_;
  assign new_n44_ = ~v15 & ~new_n43_;
  assign new_n45_ = v11 & v15;
  assign new_n46_ = ~new_n44_ & ~new_n45_;
  assign new_n47_ = ~v13 & ~new_n46_;
  assign new_n48_ = v15 & ~v16;
  assign new_n49_ = v15 & ~new_n48_;
  assign new_n50_ = v13 & ~new_n49_;
  assign new_n51_ = v11 & new_n50_;
  assign new_n52_ = ~new_n47_ & ~new_n51_;
  assign new_n53_ = ~v14 & ~new_n52_;
  assign new_n54_ = v14 & ~v15;
  assign new_n55_ = ~v13 & new_n54_;
  assign new_n56_ = v11 & new_n55_;
  assign new_n57_ = ~new_n53_ & ~new_n56_;
  assign new_n58_ = ~v12 & ~new_n57_;
  assign \v17.0  = ~v0 & new_n58_;
  assign new_n60_ = v13 & ~v14;
  assign new_n61_ = v13 & ~new_n60_;
  assign new_n62_ = v13 & new_n54_;
  assign new_n63_ = new_n61_ & ~new_n62_;
  assign new_n64_ = v13 & v14;
  assign new_n65_ = new_n48_ & new_n64_;
  assign new_n66_ = new_n63_ & ~new_n65_;
  assign new_n67_ = v12 & ~new_n66_;
  assign new_n68_ = v1 & ~v2;
  assign new_n69_ = v4 & ~v5;
  assign new_n70_ = ~v3 & new_n69_;
  assign new_n71_ = new_n68_ & new_n70_;
  assign new_n72_ = ~v12 & ~v13;
  assign new_n73_ = ~v15 & ~v16;
  assign new_n74_ = ~v14 & new_n73_;
  assign new_n75_ = new_n72_ & new_n74_;
  assign new_n76_ = new_n71_ & new_n75_;
  assign new_n77_ = ~new_n67_ & ~new_n76_;
  assign new_n78_ = ~v11 & ~new_n77_;
  assign \v17.1  = ~v0 & new_n78_;
  assign new_n80_ = v12 & v14;
  assign new_n81_ = v15 & v16;
  assign new_n82_ = new_n80_ & new_n81_;
  assign new_n83_ = v1 & v3;
  assign new_n84_ = ~v4 & v6;
  assign new_n85_ = new_n83_ & new_n84_;
  assign new_n86_ = ~v12 & ~v14;
  assign new_n87_ = new_n73_ & new_n86_;
  assign new_n88_ = new_n85_ & new_n87_;
  assign new_n89_ = ~new_n82_ & ~new_n88_;
  assign new_n90_ = ~v13 & ~new_n89_;
  assign new_n91_ = v14 & ~new_n54_;
  assign new_n92_ = v14 & new_n48_;
  assign new_n93_ = new_n91_ & ~new_n92_;
  assign new_n94_ = v13 & ~new_n93_;
  assign new_n95_ = v12 & new_n94_;
  assign new_n96_ = ~new_n90_ & ~new_n95_;
  assign new_n97_ = ~v11 & ~new_n96_;
  assign new_n98_ = ~v14 & ~new_n49_;
  assign new_n99_ = v13 & new_n98_;
  assign new_n100_ = ~v12 & new_n99_;
  assign new_n101_ = v11 & new_n100_;
  assign new_n102_ = ~new_n97_ & ~new_n101_;
  assign \v17.2  = ~v0 & ~new_n102_;
  assign new_n104_ = ~v14 & new_n81_;
  assign new_n105_ = ~new_n54_ & ~new_n104_;
  assign new_n106_ = ~v11 & v12;
  assign new_n107_ = v11 & new_n72_;
  assign new_n108_ = ~new_n106_ & ~new_n107_;
  assign new_n109_ = ~new_n105_ & ~new_n108_;
  assign new_n110_ = v12 & v15;
  assign new_n111_ = ~v7 & v10;
  assign new_n112_ = ~v13 & ~v15;
  assign new_n113_ = ~v12 & new_n112_;
  assign new_n114_ = new_n111_ & new_n113_;
  assign new_n115_ = ~new_n110_ & ~new_n114_;
  assign new_n116_ = ~v16 & ~new_n115_;
  assign new_n117_ = v14 & new_n116_;
  assign new_n118_ = ~v11 & new_n117_;
  assign new_n119_ = ~v12 & v13;
  assign new_n120_ = v11 & new_n119_;
  assign new_n121_ = new_n104_ & new_n120_;
  assign new_n122_ = ~new_n118_ & ~new_n121_;
  assign new_n123_ = ~new_n109_ & new_n122_;
  assign \v17.3  = ~v0 & ~new_n123_;
  assign new_n125_ = ~v15 & v16;
  assign new_n126_ = ~new_n48_ & ~new_n125_;
  assign new_n127_ = v11 & new_n86_;
  assign new_n128_ = ~new_n106_ & ~new_n127_;
  assign new_n129_ = ~new_n126_ & ~new_n128_;
  assign new_n130_ = v11 & v14;
  assign new_n131_ = ~v11 & ~v14;
  assign new_n132_ = ~new_n130_ & ~new_n131_;
  assign new_n133_ = v16 & ~new_n132_;
  assign new_n134_ = ~v15 & new_n133_;
  assign new_n135_ = ~v13 & new_n134_;
  assign new_n136_ = ~v12 & new_n135_;
  assign new_n137_ = ~new_n129_ & ~new_n136_;
  assign \v17.4  = ~v0 & ~new_n137_;
  assign new_n139_ = ~v3 & v4;
  assign new_n140_ = v1 & new_n139_;
  assign new_n141_ = v5 & new_n131_;
  assign new_n142_ = new_n140_ & new_n141_;
  assign new_n143_ = ~new_n130_ & ~new_n142_;
  assign new_n144_ = ~v15 & ~new_n143_;
  assign new_n145_ = ~v13 & new_n144_;
  assign new_n146_ = ~v12 & new_n145_;
  assign new_n147_ = new_n128_ & ~new_n146_;
  assign new_n148_ = ~v16 & ~new_n147_;
  assign \v17.5  = ~v0 & new_n148_;
  assign new_n150_ = v12 & v13;
  assign new_n151_ = v4 & v5;
  assign new_n152_ = v3 & v6;
  assign new_n153_ = ~new_n151_ & ~new_n152_;
  assign new_n154_ = v2 & new_n153_;
  assign new_n155_ = ~v16 & ~new_n154_;
  assign new_n156_ = v1 & new_n155_;
  assign new_n157_ = ~v16 & ~new_n156_;
  assign new_n158_ = ~v12 & ~new_n157_;
  assign new_n159_ = ~v12 & ~new_n158_;
  assign new_n160_ = ~v15 & ~new_n159_;
  assign new_n161_ = ~v12 & ~v16;
  assign new_n162_ = ~v12 & ~new_n161_;
  assign new_n163_ = v15 & ~new_n162_;
  assign new_n164_ = ~new_n160_ & ~new_n163_;
  assign new_n165_ = ~v14 & ~new_n164_;
  assign new_n166_ = ~new_n80_ & ~new_n165_;
  assign new_n167_ = ~v13 & ~new_n166_;
  assign new_n168_ = ~new_n150_ & ~new_n167_;
  assign new_n169_ = ~v11 & ~new_n168_;
  assign new_n170_ = v14 & ~new_n55_;
  assign new_n171_ = ~v13 & v14;
  assign new_n172_ = new_n48_ & new_n171_;
  assign new_n173_ = new_n170_ & ~new_n172_;
  assign new_n174_ = ~v12 & ~new_n173_;
  assign new_n175_ = v11 & new_n174_;
  assign new_n176_ = ~new_n169_ & ~new_n175_;
  assign \v17.6  = ~v0 & ~new_n176_;
  assign new_n178_ = v11 & v13;
  assign new_n179_ = v1 & new_n152_;
  assign new_n180_ = ~v13 & ~v16;
  assign new_n181_ = ~v11 & new_n180_;
  assign new_n182_ = new_n179_ & new_n181_;
  assign new_n183_ = ~new_n178_ & ~new_n182_;
  assign new_n184_ = ~v14 & ~new_n183_;
  assign new_n185_ = ~v11 & ~v13;
  assign new_n186_ = v14 & ~v16;
  assign new_n187_ = new_n185_ & new_n186_;
  assign new_n188_ = ~new_n184_ & ~new_n187_;
  assign new_n189_ = ~v15 & ~new_n188_;
  assign new_n190_ = ~v14 & v15;
  assign new_n191_ = v13 & new_n190_;
  assign new_n192_ = v11 & new_n191_;
  assign new_n193_ = ~new_n189_ & ~new_n192_;
  assign new_n194_ = ~v12 & ~new_n193_;
  assign \v17.7  = ~v0 & new_n194_;
  assign new_n196_ = ~v14 & ~new_n126_;
  assign new_n197_ = ~v13 & new_n196_;
  assign new_n198_ = ~v12 & new_n197_;
  assign new_n199_ = ~v11 & new_n198_;
  assign \v17.8  = v7 & new_n199_;
  assign new_n201_ = ~new_n126_ & ~new_n132_;
  assign new_n202_ = ~v13 & new_n201_;
  assign new_n203_ = ~v12 & new_n202_;
  assign new_n204_ = v14 & new_n73_;
  assign new_n205_ = ~new_n104_ & ~new_n204_;
  assign new_n206_ = v13 & ~new_n205_;
  assign new_n207_ = v12 & new_n206_;
  assign new_n208_ = ~v11 & new_n207_;
  assign new_n209_ = ~new_n203_ & ~new_n208_;
  assign new_n210_ = ~v7 & ~new_n209_;
  assign new_n211_ = v11 & ~v12;
  assign new_n212_ = ~new_n106_ & ~new_n211_;
  assign new_n213_ = ~v15 & ~new_n212_;
  assign new_n214_ = ~v14 & new_n213_;
  assign new_n215_ = ~v13 & new_n214_;
  assign new_n216_ = v7 & new_n215_;
  assign \v17.9  = new_n210_ | new_n216_;
  assign new_n218_ = ~new_n60_ & ~new_n171_;
  assign new_n219_ = ~new_n62_ & new_n218_;
  assign new_n220_ = ~v13 & ~v14;
  assign new_n221_ = new_n81_ & new_n220_;
  assign new_n222_ = new_n219_ & ~new_n221_;
  assign new_n223_ = v12 & ~new_n222_;
  assign \v17.10  = ~v11 & new_n223_;
  assign new_n225_ = ~v13 & new_n81_;
  assign new_n226_ = v13 & new_n73_;
  assign new_n227_ = ~new_n225_ & ~new_n226_;
  assign new_n228_ = v14 & ~new_n227_;
  assign new_n229_ = ~new_n60_ & ~new_n228_;
  assign new_n230_ = v12 & ~new_n229_;
  assign \v17.11  = ~v11 & new_n230_;
  assign new_n232_ = ~new_n54_ & ~new_n190_;
  assign new_n233_ = ~v13 & ~new_n232_;
  assign new_n234_ = ~v12 & new_n233_;
  assign new_n235_ = v11 & new_n234_;
  assign \v17.12  = v7 & new_n235_;
  assign new_n237_ = ~v8 & new_n235_;
  assign \v17.13  = v7 & new_n237_;
  assign new_n239_ = v9 & new_n235_;
  assign \v17.14  = v7 & new_n239_;
  assign new_n241_ = v7 & v11;
  assign new_n242_ = ~v12 & new_n241_;
  assign new_n243_ = v13 & new_n242_;
  assign new_n244_ = ~v14 & new_n243_;
  assign new_n245_ = v15 & new_n244_;
  assign \v17.15  = v16 & new_n245_;
endmodule


