// Benchmark "sin" written by ABC on Tue Sep  5 18:13:10 2023

module sin ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] ;
  wire new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_,
    new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_,
    new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_,
    new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_,
    new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_,
    new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_,
    new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_,
    new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_,
    new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_,
    new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_,
    new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_,
    new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_,
    new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_,
    new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_,
    new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_,
    new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_,
    new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_,
    new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_,
    new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_,
    new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_,
    new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_,
    new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_,
    new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_,
    new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_,
    new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_,
    new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_,
    new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_,
    new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_,
    new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_,
    new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_,
    new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_,
    new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_,
    new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_,
    new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_,
    new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_,
    new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_,
    new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_,
    new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_,
    new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_,
    new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_,
    new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_,
    new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_,
    new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_,
    new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_,
    new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_,
    new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_,
    new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_,
    new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_,
    new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_,
    new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_,
    new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_,
    new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_,
    new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_,
    new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_,
    new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_,
    new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_,
    new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_,
    new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_,
    new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_,
    new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_,
    new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_,
    new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_,
    new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_,
    new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_,
    new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_,
    new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_,
    new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_,
    new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_,
    new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_,
    new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_,
    new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_,
    new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_,
    new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_,
    new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_,
    new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_,
    new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_,
    new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_,
    new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_,
    new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_,
    new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_,
    new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_,
    new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_,
    new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_,
    new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_,
    new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_,
    new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_,
    new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_,
    new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_,
    new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_,
    new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_,
    new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_,
    new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_,
    new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_,
    new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_,
    new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_,
    new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_,
    new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_,
    new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_,
    new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_,
    new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_,
    new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_,
    new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_,
    new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_,
    new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_,
    new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_,
    new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_,
    new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_,
    new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_,
    new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_,
    new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_,
    new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_,
    new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_,
    new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_,
    new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4264_,
    new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_,
    new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_,
    new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_,
    new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_,
    new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_,
    new_n4427_, new_n4428_, new_n4429_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_,
    new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_,
    new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_,
    new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_,
    new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_,
    new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_,
    new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4781_, new_n4782_, new_n4783_, new_n4784_,
    new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_,
    new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_,
    new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_,
    new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_,
    new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_,
    new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_,
    new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_,
    new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_,
    new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_,
    new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_,
    new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_,
    new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_,
    new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_,
    new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_,
    new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_,
    new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_,
    new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_,
    new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_,
    new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_,
    new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_,
    new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_,
    new_n5081_, new_n5082_, new_n5083_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5274_, new_n5275_, new_n5276_,
    new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_,
    new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_,
    new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_,
    new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_,
    new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_,
    new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_,
    new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_,
    new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_,
    new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_,
    new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_,
    new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_,
    new_n5343_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_,
    new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5656_,
    new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_,
    new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_,
    new_n5669_, new_n5670_, new_n5671_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5738_,
    new_n5739_, new_n5740_, new_n5741_;
  INV_X1     g0000(.I(\a[4] ), .ZN(new_n50_));
  NOR4_X1    g0001(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[2] ), .A4(\a[3] ), .ZN(new_n51_));
  OR4_X2     g0002(.A1(\a[0] ), .A2(\a[1] ), .A3(\a[2] ), .A4(\a[3] ), .Z(new_n52_));
  NOR2_X1    g0003(.A1(new_n52_), .A2(\a[22] ), .ZN(new_n53_));
  INV_X1     g0004(.I(new_n53_), .ZN(new_n54_));
  NOR2_X1    g0005(.A1(new_n50_), .A2(\a[22] ), .ZN(new_n55_));
  AOI22_X1   g0006(.A1(new_n54_), .A2(new_n50_), .B1(new_n51_), .B2(new_n55_), .ZN(new_n56_));
  NOR2_X1    g0007(.A1(new_n51_), .A2(\a[4] ), .ZN(new_n57_));
  NOR2_X1    g0008(.A1(new_n57_), .A2(\a[22] ), .ZN(new_n58_));
  NOR2_X1    g0009(.A1(new_n58_), .A2(\a[5] ), .ZN(new_n59_));
  INV_X1     g0010(.I(\a[5] ), .ZN(new_n60_));
  NOR3_X1    g0011(.A1(new_n57_), .A2(new_n60_), .A3(\a[22] ), .ZN(new_n61_));
  NOR2_X1    g0012(.A1(new_n59_), .A2(new_n61_), .ZN(new_n62_));
  XNOR2_X1   g0013(.A1(new_n62_), .A2(new_n56_), .ZN(new_n63_));
  INV_X1     g0014(.I(\a[2] ), .ZN(new_n64_));
  NOR2_X1    g0015(.A1(\a[0] ), .A2(\a[1] ), .ZN(new_n65_));
  AOI21_X1   g0016(.A1(new_n65_), .A2(new_n64_), .B(\a[22] ), .ZN(new_n66_));
  XOR2_X1    g0017(.A1(new_n66_), .A2(\a[3] ), .Z(new_n67_));
  NOR2_X1    g0018(.A1(new_n65_), .A2(\a[22] ), .ZN(new_n68_));
  XOR2_X1    g0019(.A1(new_n68_), .A2(new_n64_), .Z(new_n69_));
  XNOR2_X1   g0020(.A1(new_n67_), .A2(new_n69_), .ZN(new_n70_));
  NOR2_X1    g0021(.A1(new_n63_), .A2(new_n70_), .ZN(new_n71_));
  INV_X1     g0022(.I(new_n71_), .ZN(new_n72_));
  INV_X1     g0023(.I(\a[15] ), .ZN(new_n73_));
  OR3_X2     g0024(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .Z(new_n74_));
  OR3_X2     g0025(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[9] ), .Z(new_n75_));
  OR3_X2     g0026(.A1(\a[10] ), .A2(\a[11] ), .A3(\a[12] ), .Z(new_n76_));
  NOR4_X1    g0027(.A1(new_n74_), .A2(new_n75_), .A3(new_n76_), .A4(new_n51_), .ZN(new_n77_));
  NOR2_X1    g0028(.A1(\a[13] ), .A2(\a[14] ), .ZN(new_n78_));
  NAND2_X1   g0029(.A1(new_n77_), .A2(new_n78_), .ZN(new_n79_));
  INV_X1     g0030(.I(\a[22] ), .ZN(new_n80_));
  NOR3_X1    g0031(.A1(\a[4] ), .A2(\a[5] ), .A3(\a[6] ), .ZN(new_n81_));
  NOR3_X1    g0032(.A1(\a[7] ), .A2(\a[8] ), .A3(\a[9] ), .ZN(new_n82_));
  NOR3_X1    g0033(.A1(\a[10] ), .A2(\a[11] ), .A3(\a[12] ), .ZN(new_n83_));
  NAND4_X1   g0034(.A1(new_n52_), .A2(new_n81_), .A3(new_n82_), .A4(new_n83_), .ZN(new_n84_));
  INV_X1     g0035(.I(new_n78_), .ZN(new_n85_));
  OAI21_X1   g0036(.A1(new_n84_), .A2(new_n85_), .B(new_n80_), .ZN(new_n86_));
  NOR2_X1    g0037(.A1(new_n73_), .A2(\a[22] ), .ZN(new_n87_));
  AOI22_X1   g0038(.A1(new_n86_), .A2(new_n73_), .B1(new_n79_), .B2(new_n87_), .ZN(new_n88_));
  NOR3_X1    g0039(.A1(\a[15] ), .A2(\a[16] ), .A3(\a[17] ), .ZN(new_n89_));
  NOR2_X1    g0040(.A1(\a[18] ), .A2(\a[19] ), .ZN(new_n90_));
  NAND4_X1   g0041(.A1(new_n77_), .A2(new_n78_), .A3(new_n89_), .A4(new_n90_), .ZN(new_n91_));
  AOI21_X1   g0042(.A1(new_n91_), .A2(new_n80_), .B(\a[20] ), .ZN(new_n92_));
  INV_X1     g0043(.I(\a[20] ), .ZN(new_n93_));
  INV_X1     g0044(.I(new_n89_), .ZN(new_n94_));
  INV_X1     g0045(.I(new_n90_), .ZN(new_n95_));
  NOR4_X1    g0046(.A1(new_n84_), .A2(new_n85_), .A3(new_n94_), .A4(new_n95_), .ZN(new_n96_));
  NOR3_X1    g0047(.A1(new_n96_), .A2(new_n93_), .A3(\a[22] ), .ZN(new_n97_));
  NOR2_X1    g0048(.A1(new_n97_), .A2(new_n92_), .ZN(new_n98_));
  NAND2_X1   g0049(.A1(new_n90_), .A2(new_n93_), .ZN(new_n99_));
  INV_X1     g0050(.I(new_n99_), .ZN(new_n100_));
  NAND4_X1   g0051(.A1(new_n77_), .A2(new_n78_), .A3(new_n89_), .A4(new_n100_), .ZN(new_n101_));
  AOI21_X1   g0052(.A1(new_n101_), .A2(new_n80_), .B(\a[21] ), .ZN(new_n102_));
  NOR4_X1    g0053(.A1(new_n84_), .A2(new_n85_), .A3(new_n94_), .A4(new_n99_), .ZN(new_n103_));
  INV_X1     g0054(.I(\a[21] ), .ZN(new_n104_));
  NOR2_X1    g0055(.A1(new_n104_), .A2(\a[22] ), .ZN(new_n105_));
  INV_X1     g0056(.I(new_n105_), .ZN(new_n106_));
  NOR2_X1    g0057(.A1(new_n103_), .A2(new_n106_), .ZN(new_n107_));
  NOR2_X1    g0058(.A1(new_n102_), .A2(new_n107_), .ZN(new_n108_));
  NOR3_X1    g0059(.A1(new_n98_), .A2(new_n108_), .A3(new_n88_), .ZN(new_n109_));
  NOR3_X1    g0060(.A1(new_n74_), .A2(new_n75_), .A3(new_n51_), .ZN(new_n110_));
  NAND4_X1   g0061(.A1(new_n110_), .A2(new_n73_), .A3(new_n83_), .A4(new_n78_), .ZN(new_n111_));
  AOI21_X1   g0062(.A1(new_n111_), .A2(new_n80_), .B(\a[16] ), .ZN(new_n112_));
  INV_X1     g0063(.I(\a[16] ), .ZN(new_n113_));
  NOR3_X1    g0064(.A1(new_n84_), .A2(\a[15] ), .A3(new_n85_), .ZN(new_n114_));
  NOR3_X1    g0065(.A1(new_n114_), .A2(new_n113_), .A3(\a[22] ), .ZN(new_n115_));
  AOI21_X1   g0066(.A1(new_n111_), .A2(new_n80_), .B(\a[17] ), .ZN(new_n116_));
  INV_X1     g0067(.I(\a[17] ), .ZN(new_n117_));
  NOR3_X1    g0068(.A1(new_n114_), .A2(new_n117_), .A3(\a[22] ), .ZN(new_n118_));
  OAI22_X1   g0069(.A1(new_n112_), .A2(new_n115_), .B1(new_n118_), .B2(new_n116_), .ZN(new_n119_));
  INV_X1     g0070(.I(\a[18] ), .ZN(new_n120_));
  NOR3_X1    g0071(.A1(new_n84_), .A2(new_n85_), .A3(new_n94_), .ZN(new_n121_));
  OAI21_X1   g0072(.A1(new_n121_), .A2(\a[22] ), .B(new_n120_), .ZN(new_n122_));
  NAND4_X1   g0073(.A1(new_n110_), .A2(new_n83_), .A3(new_n78_), .A4(new_n89_), .ZN(new_n123_));
  NAND3_X1   g0074(.A1(new_n123_), .A2(\a[18] ), .A3(new_n80_), .ZN(new_n124_));
  NAND2_X1   g0075(.A1(new_n122_), .A2(new_n124_), .ZN(new_n125_));
  AOI21_X1   g0076(.A1(new_n123_), .A2(new_n80_), .B(\a[19] ), .ZN(new_n126_));
  INV_X1     g0077(.I(\a[19] ), .ZN(new_n127_));
  NOR3_X1    g0078(.A1(new_n121_), .A2(new_n127_), .A3(\a[22] ), .ZN(new_n128_));
  NOR2_X1    g0079(.A1(new_n128_), .A2(new_n126_), .ZN(new_n129_));
  NOR3_X1    g0080(.A1(new_n119_), .A2(new_n125_), .A3(new_n129_), .ZN(new_n130_));
  NAND2_X1   g0081(.A1(new_n130_), .A2(new_n109_), .ZN(new_n131_));
  OAI21_X1   g0082(.A1(new_n114_), .A2(\a[22] ), .B(new_n113_), .ZN(new_n132_));
  NAND3_X1   g0083(.A1(new_n111_), .A2(\a[16] ), .A3(new_n80_), .ZN(new_n133_));
  NAND2_X1   g0084(.A1(new_n132_), .A2(new_n133_), .ZN(new_n134_));
  NOR2_X1    g0085(.A1(new_n118_), .A2(new_n116_), .ZN(new_n135_));
  NOR3_X1    g0086(.A1(new_n121_), .A2(new_n120_), .A3(\a[19] ), .ZN(new_n136_));
  AOI21_X1   g0087(.A1(new_n123_), .A2(new_n127_), .B(\a[18] ), .ZN(new_n137_));
  XNOR2_X1   g0088(.A1(\a[19] ), .A2(\a[22] ), .ZN(new_n138_));
  INV_X1     g0089(.I(new_n138_), .ZN(new_n139_));
  NOR3_X1    g0090(.A1(new_n136_), .A2(new_n137_), .A3(new_n139_), .ZN(new_n140_));
  NOR3_X1    g0091(.A1(new_n140_), .A2(new_n135_), .A3(new_n134_), .ZN(new_n141_));
  OAI21_X1   g0092(.A1(new_n103_), .A2(\a[22] ), .B(new_n104_), .ZN(new_n142_));
  NAND2_X1   g0093(.A1(new_n101_), .A2(new_n105_), .ZN(new_n143_));
  NAND2_X1   g0094(.A1(new_n142_), .A2(new_n143_), .ZN(new_n144_));
  NOR3_X1    g0095(.A1(new_n98_), .A2(new_n144_), .A3(new_n88_), .ZN(new_n145_));
  NAND2_X1   g0096(.A1(new_n145_), .A2(new_n141_), .ZN(new_n146_));
  NOR2_X1    g0097(.A1(new_n84_), .A2(new_n85_), .ZN(new_n147_));
  AOI21_X1   g0098(.A1(new_n77_), .A2(new_n78_), .B(\a[22] ), .ZN(new_n148_));
  INV_X1     g0099(.I(new_n87_), .ZN(new_n149_));
  OAI22_X1   g0100(.A1(new_n148_), .A2(\a[15] ), .B1(new_n147_), .B2(new_n149_), .ZN(new_n150_));
  NOR3_X1    g0101(.A1(new_n98_), .A2(new_n144_), .A3(new_n150_), .ZN(new_n151_));
  NOR4_X1    g0102(.A1(new_n134_), .A2(new_n135_), .A3(new_n129_), .A4(new_n125_), .ZN(new_n152_));
  NAND2_X1   g0103(.A1(new_n152_), .A2(new_n151_), .ZN(new_n153_));
  NAND3_X1   g0104(.A1(new_n131_), .A2(new_n153_), .A3(new_n146_), .ZN(new_n154_));
  NOR2_X1    g0105(.A1(new_n115_), .A2(new_n112_), .ZN(new_n155_));
  OAI21_X1   g0106(.A1(new_n114_), .A2(\a[22] ), .B(new_n117_), .ZN(new_n156_));
  NAND3_X1   g0107(.A1(new_n111_), .A2(\a[17] ), .A3(new_n80_), .ZN(new_n157_));
  NAND2_X1   g0108(.A1(new_n156_), .A2(new_n157_), .ZN(new_n158_));
  AOI21_X1   g0109(.A1(new_n123_), .A2(new_n80_), .B(\a[18] ), .ZN(new_n159_));
  NOR3_X1    g0110(.A1(new_n121_), .A2(new_n120_), .A3(\a[22] ), .ZN(new_n160_));
  NOR2_X1    g0111(.A1(new_n160_), .A2(new_n159_), .ZN(new_n161_));
  OAI21_X1   g0112(.A1(new_n121_), .A2(\a[22] ), .B(new_n127_), .ZN(new_n162_));
  NAND3_X1   g0113(.A1(new_n123_), .A2(\a[19] ), .A3(new_n80_), .ZN(new_n163_));
  NAND2_X1   g0114(.A1(new_n162_), .A2(new_n163_), .ZN(new_n164_));
  NAND4_X1   g0115(.A1(new_n155_), .A2(new_n158_), .A3(new_n161_), .A4(new_n164_), .ZN(new_n165_));
  OAI21_X1   g0116(.A1(new_n96_), .A2(\a[22] ), .B(new_n93_), .ZN(new_n166_));
  NAND2_X1   g0117(.A1(new_n104_), .A2(\a[22] ), .ZN(new_n167_));
  NAND2_X1   g0118(.A1(new_n106_), .A2(new_n167_), .ZN(new_n168_));
  NAND3_X1   g0119(.A1(new_n91_), .A2(\a[20] ), .A3(new_n80_), .ZN(new_n169_));
  AOI21_X1   g0120(.A1(new_n166_), .A2(new_n169_), .B(new_n168_), .ZN(new_n170_));
  NAND2_X1   g0121(.A1(new_n170_), .A2(new_n150_), .ZN(new_n171_));
  NOR2_X1    g0122(.A1(new_n165_), .A2(new_n171_), .ZN(new_n172_));
  NAND3_X1   g0123(.A1(new_n91_), .A2(\a[20] ), .A3(new_n80_), .ZN(new_n173_));
  AOI21_X1   g0124(.A1(new_n166_), .A2(new_n173_), .B(new_n150_), .ZN(new_n174_));
  NAND2_X1   g0125(.A1(new_n174_), .A2(new_n108_), .ZN(new_n175_));
  XNOR2_X1   g0126(.A1(\a[17] ), .A2(\a[22] ), .ZN(new_n176_));
  INV_X1     g0127(.I(new_n176_), .ZN(new_n177_));
  AOI21_X1   g0128(.A1(new_n132_), .A2(new_n133_), .B(new_n177_), .ZN(new_n178_));
  AOI21_X1   g0129(.A1(new_n122_), .A2(new_n124_), .B(new_n139_), .ZN(new_n179_));
  NAND2_X1   g0130(.A1(new_n178_), .A2(new_n179_), .ZN(new_n180_));
  NOR2_X1    g0131(.A1(new_n175_), .A2(new_n180_), .ZN(new_n181_));
  NOR3_X1    g0132(.A1(new_n154_), .A2(new_n172_), .A3(new_n181_), .ZN(new_n182_));
  INV_X1     g0133(.I(new_n182_), .ZN(new_n183_));
  INV_X1     g0134(.I(new_n168_), .ZN(new_n184_));
  NAND3_X1   g0135(.A1(new_n91_), .A2(\a[20] ), .A3(new_n104_), .ZN(new_n185_));
  OAI21_X1   g0136(.A1(new_n96_), .A2(\a[21] ), .B(new_n93_), .ZN(new_n186_));
  NAND3_X1   g0137(.A1(new_n186_), .A2(new_n185_), .A3(new_n184_), .ZN(new_n187_));
  NAND2_X1   g0138(.A1(new_n187_), .A2(new_n88_), .ZN(new_n188_));
  NOR2_X1    g0139(.A1(new_n165_), .A2(new_n188_), .ZN(new_n189_));
  NAND2_X1   g0140(.A1(new_n166_), .A2(new_n173_), .ZN(new_n190_));
  NAND3_X1   g0141(.A1(new_n190_), .A2(new_n144_), .A3(new_n150_), .ZN(new_n191_));
  NOR2_X1    g0142(.A1(new_n165_), .A2(new_n191_), .ZN(new_n192_));
  NOR2_X1    g0143(.A1(new_n189_), .A2(new_n192_), .ZN(new_n193_));
  INV_X1     g0144(.I(new_n193_), .ZN(new_n194_));
  NAND3_X1   g0145(.A1(new_n190_), .A2(new_n108_), .A3(new_n150_), .ZN(new_n195_));
  AOI22_X1   g0146(.A1(new_n122_), .A2(new_n124_), .B1(new_n162_), .B2(new_n163_), .ZN(new_n196_));
  NAND3_X1   g0147(.A1(new_n196_), .A2(new_n155_), .A3(new_n158_), .ZN(new_n197_));
  NOR2_X1    g0148(.A1(new_n197_), .A2(new_n195_), .ZN(new_n198_));
  NOR3_X1    g0149(.A1(new_n114_), .A2(new_n113_), .A3(\a[17] ), .ZN(new_n199_));
  AOI21_X1   g0150(.A1(new_n111_), .A2(new_n117_), .B(\a[16] ), .ZN(new_n200_));
  NOR3_X1    g0151(.A1(new_n199_), .A2(new_n200_), .A3(new_n177_), .ZN(new_n201_));
  NOR2_X1    g0152(.A1(new_n140_), .A2(new_n201_), .ZN(new_n202_));
  NAND2_X1   g0153(.A1(new_n109_), .A2(new_n202_), .ZN(new_n203_));
  INV_X1     g0154(.I(new_n203_), .ZN(new_n204_));
  NAND3_X1   g0155(.A1(new_n123_), .A2(\a[18] ), .A3(new_n127_), .ZN(new_n205_));
  OAI21_X1   g0156(.A1(new_n121_), .A2(\a[19] ), .B(new_n120_), .ZN(new_n206_));
  NAND3_X1   g0157(.A1(new_n206_), .A2(new_n205_), .A3(new_n138_), .ZN(new_n207_));
  NAND3_X1   g0158(.A1(new_n155_), .A2(new_n207_), .A3(new_n158_), .ZN(new_n208_));
  NOR2_X1    g0159(.A1(new_n191_), .A2(new_n208_), .ZN(new_n209_));
  AOI22_X1   g0160(.A1(new_n132_), .A2(new_n133_), .B1(new_n156_), .B2(new_n157_), .ZN(new_n210_));
  NAND4_X1   g0161(.A1(new_n174_), .A2(new_n210_), .A3(new_n144_), .A4(new_n179_), .ZN(new_n211_));
  INV_X1     g0162(.I(new_n211_), .ZN(new_n212_));
  NOR2_X1    g0163(.A1(new_n212_), .A2(new_n209_), .ZN(new_n213_));
  INV_X1     g0164(.I(new_n213_), .ZN(new_n214_));
  NOR4_X1    g0165(.A1(new_n194_), .A2(new_n214_), .A3(new_n198_), .A4(new_n204_), .ZN(new_n215_));
  INV_X1     g0166(.I(new_n215_), .ZN(new_n216_));
  OAI21_X1   g0167(.A1(new_n115_), .A2(new_n112_), .B(new_n176_), .ZN(new_n217_));
  OAI21_X1   g0168(.A1(new_n160_), .A2(new_n159_), .B(new_n138_), .ZN(new_n218_));
  NOR2_X1    g0169(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR3_X1    g0170(.A1(new_n96_), .A2(new_n93_), .A3(\a[22] ), .ZN(new_n220_));
  OAI21_X1   g0171(.A1(new_n220_), .A2(new_n92_), .B(new_n184_), .ZN(new_n221_));
  NOR2_X1    g0172(.A1(new_n221_), .A2(new_n150_), .ZN(new_n222_));
  NAND2_X1   g0173(.A1(new_n222_), .A2(new_n219_), .ZN(new_n223_));
  NOR2_X1    g0174(.A1(new_n221_), .A2(new_n88_), .ZN(new_n224_));
  OAI22_X1   g0175(.A1(new_n159_), .A2(new_n160_), .B1(new_n128_), .B2(new_n126_), .ZN(new_n225_));
  NOR3_X1    g0176(.A1(new_n225_), .A2(new_n134_), .A3(new_n135_), .ZN(new_n226_));
  NOR2_X1    g0177(.A1(new_n119_), .A2(new_n218_), .ZN(new_n227_));
  OAI21_X1   g0178(.A1(new_n226_), .A2(new_n227_), .B(new_n224_), .ZN(new_n228_));
  NAND3_X1   g0179(.A1(new_n111_), .A2(\a[16] ), .A3(new_n117_), .ZN(new_n229_));
  OAI21_X1   g0180(.A1(new_n114_), .A2(\a[17] ), .B(new_n113_), .ZN(new_n230_));
  NAND3_X1   g0181(.A1(new_n230_), .A2(new_n229_), .A3(new_n176_), .ZN(new_n231_));
  NAND4_X1   g0182(.A1(new_n174_), .A2(new_n196_), .A3(new_n108_), .A4(new_n231_), .ZN(new_n232_));
  NOR2_X1    g0183(.A1(new_n218_), .A2(new_n201_), .ZN(new_n233_));
  NOR2_X1    g0184(.A1(new_n119_), .A2(new_n225_), .ZN(new_n234_));
  OAI21_X1   g0185(.A1(new_n234_), .A2(new_n233_), .B(new_n224_), .ZN(new_n235_));
  NAND4_X1   g0186(.A1(new_n228_), .A2(new_n235_), .A3(new_n223_), .A4(new_n232_), .ZN(new_n236_));
  NAND2_X1   g0187(.A1(new_n170_), .A2(new_n88_), .ZN(new_n237_));
  NOR2_X1    g0188(.A1(new_n237_), .A2(new_n208_), .ZN(new_n238_));
  NOR2_X1    g0189(.A1(new_n175_), .A2(new_n208_), .ZN(new_n239_));
  NAND2_X1   g0190(.A1(new_n174_), .A2(new_n144_), .ZN(new_n240_));
  NAND3_X1   g0191(.A1(new_n178_), .A2(new_n161_), .A3(new_n164_), .ZN(new_n241_));
  NOR2_X1    g0192(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NOR3_X1    g0193(.A1(new_n88_), .A2(new_n102_), .A3(new_n107_), .ZN(new_n243_));
  NAND2_X1   g0194(.A1(new_n243_), .A2(new_n190_), .ZN(new_n244_));
  NAND3_X1   g0195(.A1(new_n161_), .A2(new_n231_), .A3(new_n164_), .ZN(new_n245_));
  NOR2_X1    g0196(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR4_X1    g0197(.A1(new_n238_), .A2(new_n239_), .A3(new_n242_), .A4(new_n246_), .ZN(new_n247_));
  NOR4_X1    g0198(.A1(new_n216_), .A2(new_n183_), .A3(new_n236_), .A4(new_n247_), .ZN(new_n248_));
  INV_X1     g0199(.I(new_n248_), .ZN(new_n249_));
  NOR2_X1    g0200(.A1(new_n165_), .A2(new_n195_), .ZN(new_n250_));
  NOR3_X1    g0201(.A1(new_n98_), .A2(new_n108_), .A3(new_n150_), .ZN(new_n251_));
  NAND2_X1   g0202(.A1(new_n251_), .A2(new_n233_), .ZN(new_n252_));
  NAND2_X1   g0203(.A1(new_n91_), .A2(new_n104_), .ZN(new_n253_));
  AOI21_X1   g0204(.A1(new_n253_), .A2(new_n93_), .B(new_n168_), .ZN(new_n254_));
  AOI21_X1   g0205(.A1(new_n254_), .A2(new_n185_), .B(new_n150_), .ZN(new_n255_));
  NAND2_X1   g0206(.A1(new_n141_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1   g0207(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  NOR3_X1    g0208(.A1(new_n249_), .A2(new_n250_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1     g0209(.I(new_n258_), .ZN(new_n259_));
  OAI22_X1   g0210(.A1(new_n92_), .A2(new_n97_), .B1(new_n102_), .B2(new_n107_), .ZN(new_n260_));
  NOR4_X1    g0211(.A1(new_n260_), .A2(new_n225_), .A3(new_n88_), .A4(new_n217_), .ZN(new_n261_));
  NAND2_X1   g0212(.A1(new_n161_), .A2(new_n164_), .ZN(new_n262_));
  NOR3_X1    g0213(.A1(new_n244_), .A2(new_n119_), .A3(new_n262_), .ZN(new_n263_));
  NOR2_X1    g0214(.A1(new_n263_), .A2(new_n261_), .ZN(new_n264_));
  NAND2_X1   g0215(.A1(new_n187_), .A2(new_n150_), .ZN(new_n265_));
  NOR2_X1    g0216(.A1(new_n265_), .A2(new_n180_), .ZN(new_n266_));
  NOR2_X1    g0217(.A1(new_n241_), .A2(new_n188_), .ZN(new_n267_));
  NOR2_X1    g0218(.A1(new_n267_), .A2(new_n266_), .ZN(new_n268_));
  NAND2_X1   g0219(.A1(new_n210_), .A2(new_n196_), .ZN(new_n269_));
  NAND3_X1   g0220(.A1(new_n190_), .A2(new_n108_), .A3(new_n88_), .ZN(new_n270_));
  OAI22_X1   g0221(.A1(new_n269_), .A2(new_n191_), .B1(new_n270_), .B2(new_n241_), .ZN(new_n271_));
  NOR2_X1    g0222(.A1(new_n165_), .A2(new_n265_), .ZN(new_n272_));
  OAI21_X1   g0223(.A1(new_n92_), .A2(new_n97_), .B(new_n88_), .ZN(new_n273_));
  NOR4_X1    g0224(.A1(new_n119_), .A2(new_n273_), .A3(new_n225_), .A4(new_n108_), .ZN(new_n274_));
  NOR2_X1    g0225(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1     g0226(.I(new_n275_), .ZN(new_n276_));
  NAND2_X1   g0227(.A1(new_n207_), .A2(new_n231_), .ZN(new_n277_));
  NOR2_X1    g0228(.A1(new_n171_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1   g0229(.A1(new_n179_), .A2(new_n155_), .A3(new_n158_), .ZN(new_n279_));
  NOR2_X1    g0230(.A1(new_n244_), .A2(new_n279_), .ZN(new_n280_));
  NOR2_X1    g0231(.A1(new_n280_), .A2(new_n278_), .ZN(new_n281_));
  INV_X1     g0232(.I(new_n281_), .ZN(new_n282_));
  NOR2_X1    g0233(.A1(new_n119_), .A2(new_n140_), .ZN(new_n283_));
  NAND2_X1   g0234(.A1(new_n283_), .A2(new_n251_), .ZN(new_n284_));
  NOR2_X1    g0235(.A1(new_n225_), .A2(new_n201_), .ZN(new_n285_));
  NAND3_X1   g0236(.A1(new_n150_), .A2(new_n142_), .A3(new_n143_), .ZN(new_n286_));
  NOR2_X1    g0237(.A1(new_n286_), .A2(new_n98_), .ZN(new_n287_));
  NAND2_X1   g0238(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1   g0239(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  NOR4_X1    g0240(.A1(new_n276_), .A2(new_n282_), .A3(new_n271_), .A4(new_n289_), .ZN(new_n290_));
  NAND4_X1   g0241(.A1(new_n196_), .A2(new_n170_), .A3(new_n150_), .A4(new_n178_), .ZN(new_n291_));
  NAND3_X1   g0242(.A1(new_n210_), .A2(new_n161_), .A3(new_n164_), .ZN(new_n292_));
  NOR2_X1    g0243(.A1(new_n292_), .A2(new_n175_), .ZN(new_n293_));
  INV_X1     g0244(.I(new_n293_), .ZN(new_n294_));
  AOI21_X1   g0245(.A1(new_n254_), .A2(new_n185_), .B(new_n88_), .ZN(new_n295_));
  NAND2_X1   g0246(.A1(new_n285_), .A2(new_n295_), .ZN(new_n296_));
  NOR3_X1    g0247(.A1(new_n96_), .A2(new_n93_), .A3(\a[21] ), .ZN(new_n297_));
  AOI21_X1   g0248(.A1(new_n91_), .A2(new_n104_), .B(\a[20] ), .ZN(new_n298_));
  NOR3_X1    g0249(.A1(new_n297_), .A2(new_n298_), .A3(new_n168_), .ZN(new_n299_));
  NOR4_X1    g0250(.A1(new_n119_), .A2(new_n299_), .A3(new_n150_), .A4(new_n140_), .ZN(new_n300_));
  NOR2_X1    g0251(.A1(new_n292_), .A2(new_n265_), .ZN(new_n301_));
  NOR2_X1    g0252(.A1(new_n301_), .A2(new_n300_), .ZN(new_n302_));
  NAND4_X1   g0253(.A1(new_n302_), .A2(new_n294_), .A3(new_n291_), .A4(new_n296_), .ZN(new_n303_));
  NAND2_X1   g0254(.A1(new_n226_), .A2(new_n295_), .ZN(new_n304_));
  INV_X1     g0255(.I(new_n304_), .ZN(new_n305_));
  NOR2_X1    g0256(.A1(new_n175_), .A2(new_n277_), .ZN(new_n306_));
  NOR2_X1    g0257(.A1(new_n244_), .A2(new_n180_), .ZN(new_n307_));
  NOR3_X1    g0258(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1   g0259(.A1(new_n109_), .A2(new_n219_), .ZN(new_n309_));
  NAND3_X1   g0260(.A1(new_n233_), .A2(new_n190_), .A3(new_n243_), .ZN(new_n310_));
  NOR2_X1    g0261(.A1(new_n191_), .A2(new_n245_), .ZN(new_n311_));
  INV_X1     g0262(.I(new_n311_), .ZN(new_n312_));
  NAND4_X1   g0263(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .A4(new_n312_), .ZN(new_n313_));
  NOR2_X1    g0264(.A1(new_n313_), .A2(new_n303_), .ZN(new_n314_));
  NAND4_X1   g0265(.A1(new_n314_), .A2(new_n264_), .A3(new_n268_), .A4(new_n290_), .ZN(new_n315_));
  NAND2_X1   g0266(.A1(new_n141_), .A2(new_n295_), .ZN(new_n316_));
  NAND3_X1   g0267(.A1(new_n226_), .A2(new_n88_), .A3(new_n187_), .ZN(new_n317_));
  NOR3_X1    g0268(.A1(new_n218_), .A2(new_n135_), .A3(new_n134_), .ZN(new_n318_));
  NAND2_X1   g0269(.A1(new_n151_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1   g0270(.A1(new_n317_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  NAND4_X1   g0271(.A1(new_n187_), .A2(new_n178_), .A3(new_n179_), .A4(new_n88_), .ZN(new_n321_));
  INV_X1     g0272(.I(new_n321_), .ZN(new_n322_));
  NAND3_X1   g0273(.A1(new_n207_), .A2(new_n231_), .A3(new_n88_), .ZN(new_n323_));
  NOR2_X1    g0274(.A1(new_n323_), .A2(new_n221_), .ZN(new_n324_));
  NAND4_X1   g0275(.A1(new_n174_), .A2(new_n108_), .A3(new_n179_), .A4(new_n231_), .ZN(new_n325_));
  INV_X1     g0276(.I(new_n325_), .ZN(new_n326_));
  NOR4_X1    g0277(.A1(new_n286_), .A2(new_n98_), .A3(new_n140_), .A4(new_n201_), .ZN(new_n327_));
  NOR4_X1    g0278(.A1(new_n326_), .A2(new_n322_), .A3(new_n324_), .A4(new_n327_), .ZN(new_n328_));
  NAND2_X1   g0279(.A1(new_n130_), .A2(new_n224_), .ZN(new_n329_));
  NAND2_X1   g0280(.A1(new_n285_), .A2(new_n224_), .ZN(new_n330_));
  NAND2_X1   g0281(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR3_X1    g0282(.A1(new_n328_), .A2(new_n320_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1     g0283(.I(new_n332_), .ZN(new_n333_));
  NAND2_X1   g0284(.A1(new_n210_), .A2(new_n207_), .ZN(new_n334_));
  NOR2_X1    g0285(.A1(new_n334_), .A2(new_n237_), .ZN(new_n335_));
  NOR2_X1    g0286(.A1(new_n244_), .A2(new_n241_), .ZN(new_n336_));
  NAND3_X1   g0287(.A1(new_n190_), .A2(new_n144_), .A3(new_n88_), .ZN(new_n337_));
  NOR2_X1    g0288(.A1(new_n337_), .A2(new_n245_), .ZN(new_n338_));
  NOR2_X1    g0289(.A1(new_n292_), .A2(new_n237_), .ZN(new_n339_));
  NOR4_X1    g0290(.A1(new_n335_), .A2(new_n339_), .A3(new_n336_), .A4(new_n338_), .ZN(new_n340_));
  NAND4_X1   g0291(.A1(new_n187_), .A2(new_n179_), .A3(new_n231_), .A4(new_n88_), .ZN(new_n341_));
  NAND4_X1   g0292(.A1(new_n210_), .A2(new_n243_), .A3(new_n190_), .A4(new_n179_), .ZN(new_n342_));
  NAND4_X1   g0293(.A1(new_n174_), .A2(new_n210_), .A3(new_n108_), .A4(new_n179_), .ZN(new_n343_));
  NAND4_X1   g0294(.A1(new_n210_), .A2(new_n187_), .A3(new_n150_), .A4(new_n207_), .ZN(new_n344_));
  NAND4_X1   g0295(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .A4(new_n341_), .ZN(new_n345_));
  NAND3_X1   g0296(.A1(new_n210_), .A2(new_n150_), .A3(new_n207_), .ZN(new_n346_));
  NAND3_X1   g0297(.A1(new_n158_), .A2(new_n132_), .A3(new_n133_), .ZN(new_n347_));
  OAI21_X1   g0298(.A1(new_n347_), .A2(new_n218_), .B(new_n150_), .ZN(new_n348_));
  AOI21_X1   g0299(.A1(new_n348_), .A2(new_n346_), .B(new_n221_), .ZN(new_n349_));
  AOI22_X1   g0300(.A1(new_n226_), .A2(new_n151_), .B1(new_n251_), .B2(new_n219_), .ZN(new_n350_));
  NAND3_X1   g0301(.A1(new_n345_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1    g0302(.A1(new_n351_), .A2(new_n340_), .ZN(new_n352_));
  INV_X1     g0303(.I(new_n352_), .ZN(new_n353_));
  NOR4_X1    g0304(.A1(new_n259_), .A2(new_n315_), .A3(new_n333_), .A4(new_n353_), .ZN(new_n354_));
  INV_X1     g0305(.I(new_n354_), .ZN(new_n355_));
  NAND2_X1   g0306(.A1(new_n283_), .A2(new_n224_), .ZN(new_n356_));
  NAND2_X1   g0307(.A1(new_n234_), .A2(new_n287_), .ZN(new_n357_));
  NAND3_X1   g0308(.A1(new_n357_), .A2(new_n356_), .A3(new_n232_), .ZN(new_n358_));
  INV_X1     g0309(.I(new_n198_), .ZN(new_n359_));
  NOR4_X1    g0310(.A1(new_n347_), .A2(new_n144_), .A3(new_n273_), .A4(new_n225_), .ZN(new_n360_));
  NOR4_X1    g0311(.A1(new_n273_), .A2(new_n225_), .A3(new_n144_), .A4(new_n217_), .ZN(new_n361_));
  NOR2_X1    g0312(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1   g0313(.A1(new_n210_), .A2(new_n174_), .A3(new_n196_), .A4(new_n108_), .ZN(new_n363_));
  NAND4_X1   g0314(.A1(new_n281_), .A2(new_n359_), .A3(new_n362_), .A4(new_n363_), .ZN(new_n364_));
  NOR2_X1    g0315(.A1(new_n364_), .A2(new_n358_), .ZN(new_n365_));
  NOR3_X1    g0316(.A1(new_n119_), .A2(new_n150_), .A3(new_n140_), .ZN(new_n366_));
  NOR2_X1    g0317(.A1(new_n217_), .A2(new_n140_), .ZN(new_n367_));
  OAI21_X1   g0318(.A1(new_n366_), .A2(new_n367_), .B(new_n170_), .ZN(new_n368_));
  NOR2_X1    g0319(.A1(new_n237_), .A2(new_n245_), .ZN(new_n369_));
  NOR3_X1    g0320(.A1(new_n201_), .A2(new_n129_), .A3(new_n125_), .ZN(new_n370_));
  NAND2_X1   g0321(.A1(new_n224_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1     g0322(.I(new_n371_), .ZN(new_n372_));
  NOR4_X1    g0323(.A1(new_n372_), .A2(new_n238_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n373_));
  NOR2_X1    g0324(.A1(new_n225_), .A2(new_n217_), .ZN(new_n374_));
  NAND2_X1   g0325(.A1(new_n374_), .A2(new_n145_), .ZN(new_n375_));
  INV_X1     g0326(.I(new_n375_), .ZN(new_n376_));
  NOR2_X1    g0327(.A1(new_n171_), .A2(new_n208_), .ZN(new_n377_));
  NOR2_X1    g0328(.A1(new_n165_), .A2(new_n237_), .ZN(new_n378_));
  NOR3_X1    g0329(.A1(new_n140_), .A2(new_n201_), .A3(new_n150_), .ZN(new_n379_));
  NAND2_X1   g0330(.A1(new_n379_), .A2(new_n170_), .ZN(new_n380_));
  NAND2_X1   g0331(.A1(new_n288_), .A2(new_n380_), .ZN(new_n381_));
  NOR4_X1    g0332(.A1(new_n381_), .A2(new_n376_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n382_));
  NAND3_X1   g0333(.A1(new_n365_), .A2(new_n373_), .A3(new_n382_), .ZN(new_n383_));
  NOR2_X1    g0334(.A1(new_n191_), .A2(new_n241_), .ZN(new_n384_));
  NOR2_X1    g0335(.A1(new_n292_), .A2(new_n240_), .ZN(new_n385_));
  NOR4_X1    g0336(.A1(new_n385_), .A2(new_n192_), .A3(new_n242_), .A4(new_n384_), .ZN(new_n386_));
  NOR2_X1    g0337(.A1(new_n240_), .A2(new_n334_), .ZN(new_n387_));
  NAND2_X1   g0338(.A1(new_n178_), .A2(new_n207_), .ZN(new_n388_));
  NOR2_X1    g0339(.A1(new_n337_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1    g0340(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NOR4_X1    g0341(.A1(new_n119_), .A2(new_n286_), .A3(new_n98_), .A4(new_n218_), .ZN(new_n391_));
  NOR2_X1    g0342(.A1(new_n307_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1    g0343(.A1(new_n269_), .A2(new_n171_), .ZN(new_n393_));
  NOR2_X1    g0344(.A1(new_n337_), .A2(new_n208_), .ZN(new_n394_));
  NOR2_X1    g0345(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1   g0346(.A1(new_n395_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n396_));
  NAND2_X1   g0347(.A1(new_n251_), .A2(new_n202_), .ZN(new_n397_));
  INV_X1     g0348(.I(new_n397_), .ZN(new_n398_));
  NOR4_X1    g0349(.A1(new_n260_), .A2(new_n88_), .A3(new_n140_), .A4(new_n217_), .ZN(new_n399_));
  NOR4_X1    g0350(.A1(new_n204_), .A2(new_n398_), .A3(new_n209_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1   g0351(.A1(new_n234_), .A2(new_n222_), .ZN(new_n401_));
  NOR4_X1    g0352(.A1(new_n273_), .A2(new_n119_), .A3(new_n144_), .A4(new_n218_), .ZN(new_n402_));
  NOR2_X1    g0353(.A1(new_n181_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1   g0354(.A1(new_n403_), .A2(new_n401_), .ZN(new_n404_));
  NOR3_X1    g0355(.A1(new_n396_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  OAI21_X1   g0356(.A1(new_n102_), .A2(new_n107_), .B(new_n88_), .ZN(new_n406_));
  NOR2_X1    g0357(.A1(new_n406_), .A2(new_n98_), .ZN(new_n407_));
  NAND2_X1   g0358(.A1(new_n407_), .A2(new_n370_), .ZN(new_n408_));
  AOI22_X1   g0359(.A1(new_n166_), .A2(new_n173_), .B1(new_n142_), .B2(new_n143_), .ZN(new_n409_));
  NOR3_X1    g0360(.A1(new_n119_), .A2(new_n88_), .A3(new_n140_), .ZN(new_n410_));
  NAND2_X1   g0361(.A1(new_n410_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1   g0362(.A1(new_n152_), .A2(new_n407_), .ZN(new_n412_));
  NAND4_X1   g0363(.A1(new_n312_), .A2(new_n408_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  NAND2_X1   g0364(.A1(new_n405_), .A2(new_n413_), .ZN(new_n414_));
  NOR3_X1    g0365(.A1(new_n414_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n415_));
  INV_X1     g0366(.I(new_n415_), .ZN(new_n416_));
  OAI22_X1   g0367(.A1(new_n208_), .A2(new_n237_), .B1(new_n171_), .B2(new_n180_), .ZN(new_n417_));
  NAND2_X1   g0368(.A1(new_n152_), .A2(new_n295_), .ZN(new_n418_));
  NAND2_X1   g0369(.A1(new_n370_), .A2(new_n295_), .ZN(new_n419_));
  NAND2_X1   g0370(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR3_X1    g0371(.A1(new_n420_), .A2(new_n257_), .A3(new_n417_), .ZN(new_n421_));
  NOR2_X1    g0372(.A1(new_n240_), .A2(new_n279_), .ZN(new_n422_));
  NAND2_X1   g0373(.A1(new_n179_), .A2(new_n231_), .ZN(new_n423_));
  NOR2_X1    g0374(.A1(new_n265_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1   g0375(.A1(new_n151_), .A2(new_n141_), .ZN(new_n425_));
  NOR2_X1    g0376(.A1(new_n265_), .A2(new_n388_), .ZN(new_n426_));
  NOR2_X1    g0377(.A1(new_n377_), .A2(new_n426_), .ZN(new_n427_));
  NOR3_X1    g0378(.A1(new_n217_), .A2(new_n129_), .A3(new_n125_), .ZN(new_n428_));
  OAI21_X1   g0379(.A1(new_n428_), .A2(new_n318_), .B(new_n295_), .ZN(new_n429_));
  NAND4_X1   g0380(.A1(new_n427_), .A2(new_n425_), .A3(new_n341_), .A4(new_n429_), .ZN(new_n430_));
  NOR4_X1    g0381(.A1(new_n430_), .A2(new_n267_), .A3(new_n422_), .A4(new_n424_), .ZN(new_n431_));
  NAND2_X1   g0382(.A1(new_n431_), .A2(new_n421_), .ZN(new_n432_));
  NAND2_X1   g0383(.A1(new_n210_), .A2(new_n179_), .ZN(new_n433_));
  NOR2_X1    g0384(.A1(new_n433_), .A2(new_n171_), .ZN(new_n434_));
  NOR2_X1    g0385(.A1(new_n292_), .A2(new_n188_), .ZN(new_n435_));
  NOR3_X1    g0386(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NOR2_X1    g0387(.A1(new_n245_), .A2(new_n188_), .ZN(new_n437_));
  NOR2_X1    g0388(.A1(new_n197_), .A2(new_n191_), .ZN(new_n438_));
  NAND2_X1   g0389(.A1(new_n152_), .A2(new_n255_), .ZN(new_n439_));
  NAND4_X1   g0390(.A1(new_n187_), .A2(new_n207_), .A3(new_n231_), .A4(new_n88_), .ZN(new_n440_));
  NAND2_X1   g0391(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1   g0392(.A1(new_n318_), .A2(new_n190_), .A3(new_n243_), .ZN(new_n442_));
  NAND2_X1   g0393(.A1(new_n442_), .A2(new_n316_), .ZN(new_n443_));
  NOR4_X1    g0394(.A1(new_n441_), .A2(new_n443_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n444_));
  NAND2_X1   g0395(.A1(new_n287_), .A2(new_n367_), .ZN(new_n445_));
  NAND2_X1   g0396(.A1(new_n151_), .A2(new_n367_), .ZN(new_n446_));
  NAND3_X1   g0397(.A1(new_n408_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1   g0398(.A1(new_n285_), .A2(new_n88_), .A3(new_n170_), .ZN(new_n448_));
  NAND2_X1   g0399(.A1(new_n285_), .A2(new_n251_), .ZN(new_n449_));
  NAND3_X1   g0400(.A1(new_n448_), .A2(new_n449_), .A3(new_n397_), .ZN(new_n450_));
  NOR2_X1    g0401(.A1(new_n450_), .A2(new_n447_), .ZN(new_n451_));
  NAND2_X1   g0402(.A1(new_n109_), .A2(new_n318_), .ZN(new_n452_));
  NAND2_X1   g0403(.A1(new_n226_), .A2(new_n407_), .ZN(new_n453_));
  NAND2_X1   g0404(.A1(new_n453_), .A2(new_n452_), .ZN(new_n454_));
  NAND2_X1   g0405(.A1(new_n219_), .A2(new_n295_), .ZN(new_n455_));
  NAND3_X1   g0406(.A1(new_n203_), .A2(new_n455_), .A3(new_n321_), .ZN(new_n456_));
  NOR2_X1    g0407(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  NAND4_X1   g0408(.A1(new_n187_), .A2(new_n178_), .A3(new_n207_), .A4(new_n88_), .ZN(new_n458_));
  NAND2_X1   g0409(.A1(new_n401_), .A2(new_n458_), .ZN(new_n459_));
  NOR3_X1    g0410(.A1(new_n459_), .A2(new_n246_), .A3(new_n300_), .ZN(new_n460_));
  NOR4_X1    g0411(.A1(new_n119_), .A2(new_n299_), .A3(new_n88_), .A4(new_n140_), .ZN(new_n461_));
  NOR2_X1    g0412(.A1(new_n391_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1   g0413(.A1(new_n222_), .A2(new_n428_), .ZN(new_n463_));
  NAND3_X1   g0414(.A1(new_n312_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NOR2_X1    g0415(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1   g0416(.A1(new_n465_), .A2(new_n444_), .A3(new_n451_), .A4(new_n457_), .ZN(new_n466_));
  INV_X1     g0417(.I(new_n278_), .ZN(new_n467_));
  NAND2_X1   g0418(.A1(new_n130_), .A2(new_n222_), .ZN(new_n468_));
  NAND2_X1   g0419(.A1(new_n234_), .A2(new_n224_), .ZN(new_n469_));
  NAND3_X1   g0420(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NOR4_X1    g0421(.A1(new_n225_), .A2(new_n286_), .A3(new_n98_), .A4(new_n201_), .ZN(new_n471_));
  NOR4_X1    g0422(.A1(new_n119_), .A2(new_n286_), .A3(new_n98_), .A4(new_n140_), .ZN(new_n472_));
  NOR2_X1    g0423(.A1(new_n237_), .A2(new_n388_), .ZN(new_n473_));
  NOR4_X1    g0424(.A1(new_n307_), .A2(new_n473_), .A3(new_n471_), .A4(new_n472_), .ZN(new_n474_));
  NAND2_X1   g0425(.A1(new_n283_), .A2(new_n151_), .ZN(new_n475_));
  NAND2_X1   g0426(.A1(new_n285_), .A2(new_n109_), .ZN(new_n476_));
  NAND2_X1   g0427(.A1(new_n476_), .A2(new_n475_), .ZN(new_n477_));
  NOR2_X1    g0428(.A1(new_n191_), .A2(new_n423_), .ZN(new_n478_));
  NOR4_X1    g0429(.A1(new_n470_), .A2(new_n474_), .A3(new_n477_), .A4(new_n478_), .ZN(new_n479_));
  NAND2_X1   g0430(.A1(new_n151_), .A2(new_n370_), .ZN(new_n480_));
  NAND2_X1   g0431(.A1(new_n318_), .A2(new_n255_), .ZN(new_n481_));
  NAND3_X1   g0432(.A1(new_n480_), .A2(new_n481_), .A3(new_n343_), .ZN(new_n482_));
  INV_X1     g0433(.I(new_n232_), .ZN(new_n483_));
  NOR2_X1    g0434(.A1(new_n346_), .A2(new_n260_), .ZN(new_n484_));
  NOR4_X1    g0435(.A1(new_n484_), .A2(new_n483_), .A3(new_n301_), .A4(new_n324_), .ZN(new_n485_));
  NOR2_X1    g0436(.A1(new_n485_), .A2(new_n482_), .ZN(new_n486_));
  NOR4_X1    g0437(.A1(new_n299_), .A2(new_n140_), .A3(new_n201_), .A4(new_n88_), .ZN(new_n487_));
  NOR4_X1    g0438(.A1(new_n119_), .A2(new_n221_), .A3(new_n150_), .A4(new_n218_), .ZN(new_n488_));
  NOR2_X1    g0439(.A1(new_n488_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1   g0440(.A1(new_n224_), .A2(new_n428_), .ZN(new_n490_));
  AND4_X2    g0441(.A1(new_n329_), .A2(new_n489_), .A3(new_n412_), .A4(new_n490_), .Z(new_n491_));
  NAND4_X1   g0442(.A1(new_n479_), .A2(new_n486_), .A3(new_n182_), .A4(new_n491_), .ZN(new_n492_));
  NOR2_X1    g0443(.A1(new_n466_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1   g0444(.A1(new_n436_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1    g0445(.A1(new_n240_), .A2(new_n423_), .ZN(new_n495_));
  NOR4_X1    g0446(.A1(new_n495_), .A2(new_n280_), .A3(new_n437_), .A4(new_n307_), .ZN(new_n496_));
  OAI21_X1   g0447(.A1(new_n226_), .A2(new_n227_), .B(new_n255_), .ZN(new_n497_));
  NAND2_X1   g0448(.A1(new_n395_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1   g0449(.A1(new_n196_), .A2(new_n231_), .ZN(new_n499_));
  NOR2_X1    g0450(.A1(new_n499_), .A2(new_n265_), .ZN(new_n500_));
  NOR2_X1    g0451(.A1(new_n208_), .A2(new_n265_), .ZN(new_n501_));
  NOR3_X1    g0452(.A1(new_n420_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1   g0453(.A1(new_n151_), .A2(new_n219_), .ZN(new_n503_));
  NAND2_X1   g0454(.A1(new_n227_), .A2(new_n295_), .ZN(new_n504_));
  NAND2_X1   g0455(.A1(new_n224_), .A2(new_n233_), .ZN(new_n505_));
  NAND4_X1   g0456(.A1(new_n503_), .A2(new_n309_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  NOR2_X1    g0457(.A1(new_n237_), .A2(new_n423_), .ZN(new_n507_));
  NOR2_X1    g0458(.A1(new_n172_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1   g0459(.A1(new_n196_), .A2(new_n178_), .ZN(new_n509_));
  AOI21_X1   g0460(.A1(new_n509_), .A2(new_n208_), .B(new_n188_), .ZN(new_n510_));
  INV_X1     g0461(.I(new_n510_), .ZN(new_n511_));
  NAND3_X1   g0462(.A1(new_n506_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n512_));
  NOR4_X1    g0463(.A1(new_n512_), .A2(new_n496_), .A3(new_n498_), .A4(new_n502_), .ZN(new_n513_));
  NOR2_X1    g0464(.A1(new_n292_), .A2(new_n191_), .ZN(new_n514_));
  INV_X1     g0465(.I(new_n440_), .ZN(new_n515_));
  NOR2_X1    g0466(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1   g0467(.A1(new_n241_), .A2(new_n279_), .B(new_n265_), .ZN(new_n517_));
  INV_X1     g0468(.I(new_n452_), .ZN(new_n518_));
  NOR2_X1    g0469(.A1(new_n279_), .A2(new_n188_), .ZN(new_n519_));
  NOR2_X1    g0470(.A1(new_n171_), .A2(new_n279_), .ZN(new_n520_));
  NOR4_X1    g0471(.A1(new_n518_), .A2(new_n339_), .A3(new_n519_), .A4(new_n520_), .ZN(new_n521_));
  OAI21_X1   g0472(.A1(new_n188_), .A2(new_n241_), .B(new_n401_), .ZN(new_n522_));
  NOR4_X1    g0473(.A1(new_n521_), .A2(new_n214_), .A3(new_n517_), .A4(new_n522_), .ZN(new_n523_));
  NOR4_X1    g0474(.A1(new_n299_), .A2(new_n218_), .A3(new_n201_), .A4(new_n150_), .ZN(new_n524_));
  NOR2_X1    g0475(.A1(new_n237_), .A2(new_n241_), .ZN(new_n525_));
  NOR4_X1    g0476(.A1(new_n119_), .A2(new_n225_), .A3(new_n299_), .A4(new_n150_), .ZN(new_n526_));
  NOR4_X1    g0477(.A1(new_n525_), .A2(new_n266_), .A3(new_n524_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1     g0478(.I(new_n301_), .ZN(new_n528_));
  NOR2_X1    g0479(.A1(new_n509_), .A2(new_n265_), .ZN(new_n529_));
  INV_X1     g0480(.I(new_n529_), .ZN(new_n530_));
  NAND3_X1   g0481(.A1(new_n528_), .A2(new_n530_), .A3(new_n329_), .ZN(new_n531_));
  NAND2_X1   g0482(.A1(new_n251_), .A2(new_n219_), .ZN(new_n532_));
  INV_X1     g0483(.I(new_n532_), .ZN(new_n533_));
  NOR4_X1    g0484(.A1(new_n119_), .A2(new_n273_), .A3(new_n225_), .A4(new_n144_), .ZN(new_n534_));
  NOR2_X1    g0485(.A1(new_n433_), .A2(new_n191_), .ZN(new_n535_));
  NOR4_X1    g0486(.A1(new_n533_), .A2(new_n535_), .A3(new_n402_), .A4(new_n534_), .ZN(new_n536_));
  NOR4_X1    g0487(.A1(new_n536_), .A2(new_n531_), .A3(new_n289_), .A4(new_n527_), .ZN(new_n537_));
  AND4_X2    g0488(.A1(new_n513_), .A2(new_n516_), .A3(new_n523_), .A4(new_n537_), .Z(new_n538_));
  NAND4_X1   g0489(.A1(new_n174_), .A2(new_n196_), .A3(new_n108_), .A4(new_n178_), .ZN(new_n539_));
  NAND3_X1   g0490(.A1(new_n359_), .A2(new_n304_), .A3(new_n439_), .ZN(new_n540_));
  NOR4_X1    g0491(.A1(new_n398_), .A2(new_n422_), .A3(new_n322_), .A4(new_n426_), .ZN(new_n541_));
  NAND2_X1   g0492(.A1(new_n151_), .A2(new_n202_), .ZN(new_n542_));
  NAND2_X1   g0493(.A1(new_n375_), .A2(new_n542_), .ZN(new_n543_));
  NOR3_X1    g0494(.A1(new_n541_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  NAND3_X1   g0495(.A1(new_n285_), .A2(new_n88_), .A3(new_n187_), .ZN(new_n545_));
  NAND3_X1   g0496(.A1(new_n544_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n546_));
  NAND4_X1   g0497(.A1(new_n210_), .A2(new_n187_), .A3(new_n88_), .A4(new_n207_), .ZN(new_n547_));
  NOR2_X1    g0498(.A1(new_n135_), .A2(new_n134_), .ZN(new_n548_));
  NAND3_X1   g0499(.A1(new_n151_), .A2(new_n548_), .A3(new_n196_), .ZN(new_n549_));
  NAND4_X1   g0500(.A1(new_n187_), .A2(new_n207_), .A3(new_n231_), .A4(new_n150_), .ZN(new_n550_));
  NAND2_X1   g0501(.A1(new_n222_), .A2(new_n318_), .ZN(new_n551_));
  NAND4_X1   g0502(.A1(new_n549_), .A2(new_n551_), .A3(new_n547_), .A4(new_n550_), .ZN(new_n552_));
  NOR4_X1    g0503(.A1(new_n119_), .A2(new_n225_), .A3(new_n299_), .A4(new_n88_), .ZN(new_n553_));
  NOR2_X1    g0504(.A1(new_n553_), .A2(new_n327_), .ZN(new_n554_));
  NAND4_X1   g0505(.A1(new_n552_), .A2(new_n458_), .A3(new_n490_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1   g0506(.A1(new_n407_), .A2(new_n367_), .ZN(new_n556_));
  NAND2_X1   g0507(.A1(new_n233_), .A2(new_n295_), .ZN(new_n557_));
  NOR2_X1    g0508(.A1(new_n129_), .A2(new_n125_), .ZN(new_n558_));
  NAND3_X1   g0509(.A1(new_n255_), .A2(new_n558_), .A3(new_n210_), .ZN(new_n559_));
  NAND3_X1   g0510(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1    g0511(.A1(new_n237_), .A2(new_n180_), .ZN(new_n561_));
  NOR4_X1    g0512(.A1(new_n204_), .A2(new_n561_), .A3(new_n483_), .A4(new_n478_), .ZN(new_n562_));
  NOR2_X1    g0513(.A1(new_n269_), .A2(new_n244_), .ZN(new_n563_));
  NOR2_X1    g0514(.A1(new_n563_), .A2(new_n399_), .ZN(new_n564_));
  NAND4_X1   g0515(.A1(new_n562_), .A2(new_n462_), .A3(new_n560_), .A4(new_n564_), .ZN(new_n565_));
  NOR3_X1    g0516(.A1(new_n546_), .A2(new_n555_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1   g0517(.A1(new_n538_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1   g0518(.A1(new_n567_), .A2(new_n494_), .ZN(new_n568_));
  NAND2_X1   g0519(.A1(new_n568_), .A2(new_n416_), .ZN(new_n569_));
  INV_X1     g0520(.I(\a[11] ), .ZN(new_n570_));
  INV_X1     g0521(.I(new_n110_), .ZN(new_n571_));
  NOR2_X1    g0522(.A1(new_n571_), .A2(\a[10] ), .ZN(new_n572_));
  OAI21_X1   g0523(.A1(new_n572_), .A2(\a[22] ), .B(new_n570_), .ZN(new_n573_));
  INV_X1     g0524(.I(new_n572_), .ZN(new_n574_));
  NAND3_X1   g0525(.A1(new_n574_), .A2(\a[11] ), .A3(new_n80_), .ZN(new_n575_));
  NAND2_X1   g0526(.A1(new_n575_), .A2(new_n573_), .ZN(new_n576_));
  AOI21_X1   g0527(.A1(new_n574_), .A2(\a[11] ), .B(\a[22] ), .ZN(new_n577_));
  NOR2_X1    g0528(.A1(new_n577_), .A2(\a[12] ), .ZN(new_n578_));
  NAND2_X1   g0529(.A1(new_n577_), .A2(\a[12] ), .ZN(new_n579_));
  INV_X1     g0530(.I(new_n579_), .ZN(new_n580_));
  NOR2_X1    g0531(.A1(new_n580_), .A2(new_n578_), .ZN(new_n581_));
  INV_X1     g0532(.I(new_n581_), .ZN(new_n582_));
  NOR2_X1    g0533(.A1(new_n582_), .A2(new_n576_), .ZN(new_n583_));
  NOR2_X1    g0534(.A1(new_n433_), .A2(new_n265_), .ZN(new_n584_));
  NOR4_X1    g0535(.A1(new_n336_), .A2(new_n584_), .A3(new_n519_), .A4(new_n424_), .ZN(new_n585_));
  INV_X1     g0536(.I(new_n585_), .ZN(new_n586_));
  NOR2_X1    g0537(.A1(new_n293_), .A2(new_n524_), .ZN(new_n587_));
  NOR2_X1    g0538(.A1(new_n270_), .A2(new_n241_), .ZN(new_n588_));
  NOR2_X1    g0539(.A1(new_n433_), .A2(new_n188_), .ZN(new_n589_));
  NOR3_X1    g0540(.A1(new_n263_), .A2(new_n589_), .A3(new_n588_), .ZN(new_n590_));
  NAND3_X1   g0541(.A1(new_n586_), .A2(new_n590_), .A3(new_n587_), .ZN(new_n591_));
  INV_X1     g0542(.I(new_n591_), .ZN(new_n592_));
  NOR2_X1    g0543(.A1(new_n244_), .A2(new_n388_), .ZN(new_n593_));
  NOR2_X1    g0544(.A1(new_n245_), .A2(new_n265_), .ZN(new_n594_));
  NOR3_X1    g0545(.A1(new_n499_), .A2(new_n150_), .A3(new_n299_), .ZN(new_n595_));
  NOR3_X1    g0546(.A1(new_n595_), .A2(new_n189_), .A3(new_n594_), .ZN(new_n596_));
  NOR2_X1    g0547(.A1(new_n175_), .A2(new_n334_), .ZN(new_n597_));
  NOR2_X1    g0548(.A1(new_n597_), .A2(new_n500_), .ZN(new_n598_));
  NAND4_X1   g0549(.A1(new_n596_), .A2(new_n418_), .A3(new_n598_), .A4(new_n446_), .ZN(new_n599_));
  NOR3_X1    g0550(.A1(new_n599_), .A2(new_n593_), .A3(new_n472_), .ZN(new_n600_));
  NOR2_X1    g0551(.A1(new_n306_), .A2(new_n501_), .ZN(new_n601_));
  NOR2_X1    g0552(.A1(new_n267_), .A2(new_n553_), .ZN(new_n602_));
  NOR4_X1    g0553(.A1(new_n299_), .A2(new_n140_), .A3(new_n217_), .A4(new_n150_), .ZN(new_n603_));
  NOR4_X1    g0554(.A1(new_n529_), .A2(new_n426_), .A3(new_n603_), .A4(new_n526_), .ZN(new_n604_));
  AOI21_X1   g0555(.A1(new_n601_), .A2(new_n602_), .B(new_n604_), .ZN(new_n605_));
  NAND3_X1   g0556(.A1(new_n592_), .A2(new_n600_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1     g0557(.I(new_n606_), .ZN(new_n607_));
  INV_X1     g0558(.I(new_n480_), .ZN(new_n608_));
  NOR2_X1    g0559(.A1(new_n98_), .A2(new_n144_), .ZN(new_n609_));
  NAND2_X1   g0560(.A1(new_n152_), .A2(new_n609_), .ZN(new_n610_));
  NOR4_X1    g0561(.A1(new_n608_), .A2(new_n266_), .A3(new_n435_), .A4(new_n610_), .ZN(new_n611_));
  NAND2_X1   g0562(.A1(new_n325_), .A2(new_n321_), .ZN(new_n612_));
  NAND2_X1   g0563(.A1(new_n287_), .A2(new_n370_), .ZN(new_n613_));
  NAND2_X1   g0564(.A1(new_n528_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1   g0565(.A1(new_n319_), .A2(new_n310_), .ZN(new_n615_));
  NOR4_X1    g0566(.A1(new_n614_), .A2(new_n615_), .A3(new_n517_), .A4(new_n612_), .ZN(new_n616_));
  NAND2_X1   g0567(.A1(new_n616_), .A2(new_n611_), .ZN(new_n617_));
  INV_X1     g0568(.I(new_n617_), .ZN(new_n618_));
  NAND4_X1   g0569(.A1(new_n243_), .A2(new_n190_), .A3(new_n207_), .A4(new_n231_), .ZN(new_n619_));
  NOR2_X1    g0570(.A1(new_n195_), .A2(new_n208_), .ZN(new_n620_));
  NOR2_X1    g0571(.A1(new_n620_), .A2(new_n437_), .ZN(new_n621_));
  NAND3_X1   g0572(.A1(new_n621_), .A2(new_n619_), .A3(new_n344_), .ZN(new_n622_));
  NOR2_X1    g0573(.A1(new_n239_), .A2(new_n300_), .ZN(new_n623_));
  NAND2_X1   g0574(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1    g0575(.A1(new_n226_), .A2(new_n202_), .ZN(new_n625_));
  NOR4_X1    g0576(.A1(new_n624_), .A2(new_n299_), .A3(new_n510_), .A4(new_n625_), .ZN(new_n626_));
  NAND3_X1   g0577(.A1(new_n607_), .A2(new_n618_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1     g0578(.I(new_n627_), .ZN(new_n628_));
  AOI21_X1   g0579(.A1(new_n576_), .A2(new_n582_), .B(new_n628_), .ZN(new_n629_));
  OAI21_X1   g0580(.A1(new_n569_), .A2(new_n583_), .B(new_n629_), .ZN(new_n630_));
  NOR2_X1    g0581(.A1(new_n171_), .A2(new_n180_), .ZN(new_n631_));
  OAI22_X1   g0582(.A1(new_n165_), .A2(new_n171_), .B1(new_n237_), .B2(new_n423_), .ZN(new_n632_));
  NAND4_X1   g0583(.A1(new_n463_), .A2(new_n490_), .A3(new_n551_), .A4(new_n505_), .ZN(new_n633_));
  NAND2_X1   g0584(.A1(new_n224_), .A2(new_n318_), .ZN(new_n634_));
  NAND4_X1   g0585(.A1(new_n329_), .A2(new_n468_), .A3(new_n634_), .A4(new_n223_), .ZN(new_n635_));
  NOR3_X1    g0586(.A1(new_n635_), .A2(new_n633_), .A3(new_n632_), .ZN(new_n636_));
  NAND3_X1   g0587(.A1(new_n636_), .A2(new_n392_), .A3(new_n403_), .ZN(new_n637_));
  NOR2_X1    g0588(.A1(new_n499_), .A2(new_n171_), .ZN(new_n638_));
  NAND2_X1   g0589(.A1(new_n227_), .A2(new_n222_), .ZN(new_n639_));
  NAND2_X1   g0590(.A1(new_n639_), .A2(new_n291_), .ZN(new_n640_));
  NAND3_X1   g0591(.A1(new_n224_), .A2(new_n548_), .A3(new_n196_), .ZN(new_n641_));
  INV_X1     g0592(.I(new_n641_), .ZN(new_n642_));
  NOR4_X1    g0593(.A1(new_n225_), .A2(new_n221_), .A3(new_n150_), .A4(new_n217_), .ZN(new_n643_));
  NOR4_X1    g0594(.A1(new_n640_), .A2(new_n642_), .A3(new_n638_), .A4(new_n643_), .ZN(new_n644_));
  INV_X1     g0595(.I(new_n434_), .ZN(new_n645_));
  NAND4_X1   g0596(.A1(new_n548_), .A2(new_n88_), .A3(new_n170_), .A4(new_n196_), .ZN(new_n646_));
  NAND3_X1   g0597(.A1(new_n645_), .A2(new_n448_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1     g0598(.I(new_n647_), .ZN(new_n648_));
  NAND2_X1   g0599(.A1(new_n648_), .A2(new_n644_), .ZN(new_n649_));
  NOR4_X1    g0600(.A1(new_n383_), .A2(new_n631_), .A3(new_n637_), .A4(new_n649_), .ZN(new_n650_));
  XNOR2_X1   g0601(.A1(new_n650_), .A2(new_n415_), .ZN(new_n651_));
  NOR2_X1    g0602(.A1(new_n650_), .A2(new_n415_), .ZN(new_n652_));
  XNOR2_X1   g0603(.A1(new_n627_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1   g0604(.A1(new_n84_), .A2(\a[13] ), .B(\a[22] ), .ZN(new_n654_));
  NOR2_X1    g0605(.A1(new_n654_), .A2(\a[14] ), .ZN(new_n655_));
  NAND2_X1   g0606(.A1(new_n654_), .A2(\a[14] ), .ZN(new_n656_));
  INV_X1     g0607(.I(new_n656_), .ZN(new_n657_));
  NOR2_X1    g0608(.A1(new_n657_), .A2(new_n655_), .ZN(new_n658_));
  INV_X1     g0609(.I(new_n658_), .ZN(new_n659_));
  NOR2_X1    g0610(.A1(new_n627_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1    g0611(.A1(new_n628_), .A2(new_n658_), .ZN(new_n661_));
  NOR2_X1    g0612(.A1(new_n661_), .A2(new_n660_), .ZN(new_n662_));
  AOI21_X1   g0613(.A1(new_n651_), .A2(new_n662_), .B(new_n653_), .ZN(new_n663_));
  AOI21_X1   g0614(.A1(new_n84_), .A2(new_n80_), .B(\a[13] ), .ZN(new_n664_));
  INV_X1     g0615(.I(\a[13] ), .ZN(new_n665_));
  NOR2_X1    g0616(.A1(new_n665_), .A2(\a[22] ), .ZN(new_n666_));
  AOI21_X1   g0617(.A1(new_n84_), .A2(new_n666_), .B(new_n664_), .ZN(new_n667_));
  NAND2_X1   g0618(.A1(new_n627_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1   g0619(.A1(new_n663_), .A2(new_n668_), .ZN(new_n669_));
  XOR2_X1    g0620(.A1(new_n669_), .A2(new_n630_), .Z(new_n670_));
  NOR2_X1    g0621(.A1(new_n651_), .A2(new_n627_), .ZN(new_n671_));
  NAND2_X1   g0622(.A1(new_n650_), .A2(new_n415_), .ZN(new_n672_));
  NOR2_X1    g0623(.A1(new_n650_), .A2(new_n415_), .ZN(new_n673_));
  INV_X1     g0624(.I(new_n673_), .ZN(new_n674_));
  NAND3_X1   g0625(.A1(new_n674_), .A2(new_n627_), .A3(new_n672_), .ZN(new_n675_));
  INV_X1     g0626(.I(new_n675_), .ZN(new_n676_));
  NOR3_X1    g0627(.A1(new_n676_), .A2(new_n671_), .A3(new_n658_), .ZN(new_n677_));
  INV_X1     g0628(.I(new_n667_), .ZN(new_n678_));
  OAI21_X1   g0629(.A1(new_n628_), .A2(new_n674_), .B(new_n672_), .ZN(new_n679_));
  NOR2_X1    g0630(.A1(new_n679_), .A2(new_n678_), .ZN(new_n680_));
  NOR2_X1    g0631(.A1(new_n627_), .A2(new_n672_), .ZN(new_n681_));
  NOR2_X1    g0632(.A1(new_n681_), .A2(new_n673_), .ZN(new_n682_));
  AOI21_X1   g0633(.A1(new_n678_), .A2(new_n682_), .B(new_n680_), .ZN(new_n683_));
  NAND2_X1   g0634(.A1(new_n683_), .A2(new_n677_), .ZN(new_n684_));
  XOR2_X1    g0635(.A1(new_n581_), .A2(new_n576_), .Z(new_n685_));
  INV_X1     g0636(.I(new_n685_), .ZN(new_n686_));
  NAND2_X1   g0637(.A1(new_n627_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1   g0638(.A1(new_n569_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X2    g0639(.A1(new_n684_), .A2(new_n688_), .Z(new_n689_));
  XNOR2_X1   g0640(.A1(new_n567_), .A2(new_n494_), .ZN(new_n690_));
  NAND2_X1   g0641(.A1(new_n567_), .A2(new_n494_), .ZN(new_n691_));
  XOR2_X1    g0642(.A1(new_n691_), .A2(new_n416_), .Z(new_n692_));
  XOR2_X1    g0643(.A1(new_n415_), .A2(new_n658_), .Z(new_n693_));
  AOI21_X1   g0644(.A1(new_n690_), .A2(new_n693_), .B(new_n692_), .ZN(new_n694_));
  NOR3_X1    g0645(.A1(new_n694_), .A2(new_n576_), .A3(new_n628_), .ZN(new_n695_));
  INV_X1     g0646(.I(new_n671_), .ZN(new_n696_));
  NOR2_X1    g0647(.A1(new_n679_), .A2(new_n582_), .ZN(new_n697_));
  AOI21_X1   g0648(.A1(new_n582_), .A2(new_n682_), .B(new_n697_), .ZN(new_n698_));
  NAND4_X1   g0649(.A1(new_n698_), .A2(new_n678_), .A3(new_n696_), .A4(new_n675_), .ZN(new_n699_));
  INV_X1     g0650(.I(new_n694_), .ZN(new_n700_));
  NOR2_X1    g0651(.A1(new_n628_), .A2(new_n576_), .ZN(new_n701_));
  NOR2_X1    g0652(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1     g0653(.I(new_n702_), .ZN(new_n703_));
  AOI21_X1   g0654(.A1(new_n703_), .A2(new_n699_), .B(new_n695_), .ZN(new_n704_));
  NOR2_X1    g0655(.A1(new_n684_), .A2(new_n688_), .ZN(new_n705_));
  NOR2_X1    g0656(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1    g0657(.A1(new_n706_), .A2(new_n689_), .ZN(new_n707_));
  XOR2_X1    g0658(.A1(new_n707_), .A2(new_n670_), .Z(new_n708_));
  NAND2_X1   g0659(.A1(new_n708_), .A2(new_n670_), .ZN(new_n709_));
  NAND2_X1   g0660(.A1(new_n407_), .A2(new_n141_), .ZN(new_n710_));
  NAND4_X1   g0661(.A1(new_n196_), .A2(new_n170_), .A3(new_n88_), .A4(new_n178_), .ZN(new_n711_));
  NAND4_X1   g0662(.A1(new_n131_), .A2(new_n490_), .A3(new_n634_), .A4(new_n711_), .ZN(new_n712_));
  NAND3_X1   g0663(.A1(new_n712_), .A2(new_n528_), .A3(new_n710_), .ZN(new_n713_));
  NAND2_X1   g0664(.A1(new_n428_), .A2(new_n295_), .ZN(new_n714_));
  INV_X1     g0665(.I(new_n714_), .ZN(new_n715_));
  OR3_X2     g0666(.A1(new_n404_), .A2(new_n209_), .A3(new_n715_), .Z(new_n716_));
  NOR4_X1    g0667(.A1(new_n406_), .A2(new_n225_), .A3(new_n98_), .A4(new_n217_), .ZN(new_n717_));
  NOR4_X1    g0668(.A1(new_n608_), .A2(new_n172_), .A3(new_n588_), .A4(new_n717_), .ZN(new_n718_));
  INV_X1     g0669(.I(new_n335_), .ZN(new_n719_));
  INV_X1     g0670(.I(new_n507_), .ZN(new_n720_));
  NAND4_X1   g0671(.A1(new_n719_), .A2(new_n720_), .A3(new_n453_), .A4(new_n646_), .ZN(new_n721_));
  INV_X1     g0672(.I(new_n721_), .ZN(new_n722_));
  NOR4_X1    g0673(.A1(new_n716_), .A2(new_n713_), .A3(new_n718_), .A4(new_n722_), .ZN(new_n723_));
  NOR4_X1    g0674(.A1(new_n250_), .A2(new_n280_), .A3(new_n631_), .A4(new_n472_), .ZN(new_n724_));
  NOR3_X1    g0675(.A1(new_n724_), .A2(new_n424_), .A3(new_n435_), .ZN(new_n725_));
  NAND2_X1   g0676(.A1(new_n224_), .A2(new_n141_), .ZN(new_n726_));
  INV_X1     g0677(.I(new_n384_), .ZN(new_n727_));
  NOR2_X1    g0678(.A1(new_n339_), .A2(new_n422_), .ZN(new_n728_));
  NOR2_X1    g0679(.A1(new_n324_), .A2(new_n399_), .ZN(new_n729_));
  NAND4_X1   g0680(.A1(new_n728_), .A2(new_n726_), .A3(new_n727_), .A4(new_n729_), .ZN(new_n730_));
  NOR2_X1    g0681(.A1(new_n212_), .A2(new_n391_), .ZN(new_n731_));
  NAND2_X1   g0682(.A1(new_n731_), .A2(new_n532_), .ZN(new_n732_));
  NAND2_X1   g0683(.A1(new_n130_), .A2(new_n287_), .ZN(new_n733_));
  NAND2_X1   g0684(.A1(new_n733_), .A2(new_n296_), .ZN(new_n734_));
  NOR4_X1    g0685(.A1(new_n730_), .A2(new_n478_), .A3(new_n732_), .A4(new_n734_), .ZN(new_n735_));
  NAND2_X1   g0686(.A1(new_n735_), .A2(new_n725_), .ZN(new_n736_));
  INV_X1     g0687(.I(new_n736_), .ZN(new_n737_));
  INV_X1     g0688(.I(new_n551_), .ZN(new_n738_));
  NOR3_X1    g0689(.A1(new_n738_), .A2(new_n526_), .A3(new_n589_), .ZN(new_n739_));
  NAND4_X1   g0690(.A1(new_n146_), .A2(new_n449_), .A3(new_n504_), .A4(new_n425_), .ZN(new_n740_));
  INV_X1     g0691(.I(new_n446_), .ZN(new_n741_));
  NOR3_X1    g0692(.A1(new_n376_), .A2(new_n741_), .A3(new_n360_), .ZN(new_n742_));
  NAND3_X1   g0693(.A1(new_n742_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n743_));
  NOR4_X1    g0694(.A1(new_n398_), .A2(new_n326_), .A3(new_n638_), .A4(new_n369_), .ZN(new_n744_));
  NOR3_X1    g0695(.A1(new_n744_), .A2(new_n311_), .A3(new_n524_), .ZN(new_n745_));
  NOR4_X1    g0696(.A1(new_n484_), .A2(new_n192_), .A3(new_n434_), .A4(new_n553_), .ZN(new_n746_));
  NOR2_X1    g0697(.A1(new_n171_), .A2(new_n388_), .ZN(new_n747_));
  NOR4_X1    g0698(.A1(new_n595_), .A2(new_n529_), .A3(new_n747_), .A4(new_n274_), .ZN(new_n748_));
  NOR2_X1    g0699(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1   g0700(.A1(new_n745_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1    g0701(.A1(new_n750_), .A2(new_n743_), .ZN(new_n751_));
  NAND3_X1   g0702(.A1(new_n737_), .A2(new_n723_), .A3(new_n751_), .ZN(new_n752_));
  AND2_X2    g0703(.A1(new_n513_), .A2(new_n516_), .Z(new_n753_));
  NOR3_X1    g0704(.A1(new_n540_), .A2(new_n209_), .A3(new_n239_), .ZN(new_n754_));
  NOR2_X1    g0705(.A1(new_n250_), .A2(new_n638_), .ZN(new_n755_));
  NAND3_X1   g0706(.A1(new_n755_), .A2(new_n445_), .A3(new_n545_), .ZN(new_n756_));
  NOR3_X1    g0707(.A1(new_n267_), .A2(new_n324_), .A3(new_n461_), .ZN(new_n757_));
  NOR4_X1    g0708(.A1(new_n597_), .A2(new_n242_), .A3(new_n525_), .A4(new_n278_), .ZN(new_n758_));
  NAND3_X1   g0709(.A1(new_n411_), .A2(new_n356_), .A3(new_n458_), .ZN(new_n759_));
  NOR2_X1    g0710(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1   g0711(.A1(new_n754_), .A2(new_n760_), .A3(new_n756_), .A4(new_n757_), .ZN(new_n761_));
  OAI22_X1   g0712(.A1(new_n175_), .A2(new_n197_), .B1(new_n240_), .B2(new_n180_), .ZN(new_n762_));
  NOR3_X1    g0713(.A1(new_n417_), .A2(new_n192_), .A3(new_n261_), .ZN(new_n763_));
  NAND2_X1   g0714(.A1(new_n476_), .A2(new_n539_), .ZN(new_n764_));
  NOR3_X1    g0715(.A1(new_n763_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1   g0716(.A1(new_n765_), .A2(new_n719_), .A3(new_n646_), .ZN(new_n766_));
  NOR2_X1    g0717(.A1(new_n741_), .A2(new_n336_), .ZN(new_n767_));
  NOR2_X1    g0718(.A1(new_n588_), .A2(new_n300_), .ZN(new_n768_));
  NOR2_X1    g0719(.A1(new_n293_), .A2(new_n426_), .ZN(new_n769_));
  NAND4_X1   g0720(.A1(new_n767_), .A2(new_n489_), .A3(new_n768_), .A4(new_n769_), .ZN(new_n770_));
  INV_X1     g0721(.I(new_n747_), .ZN(new_n771_));
  NAND4_X1   g0722(.A1(new_n771_), .A2(new_n146_), .A3(new_n556_), .A4(new_n449_), .ZN(new_n772_));
  AOI21_X1   g0723(.A1(new_n142_), .A2(new_n143_), .B(new_n150_), .ZN(new_n773_));
  NAND4_X1   g0724(.A1(new_n773_), .A2(new_n196_), .A3(new_n190_), .A4(new_n178_), .ZN(new_n774_));
  NAND4_X1   g0725(.A1(new_n401_), .A2(new_n408_), .A3(new_n641_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1   g0726(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  NOR4_X1    g0727(.A1(new_n761_), .A2(new_n766_), .A3(new_n770_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1   g0728(.A1(new_n777_), .A2(new_n753_), .ZN(new_n778_));
  NAND2_X1   g0729(.A1(new_n778_), .A2(new_n752_), .ZN(new_n779_));
  NAND2_X1   g0730(.A1(new_n779_), .A2(new_n494_), .ZN(new_n780_));
  INV_X1     g0731(.I(new_n780_), .ZN(new_n781_));
  NOR2_X1    g0732(.A1(new_n778_), .A2(new_n752_), .ZN(new_n782_));
  INV_X1     g0733(.I(new_n782_), .ZN(new_n783_));
  NAND2_X1   g0734(.A1(new_n783_), .A2(new_n779_), .ZN(new_n784_));
  NOR2_X1    g0735(.A1(new_n784_), .A2(new_n781_), .ZN(new_n785_));
  NOR2_X1    g0736(.A1(new_n782_), .A2(new_n494_), .ZN(new_n786_));
  NOR2_X1    g0737(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NOR3_X1    g0738(.A1(new_n785_), .A2(new_n787_), .A3(new_n581_), .ZN(new_n788_));
  INV_X1     g0739(.I(new_n788_), .ZN(new_n789_));
  INV_X1     g0740(.I(new_n576_), .ZN(new_n790_));
  INV_X1     g0741(.I(new_n779_), .ZN(new_n791_));
  NOR2_X1    g0742(.A1(new_n791_), .A2(new_n782_), .ZN(new_n792_));
  NOR2_X1    g0743(.A1(new_n792_), .A2(new_n781_), .ZN(new_n793_));
  NOR2_X1    g0744(.A1(new_n793_), .A2(new_n790_), .ZN(new_n794_));
  NOR2_X1    g0745(.A1(new_n792_), .A2(new_n786_), .ZN(new_n795_));
  NOR2_X1    g0746(.A1(new_n795_), .A2(new_n576_), .ZN(new_n796_));
  NOR3_X1    g0747(.A1(new_n789_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1     g0748(.I(new_n797_), .ZN(new_n798_));
  NAND2_X1   g0749(.A1(new_n411_), .A2(new_n613_), .ZN(new_n799_));
  NOR4_X1    g0750(.A1(new_n799_), .A2(new_n250_), .A3(new_n274_), .A4(new_n529_), .ZN(new_n800_));
  INV_X1     g0751(.I(new_n453_), .ZN(new_n801_));
  NOR4_X1    g0752(.A1(new_n377_), .A2(new_n747_), .A3(new_n426_), .A4(new_n534_), .ZN(new_n802_));
  NOR4_X1    g0753(.A1(new_n802_), .A2(new_n338_), .A3(new_n801_), .A4(new_n478_), .ZN(new_n803_));
  NOR2_X1    g0754(.A1(new_n318_), .A2(new_n88_), .ZN(new_n804_));
  OAI21_X1   g0755(.A1(new_n804_), .A2(new_n410_), .B(new_n170_), .ZN(new_n805_));
  NOR4_X1    g0756(.A1(new_n597_), .A2(new_n487_), .A3(new_n507_), .A4(new_n643_), .ZN(new_n806_));
  NOR4_X1    g0757(.A1(new_n806_), .A2(new_n495_), .A3(new_n805_), .A4(new_n594_), .ZN(new_n807_));
  NAND4_X1   g0758(.A1(new_n803_), .A2(new_n807_), .A3(new_n332_), .A4(new_n800_), .ZN(new_n808_));
  NAND2_X1   g0759(.A1(new_n152_), .A2(new_n224_), .ZN(new_n809_));
  NAND4_X1   g0760(.A1(new_n809_), .A2(new_n439_), .A3(new_n476_), .A4(new_n203_), .ZN(new_n810_));
  NAND3_X1   g0761(.A1(new_n810_), .A2(new_n733_), .A3(new_n587_), .ZN(new_n811_));
  INV_X1     g0762(.I(new_n811_), .ZN(new_n812_));
  NAND2_X1   g0763(.A1(new_n224_), .A2(new_n219_), .ZN(new_n813_));
  NAND3_X1   g0764(.A1(new_n545_), .A2(new_n490_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1   g0765(.A1(new_n310_), .A2(new_n714_), .ZN(new_n815_));
  NOR4_X1    g0766(.A1(new_n814_), .A2(new_n336_), .A3(new_n815_), .A4(new_n603_), .ZN(new_n816_));
  NOR4_X1    g0767(.A1(new_n385_), .A2(new_n198_), .A3(new_n384_), .A4(new_n278_), .ZN(new_n817_));
  NOR2_X1    g0768(.A1(new_n817_), .A2(new_n450_), .ZN(new_n818_));
  NAND3_X1   g0769(.A1(new_n812_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1   g0770(.A1(new_n227_), .A2(new_n255_), .ZN(new_n820_));
  NAND3_X1   g0771(.A1(new_n131_), .A2(new_n820_), .A3(new_n256_), .ZN(new_n821_));
  NOR4_X1    g0772(.A1(new_n438_), .A2(new_n306_), .A3(new_n360_), .A4(new_n261_), .ZN(new_n822_));
  NAND3_X1   g0773(.A1(new_n710_), .A2(new_n371_), .A3(new_n440_), .ZN(new_n823_));
  OR3_X2     g0774(.A1(new_n822_), .A2(new_n821_), .A3(new_n823_), .Z(new_n824_));
  NOR2_X1    g0775(.A1(new_n175_), .A2(new_n165_), .ZN(new_n825_));
  NOR4_X1    g0776(.A1(new_n825_), .A2(new_n239_), .A3(new_n391_), .A4(new_n526_), .ZN(new_n826_));
  NOR4_X1    g0777(.A1(new_n826_), .A2(new_n387_), .A3(new_n472_), .A4(new_n717_), .ZN(new_n827_));
  NOR3_X1    g0778(.A1(new_n482_), .A2(new_n640_), .A3(new_n271_), .ZN(new_n828_));
  NAND2_X1   g0779(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NOR4_X1    g0780(.A1(new_n819_), .A2(new_n808_), .A3(new_n824_), .A4(new_n829_), .ZN(new_n830_));
  NOR4_X1    g0781(.A1(new_n280_), .A2(new_n336_), .A3(new_n478_), .A4(new_n717_), .ZN(new_n831_));
  NOR4_X1    g0782(.A1(new_n225_), .A2(new_n299_), .A3(new_n150_), .A4(new_n217_), .ZN(new_n832_));
  NOR4_X1    g0783(.A1(new_n526_), .A2(new_n553_), .A3(new_n832_), .A4(new_n327_), .ZN(new_n833_));
  NOR3_X1    g0784(.A1(new_n831_), .A2(new_n799_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1   g0785(.A1(new_n503_), .A2(new_n343_), .ZN(new_n835_));
  NOR2_X1    g0786(.A1(new_n447_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1   g0787(.A1(new_n409_), .A2(new_n196_), .A3(new_n150_), .A4(new_n178_), .ZN(new_n837_));
  NAND4_X1   g0788(.A1(new_n480_), .A2(new_n252_), .A3(new_n211_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1   g0789(.A1(new_n152_), .A2(new_n109_), .ZN(new_n839_));
  NAND3_X1   g0790(.A1(new_n733_), .A2(new_n839_), .A3(new_n425_), .ZN(new_n840_));
  OAI22_X1   g0791(.A1(new_n88_), .A2(new_n260_), .B1(new_n273_), .B2(new_n108_), .ZN(new_n841_));
  AOI22_X1   g0792(.A1(new_n841_), .A2(new_n234_), .B1(new_n130_), .B2(new_n151_), .ZN(new_n842_));
  NOR2_X1    g0793(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1   g0794(.A1(new_n834_), .A2(new_n836_), .A3(new_n843_), .A4(new_n838_), .ZN(new_n844_));
  NOR3_X1    g0795(.A1(new_n435_), .A2(new_n389_), .A3(new_n424_), .ZN(new_n845_));
  NOR2_X1    g0796(.A1(new_n845_), .A2(new_n821_), .ZN(new_n846_));
  NOR4_X1    g0797(.A1(new_n272_), .A2(new_n525_), .A3(new_n501_), .A4(new_n487_), .ZN(new_n847_));
  NOR4_X1    g0798(.A1(new_n165_), .A2(new_n98_), .A3(new_n144_), .A4(new_n221_), .ZN(new_n848_));
  OAI21_X1   g0799(.A1(new_n165_), .A2(new_n150_), .B(new_n245_), .ZN(new_n849_));
  NAND4_X1   g0800(.A1(new_n848_), .A2(new_n849_), .A3(new_n710_), .A4(new_n639_), .ZN(new_n850_));
  NOR2_X1    g0801(.A1(new_n850_), .A2(new_n847_), .ZN(new_n851_));
  OAI21_X1   g0802(.A1(new_n241_), .A2(new_n270_), .B(new_n547_), .ZN(new_n852_));
  NOR4_X1    g0803(.A1(new_n515_), .A2(new_n519_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n853_));
  AOI22_X1   g0804(.A1(new_n109_), .A2(new_n227_), .B1(new_n251_), .B2(new_n428_), .ZN(new_n854_));
  NOR3_X1    g0805(.A1(new_n853_), .A2(new_n852_), .A3(new_n854_), .ZN(new_n855_));
  NOR2_X1    g0806(.A1(new_n191_), .A2(new_n180_), .ZN(new_n856_));
  NOR4_X1    g0807(.A1(new_n612_), .A2(new_n563_), .A3(new_n856_), .A4(new_n638_), .ZN(new_n857_));
  NAND4_X1   g0808(.A1(new_n851_), .A2(new_n855_), .A3(new_n846_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1   g0809(.A1(new_n197_), .A2(new_n433_), .B(new_n171_), .ZN(new_n859_));
  AOI21_X1   g0810(.A1(new_n269_), .A2(new_n423_), .B(new_n171_), .ZN(new_n860_));
  NOR4_X1    g0811(.A1(new_n860_), .A2(new_n859_), .A3(new_n483_), .A4(new_n561_), .ZN(new_n861_));
  OAI22_X1   g0812(.A1(new_n191_), .A2(new_n388_), .B1(new_n323_), .B2(new_n221_), .ZN(new_n862_));
  NOR4_X1    g0813(.A1(new_n632_), .A2(new_n862_), .A3(new_n368_), .A4(new_n517_), .ZN(new_n863_));
  NAND4_X1   g0814(.A1(new_n356_), .A2(new_n726_), .A3(new_n504_), .A4(new_n455_), .ZN(new_n864_));
  NOR4_X1    g0815(.A1(new_n225_), .A2(new_n221_), .A3(new_n88_), .A4(new_n217_), .ZN(new_n865_));
  NOR3_X1    g0816(.A1(new_n595_), .A2(new_n594_), .A3(new_n865_), .ZN(new_n866_));
  NAND4_X1   g0817(.A1(new_n863_), .A2(new_n861_), .A3(new_n864_), .A4(new_n866_), .ZN(new_n867_));
  NOR3_X1    g0818(.A1(new_n858_), .A2(new_n844_), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1   g0819(.A1(new_n227_), .A2(new_n374_), .B(new_n295_), .ZN(new_n869_));
  OAI21_X1   g0820(.A1(new_n292_), .A2(new_n188_), .B(new_n440_), .ZN(new_n870_));
  NOR4_X1    g0821(.A1(new_n870_), .A2(new_n417_), .A3(new_n869_), .A4(new_n593_), .ZN(new_n871_));
  NOR3_X1    g0822(.A1(new_n423_), .A2(new_n98_), .A3(new_n286_), .ZN(new_n872_));
  NOR3_X1    g0823(.A1(new_n337_), .A2(new_n262_), .A3(new_n347_), .ZN(new_n873_));
  NOR4_X1    g0824(.A1(new_n873_), .A2(new_n872_), .A3(new_n324_), .A4(new_n487_), .ZN(new_n874_));
  NAND4_X1   g0825(.A1(new_n548_), .A2(new_n150_), .A3(new_n409_), .A4(new_n196_), .ZN(new_n875_));
  NAND3_X1   g0826(.A1(new_n146_), .A2(new_n875_), .A3(new_n363_), .ZN(new_n876_));
  NOR2_X1    g0827(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NOR4_X1    g0828(.A1(new_n262_), .A2(new_n88_), .A3(new_n221_), .A4(new_n217_), .ZN(new_n878_));
  NOR4_X1    g0829(.A1(new_n878_), .A2(new_n471_), .A3(new_n399_), .A4(new_n300_), .ZN(new_n879_));
  NAND3_X1   g0830(.A1(new_n442_), .A2(new_n291_), .A3(new_n711_), .ZN(new_n880_));
  NOR2_X1    g0831(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1   g0832(.A1(new_n877_), .A2(new_n881_), .A3(new_n871_), .ZN(new_n882_));
  NAND3_X1   g0833(.A1(new_n152_), .A2(new_n609_), .A3(new_n170_), .ZN(new_n883_));
  AOI21_X1   g0834(.A1(new_n152_), .A2(new_n88_), .B(new_n370_), .ZN(new_n884_));
  NOR4_X1    g0835(.A1(new_n884_), .A2(new_n883_), .A3(new_n394_), .A4(new_n488_), .ZN(new_n885_));
  OAI22_X1   g0836(.A1(new_n175_), .A2(new_n208_), .B1(new_n279_), .B2(new_n265_), .ZN(new_n886_));
  OAI22_X1   g0837(.A1(new_n292_), .A2(new_n175_), .B1(new_n171_), .B2(new_n388_), .ZN(new_n887_));
  NOR4_X1    g0838(.A1(new_n271_), .A2(new_n854_), .A3(new_n887_), .A4(new_n886_), .ZN(new_n888_));
  AOI21_X1   g0839(.A1(new_n197_), .A2(new_n433_), .B(new_n188_), .ZN(new_n889_));
  NOR3_X1    g0840(.A1(new_n197_), .A2(new_n150_), .A3(new_n221_), .ZN(new_n890_));
  NOR4_X1    g0841(.A1(new_n889_), .A2(new_n890_), .A3(new_n500_), .A4(new_n478_), .ZN(new_n891_));
  NAND4_X1   g0842(.A1(new_n888_), .A2(new_n457_), .A3(new_n885_), .A4(new_n891_), .ZN(new_n892_));
  NAND2_X1   g0843(.A1(new_n287_), .A2(new_n428_), .ZN(new_n893_));
  NAND4_X1   g0844(.A1(new_n719_), .A2(new_n468_), .A3(new_n408_), .A4(new_n893_), .ZN(new_n894_));
  NOR4_X1    g0845(.A1(new_n402_), .A2(new_n391_), .A3(new_n461_), .A4(new_n524_), .ZN(new_n895_));
  NOR3_X1    g0846(.A1(new_n895_), .A2(new_n805_), .A3(new_n762_), .ZN(new_n896_));
  NOR4_X1    g0847(.A1(new_n274_), .A2(new_n526_), .A3(new_n472_), .A4(new_n603_), .ZN(new_n897_));
  OAI22_X1   g0848(.A1(new_n197_), .A2(new_n195_), .B1(new_n237_), .B2(new_n423_), .ZN(new_n898_));
  NAND2_X1   g0849(.A1(new_n130_), .A2(new_n251_), .ZN(new_n899_));
  NAND3_X1   g0850(.A1(new_n899_), .A2(new_n641_), .A3(new_n232_), .ZN(new_n900_));
  NOR3_X1    g0851(.A1(new_n900_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n901_));
  NAND3_X1   g0852(.A1(new_n901_), .A2(new_n896_), .A3(new_n894_), .ZN(new_n902_));
  NOR3_X1    g0853(.A1(new_n892_), .A2(new_n902_), .A3(new_n882_), .ZN(new_n903_));
  NOR2_X1    g0854(.A1(new_n868_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1    g0855(.A1(new_n904_), .A2(new_n830_), .ZN(new_n905_));
  AOI22_X1   g0856(.A1(new_n141_), .A2(new_n222_), .B1(new_n224_), .B2(new_n219_), .ZN(new_n906_));
  AOI21_X1   g0857(.A1(new_n433_), .A2(new_n509_), .B(new_n265_), .ZN(new_n907_));
  AOI22_X1   g0858(.A1(new_n130_), .A2(new_n255_), .B1(new_n379_), .B2(new_n187_), .ZN(new_n908_));
  NAND4_X1   g0859(.A1(new_n908_), .A2(new_n906_), .A3(new_n907_), .A4(new_n445_), .ZN(new_n909_));
  NAND4_X1   g0860(.A1(new_n412_), .A2(new_n310_), .A3(new_n380_), .A4(new_n550_), .ZN(new_n910_));
  NOR3_X1    g0861(.A1(new_n438_), .A2(new_n620_), .A3(new_n534_), .ZN(new_n911_));
  NAND2_X1   g0862(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1   g0863(.A1(new_n367_), .A2(new_n150_), .A3(new_n409_), .ZN(new_n913_));
  NAND4_X1   g0864(.A1(new_n288_), .A2(new_n490_), .A3(new_n913_), .A4(new_n547_), .ZN(new_n914_));
  NOR3_X1    g0865(.A1(new_n280_), .A2(new_n865_), .A3(new_n643_), .ZN(new_n915_));
  NAND2_X1   g0866(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NOR3_X1    g0867(.A1(new_n912_), .A2(new_n916_), .A3(new_n909_), .ZN(new_n917_));
  AOI22_X1   g0868(.A1(new_n226_), .A2(new_n407_), .B1(new_n109_), .B2(new_n318_), .ZN(new_n918_));
  NAND4_X1   g0869(.A1(new_n918_), .A2(new_n203_), .A3(new_n455_), .A4(new_n321_), .ZN(new_n919_));
  NOR3_X1    g0870(.A1(new_n98_), .A2(new_n144_), .A3(new_n150_), .ZN(new_n920_));
  AOI22_X1   g0871(.A1(new_n234_), .A2(new_n109_), .B1(new_n920_), .B2(new_n428_), .ZN(new_n921_));
  OAI22_X1   g0872(.A1(new_n240_), .A2(new_n241_), .B1(new_n433_), .B2(new_n191_), .ZN(new_n922_));
  AOI22_X1   g0873(.A1(new_n151_), .A2(new_n141_), .B1(new_n318_), .B2(new_n295_), .ZN(new_n923_));
  AOI22_X1   g0874(.A1(new_n130_), .A2(new_n151_), .B1(new_n224_), .B2(new_n367_), .ZN(new_n924_));
  NAND4_X1   g0875(.A1(new_n921_), .A2(new_n922_), .A3(new_n924_), .A4(new_n923_), .ZN(new_n925_));
  NAND4_X1   g0876(.A1(new_n409_), .A2(new_n150_), .A3(new_n179_), .A4(new_n231_), .ZN(new_n926_));
  NAND4_X1   g0877(.A1(new_n497_), .A2(new_n296_), .A3(new_n926_), .A4(new_n646_), .ZN(new_n927_));
  NOR4_X1    g0878(.A1(new_n925_), .A2(new_n919_), .A3(new_n850_), .A4(new_n927_), .ZN(new_n928_));
  NAND4_X1   g0879(.A1(new_n210_), .A2(new_n174_), .A3(new_n196_), .A4(new_n144_), .ZN(new_n929_));
  NAND4_X1   g0880(.A1(new_n210_), .A2(new_n243_), .A3(new_n190_), .A4(new_n207_), .ZN(new_n930_));
  NAND4_X1   g0881(.A1(new_n210_), .A2(new_n196_), .A3(new_n187_), .A4(new_n88_), .ZN(new_n931_));
  NAND4_X1   g0882(.A1(new_n929_), .A2(new_n931_), .A3(new_n930_), .A4(new_n458_), .ZN(new_n932_));
  AOI22_X1   g0883(.A1(new_n226_), .A2(new_n145_), .B1(new_n222_), .B2(new_n233_), .ZN(new_n933_));
  AOI22_X1   g0884(.A1(new_n130_), .A2(new_n251_), .B1(new_n285_), .B2(new_n151_), .ZN(new_n934_));
  NAND4_X1   g0885(.A1(new_n932_), .A2(new_n934_), .A3(new_n933_), .A4(new_n641_), .ZN(new_n935_));
  NOR3_X1    g0886(.A1(new_n935_), .A2(new_n351_), .A3(new_n340_), .ZN(new_n936_));
  NAND3_X1   g0887(.A1(new_n917_), .A2(new_n928_), .A3(new_n936_), .ZN(new_n937_));
  OAI21_X1   g0888(.A1(new_n57_), .A2(new_n60_), .B(new_n80_), .ZN(new_n938_));
  XNOR2_X1   g0889(.A1(new_n938_), .A2(\a[6] ), .ZN(new_n939_));
  NAND2_X1   g0890(.A1(new_n627_), .A2(new_n939_), .ZN(new_n940_));
  XOR2_X1    g0891(.A1(new_n940_), .A2(new_n937_), .Z(new_n941_));
  XOR2_X1    g0892(.A1(new_n941_), .A2(new_n905_), .Z(new_n942_));
  INV_X1     g0893(.I(new_n62_), .ZN(new_n943_));
  NOR2_X1    g0894(.A1(new_n628_), .A2(new_n943_), .ZN(new_n944_));
  XOR2_X1    g0895(.A1(new_n944_), .A2(new_n903_), .Z(new_n945_));
  NAND2_X1   g0896(.A1(new_n944_), .A2(new_n903_), .ZN(new_n946_));
  NOR2_X1    g0897(.A1(new_n484_), .A2(new_n246_), .ZN(new_n947_));
  NAND4_X1   g0898(.A1(new_n893_), .A2(new_n442_), .A3(new_n926_), .A4(new_n774_), .ZN(new_n948_));
  NAND4_X1   g0899(.A1(new_n210_), .A2(new_n196_), .A3(new_n187_), .A4(new_n150_), .ZN(new_n949_));
  NAND4_X1   g0900(.A1(new_n196_), .A2(new_n187_), .A3(new_n88_), .A4(new_n178_), .ZN(new_n950_));
  NAND4_X1   g0901(.A1(new_n931_), .A2(new_n949_), .A3(new_n950_), .A4(new_n619_), .ZN(new_n951_));
  NAND3_X1   g0902(.A1(new_n948_), .A2(new_n947_), .A3(new_n951_), .ZN(new_n952_));
  NAND4_X1   g0903(.A1(new_n403_), .A2(new_n408_), .A3(new_n445_), .A4(new_n446_), .ZN(new_n953_));
  NOR3_X1    g0904(.A1(new_n192_), .A2(new_n239_), .A3(new_n263_), .ZN(new_n954_));
  AOI22_X1   g0905(.A1(new_n409_), .A2(new_n150_), .B1(new_n174_), .B2(new_n144_), .ZN(new_n955_));
  OAI22_X1   g0906(.A1(new_n955_), .A2(new_n269_), .B1(new_n292_), .B2(new_n175_), .ZN(new_n956_));
  NAND3_X1   g0907(.A1(new_n954_), .A2(new_n838_), .A3(new_n956_), .ZN(new_n957_));
  NOR3_X1    g0908(.A1(new_n957_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n958_));
  AOI22_X1   g0909(.A1(new_n130_), .A2(new_n109_), .B1(new_n141_), .B2(new_n255_), .ZN(new_n959_));
  NAND3_X1   g0910(.A1(new_n560_), .A2(new_n820_), .A3(new_n959_), .ZN(new_n960_));
  NAND4_X1   g0911(.A1(new_n418_), .A2(new_n463_), .A3(new_n316_), .A4(new_n550_), .ZN(new_n961_));
  NOR2_X1    g0912(.A1(new_n883_), .A2(new_n394_), .ZN(new_n962_));
  NAND3_X1   g0913(.A1(new_n558_), .A2(new_n548_), .A3(new_n88_), .ZN(new_n963_));
  AOI21_X1   g0914(.A1(new_n963_), .A2(new_n245_), .B(new_n488_), .ZN(new_n964_));
  NAND3_X1   g0915(.A1(new_n961_), .A2(new_n962_), .A3(new_n964_), .ZN(new_n965_));
  NAND4_X1   g0916(.A1(new_n549_), .A2(new_n481_), .A3(new_n539_), .A4(new_n440_), .ZN(new_n966_));
  NAND3_X1   g0917(.A1(new_n966_), .A2(new_n768_), .A3(new_n922_), .ZN(new_n967_));
  AOI22_X1   g0918(.A1(new_n151_), .A2(new_n233_), .B1(new_n219_), .B2(new_n255_), .ZN(new_n968_));
  NAND4_X1   g0919(.A1(new_n968_), .A2(new_n309_), .A3(new_n357_), .A4(new_n330_), .ZN(new_n969_));
  NOR4_X1    g0920(.A1(new_n965_), .A2(new_n967_), .A3(new_n960_), .A4(new_n969_), .ZN(new_n970_));
  NAND3_X1   g0921(.A1(new_n210_), .A2(new_n88_), .A3(new_n207_), .ZN(new_n971_));
  AOI21_X1   g0922(.A1(new_n971_), .A2(new_n388_), .B(new_n221_), .ZN(new_n972_));
  NAND4_X1   g0923(.A1(new_n508_), .A2(new_n972_), .A3(new_n729_), .A4(new_n429_), .ZN(new_n973_));
  NOR2_X1    g0924(.A1(new_n334_), .A2(new_n171_), .ZN(new_n974_));
  NOR4_X1    g0925(.A1(new_n974_), .A2(new_n377_), .A3(new_n584_), .A4(new_n266_), .ZN(new_n975_));
  NAND3_X1   g0926(.A1(new_n545_), .A2(new_n291_), .A3(new_n419_), .ZN(new_n976_));
  NOR4_X1    g0927(.A1(new_n973_), .A2(new_n236_), .A3(new_n975_), .A4(new_n976_), .ZN(new_n977_));
  NAND3_X1   g0928(.A1(new_n970_), .A2(new_n958_), .A3(new_n977_), .ZN(new_n978_));
  NOR2_X1    g0929(.A1(new_n978_), .A2(new_n903_), .ZN(new_n979_));
  NOR2_X1    g0930(.A1(new_n868_), .A2(new_n937_), .ZN(new_n980_));
  NOR2_X1    g0931(.A1(new_n980_), .A2(new_n979_), .ZN(new_n981_));
  NOR2_X1    g0932(.A1(new_n868_), .A2(new_n903_), .ZN(new_n982_));
  XOR2_X1    g0933(.A1(new_n982_), .A2(new_n830_), .Z(new_n983_));
  NAND2_X1   g0934(.A1(new_n830_), .A2(new_n658_), .ZN(new_n984_));
  INV_X1     g0935(.I(new_n808_), .ZN(new_n985_));
  NAND2_X1   g0936(.A1(new_n816_), .A2(new_n818_), .ZN(new_n986_));
  NOR4_X1    g0937(.A1(new_n829_), .A2(new_n986_), .A3(new_n811_), .A4(new_n824_), .ZN(new_n987_));
  NAND2_X1   g0938(.A1(new_n987_), .A2(new_n985_), .ZN(new_n988_));
  NAND2_X1   g0939(.A1(new_n988_), .A2(new_n659_), .ZN(new_n989_));
  AND2_X2    g0940(.A1(new_n989_), .A2(new_n984_), .Z(new_n990_));
  AOI21_X1   g0941(.A1(new_n990_), .A2(new_n981_), .B(new_n983_), .ZN(new_n991_));
  OAI21_X1   g0942(.A1(new_n945_), .A2(new_n991_), .B(new_n946_), .ZN(new_n992_));
  INV_X1     g0943(.I(new_n992_), .ZN(new_n993_));
  NOR2_X1    g0944(.A1(new_n993_), .A2(new_n942_), .ZN(new_n994_));
  INV_X1     g0945(.I(new_n942_), .ZN(new_n995_));
  NOR2_X1    g0946(.A1(new_n995_), .A2(new_n992_), .ZN(new_n996_));
  NOR2_X1    g0947(.A1(new_n996_), .A2(new_n994_), .ZN(new_n997_));
  NOR2_X1    g0948(.A1(new_n997_), .A2(new_n798_), .ZN(new_n998_));
  XOR2_X1    g0949(.A1(new_n942_), .A2(new_n992_), .Z(new_n999_));
  NOR2_X1    g0950(.A1(new_n999_), .A2(new_n797_), .ZN(new_n1000_));
  NOR2_X1    g0951(.A1(new_n998_), .A2(new_n1000_), .ZN(new_n1001_));
  NOR3_X1    g0952(.A1(new_n676_), .A2(new_n671_), .A3(new_n939_), .ZN(new_n1002_));
  INV_X1     g0953(.I(new_n1002_), .ZN(new_n1003_));
  NOR2_X1    g0954(.A1(new_n679_), .A2(new_n943_), .ZN(new_n1004_));
  INV_X1     g0955(.I(new_n682_), .ZN(new_n1005_));
  NOR2_X1    g0956(.A1(new_n1005_), .A2(new_n62_), .ZN(new_n1006_));
  NOR3_X1    g0957(.A1(new_n1003_), .A2(new_n1004_), .A3(new_n1006_), .ZN(new_n1007_));
  INV_X1     g0958(.I(new_n1007_), .ZN(new_n1008_));
  NOR2_X1    g0959(.A1(new_n239_), .A2(new_n263_), .ZN(new_n1009_));
  NAND4_X1   g0960(.A1(new_n1009_), .A2(new_n564_), .A3(new_n203_), .A4(new_n445_), .ZN(new_n1010_));
  NAND2_X1   g0961(.A1(new_n755_), .A2(new_n481_), .ZN(new_n1011_));
  NAND4_X1   g0962(.A1(new_n511_), .A2(new_n528_), .A3(new_n448_), .A4(new_n931_), .ZN(new_n1012_));
  NOR4_X1    g0963(.A1(new_n1010_), .A2(new_n1012_), .A3(new_n474_), .A4(new_n1011_), .ZN(new_n1013_));
  INV_X1     g0964(.I(new_n1013_), .ZN(new_n1014_));
  NAND4_X1   g0965(.A1(new_n639_), .A2(new_n532_), .A3(new_n455_), .A4(new_n344_), .ZN(new_n1015_));
  NOR2_X1    g0966(.A1(new_n535_), .A2(new_n561_), .ZN(new_n1016_));
  NAND4_X1   g0967(.A1(new_n1015_), .A2(new_n213_), .A3(new_n1016_), .A4(new_n837_), .ZN(new_n1017_));
  OR2_X2     g0968(.A1(new_n1017_), .A2(new_n599_), .Z(new_n1018_));
  NAND2_X1   g0969(.A1(new_n234_), .A2(new_n109_), .ZN(new_n1019_));
  NAND4_X1   g0970(.A1(new_n809_), .A2(new_n1019_), .A3(new_n469_), .A4(new_n284_), .ZN(new_n1020_));
  NOR2_X1    g0971(.A1(new_n269_), .A2(new_n237_), .ZN(new_n1021_));
  NOR3_X1    g0972(.A1(new_n483_), .A2(new_n1021_), .A3(new_n878_), .ZN(new_n1022_));
  NAND4_X1   g0973(.A1(new_n1020_), .A2(new_n252_), .A3(new_n1022_), .A4(new_n363_), .ZN(new_n1023_));
  NOR4_X1    g0974(.A1(new_n438_), .A2(new_n278_), .A3(new_n360_), .A4(new_n478_), .ZN(new_n1024_));
  NOR4_X1    g0975(.A1(new_n246_), .A2(new_n588_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n1025_));
  OR3_X2     g0976(.A1(new_n1024_), .A2(new_n1025_), .A3(new_n764_), .Z(new_n1026_));
  NOR4_X1    g0977(.A1(new_n1014_), .A2(new_n1018_), .A3(new_n1023_), .A4(new_n1026_), .ZN(new_n1027_));
  AOI21_X1   g0978(.A1(new_n1027_), .A2(new_n658_), .B(new_n903_), .ZN(new_n1028_));
  INV_X1     g0979(.I(new_n1028_), .ZN(new_n1029_));
  NOR2_X1    g0980(.A1(new_n978_), .A2(new_n937_), .ZN(new_n1030_));
  AOI21_X1   g0981(.A1(new_n830_), .A2(new_n1030_), .B(new_n904_), .ZN(new_n1031_));
  INV_X1     g0982(.I(new_n1031_), .ZN(new_n1032_));
  AOI21_X1   g0983(.A1(new_n988_), .A2(new_n904_), .B(new_n1030_), .ZN(new_n1033_));
  INV_X1     g0984(.I(new_n1033_), .ZN(new_n1034_));
  OAI21_X1   g0985(.A1(new_n980_), .A2(new_n979_), .B(new_n830_), .ZN(new_n1035_));
  NAND2_X1   g0986(.A1(new_n1035_), .A2(new_n678_), .ZN(new_n1036_));
  NOR2_X1    g0987(.A1(new_n981_), .A2(new_n830_), .ZN(new_n1037_));
  OAI21_X1   g0988(.A1(new_n678_), .A2(new_n1037_), .B(new_n1036_), .ZN(new_n1038_));
  NOR4_X1    g0989(.A1(new_n1038_), .A2(new_n581_), .A3(new_n1032_), .A4(new_n1034_), .ZN(new_n1039_));
  XOR2_X1    g0990(.A1(new_n1039_), .A2(new_n1029_), .Z(new_n1040_));
  NAND2_X1   g0991(.A1(new_n627_), .A2(new_n67_), .ZN(new_n1041_));
  AOI21_X1   g0992(.A1(new_n1028_), .A2(new_n1041_), .B(new_n1040_), .ZN(new_n1042_));
  NAND2_X1   g0993(.A1(new_n1042_), .A2(new_n1008_), .ZN(new_n1043_));
  INV_X1     g0994(.I(new_n568_), .ZN(new_n1044_));
  NOR2_X1    g0995(.A1(new_n567_), .A2(new_n494_), .ZN(new_n1045_));
  NOR2_X1    g0996(.A1(new_n1044_), .A2(new_n1045_), .ZN(new_n1046_));
  NAND2_X1   g0997(.A1(new_n1046_), .A2(new_n569_), .ZN(new_n1047_));
  INV_X1     g0998(.I(\a[7] ), .ZN(new_n1048_));
  NOR2_X1    g0999(.A1(new_n74_), .A2(new_n51_), .ZN(new_n1049_));
  INV_X1     g1000(.I(new_n1049_), .ZN(new_n1050_));
  NAND2_X1   g1001(.A1(new_n1050_), .A2(new_n80_), .ZN(new_n1051_));
  NOR2_X1    g1002(.A1(new_n1048_), .A2(\a[22] ), .ZN(new_n1052_));
  AOI22_X1   g1003(.A1(new_n1051_), .A2(new_n1048_), .B1(new_n1050_), .B2(new_n1052_), .ZN(new_n1053_));
  NOR2_X1    g1004(.A1(new_n1047_), .A2(new_n1053_), .ZN(new_n1054_));
  XOR2_X1    g1005(.A1(new_n567_), .A2(new_n415_), .Z(new_n1055_));
  XOR2_X1    g1006(.A1(new_n494_), .A2(new_n939_), .Z(new_n1056_));
  NOR2_X1    g1007(.A1(new_n1055_), .A2(new_n1056_), .ZN(new_n1057_));
  INV_X1     g1008(.I(new_n1045_), .ZN(new_n1058_));
  NAND2_X1   g1009(.A1(new_n1058_), .A2(new_n568_), .ZN(new_n1059_));
  NOR2_X1    g1010(.A1(new_n1045_), .A2(new_n416_), .ZN(new_n1060_));
  NOR2_X1    g1011(.A1(new_n1059_), .A2(new_n1060_), .ZN(new_n1061_));
  INV_X1     g1012(.I(new_n1053_), .ZN(new_n1062_));
  NAND2_X1   g1013(.A1(new_n690_), .A2(new_n1062_), .ZN(new_n1063_));
  NOR4_X1    g1014(.A1(new_n1054_), .A2(new_n1057_), .A3(new_n1061_), .A4(new_n1063_), .ZN(new_n1064_));
  INV_X1     g1015(.I(new_n723_), .ZN(new_n1065_));
  NOR4_X1    g1016(.A1(new_n1065_), .A2(new_n736_), .A3(new_n743_), .A4(new_n750_), .ZN(new_n1066_));
  NAND3_X1   g1017(.A1(new_n908_), .A2(new_n907_), .A3(new_n445_), .ZN(new_n1067_));
  NOR2_X1    g1018(.A1(new_n459_), .A2(new_n543_), .ZN(new_n1068_));
  NAND2_X1   g1019(.A1(new_n771_), .A2(new_n146_), .ZN(new_n1069_));
  OR3_X2     g1020(.A1(new_n1068_), .A2(new_n1067_), .A3(new_n1069_), .Z(new_n1070_));
  NOR4_X1    g1021(.A1(new_n817_), .A2(new_n242_), .A3(new_n305_), .A4(new_n519_), .ZN(new_n1071_));
  NAND3_X1   g1022(.A1(new_n302_), .A2(new_n131_), .A3(new_n926_), .ZN(new_n1072_));
  INV_X1     g1023(.I(new_n473_), .ZN(new_n1073_));
  NAND4_X1   g1024(.A1(new_n1073_), .A2(new_n316_), .A3(new_n344_), .A4(new_n550_), .ZN(new_n1074_));
  NAND3_X1   g1025(.A1(new_n1071_), .A2(new_n1072_), .A3(new_n1074_), .ZN(new_n1075_));
  NOR2_X1    g1026(.A1(new_n1075_), .A2(new_n1070_), .ZN(new_n1076_));
  NOR2_X1    g1027(.A1(new_n372_), .A2(new_n738_), .ZN(new_n1077_));
  NAND4_X1   g1028(.A1(new_n1077_), .A2(new_n613_), .A3(new_n312_), .A4(new_n343_), .ZN(new_n1078_));
  NAND2_X1   g1029(.A1(new_n469_), .A2(new_n710_), .ZN(new_n1079_));
  NOR3_X1    g1030(.A1(new_n496_), .A2(new_n1079_), .A3(new_n889_), .ZN(new_n1080_));
  NOR4_X1    g1031(.A1(new_n204_), .A2(new_n336_), .A3(new_n517_), .A4(new_n878_), .ZN(new_n1081_));
  NAND2_X1   g1032(.A1(new_n1080_), .A2(new_n1081_), .ZN(new_n1082_));
  INV_X1     g1033(.I(new_n426_), .ZN(new_n1083_));
  NAND4_X1   g1034(.A1(new_n1083_), .A2(new_n310_), .A3(new_n330_), .A4(new_n363_), .ZN(new_n1084_));
  NAND2_X1   g1035(.A1(new_n412_), .A2(new_n397_), .ZN(new_n1085_));
  INV_X1     g1036(.I(new_n1085_), .ZN(new_n1086_));
  NAND3_X1   g1037(.A1(new_n1086_), .A2(new_n1084_), .A3(new_n954_), .ZN(new_n1087_));
  NOR3_X1    g1038(.A1(new_n483_), .A2(new_n369_), .A3(new_n525_), .ZN(new_n1088_));
  NOR2_X1    g1039(.A1(new_n208_), .A2(new_n188_), .ZN(new_n1089_));
  NOR3_X1    g1040(.A1(new_n499_), .A2(new_n150_), .A3(new_n221_), .ZN(new_n1090_));
  NOR2_X1    g1041(.A1(new_n171_), .A2(new_n423_), .ZN(new_n1091_));
  NOR4_X1    g1042(.A1(new_n1090_), .A2(new_n250_), .A3(new_n434_), .A4(new_n1091_), .ZN(new_n1092_));
  NOR3_X1    g1043(.A1(new_n1092_), .A2(new_n1089_), .A3(new_n472_), .ZN(new_n1093_));
  NAND2_X1   g1044(.A1(new_n1093_), .A2(new_n1088_), .ZN(new_n1094_));
  NOR4_X1    g1045(.A1(new_n1094_), .A2(new_n1082_), .A3(new_n1078_), .A4(new_n1087_), .ZN(new_n1095_));
  NAND2_X1   g1046(.A1(new_n1095_), .A2(new_n1076_), .ZN(new_n1096_));
  XOR2_X1    g1047(.A1(new_n1096_), .A2(new_n988_), .Z(new_n1097_));
  NAND2_X1   g1048(.A1(new_n1097_), .A2(new_n1066_), .ZN(new_n1098_));
  XOR2_X1    g1049(.A1(new_n1096_), .A2(new_n830_), .Z(new_n1099_));
  NOR2_X1    g1050(.A1(new_n1099_), .A2(new_n1066_), .ZN(new_n1100_));
  NOR2_X1    g1051(.A1(new_n1100_), .A2(new_n576_), .ZN(new_n1101_));
  AOI21_X1   g1052(.A1(new_n576_), .A2(new_n1098_), .B(new_n1101_), .ZN(new_n1102_));
  AOI21_X1   g1053(.A1(new_n571_), .A2(new_n80_), .B(\a[10] ), .ZN(new_n1103_));
  NAND3_X1   g1054(.A1(new_n571_), .A2(\a[10] ), .A3(new_n80_), .ZN(new_n1104_));
  INV_X1     g1055(.I(new_n1104_), .ZN(new_n1105_));
  NOR2_X1    g1056(.A1(new_n1105_), .A2(new_n1103_), .ZN(new_n1106_));
  NAND2_X1   g1057(.A1(new_n1096_), .A2(new_n988_), .ZN(new_n1107_));
  AND2_X2    g1058(.A1(new_n1095_), .A2(new_n1076_), .Z(new_n1108_));
  NAND2_X1   g1059(.A1(new_n1108_), .A2(new_n830_), .ZN(new_n1109_));
  OAI21_X1   g1060(.A1(new_n1109_), .A2(new_n752_), .B(new_n1107_), .ZN(new_n1110_));
  NOR2_X1    g1061(.A1(new_n1110_), .A2(new_n1106_), .ZN(new_n1111_));
  NOR2_X1    g1062(.A1(new_n1096_), .A2(new_n988_), .ZN(new_n1112_));
  NOR2_X1    g1063(.A1(new_n1107_), .A2(new_n1066_), .ZN(new_n1113_));
  NOR2_X1    g1064(.A1(new_n1113_), .A2(new_n1112_), .ZN(new_n1114_));
  AOI21_X1   g1065(.A1(new_n1106_), .A2(new_n1114_), .B(new_n1111_), .ZN(new_n1115_));
  NAND2_X1   g1066(.A1(new_n1102_), .A2(new_n1115_), .ZN(new_n1116_));
  INV_X1     g1067(.I(new_n1116_), .ZN(new_n1117_));
  NOR2_X1    g1068(.A1(new_n1117_), .A2(new_n1064_), .ZN(new_n1118_));
  NAND2_X1   g1069(.A1(new_n792_), .A2(new_n780_), .ZN(new_n1119_));
  INV_X1     g1070(.I(new_n494_), .ZN(new_n1120_));
  NAND2_X1   g1071(.A1(new_n783_), .A2(new_n1120_), .ZN(new_n1121_));
  NAND2_X1   g1072(.A1(new_n792_), .A2(new_n1121_), .ZN(new_n1122_));
  OR2_X2     g1073(.A1(\a[7] ), .A2(\a[8] ), .Z(new_n1123_));
  AOI21_X1   g1074(.A1(new_n1050_), .A2(new_n1123_), .B(\a[22] ), .ZN(new_n1124_));
  XNOR2_X1   g1075(.A1(new_n1124_), .A2(\a[9] ), .ZN(new_n1125_));
  INV_X1     g1076(.I(new_n1125_), .ZN(new_n1126_));
  NAND3_X1   g1077(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n1126_), .ZN(new_n1127_));
  AOI21_X1   g1078(.A1(new_n1050_), .A2(\a[7] ), .B(\a[22] ), .ZN(new_n1128_));
  NOR2_X1    g1079(.A1(new_n1128_), .A2(\a[8] ), .ZN(new_n1129_));
  NAND2_X1   g1080(.A1(new_n1128_), .A2(\a[8] ), .ZN(new_n1130_));
  INV_X1     g1081(.I(new_n1130_), .ZN(new_n1131_));
  NOR2_X1    g1082(.A1(new_n1131_), .A2(new_n1129_), .ZN(new_n1132_));
  NOR2_X1    g1083(.A1(new_n793_), .A2(new_n1132_), .ZN(new_n1133_));
  INV_X1     g1084(.I(new_n1132_), .ZN(new_n1134_));
  NOR2_X1    g1085(.A1(new_n795_), .A2(new_n1134_), .ZN(new_n1135_));
  NOR3_X1    g1086(.A1(new_n1127_), .A2(new_n1133_), .A3(new_n1135_), .ZN(new_n1136_));
  INV_X1     g1087(.I(new_n1136_), .ZN(new_n1137_));
  NAND2_X1   g1088(.A1(new_n1117_), .A2(new_n1064_), .ZN(new_n1138_));
  AOI21_X1   g1089(.A1(new_n1137_), .A2(new_n1138_), .B(new_n1118_), .ZN(new_n1139_));
  NOR2_X1    g1090(.A1(new_n1042_), .A2(new_n1008_), .ZN(new_n1140_));
  OAI21_X1   g1091(.A1(new_n1139_), .A2(new_n1140_), .B(new_n1043_), .ZN(new_n1141_));
  INV_X1     g1092(.I(new_n1141_), .ZN(new_n1142_));
  XOR2_X1    g1093(.A1(new_n945_), .A2(new_n991_), .Z(new_n1143_));
  INV_X1     g1094(.I(new_n1143_), .ZN(new_n1144_));
  INV_X1     g1095(.I(new_n1047_), .ZN(new_n1145_));
  NAND2_X1   g1096(.A1(new_n1059_), .A2(new_n569_), .ZN(new_n1146_));
  NAND2_X1   g1097(.A1(new_n1146_), .A2(new_n1134_), .ZN(new_n1147_));
  NOR2_X1    g1098(.A1(new_n1046_), .A2(new_n1060_), .ZN(new_n1148_));
  OAI21_X1   g1099(.A1(new_n1134_), .A2(new_n1148_), .B(new_n1147_), .ZN(new_n1149_));
  NOR4_X1    g1100(.A1(new_n1149_), .A2(new_n1145_), .A3(new_n1061_), .A4(new_n1125_), .ZN(new_n1150_));
  NAND3_X1   g1101(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n576_), .ZN(new_n1151_));
  NOR2_X1    g1102(.A1(new_n793_), .A2(new_n1106_), .ZN(new_n1152_));
  INV_X1     g1103(.I(new_n1106_), .ZN(new_n1153_));
  NOR2_X1    g1104(.A1(new_n795_), .A2(new_n1153_), .ZN(new_n1154_));
  NOR3_X1    g1105(.A1(new_n1151_), .A2(new_n1152_), .A3(new_n1154_), .ZN(new_n1155_));
  NOR2_X1    g1106(.A1(new_n1100_), .A2(new_n678_), .ZN(new_n1156_));
  AOI21_X1   g1107(.A1(new_n678_), .A2(new_n1098_), .B(new_n1156_), .ZN(new_n1157_));
  NOR2_X1    g1108(.A1(new_n1110_), .A2(new_n581_), .ZN(new_n1158_));
  AOI21_X1   g1109(.A1(new_n581_), .A2(new_n1114_), .B(new_n1158_), .ZN(new_n1159_));
  NAND2_X1   g1110(.A1(new_n1157_), .A2(new_n1159_), .ZN(new_n1160_));
  XNOR2_X1   g1111(.A1(new_n1160_), .A2(new_n1155_), .ZN(new_n1161_));
  NAND2_X1   g1112(.A1(new_n1161_), .A2(new_n1150_), .ZN(new_n1162_));
  INV_X1     g1113(.I(new_n1150_), .ZN(new_n1163_));
  AOI21_X1   g1114(.A1(new_n1157_), .A2(new_n1159_), .B(new_n1155_), .ZN(new_n1164_));
  NOR4_X1    g1115(.A1(new_n1160_), .A2(new_n1151_), .A3(new_n1152_), .A4(new_n1154_), .ZN(new_n1165_));
  OAI21_X1   g1116(.A1(new_n1164_), .A2(new_n1165_), .B(new_n1163_), .ZN(new_n1166_));
  NAND2_X1   g1117(.A1(new_n1162_), .A2(new_n1166_), .ZN(new_n1167_));
  OAI21_X1   g1118(.A1(new_n1141_), .A2(new_n1144_), .B(new_n1167_), .ZN(new_n1168_));
  OAI21_X1   g1119(.A1(new_n1142_), .A2(new_n1143_), .B(new_n1168_), .ZN(new_n1169_));
  NAND2_X1   g1120(.A1(new_n1169_), .A2(new_n1001_), .ZN(new_n1170_));
  INV_X1     g1121(.I(new_n939_), .ZN(new_n1171_));
  NOR2_X1    g1122(.A1(new_n679_), .A2(new_n1171_), .ZN(new_n1172_));
  NOR2_X1    g1123(.A1(new_n1005_), .A2(new_n939_), .ZN(new_n1173_));
  NOR2_X1    g1124(.A1(new_n1173_), .A2(new_n1172_), .ZN(new_n1174_));
  AND4_X2    g1125(.A1(new_n696_), .A2(new_n1174_), .A3(new_n675_), .A4(new_n1062_), .Z(new_n1175_));
  INV_X1     g1126(.I(new_n56_), .ZN(new_n1176_));
  NOR2_X1    g1127(.A1(new_n628_), .A2(new_n1176_), .ZN(new_n1177_));
  NAND2_X1   g1128(.A1(new_n1177_), .A2(new_n903_), .ZN(new_n1178_));
  XOR2_X1    g1129(.A1(new_n1177_), .A2(new_n937_), .Z(new_n1179_));
  NOR3_X1    g1130(.A1(new_n1032_), .A2(new_n1034_), .A3(new_n667_), .ZN(new_n1180_));
  NAND2_X1   g1131(.A1(new_n1035_), .A2(new_n659_), .ZN(new_n1181_));
  NOR3_X1    g1132(.A1(new_n514_), .A2(new_n589_), .A3(new_n1089_), .ZN(new_n1182_));
  NAND4_X1   g1133(.A1(new_n885_), .A2(new_n1182_), .A3(new_n961_), .A4(new_n560_), .ZN(new_n1183_));
  NAND4_X1   g1134(.A1(new_n857_), .A2(new_n768_), .A3(new_n966_), .A4(new_n922_), .ZN(new_n1184_));
  NOR3_X1    g1135(.A1(new_n867_), .A2(new_n1183_), .A3(new_n1184_), .ZN(new_n1185_));
  NAND3_X1   g1136(.A1(new_n937_), .A2(new_n958_), .A3(new_n1185_), .ZN(new_n1186_));
  NAND2_X1   g1137(.A1(new_n978_), .A2(new_n903_), .ZN(new_n1187_));
  NAND2_X1   g1138(.A1(new_n1187_), .A2(new_n1186_), .ZN(new_n1188_));
  NAND2_X1   g1139(.A1(new_n1188_), .A2(new_n988_), .ZN(new_n1189_));
  NAND2_X1   g1140(.A1(new_n1189_), .A2(new_n658_), .ZN(new_n1190_));
  NAND3_X1   g1141(.A1(new_n1180_), .A2(new_n1181_), .A3(new_n1190_), .ZN(new_n1191_));
  NAND2_X1   g1142(.A1(new_n1179_), .A2(new_n1191_), .ZN(new_n1192_));
  NAND2_X1   g1143(.A1(new_n1192_), .A2(new_n1178_), .ZN(new_n1193_));
  INV_X1     g1144(.I(new_n1193_), .ZN(new_n1194_));
  NOR2_X1    g1145(.A1(new_n1194_), .A2(new_n1175_), .ZN(new_n1195_));
  INV_X1     g1146(.I(new_n1195_), .ZN(new_n1196_));
  NAND3_X1   g1147(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n1153_), .ZN(new_n1197_));
  NOR2_X1    g1148(.A1(new_n793_), .A2(new_n1125_), .ZN(new_n1198_));
  NOR2_X1    g1149(.A1(new_n795_), .A2(new_n1126_), .ZN(new_n1199_));
  NOR3_X1    g1150(.A1(new_n1197_), .A2(new_n1198_), .A3(new_n1199_), .ZN(new_n1200_));
  INV_X1     g1151(.I(new_n1200_), .ZN(new_n1201_));
  NOR2_X1    g1152(.A1(new_n1100_), .A2(new_n582_), .ZN(new_n1202_));
  AOI21_X1   g1153(.A1(new_n582_), .A2(new_n1098_), .B(new_n1202_), .ZN(new_n1203_));
  NOR2_X1    g1154(.A1(new_n1110_), .A2(new_n790_), .ZN(new_n1204_));
  AOI21_X1   g1155(.A1(new_n790_), .A2(new_n1114_), .B(new_n1204_), .ZN(new_n1205_));
  NAND2_X1   g1156(.A1(new_n1203_), .A2(new_n1205_), .ZN(new_n1206_));
  NAND2_X1   g1157(.A1(new_n1201_), .A2(new_n1206_), .ZN(new_n1207_));
  INV_X1     g1158(.I(new_n1207_), .ZN(new_n1208_));
  NAND2_X1   g1159(.A1(new_n1146_), .A2(new_n1062_), .ZN(new_n1209_));
  OAI21_X1   g1160(.A1(new_n1062_), .A2(new_n1148_), .B(new_n1209_), .ZN(new_n1210_));
  NOR4_X1    g1161(.A1(new_n1210_), .A2(new_n1145_), .A3(new_n1061_), .A4(new_n1132_), .ZN(new_n1211_));
  INV_X1     g1162(.I(new_n1211_), .ZN(new_n1212_));
  NAND3_X1   g1163(.A1(new_n1200_), .A2(new_n1203_), .A3(new_n1205_), .ZN(new_n1213_));
  AOI21_X1   g1164(.A1(new_n1212_), .A2(new_n1213_), .B(new_n1208_), .ZN(new_n1214_));
  NAND2_X1   g1165(.A1(new_n1194_), .A2(new_n1175_), .ZN(new_n1215_));
  INV_X1     g1166(.I(new_n1215_), .ZN(new_n1216_));
  OAI21_X1   g1167(.A1(new_n1214_), .A2(new_n1216_), .B(new_n1196_), .ZN(new_n1217_));
  NOR3_X1    g1168(.A1(new_n1145_), .A2(new_n1061_), .A3(new_n1106_), .ZN(new_n1218_));
  INV_X1     g1169(.I(new_n1218_), .ZN(new_n1219_));
  INV_X1     g1170(.I(new_n1146_), .ZN(new_n1220_));
  NOR2_X1    g1171(.A1(new_n1220_), .A2(new_n1125_), .ZN(new_n1221_));
  NOR2_X1    g1172(.A1(new_n1148_), .A2(new_n1126_), .ZN(new_n1222_));
  OR3_X2     g1173(.A1(new_n1219_), .A2(new_n1221_), .A3(new_n1222_), .Z(new_n1223_));
  NOR3_X1    g1174(.A1(new_n676_), .A2(new_n671_), .A3(new_n1132_), .ZN(new_n1224_));
  INV_X1     g1175(.I(new_n1224_), .ZN(new_n1225_));
  NOR2_X1    g1176(.A1(new_n679_), .A2(new_n1062_), .ZN(new_n1226_));
  NOR2_X1    g1177(.A1(new_n1005_), .A2(new_n1053_), .ZN(new_n1227_));
  NOR3_X1    g1178(.A1(new_n1225_), .A2(new_n1226_), .A3(new_n1227_), .ZN(new_n1228_));
  INV_X1     g1179(.I(new_n1228_), .ZN(new_n1229_));
  NAND2_X1   g1180(.A1(new_n1097_), .A2(new_n752_), .ZN(new_n1230_));
  NOR2_X1    g1181(.A1(new_n1099_), .A2(new_n752_), .ZN(new_n1231_));
  NOR2_X1    g1182(.A1(new_n1231_), .A2(new_n658_), .ZN(new_n1232_));
  AOI21_X1   g1183(.A1(new_n658_), .A2(new_n1230_), .B(new_n1232_), .ZN(new_n1233_));
  NOR2_X1    g1184(.A1(new_n1110_), .A2(new_n667_), .ZN(new_n1234_));
  AOI21_X1   g1185(.A1(new_n667_), .A2(new_n1114_), .B(new_n1234_), .ZN(new_n1235_));
  NAND2_X1   g1186(.A1(new_n1233_), .A2(new_n1235_), .ZN(new_n1236_));
  NAND2_X1   g1187(.A1(new_n1229_), .A2(new_n1236_), .ZN(new_n1237_));
  NAND3_X1   g1188(.A1(new_n1228_), .A2(new_n1233_), .A3(new_n1235_), .ZN(new_n1238_));
  AOI21_X1   g1189(.A1(new_n1238_), .A2(new_n1237_), .B(new_n1223_), .ZN(new_n1239_));
  NOR3_X1    g1190(.A1(new_n1219_), .A2(new_n1221_), .A3(new_n1222_), .ZN(new_n1240_));
  XOR2_X1    g1191(.A1(new_n1236_), .A2(new_n1228_), .Z(new_n1241_));
  NOR2_X1    g1192(.A1(new_n1241_), .A2(new_n1240_), .ZN(new_n1242_));
  NOR2_X1    g1193(.A1(new_n1239_), .A2(new_n1242_), .ZN(new_n1243_));
  NOR2_X1    g1194(.A1(new_n1165_), .A2(new_n1150_), .ZN(new_n1244_));
  OR2_X2     g1195(.A1(new_n1244_), .A2(new_n1164_), .Z(new_n1245_));
  XOR2_X1    g1196(.A1(new_n1243_), .A2(new_n1245_), .Z(new_n1246_));
  AND2_X2    g1197(.A1(new_n1246_), .A2(new_n1217_), .Z(new_n1247_));
  NAND2_X1   g1198(.A1(new_n1243_), .A2(new_n1245_), .ZN(new_n1248_));
  OR2_X2     g1199(.A1(new_n1243_), .A2(new_n1245_), .Z(new_n1249_));
  AOI21_X1   g1200(.A1(new_n1249_), .A2(new_n1248_), .B(new_n1217_), .ZN(new_n1250_));
  NOR2_X1    g1201(.A1(new_n1247_), .A2(new_n1250_), .ZN(new_n1251_));
  OAI21_X1   g1202(.A1(new_n1169_), .A2(new_n1001_), .B(new_n1251_), .ZN(new_n1252_));
  NAND2_X1   g1203(.A1(new_n1252_), .A2(new_n1170_), .ZN(new_n1253_));
  INV_X1     g1204(.I(new_n1253_), .ZN(new_n1254_));
  NAND2_X1   g1205(.A1(new_n1249_), .A2(new_n1217_), .ZN(new_n1255_));
  NAND2_X1   g1206(.A1(new_n1255_), .A2(new_n1248_), .ZN(new_n1256_));
  INV_X1     g1207(.I(new_n1256_), .ZN(new_n1257_));
  NAND2_X1   g1208(.A1(new_n1223_), .A2(new_n1238_), .ZN(new_n1258_));
  NAND2_X1   g1209(.A1(new_n1258_), .A2(new_n1237_), .ZN(new_n1259_));
  NOR3_X1    g1210(.A1(new_n676_), .A2(new_n671_), .A3(new_n1125_), .ZN(new_n1260_));
  INV_X1     g1211(.I(new_n1260_), .ZN(new_n1261_));
  NOR2_X1    g1212(.A1(new_n679_), .A2(new_n1134_), .ZN(new_n1262_));
  NOR2_X1    g1213(.A1(new_n1005_), .A2(new_n1132_), .ZN(new_n1263_));
  NOR3_X1    g1214(.A1(new_n1261_), .A2(new_n1262_), .A3(new_n1263_), .ZN(new_n1264_));
  NAND2_X1   g1215(.A1(new_n1146_), .A2(new_n1153_), .ZN(new_n1265_));
  OAI21_X1   g1216(.A1(new_n1153_), .A2(new_n1148_), .B(new_n1265_), .ZN(new_n1266_));
  NOR4_X1    g1217(.A1(new_n1266_), .A2(new_n790_), .A3(new_n1145_), .A4(new_n1061_), .ZN(new_n1267_));
  NOR2_X1    g1218(.A1(new_n1267_), .A2(new_n1264_), .ZN(new_n1268_));
  AND2_X2    g1219(.A1(new_n1267_), .A2(new_n1264_), .Z(new_n1269_));
  NAND2_X1   g1220(.A1(new_n784_), .A2(new_n780_), .ZN(new_n1270_));
  NAND2_X1   g1221(.A1(new_n1270_), .A2(new_n582_), .ZN(new_n1271_));
  OAI21_X1   g1222(.A1(new_n582_), .A2(new_n795_), .B(new_n1271_), .ZN(new_n1272_));
  NOR4_X1    g1223(.A1(new_n1272_), .A2(new_n667_), .A3(new_n785_), .A4(new_n787_), .ZN(new_n1273_));
  NAND2_X1   g1224(.A1(new_n1096_), .A2(new_n988_), .ZN(new_n1274_));
  XOR2_X1    g1225(.A1(new_n1274_), .A2(new_n752_), .Z(new_n1275_));
  NOR2_X1    g1226(.A1(new_n752_), .A2(new_n659_), .ZN(new_n1276_));
  NOR2_X1    g1227(.A1(new_n1066_), .A2(new_n658_), .ZN(new_n1277_));
  NOR3_X1    g1228(.A1(new_n1097_), .A2(new_n1276_), .A3(new_n1277_), .ZN(new_n1278_));
  NOR2_X1    g1229(.A1(new_n1278_), .A2(new_n1275_), .ZN(new_n1279_));
  NOR2_X1    g1230(.A1(new_n628_), .A2(new_n1062_), .ZN(new_n1280_));
  INV_X1     g1231(.I(new_n1280_), .ZN(new_n1281_));
  NOR2_X1    g1232(.A1(new_n1279_), .A2(new_n1281_), .ZN(new_n1282_));
  NOR3_X1    g1233(.A1(new_n1278_), .A2(new_n1275_), .A3(new_n1280_), .ZN(new_n1283_));
  OAI21_X1   g1234(.A1(new_n1282_), .A2(new_n1283_), .B(new_n1273_), .ZN(new_n1284_));
  XOR2_X1    g1235(.A1(new_n1279_), .A2(new_n1280_), .Z(new_n1285_));
  OR2_X2     g1236(.A1(new_n1273_), .A2(new_n1285_), .Z(new_n1286_));
  NAND2_X1   g1237(.A1(new_n1286_), .A2(new_n1284_), .ZN(new_n1287_));
  NOR3_X1    g1238(.A1(new_n1287_), .A2(new_n1268_), .A3(new_n1269_), .ZN(new_n1288_));
  NOR2_X1    g1239(.A1(new_n1269_), .A2(new_n1268_), .ZN(new_n1289_));
  AOI21_X1   g1240(.A1(new_n1284_), .A2(new_n1286_), .B(new_n1289_), .ZN(new_n1290_));
  OAI21_X1   g1241(.A1(new_n1290_), .A2(new_n1288_), .B(new_n1259_), .ZN(new_n1291_));
  INV_X1     g1242(.I(new_n1259_), .ZN(new_n1292_));
  XNOR2_X1   g1243(.A1(new_n1289_), .A2(new_n1287_), .ZN(new_n1293_));
  NAND2_X1   g1244(.A1(new_n1293_), .A2(new_n1292_), .ZN(new_n1294_));
  INV_X1     g1245(.I(new_n996_), .ZN(new_n1295_));
  AOI21_X1   g1246(.A1(new_n1295_), .A2(new_n798_), .B(new_n994_), .ZN(new_n1296_));
  AOI21_X1   g1247(.A1(new_n1294_), .A2(new_n1291_), .B(new_n1296_), .ZN(new_n1297_));
  NAND2_X1   g1248(.A1(new_n1294_), .A2(new_n1291_), .ZN(new_n1298_));
  INV_X1     g1249(.I(new_n1296_), .ZN(new_n1299_));
  NOR2_X1    g1250(.A1(new_n1298_), .A2(new_n1299_), .ZN(new_n1300_));
  NOR2_X1    g1251(.A1(new_n1300_), .A2(new_n1297_), .ZN(new_n1301_));
  NOR2_X1    g1252(.A1(new_n1301_), .A2(new_n1257_), .ZN(new_n1302_));
  NAND3_X1   g1253(.A1(new_n1294_), .A2(new_n1291_), .A3(new_n1299_), .ZN(new_n1303_));
  NAND2_X1   g1254(.A1(new_n1298_), .A2(new_n1296_), .ZN(new_n1304_));
  AOI21_X1   g1255(.A1(new_n1304_), .A2(new_n1303_), .B(new_n1256_), .ZN(new_n1305_));
  NOR2_X1    g1256(.A1(new_n1302_), .A2(new_n1305_), .ZN(new_n1306_));
  INV_X1     g1257(.I(new_n1306_), .ZN(new_n1307_));
  NAND2_X1   g1258(.A1(new_n1307_), .A2(new_n1254_), .ZN(new_n1308_));
  XOR2_X1    g1259(.A1(new_n1041_), .A2(new_n1028_), .Z(new_n1309_));
  XNOR2_X1   g1260(.A1(new_n1039_), .A2(new_n1309_), .ZN(new_n1310_));
  INV_X1     g1261(.I(new_n1310_), .ZN(new_n1311_));
  NOR2_X1    g1262(.A1(new_n1116_), .A2(new_n1064_), .ZN(new_n1312_));
  NAND2_X1   g1263(.A1(new_n1116_), .A2(new_n1064_), .ZN(new_n1313_));
  INV_X1     g1264(.I(new_n1313_), .ZN(new_n1314_));
  OAI21_X1   g1265(.A1(new_n1314_), .A2(new_n1312_), .B(new_n1136_), .ZN(new_n1315_));
  INV_X1     g1266(.I(new_n1064_), .ZN(new_n1316_));
  NOR2_X1    g1267(.A1(new_n1316_), .A2(new_n1116_), .ZN(new_n1317_));
  OAI21_X1   g1268(.A1(new_n1118_), .A2(new_n1317_), .B(new_n1137_), .ZN(new_n1318_));
  AOI21_X1   g1269(.A1(new_n1318_), .A2(new_n1315_), .B(new_n1311_), .ZN(new_n1319_));
  NOR4_X1    g1270(.A1(new_n1026_), .A2(new_n599_), .A3(new_n1017_), .A4(new_n1023_), .ZN(new_n1320_));
  NAND2_X1   g1271(.A1(new_n1320_), .A2(new_n1013_), .ZN(new_n1321_));
  NAND2_X1   g1272(.A1(new_n1321_), .A2(new_n658_), .ZN(new_n1322_));
  OAI21_X1   g1273(.A1(new_n1321_), .A2(new_n678_), .B(new_n937_), .ZN(new_n1323_));
  XNOR2_X1   g1274(.A1(new_n1323_), .A2(new_n1322_), .ZN(new_n1324_));
  OR3_X2     g1275(.A1(new_n416_), .A2(new_n67_), .A3(new_n650_), .Z(new_n1325_));
  INV_X1     g1276(.I(new_n67_), .ZN(new_n1326_));
  OAI21_X1   g1277(.A1(new_n415_), .A2(new_n1326_), .B(new_n650_), .ZN(new_n1327_));
  AOI21_X1   g1278(.A1(new_n1325_), .A2(new_n1327_), .B(new_n628_), .ZN(new_n1328_));
  XOR2_X1    g1279(.A1(new_n1328_), .A2(new_n1324_), .Z(new_n1329_));
  INV_X1     g1280(.I(new_n1329_), .ZN(new_n1330_));
  NOR3_X1    g1281(.A1(new_n1032_), .A2(new_n1034_), .A3(new_n790_), .ZN(new_n1331_));
  INV_X1     g1282(.I(new_n1035_), .ZN(new_n1332_));
  NOR2_X1    g1283(.A1(new_n1332_), .A2(new_n581_), .ZN(new_n1333_));
  AOI21_X1   g1284(.A1(new_n581_), .A2(new_n1189_), .B(new_n1333_), .ZN(new_n1334_));
  NAND2_X1   g1285(.A1(new_n1334_), .A2(new_n1331_), .ZN(new_n1335_));
  INV_X1     g1286(.I(new_n1335_), .ZN(new_n1336_));
  NOR2_X1    g1287(.A1(new_n1330_), .A2(new_n1336_), .ZN(new_n1337_));
  NOR3_X1    g1288(.A1(new_n676_), .A2(new_n671_), .A3(new_n56_), .ZN(new_n1338_));
  INV_X1     g1289(.I(new_n1338_), .ZN(new_n1339_));
  NOR2_X1    g1290(.A1(new_n679_), .A2(new_n1326_), .ZN(new_n1340_));
  NOR2_X1    g1291(.A1(new_n1005_), .A2(new_n67_), .ZN(new_n1341_));
  NOR3_X1    g1292(.A1(new_n1339_), .A2(new_n1340_), .A3(new_n1341_), .ZN(new_n1342_));
  INV_X1     g1293(.I(new_n1342_), .ZN(new_n1343_));
  NOR2_X1    g1294(.A1(new_n1329_), .A2(new_n1335_), .ZN(new_n1344_));
  INV_X1     g1295(.I(new_n1344_), .ZN(new_n1345_));
  AOI21_X1   g1296(.A1(new_n1343_), .A2(new_n1345_), .B(new_n1337_), .ZN(new_n1346_));
  INV_X1     g1297(.I(new_n1346_), .ZN(new_n1347_));
  NAND3_X1   g1298(.A1(new_n1318_), .A2(new_n1315_), .A3(new_n1311_), .ZN(new_n1348_));
  AOI21_X1   g1299(.A1(new_n1347_), .A2(new_n1348_), .B(new_n1319_), .ZN(new_n1349_));
  XOR2_X1    g1300(.A1(new_n1042_), .A2(new_n1007_), .Z(new_n1350_));
  NOR2_X1    g1301(.A1(new_n1350_), .A2(new_n1139_), .ZN(new_n1351_));
  INV_X1     g1302(.I(new_n1139_), .ZN(new_n1352_));
  INV_X1     g1303(.I(new_n1140_), .ZN(new_n1353_));
  AOI21_X1   g1304(.A1(new_n1043_), .A2(new_n1353_), .B(new_n1352_), .ZN(new_n1354_));
  NOR2_X1    g1305(.A1(new_n1354_), .A2(new_n1351_), .ZN(new_n1355_));
  INV_X1     g1306(.I(new_n1355_), .ZN(new_n1356_));
  NOR2_X1    g1307(.A1(new_n1356_), .A2(new_n1349_), .ZN(new_n1357_));
  XOR2_X1    g1308(.A1(new_n1206_), .A2(new_n1200_), .Z(new_n1358_));
  NOR2_X1    g1309(.A1(new_n1358_), .A2(new_n1212_), .ZN(new_n1359_));
  AOI21_X1   g1310(.A1(new_n1207_), .A2(new_n1213_), .B(new_n1211_), .ZN(new_n1360_));
  NOR2_X1    g1311(.A1(new_n1359_), .A2(new_n1360_), .ZN(new_n1361_));
  INV_X1     g1312(.I(new_n1361_), .ZN(new_n1362_));
  XOR2_X1    g1313(.A1(new_n1179_), .A2(new_n1191_), .Z(new_n1363_));
  NAND2_X1   g1314(.A1(new_n675_), .A2(new_n62_), .ZN(new_n1364_));
  OAI21_X1   g1315(.A1(new_n671_), .A2(new_n62_), .B(new_n1364_), .ZN(new_n1365_));
  NAND2_X1   g1316(.A1(new_n682_), .A2(new_n1176_), .ZN(new_n1366_));
  OAI21_X1   g1317(.A1(new_n1176_), .A2(new_n679_), .B(new_n1366_), .ZN(new_n1367_));
  NAND2_X1   g1318(.A1(new_n1367_), .A2(new_n1365_), .ZN(new_n1368_));
  INV_X1     g1319(.I(new_n1368_), .ZN(new_n1369_));
  INV_X1     g1320(.I(new_n1328_), .ZN(new_n1370_));
  NOR2_X1    g1321(.A1(new_n1370_), .A2(new_n1324_), .ZN(new_n1371_));
  NAND2_X1   g1322(.A1(new_n1369_), .A2(new_n1371_), .ZN(new_n1372_));
  NAND2_X1   g1323(.A1(new_n1368_), .A2(new_n1371_), .ZN(new_n1373_));
  INV_X1     g1324(.I(new_n1373_), .ZN(new_n1374_));
  NOR2_X1    g1325(.A1(new_n1368_), .A2(new_n1371_), .ZN(new_n1375_));
  NOR2_X1    g1326(.A1(new_n1374_), .A2(new_n1375_), .ZN(new_n1376_));
  INV_X1     g1327(.I(new_n1376_), .ZN(new_n1377_));
  NOR2_X1    g1328(.A1(new_n1047_), .A2(new_n939_), .ZN(new_n1378_));
  XOR2_X1    g1329(.A1(new_n494_), .A2(new_n62_), .Z(new_n1379_));
  NOR2_X1    g1330(.A1(new_n1055_), .A2(new_n1379_), .ZN(new_n1380_));
  NAND2_X1   g1331(.A1(new_n690_), .A2(new_n1171_), .ZN(new_n1381_));
  NOR4_X1    g1332(.A1(new_n1378_), .A2(new_n1061_), .A3(new_n1380_), .A4(new_n1381_), .ZN(new_n1382_));
  NOR3_X1    g1333(.A1(new_n785_), .A2(new_n787_), .A3(new_n1132_), .ZN(new_n1383_));
  NAND2_X1   g1334(.A1(new_n1270_), .A2(new_n1062_), .ZN(new_n1384_));
  OAI21_X1   g1335(.A1(new_n792_), .A2(new_n786_), .B(new_n1053_), .ZN(new_n1385_));
  NAND3_X1   g1336(.A1(new_n1383_), .A2(new_n1385_), .A3(new_n1384_), .ZN(new_n1386_));
  NOR2_X1    g1337(.A1(new_n1231_), .A2(new_n1106_), .ZN(new_n1387_));
  AOI21_X1   g1338(.A1(new_n1230_), .A2(new_n1106_), .B(new_n1387_), .ZN(new_n1388_));
  NOR2_X1    g1339(.A1(new_n1110_), .A2(new_n1125_), .ZN(new_n1389_));
  AOI21_X1   g1340(.A1(new_n1114_), .A2(new_n1125_), .B(new_n1389_), .ZN(new_n1390_));
  NAND2_X1   g1341(.A1(new_n1388_), .A2(new_n1390_), .ZN(new_n1391_));
  XOR2_X1    g1342(.A1(new_n1391_), .A2(new_n1386_), .Z(new_n1392_));
  NAND2_X1   g1343(.A1(new_n1392_), .A2(new_n1382_), .ZN(new_n1393_));
  NAND3_X1   g1344(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n1134_), .ZN(new_n1394_));
  NOR2_X1    g1345(.A1(new_n793_), .A2(new_n1053_), .ZN(new_n1395_));
  INV_X1     g1346(.I(new_n1385_), .ZN(new_n1396_));
  NOR3_X1    g1347(.A1(new_n1394_), .A2(new_n1395_), .A3(new_n1396_), .ZN(new_n1397_));
  INV_X1     g1348(.I(new_n1391_), .ZN(new_n1398_));
  NAND2_X1   g1349(.A1(new_n1398_), .A2(new_n1397_), .ZN(new_n1399_));
  XOR2_X1    g1350(.A1(new_n1393_), .A2(new_n1399_), .Z(new_n1400_));
  NAND2_X1   g1351(.A1(new_n1400_), .A2(new_n1377_), .ZN(new_n1401_));
  NAND2_X1   g1352(.A1(new_n1401_), .A2(new_n1372_), .ZN(new_n1402_));
  XOR2_X1    g1353(.A1(new_n1402_), .A2(new_n1363_), .Z(new_n1403_));
  XOR2_X1    g1354(.A1(new_n1403_), .A2(new_n1362_), .Z(new_n1404_));
  NAND2_X1   g1355(.A1(new_n1356_), .A2(new_n1349_), .ZN(new_n1405_));
  AOI21_X1   g1356(.A1(new_n1404_), .A2(new_n1405_), .B(new_n1357_), .ZN(new_n1406_));
  XOR2_X1    g1357(.A1(new_n1175_), .A2(new_n1193_), .Z(new_n1407_));
  NOR2_X1    g1358(.A1(new_n1214_), .A2(new_n1407_), .ZN(new_n1408_));
  INV_X1     g1359(.I(new_n1214_), .ZN(new_n1409_));
  AOI21_X1   g1360(.A1(new_n1196_), .A2(new_n1215_), .B(new_n1409_), .ZN(new_n1410_));
  NOR2_X1    g1361(.A1(new_n1410_), .A2(new_n1408_), .ZN(new_n1411_));
  INV_X1     g1362(.I(new_n1411_), .ZN(new_n1412_));
  XOR2_X1    g1363(.A1(new_n1167_), .A2(new_n1144_), .Z(new_n1413_));
  NAND2_X1   g1364(.A1(new_n1362_), .A2(new_n1363_), .ZN(new_n1414_));
  XOR2_X1    g1365(.A1(new_n1361_), .A2(new_n1363_), .Z(new_n1415_));
  NAND3_X1   g1366(.A1(new_n1415_), .A2(new_n1401_), .A3(new_n1372_), .ZN(new_n1416_));
  NAND2_X1   g1367(.A1(new_n1416_), .A2(new_n1414_), .ZN(new_n1417_));
  NAND2_X1   g1368(.A1(new_n1417_), .A2(new_n1413_), .ZN(new_n1418_));
  XOR2_X1    g1369(.A1(new_n1167_), .A2(new_n1143_), .Z(new_n1419_));
  INV_X1     g1370(.I(new_n1417_), .ZN(new_n1420_));
  NAND2_X1   g1371(.A1(new_n1420_), .A2(new_n1419_), .ZN(new_n1421_));
  AOI21_X1   g1372(.A1(new_n1421_), .A2(new_n1418_), .B(new_n1141_), .ZN(new_n1422_));
  INV_X1     g1373(.I(new_n1422_), .ZN(new_n1423_));
  NAND3_X1   g1374(.A1(new_n1421_), .A2(new_n1141_), .A3(new_n1418_), .ZN(new_n1424_));
  AOI21_X1   g1375(.A1(new_n1423_), .A2(new_n1424_), .B(new_n1412_), .ZN(new_n1425_));
  INV_X1     g1376(.I(new_n1424_), .ZN(new_n1426_));
  NOR3_X1    g1377(.A1(new_n1426_), .A2(new_n1411_), .A3(new_n1422_), .ZN(new_n1427_));
  NOR3_X1    g1378(.A1(new_n1427_), .A2(new_n1425_), .A3(new_n1406_), .ZN(new_n1428_));
  NOR2_X1    g1379(.A1(new_n1307_), .A2(new_n1254_), .ZN(new_n1429_));
  NOR2_X1    g1380(.A1(new_n1306_), .A2(new_n1253_), .ZN(new_n1430_));
  XOR2_X1    g1381(.A1(new_n1419_), .A2(new_n1141_), .Z(new_n1431_));
  XOR2_X1    g1382(.A1(new_n1431_), .A2(new_n1411_), .Z(new_n1432_));
  AOI21_X1   g1383(.A1(new_n1417_), .A2(new_n1431_), .B(new_n1432_), .ZN(new_n1433_));
  XNOR2_X1   g1384(.A1(new_n1169_), .A2(new_n1001_), .ZN(new_n1434_));
  INV_X1     g1385(.I(new_n1434_), .ZN(new_n1435_));
  NOR2_X1    g1386(.A1(new_n1435_), .A2(new_n1251_), .ZN(new_n1436_));
  INV_X1     g1387(.I(new_n1251_), .ZN(new_n1437_));
  NOR2_X1    g1388(.A1(new_n1437_), .A2(new_n1434_), .ZN(new_n1438_));
  NOR2_X1    g1389(.A1(new_n1436_), .A2(new_n1438_), .ZN(new_n1439_));
  OAI22_X1   g1390(.A1(new_n1429_), .A2(new_n1430_), .B1(new_n1439_), .B2(new_n1433_), .ZN(new_n1440_));
  OAI21_X1   g1391(.A1(new_n1440_), .A2(new_n1428_), .B(new_n1308_), .ZN(new_n1441_));
  NOR2_X1    g1392(.A1(new_n1300_), .A2(new_n1257_), .ZN(new_n1442_));
  NOR2_X1    g1393(.A1(new_n1442_), .A2(new_n1297_), .ZN(new_n1443_));
  INV_X1     g1394(.I(new_n1443_), .ZN(new_n1444_));
  NOR2_X1    g1395(.A1(new_n1290_), .A2(new_n1292_), .ZN(new_n1445_));
  NOR2_X1    g1396(.A1(new_n1445_), .A2(new_n1288_), .ZN(new_n1446_));
  INV_X1     g1397(.I(new_n1268_), .ZN(new_n1447_));
  NOR2_X1    g1398(.A1(new_n1273_), .A2(new_n1283_), .ZN(new_n1448_));
  NOR2_X1    g1399(.A1(new_n1448_), .A2(new_n1282_), .ZN(new_n1449_));
  NAND2_X1   g1400(.A1(new_n1107_), .A2(new_n752_), .ZN(new_n1450_));
  XOR2_X1    g1401(.A1(new_n1132_), .A2(new_n1062_), .Z(new_n1451_));
  NOR2_X1    g1402(.A1(new_n628_), .A2(new_n1451_), .ZN(new_n1452_));
  XOR2_X1    g1403(.A1(new_n1452_), .A2(new_n1450_), .Z(new_n1453_));
  NOR2_X1    g1404(.A1(new_n1449_), .A2(new_n1453_), .ZN(new_n1454_));
  INV_X1     g1405(.I(new_n1454_), .ZN(new_n1455_));
  NAND2_X1   g1406(.A1(new_n1449_), .A2(new_n1453_), .ZN(new_n1456_));
  AOI21_X1   g1407(.A1(new_n1455_), .A2(new_n1456_), .B(new_n1447_), .ZN(new_n1457_));
  XOR2_X1    g1408(.A1(new_n1449_), .A2(new_n1453_), .Z(new_n1458_));
  AOI21_X1   g1409(.A1(new_n1447_), .A2(new_n1458_), .B(new_n1457_), .ZN(new_n1459_));
  INV_X1     g1410(.I(new_n1061_), .ZN(new_n1460_));
  NAND3_X1   g1411(.A1(new_n1460_), .A2(new_n1047_), .A3(new_n582_), .ZN(new_n1461_));
  NAND2_X1   g1412(.A1(new_n1146_), .A2(new_n576_), .ZN(new_n1462_));
  OAI21_X1   g1413(.A1(new_n576_), .A2(new_n1148_), .B(new_n1462_), .ZN(new_n1463_));
  NOR2_X1    g1414(.A1(new_n1463_), .A2(new_n1461_), .ZN(new_n1464_));
  INV_X1     g1415(.I(new_n1464_), .ZN(new_n1465_));
  NAND3_X1   g1416(.A1(new_n696_), .A2(new_n675_), .A3(new_n1153_), .ZN(new_n1466_));
  NOR2_X1    g1417(.A1(new_n679_), .A2(new_n1126_), .ZN(new_n1467_));
  NOR2_X1    g1418(.A1(new_n1005_), .A2(new_n1125_), .ZN(new_n1468_));
  NOR3_X1    g1419(.A1(new_n1466_), .A2(new_n1467_), .A3(new_n1468_), .ZN(new_n1469_));
  INV_X1     g1420(.I(new_n1469_), .ZN(new_n1470_));
  NAND3_X1   g1421(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n659_), .ZN(new_n1471_));
  NAND2_X1   g1422(.A1(new_n1270_), .A2(new_n678_), .ZN(new_n1472_));
  OAI21_X1   g1423(.A1(new_n678_), .A2(new_n795_), .B(new_n1472_), .ZN(new_n1473_));
  NOR2_X1    g1424(.A1(new_n1473_), .A2(new_n1471_), .ZN(new_n1474_));
  XOR2_X1    g1425(.A1(new_n1474_), .A2(new_n1470_), .Z(new_n1475_));
  NOR2_X1    g1426(.A1(new_n1475_), .A2(new_n1465_), .ZN(new_n1476_));
  OAI21_X1   g1427(.A1(new_n1473_), .A2(new_n1471_), .B(new_n1470_), .ZN(new_n1477_));
  NAND2_X1   g1428(.A1(new_n1474_), .A2(new_n1469_), .ZN(new_n1478_));
  AOI21_X1   g1429(.A1(new_n1478_), .A2(new_n1477_), .B(new_n1464_), .ZN(new_n1479_));
  NOR2_X1    g1430(.A1(new_n1476_), .A2(new_n1479_), .ZN(new_n1480_));
  NOR2_X1    g1431(.A1(new_n1459_), .A2(new_n1480_), .ZN(new_n1481_));
  INV_X1     g1432(.I(new_n1481_), .ZN(new_n1482_));
  NAND2_X1   g1433(.A1(new_n1459_), .A2(new_n1480_), .ZN(new_n1483_));
  AOI21_X1   g1434(.A1(new_n1482_), .A2(new_n1483_), .B(new_n1446_), .ZN(new_n1484_));
  XOR2_X1    g1435(.A1(new_n1459_), .A2(new_n1480_), .Z(new_n1485_));
  AOI21_X1   g1436(.A1(new_n1446_), .A2(new_n1485_), .B(new_n1484_), .ZN(new_n1486_));
  INV_X1     g1437(.I(new_n1486_), .ZN(new_n1487_));
  NOR2_X1    g1438(.A1(new_n1487_), .A2(new_n1444_), .ZN(new_n1488_));
  INV_X1     g1439(.I(new_n1488_), .ZN(new_n1489_));
  NAND2_X1   g1440(.A1(new_n1441_), .A2(new_n1489_), .ZN(new_n1490_));
  NOR3_X1    g1441(.A1(new_n1145_), .A2(new_n1061_), .A3(new_n667_), .ZN(new_n1491_));
  NOR2_X1    g1442(.A1(new_n1148_), .A2(new_n582_), .ZN(new_n1492_));
  AOI21_X1   g1443(.A1(new_n582_), .A2(new_n1146_), .B(new_n1492_), .ZN(new_n1493_));
  NAND2_X1   g1444(.A1(new_n1493_), .A2(new_n1491_), .ZN(new_n1494_));
  NAND2_X1   g1445(.A1(new_n778_), .A2(new_n752_), .ZN(new_n1495_));
  XOR2_X1    g1446(.A1(new_n1495_), .A2(new_n494_), .Z(new_n1496_));
  XOR2_X1    g1447(.A1(new_n778_), .A2(new_n752_), .Z(new_n1497_));
  INV_X1     g1448(.I(new_n1497_), .ZN(new_n1498_));
  OAI21_X1   g1449(.A1(new_n494_), .A2(new_n659_), .B(new_n1498_), .ZN(new_n1499_));
  AOI21_X1   g1450(.A1(new_n494_), .A2(new_n659_), .B(new_n1499_), .ZN(new_n1500_));
  NOR2_X1    g1451(.A1(new_n1500_), .A2(new_n1496_), .ZN(new_n1501_));
  NOR2_X1    g1452(.A1(new_n628_), .A2(new_n1126_), .ZN(new_n1502_));
  INV_X1     g1453(.I(new_n1502_), .ZN(new_n1503_));
  XOR2_X1    g1454(.A1(new_n1501_), .A2(new_n1503_), .Z(new_n1504_));
  AOI21_X1   g1455(.A1(new_n1268_), .A2(new_n1456_), .B(new_n1454_), .ZN(new_n1505_));
  NAND2_X1   g1456(.A1(new_n1478_), .A2(new_n1465_), .ZN(new_n1506_));
  NAND2_X1   g1457(.A1(new_n1506_), .A2(new_n1477_), .ZN(new_n1507_));
  NOR2_X1    g1458(.A1(new_n679_), .A2(new_n1153_), .ZN(new_n1508_));
  AOI21_X1   g1459(.A1(new_n682_), .A2(new_n1153_), .B(new_n1508_), .ZN(new_n1509_));
  NAND4_X1   g1460(.A1(new_n1509_), .A2(new_n576_), .A3(new_n696_), .A4(new_n675_), .ZN(new_n1510_));
  NOR2_X1    g1461(.A1(new_n1134_), .A2(new_n1062_), .ZN(new_n1511_));
  AOI21_X1   g1462(.A1(new_n1062_), .A2(new_n1134_), .B(new_n628_), .ZN(new_n1512_));
  OAI21_X1   g1463(.A1(new_n1450_), .A2(new_n1511_), .B(new_n1512_), .ZN(new_n1513_));
  NAND2_X1   g1464(.A1(new_n1510_), .A2(new_n1513_), .ZN(new_n1514_));
  INV_X1     g1465(.I(new_n1514_), .ZN(new_n1515_));
  NOR2_X1    g1466(.A1(new_n1510_), .A2(new_n1513_), .ZN(new_n1516_));
  OAI21_X1   g1467(.A1(new_n1515_), .A2(new_n1516_), .B(new_n1507_), .ZN(new_n1517_));
  INV_X1     g1468(.I(new_n1507_), .ZN(new_n1518_));
  XOR2_X1    g1469(.A1(new_n1510_), .A2(new_n1513_), .Z(new_n1519_));
  NAND2_X1   g1470(.A1(new_n1518_), .A2(new_n1519_), .ZN(new_n1520_));
  NAND2_X1   g1471(.A1(new_n1520_), .A2(new_n1517_), .ZN(new_n1521_));
  XOR2_X1    g1472(.A1(new_n1521_), .A2(new_n1505_), .Z(new_n1522_));
  XNOR2_X1   g1473(.A1(new_n1522_), .A2(new_n1504_), .ZN(new_n1523_));
  XOR2_X1    g1474(.A1(new_n1523_), .A2(new_n1494_), .Z(new_n1524_));
  INV_X1     g1475(.I(new_n1446_), .ZN(new_n1525_));
  AOI21_X1   g1476(.A1(new_n1525_), .A2(new_n1483_), .B(new_n1481_), .ZN(new_n1526_));
  NAND2_X1   g1477(.A1(new_n1524_), .A2(new_n1526_), .ZN(new_n1527_));
  INV_X1     g1478(.I(new_n1527_), .ZN(new_n1528_));
  NOR2_X1    g1479(.A1(new_n1524_), .A2(new_n1526_), .ZN(new_n1529_));
  NOR2_X1    g1480(.A1(new_n1486_), .A2(new_n1443_), .ZN(new_n1530_));
  NOR3_X1    g1481(.A1(new_n1528_), .A2(new_n1529_), .A3(new_n1530_), .ZN(new_n1531_));
  NAND2_X1   g1482(.A1(new_n1490_), .A2(new_n1531_), .ZN(new_n1532_));
  XNOR2_X1   g1483(.A1(new_n1306_), .A2(new_n1253_), .ZN(new_n1533_));
  INV_X1     g1484(.I(new_n1357_), .ZN(new_n1534_));
  XNOR2_X1   g1485(.A1(new_n1402_), .A2(new_n1363_), .ZN(new_n1535_));
  NAND2_X1   g1486(.A1(new_n1535_), .A2(new_n1361_), .ZN(new_n1536_));
  NAND2_X1   g1487(.A1(new_n1403_), .A2(new_n1362_), .ZN(new_n1537_));
  NAND2_X1   g1488(.A1(new_n1536_), .A2(new_n1537_), .ZN(new_n1538_));
  INV_X1     g1489(.I(new_n1405_), .ZN(new_n1539_));
  OAI21_X1   g1490(.A1(new_n1538_), .A2(new_n1539_), .B(new_n1534_), .ZN(new_n1540_));
  OAI21_X1   g1491(.A1(new_n1426_), .A2(new_n1422_), .B(new_n1411_), .ZN(new_n1541_));
  NAND3_X1   g1492(.A1(new_n1423_), .A2(new_n1412_), .A3(new_n1424_), .ZN(new_n1542_));
  NAND3_X1   g1493(.A1(new_n1542_), .A2(new_n1541_), .A3(new_n1540_), .ZN(new_n1543_));
  XOR2_X1    g1494(.A1(new_n1413_), .A2(new_n1141_), .Z(new_n1544_));
  XOR2_X1    g1495(.A1(new_n1544_), .A2(new_n1411_), .Z(new_n1545_));
  OAI21_X1   g1496(.A1(new_n1420_), .A2(new_n1544_), .B(new_n1545_), .ZN(new_n1546_));
  INV_X1     g1497(.I(new_n1439_), .ZN(new_n1547_));
  NAND2_X1   g1498(.A1(new_n1547_), .A2(new_n1546_), .ZN(new_n1548_));
  NAND3_X1   g1499(.A1(new_n1543_), .A2(new_n1533_), .A3(new_n1548_), .ZN(new_n1549_));
  AOI21_X1   g1500(.A1(new_n1549_), .A2(new_n1308_), .B(new_n1488_), .ZN(new_n1550_));
  INV_X1     g1501(.I(new_n1529_), .ZN(new_n1551_));
  INV_X1     g1502(.I(new_n1530_), .ZN(new_n1552_));
  NAND3_X1   g1503(.A1(new_n1551_), .A2(new_n1527_), .A3(new_n1552_), .ZN(new_n1553_));
  OAI21_X1   g1504(.A1(new_n1518_), .A2(new_n1516_), .B(new_n1514_), .ZN(new_n1554_));
  NAND2_X1   g1505(.A1(new_n1501_), .A2(new_n1503_), .ZN(new_n1555_));
  NAND2_X1   g1506(.A1(new_n1555_), .A2(new_n1494_), .ZN(new_n1556_));
  OAI21_X1   g1507(.A1(new_n1501_), .A2(new_n1503_), .B(new_n1556_), .ZN(new_n1557_));
  NOR3_X1    g1508(.A1(new_n1145_), .A2(new_n1061_), .A3(new_n658_), .ZN(new_n1558_));
  NOR2_X1    g1509(.A1(new_n1148_), .A2(new_n678_), .ZN(new_n1559_));
  AOI21_X1   g1510(.A1(new_n678_), .A2(new_n1146_), .B(new_n1559_), .ZN(new_n1560_));
  NAND2_X1   g1511(.A1(new_n1560_), .A2(new_n1558_), .ZN(new_n1561_));
  NOR3_X1    g1512(.A1(new_n676_), .A2(new_n671_), .A3(new_n581_), .ZN(new_n1562_));
  INV_X1     g1513(.I(new_n1562_), .ZN(new_n1563_));
  NOR2_X1    g1514(.A1(new_n679_), .A2(new_n576_), .ZN(new_n1564_));
  NOR2_X1    g1515(.A1(new_n1005_), .A2(new_n790_), .ZN(new_n1565_));
  NOR3_X1    g1516(.A1(new_n1563_), .A2(new_n1564_), .A3(new_n1565_), .ZN(new_n1566_));
  INV_X1     g1517(.I(new_n1566_), .ZN(new_n1567_));
  XOR2_X1    g1518(.A1(new_n1561_), .A2(new_n1567_), .Z(new_n1568_));
  NAND2_X1   g1519(.A1(new_n1557_), .A2(new_n1568_), .ZN(new_n1569_));
  INV_X1     g1520(.I(new_n1557_), .ZN(new_n1570_));
  AOI21_X1   g1521(.A1(new_n1560_), .A2(new_n1558_), .B(new_n1566_), .ZN(new_n1571_));
  NOR2_X1    g1522(.A1(new_n1561_), .A2(new_n1567_), .ZN(new_n1572_));
  OAI21_X1   g1523(.A1(new_n1571_), .A2(new_n1572_), .B(new_n1570_), .ZN(new_n1573_));
  NAND2_X1   g1524(.A1(new_n1573_), .A2(new_n1569_), .ZN(new_n1574_));
  NOR2_X1    g1525(.A1(new_n1153_), .A2(new_n1125_), .ZN(new_n1575_));
  NOR2_X1    g1526(.A1(new_n1126_), .A2(new_n1106_), .ZN(new_n1576_));
  OAI21_X1   g1527(.A1(new_n1575_), .A2(new_n1576_), .B(new_n627_), .ZN(new_n1577_));
  XNOR2_X1   g1528(.A1(new_n780_), .A2(new_n1577_), .ZN(new_n1578_));
  INV_X1     g1529(.I(new_n1578_), .ZN(new_n1579_));
  XOR2_X1    g1530(.A1(new_n1574_), .A2(new_n1579_), .Z(new_n1580_));
  AND2_X2    g1531(.A1(new_n1580_), .A2(new_n1554_), .Z(new_n1581_));
  NAND2_X1   g1532(.A1(new_n1574_), .A2(new_n1579_), .ZN(new_n1582_));
  NAND3_X1   g1533(.A1(new_n1573_), .A2(new_n1569_), .A3(new_n1578_), .ZN(new_n1583_));
  AOI21_X1   g1534(.A1(new_n1582_), .A2(new_n1583_), .B(new_n1554_), .ZN(new_n1584_));
  NOR2_X1    g1535(.A1(new_n1581_), .A2(new_n1584_), .ZN(new_n1585_));
  OAI21_X1   g1536(.A1(new_n1550_), .A2(new_n1553_), .B(new_n1585_), .ZN(new_n1586_));
  INV_X1     g1537(.I(new_n1585_), .ZN(new_n1587_));
  NAND3_X1   g1538(.A1(new_n1490_), .A2(new_n1531_), .A3(new_n1587_), .ZN(new_n1588_));
  AOI21_X1   g1539(.A1(new_n1517_), .A2(new_n1520_), .B(new_n1505_), .ZN(new_n1589_));
  XOR2_X1    g1540(.A1(new_n1504_), .A2(new_n1494_), .Z(new_n1590_));
  NOR2_X1    g1541(.A1(new_n1521_), .A2(new_n1590_), .ZN(new_n1591_));
  AOI21_X1   g1542(.A1(new_n1591_), .A2(new_n1505_), .B(new_n1589_), .ZN(new_n1592_));
  INV_X1     g1543(.I(new_n1592_), .ZN(new_n1593_));
  AOI22_X1   g1544(.A1(new_n1588_), .A2(new_n1586_), .B1(new_n1532_), .B2(new_n1593_), .ZN(new_n1594_));
  NAND2_X1   g1545(.A1(new_n1582_), .A2(new_n1554_), .ZN(new_n1595_));
  NAND2_X1   g1546(.A1(new_n1595_), .A2(new_n1583_), .ZN(new_n1596_));
  INV_X1     g1547(.I(new_n699_), .ZN(new_n1597_));
  OAI21_X1   g1548(.A1(new_n702_), .A2(new_n695_), .B(new_n1597_), .ZN(new_n1598_));
  XOR2_X1    g1549(.A1(new_n694_), .A2(new_n701_), .Z(new_n1599_));
  OAI21_X1   g1550(.A1(new_n1597_), .A2(new_n1599_), .B(new_n1598_), .ZN(new_n1600_));
  NOR2_X1    g1551(.A1(new_n1126_), .A2(new_n1153_), .ZN(new_n1601_));
  AOI21_X1   g1552(.A1(new_n1153_), .A2(new_n1126_), .B(new_n628_), .ZN(new_n1602_));
  OAI21_X1   g1553(.A1(new_n780_), .A2(new_n1601_), .B(new_n1602_), .ZN(new_n1603_));
  INV_X1     g1554(.I(new_n1603_), .ZN(new_n1604_));
  NOR2_X1    g1555(.A1(new_n1600_), .A2(new_n1604_), .ZN(new_n1605_));
  NOR2_X1    g1556(.A1(new_n1570_), .A2(new_n1572_), .ZN(new_n1606_));
  NOR2_X1    g1557(.A1(new_n1606_), .A2(new_n1571_), .ZN(new_n1607_));
  NAND2_X1   g1558(.A1(new_n1600_), .A2(new_n1604_), .ZN(new_n1608_));
  INV_X1     g1559(.I(new_n1608_), .ZN(new_n1609_));
  NOR2_X1    g1560(.A1(new_n1607_), .A2(new_n1609_), .ZN(new_n1610_));
  NOR2_X1    g1561(.A1(new_n1610_), .A2(new_n1605_), .ZN(new_n1611_));
  XNOR2_X1   g1562(.A1(new_n684_), .A2(new_n688_), .ZN(new_n1612_));
  OAI21_X1   g1563(.A1(new_n689_), .A2(new_n705_), .B(new_n704_), .ZN(new_n1613_));
  OAI21_X1   g1564(.A1(new_n704_), .A2(new_n1612_), .B(new_n1613_), .ZN(new_n1614_));
  INV_X1     g1565(.I(new_n1614_), .ZN(new_n1615_));
  XOR2_X1    g1566(.A1(new_n1611_), .A2(new_n1615_), .Z(new_n1616_));
  OAI22_X1   g1567(.A1(new_n1606_), .A2(new_n1571_), .B1(new_n1609_), .B2(new_n1605_), .ZN(new_n1617_));
  XOR2_X1    g1568(.A1(new_n1600_), .A2(new_n1604_), .Z(new_n1618_));
  NAND2_X1   g1569(.A1(new_n1607_), .A2(new_n1618_), .ZN(new_n1619_));
  NAND2_X1   g1570(.A1(new_n1619_), .A2(new_n1617_), .ZN(new_n1620_));
  NAND2_X1   g1571(.A1(new_n1616_), .A2(new_n1620_), .ZN(new_n1621_));
  NAND3_X1   g1572(.A1(new_n1594_), .A2(new_n1596_), .A3(new_n1621_), .ZN(new_n1622_));
  NAND2_X1   g1573(.A1(new_n1611_), .A2(new_n1614_), .ZN(new_n1623_));
  NAND3_X1   g1574(.A1(new_n1622_), .A2(new_n708_), .A3(new_n1623_), .ZN(new_n1624_));
  NOR2_X1    g1575(.A1(new_n669_), .A2(new_n630_), .ZN(new_n1625_));
  NOR2_X1    g1576(.A1(new_n669_), .A2(new_n668_), .ZN(new_n1626_));
  NOR2_X1    g1577(.A1(new_n1625_), .A2(new_n1626_), .ZN(new_n1627_));
  XOR2_X1    g1578(.A1(new_n658_), .A2(new_n667_), .Z(new_n1628_));
  AOI21_X1   g1579(.A1(new_n674_), .A2(new_n1628_), .B(new_n628_), .ZN(new_n1629_));
  OAI21_X1   g1580(.A1(new_n674_), .A2(new_n1628_), .B(new_n1629_), .ZN(new_n1630_));
  XOR2_X1    g1581(.A1(new_n1627_), .A2(new_n1630_), .Z(new_n1631_));
  AOI21_X1   g1582(.A1(new_n1624_), .A2(new_n709_), .B(new_n1631_), .ZN(new_n1632_));
  XOR2_X1    g1583(.A1(new_n1627_), .A2(new_n1630_), .Z(new_n1633_));
  AND3_X2    g1584(.A1(new_n1624_), .A2(new_n709_), .A3(new_n1633_), .Z(new_n1634_));
  NOR2_X1    g1585(.A1(new_n1634_), .A2(new_n1632_), .ZN(new_n1635_));
  INV_X1     g1586(.I(new_n1635_), .ZN(new_n1636_));
  NAND2_X1   g1587(.A1(new_n1636_), .A2(new_n355_), .ZN(new_n1637_));
  XOR2_X1    g1588(.A1(new_n1635_), .A2(new_n355_), .Z(new_n1638_));
  NOR4_X1    g1589(.A1(new_n974_), .A2(new_n631_), .A3(new_n747_), .A4(new_n534_), .ZN(new_n1639_));
  NOR4_X1    g1590(.A1(new_n1639_), .A2(new_n369_), .A3(new_n376_), .A4(new_n801_), .ZN(new_n1640_));
  NOR4_X1    g1591(.A1(new_n588_), .A2(new_n437_), .A3(new_n593_), .A4(new_n717_), .ZN(new_n1641_));
  NOR2_X1    g1592(.A1(new_n1641_), .A2(new_n527_), .ZN(new_n1642_));
  AND3_X2    g1593(.A1(new_n1640_), .A2(new_n491_), .A3(new_n1642_), .Z(new_n1643_));
  NOR4_X1    g1594(.A1(new_n239_), .A2(new_n263_), .A3(new_n377_), .A4(new_n561_), .ZN(new_n1644_));
  NAND2_X1   g1595(.A1(new_n308_), .A2(new_n1644_), .ZN(new_n1645_));
  NOR3_X1    g1596(.A1(new_n385_), .A2(new_n595_), .A3(new_n267_), .ZN(new_n1646_));
  INV_X1     g1597(.I(new_n1646_), .ZN(new_n1647_));
  NOR2_X1    g1598(.A1(new_n741_), .A2(new_n322_), .ZN(new_n1648_));
  INV_X1     g1599(.I(new_n1648_), .ZN(new_n1649_));
  NOR3_X1    g1600(.A1(new_n1649_), .A2(new_n515_), .A3(new_n890_), .ZN(new_n1650_));
  NOR2_X1    g1601(.A1(new_n1090_), .A2(new_n394_), .ZN(new_n1651_));
  NAND4_X1   g1602(.A1(new_n182_), .A2(new_n350_), .A3(new_n554_), .A4(new_n1651_), .ZN(new_n1652_));
  NOR4_X1    g1603(.A1(new_n1652_), .A2(new_n1645_), .A3(new_n1647_), .A4(new_n1650_), .ZN(new_n1653_));
  INV_X1     g1604(.I(new_n486_), .ZN(new_n1654_));
  NOR3_X1    g1605(.A1(new_n257_), .A2(new_n326_), .A3(new_n518_), .ZN(new_n1655_));
  NAND3_X1   g1606(.A1(new_n1655_), .A2(new_n390_), .A3(new_n564_), .ZN(new_n1656_));
  NOR3_X1    g1607(.A1(new_n398_), .A2(new_n520_), .A3(new_n461_), .ZN(new_n1657_));
  INV_X1     g1608(.I(new_n1657_), .ZN(new_n1658_));
  NAND4_X1   g1609(.A1(new_n317_), .A2(new_n294_), .A3(new_n727_), .A4(new_n551_), .ZN(new_n1659_));
  NOR4_X1    g1610(.A1(new_n1654_), .A2(new_n1656_), .A3(new_n1658_), .A4(new_n1659_), .ZN(new_n1660_));
  NAND3_X1   g1611(.A1(new_n1653_), .A2(new_n1643_), .A3(new_n1660_), .ZN(new_n1661_));
  INV_X1     g1612(.I(new_n1661_), .ZN(new_n1662_));
  XOR2_X1    g1613(.A1(new_n1596_), .A2(new_n1620_), .Z(new_n1663_));
  NAND2_X1   g1614(.A1(new_n1594_), .A2(new_n1663_), .ZN(new_n1664_));
  INV_X1     g1615(.I(new_n1664_), .ZN(new_n1665_));
  XOR2_X1    g1616(.A1(new_n1596_), .A2(new_n1620_), .Z(new_n1666_));
  NOR2_X1    g1617(.A1(new_n1594_), .A2(new_n1666_), .ZN(new_n1667_));
  NOR2_X1    g1618(.A1(new_n1665_), .A2(new_n1667_), .ZN(new_n1668_));
  NOR2_X1    g1619(.A1(new_n1668_), .A2(new_n1662_), .ZN(new_n1669_));
  INV_X1     g1620(.I(new_n1669_), .ZN(new_n1670_));
  NAND2_X1   g1621(.A1(new_n1551_), .A2(new_n1527_), .ZN(new_n1671_));
  NAND2_X1   g1622(.A1(new_n1441_), .A2(new_n1444_), .ZN(new_n1672_));
  XOR2_X1    g1623(.A1(new_n1672_), .A2(new_n1671_), .Z(new_n1673_));
  NAND3_X1   g1624(.A1(new_n1549_), .A2(new_n1308_), .A3(new_n1444_), .ZN(new_n1674_));
  NAND2_X1   g1625(.A1(new_n1441_), .A2(new_n1443_), .ZN(new_n1675_));
  AOI21_X1   g1626(.A1(new_n1675_), .A2(new_n1674_), .B(new_n1486_), .ZN(new_n1676_));
  NAND2_X1   g1627(.A1(new_n1673_), .A2(new_n1676_), .ZN(new_n1677_));
  INV_X1     g1628(.I(new_n1677_), .ZN(new_n1678_));
  NOR2_X1    g1629(.A1(new_n1673_), .A2(new_n1676_), .ZN(new_n1679_));
  NOR3_X1    g1630(.A1(new_n808_), .A2(new_n209_), .A3(new_n856_), .ZN(new_n1680_));
  INV_X1     g1631(.I(new_n827_), .ZN(new_n1681_));
  NOR4_X1    g1632(.A1(new_n301_), .A2(new_n369_), .A3(new_n278_), .A4(new_n361_), .ZN(new_n1682_));
  NAND4_X1   g1633(.A1(new_n193_), .A2(new_n564_), .A3(new_n429_), .A4(new_n922_), .ZN(new_n1683_));
  NOR3_X1    g1634(.A1(new_n1681_), .A2(new_n1683_), .A3(new_n1682_), .ZN(new_n1684_));
  NOR4_X1    g1635(.A1(new_n1090_), .A2(new_n172_), .A3(new_n1091_), .A4(new_n424_), .ZN(new_n1685_));
  NOR4_X1    g1636(.A1(new_n588_), .A2(new_n1021_), .A3(new_n311_), .A4(new_n437_), .ZN(new_n1686_));
  NOR2_X1    g1637(.A1(new_n1686_), .A2(new_n1685_), .ZN(new_n1687_));
  INV_X1     g1638(.I(new_n1687_), .ZN(new_n1688_));
  NAND2_X1   g1639(.A1(new_n532_), .A2(new_n559_), .ZN(new_n1689_));
  NOR4_X1    g1640(.A1(new_n1689_), .A2(new_n181_), .A3(new_n238_), .A4(new_n873_), .ZN(new_n1690_));
  INV_X1     g1641(.I(new_n1690_), .ZN(new_n1691_));
  NOR4_X1    g1642(.A1(new_n595_), .A2(new_n335_), .A3(new_n473_), .A4(new_n832_), .ZN(new_n1692_));
  NOR4_X1    g1643(.A1(new_n305_), .A2(new_n339_), .A3(new_n584_), .A4(new_n384_), .ZN(new_n1693_));
  NOR4_X1    g1644(.A1(new_n1688_), .A2(new_n1691_), .A3(new_n1692_), .A4(new_n1693_), .ZN(new_n1694_));
  NAND3_X1   g1645(.A1(new_n1680_), .A2(new_n1684_), .A3(new_n1694_), .ZN(new_n1695_));
  INV_X1     g1646(.I(new_n1695_), .ZN(new_n1696_));
  NOR3_X1    g1647(.A1(new_n1678_), .A2(new_n1679_), .A3(new_n1696_), .ZN(new_n1697_));
  NOR2_X1    g1648(.A1(new_n238_), .A2(new_n424_), .ZN(new_n1698_));
  INV_X1     g1649(.I(new_n1698_), .ZN(new_n1699_));
  NOR3_X1    g1650(.A1(new_n1699_), .A2(new_n289_), .A3(new_n612_), .ZN(new_n1700_));
  NOR2_X1    g1651(.A1(new_n520_), .A2(new_n717_), .ZN(new_n1701_));
  INV_X1     g1652(.I(new_n1701_), .ZN(new_n1702_));
  NAND2_X1   g1653(.A1(new_n223_), .A2(new_n929_), .ZN(new_n1703_));
  NOR4_X1    g1654(.A1(new_n1702_), .A2(new_n1703_), .A3(new_n563_), .A4(new_n1091_), .ZN(new_n1704_));
  NAND4_X1   g1655(.A1(new_n812_), .A2(new_n1071_), .A3(new_n1704_), .A4(new_n1700_), .ZN(new_n1705_));
  INV_X1     g1656(.I(new_n329_), .ZN(new_n1706_));
  NOR4_X1    g1657(.A1(new_n1706_), .A2(new_n873_), .A3(new_n525_), .A4(new_n856_), .ZN(new_n1707_));
  NOR4_X1    g1658(.A1(new_n1707_), .A2(new_n732_), .A3(new_n805_), .A4(new_n815_), .ZN(new_n1708_));
  INV_X1     g1659(.I(new_n1708_), .ZN(new_n1709_));
  NOR3_X1    g1660(.A1(new_n510_), .A2(new_n394_), .A3(new_n488_), .ZN(new_n1710_));
  NOR4_X1    g1661(.A1(new_n610_), .A2(new_n181_), .A3(new_n594_), .A4(new_n643_), .ZN(new_n1711_));
  NOR3_X1    g1662(.A1(new_n801_), .A2(new_n209_), .A3(new_n280_), .ZN(new_n1712_));
  NAND4_X1   g1663(.A1(new_n1712_), .A2(new_n1074_), .A3(new_n1710_), .A4(new_n1711_), .ZN(new_n1713_));
  NOR4_X1    g1664(.A1(new_n1705_), .A2(new_n1070_), .A3(new_n1709_), .A4(new_n1713_), .ZN(new_n1714_));
  INV_X1     g1665(.I(new_n1714_), .ZN(new_n1715_));
  XNOR2_X1   g1666(.A1(new_n1486_), .A2(new_n1443_), .ZN(new_n1716_));
  AOI21_X1   g1667(.A1(new_n1549_), .A2(new_n1308_), .B(new_n1716_), .ZN(new_n1717_));
  AOI21_X1   g1668(.A1(new_n1489_), .A2(new_n1552_), .B(new_n1441_), .ZN(new_n1718_));
  NOR2_X1    g1669(.A1(new_n1718_), .A2(new_n1717_), .ZN(new_n1719_));
  INV_X1     g1670(.I(new_n1719_), .ZN(new_n1720_));
  INV_X1     g1671(.I(new_n567_), .ZN(new_n1721_));
  NAND3_X1   g1672(.A1(new_n1721_), .A2(new_n1326_), .A3(new_n494_), .ZN(new_n1722_));
  OAI21_X1   g1673(.A1(new_n1721_), .A2(new_n1326_), .B(new_n1120_), .ZN(new_n1723_));
  NAND2_X1   g1674(.A1(new_n1723_), .A2(new_n1722_), .ZN(new_n1724_));
  NAND2_X1   g1675(.A1(new_n1321_), .A2(new_n581_), .ZN(new_n1725_));
  OAI21_X1   g1676(.A1(new_n1321_), .A2(new_n576_), .B(new_n937_), .ZN(new_n1726_));
  XOR2_X1    g1677(.A1(new_n1726_), .A2(new_n1725_), .Z(new_n1727_));
  NAND3_X1   g1678(.A1(new_n1724_), .A2(new_n1727_), .A3(new_n416_), .ZN(new_n1728_));
  NOR2_X1    g1679(.A1(new_n1231_), .A2(new_n1125_), .ZN(new_n1729_));
  NOR2_X1    g1680(.A1(new_n1100_), .A2(new_n1126_), .ZN(new_n1730_));
  NOR2_X1    g1681(.A1(new_n1729_), .A2(new_n1730_), .ZN(new_n1731_));
  INV_X1     g1682(.I(new_n1110_), .ZN(new_n1732_));
  NAND2_X1   g1683(.A1(new_n1732_), .A2(new_n1134_), .ZN(new_n1733_));
  NAND2_X1   g1684(.A1(new_n1114_), .A2(new_n1132_), .ZN(new_n1734_));
  NAND3_X1   g1685(.A1(new_n1731_), .A2(new_n1733_), .A3(new_n1734_), .ZN(new_n1735_));
  NAND2_X1   g1686(.A1(new_n1735_), .A2(new_n1728_), .ZN(new_n1736_));
  NAND3_X1   g1687(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n1062_), .ZN(new_n1737_));
  NOR2_X1    g1688(.A1(new_n793_), .A2(new_n939_), .ZN(new_n1738_));
  NOR2_X1    g1689(.A1(new_n795_), .A2(new_n1171_), .ZN(new_n1739_));
  NOR3_X1    g1690(.A1(new_n1737_), .A2(new_n1738_), .A3(new_n1739_), .ZN(new_n1740_));
  NOR2_X1    g1691(.A1(new_n1735_), .A2(new_n1728_), .ZN(new_n1741_));
  OAI21_X1   g1692(.A1(new_n1740_), .A2(new_n1741_), .B(new_n1736_), .ZN(new_n1742_));
  INV_X1     g1693(.I(new_n1742_), .ZN(new_n1743_));
  NOR3_X1    g1694(.A1(new_n1032_), .A2(new_n1034_), .A3(new_n1106_), .ZN(new_n1744_));
  INV_X1     g1695(.I(new_n1744_), .ZN(new_n1745_));
  NAND2_X1   g1696(.A1(new_n1035_), .A2(new_n576_), .ZN(new_n1746_));
  OAI21_X1   g1697(.A1(new_n576_), .A2(new_n1037_), .B(new_n1746_), .ZN(new_n1747_));
  NOR2_X1    g1698(.A1(new_n1745_), .A2(new_n1747_), .ZN(new_n1748_));
  NOR2_X1    g1699(.A1(new_n1027_), .A2(new_n678_), .ZN(new_n1749_));
  OAI21_X1   g1700(.A1(new_n1321_), .A2(new_n582_), .B(new_n937_), .ZN(new_n1750_));
  XOR2_X1    g1701(.A1(new_n1749_), .A2(new_n1750_), .Z(new_n1751_));
  INV_X1     g1702(.I(new_n1751_), .ZN(new_n1752_));
  NOR2_X1    g1703(.A1(new_n1748_), .A2(new_n1752_), .ZN(new_n1753_));
  NOR2_X1    g1704(.A1(new_n1047_), .A2(new_n62_), .ZN(new_n1754_));
  XOR2_X1    g1705(.A1(new_n494_), .A2(new_n56_), .Z(new_n1755_));
  NOR2_X1    g1706(.A1(new_n1055_), .A2(new_n1755_), .ZN(new_n1756_));
  NAND2_X1   g1707(.A1(new_n690_), .A2(new_n943_), .ZN(new_n1757_));
  NOR4_X1    g1708(.A1(new_n1754_), .A2(new_n1061_), .A3(new_n1756_), .A4(new_n1757_), .ZN(new_n1758_));
  NOR3_X1    g1709(.A1(new_n1747_), .A2(new_n1751_), .A3(new_n1745_), .ZN(new_n1759_));
  NOR2_X1    g1710(.A1(new_n1758_), .A2(new_n1759_), .ZN(new_n1760_));
  NOR2_X1    g1711(.A1(new_n1760_), .A2(new_n1753_), .ZN(new_n1761_));
  INV_X1     g1712(.I(new_n1761_), .ZN(new_n1762_));
  NOR2_X1    g1713(.A1(new_n1391_), .A2(new_n1382_), .ZN(new_n1763_));
  INV_X1     g1714(.I(new_n1763_), .ZN(new_n1764_));
  NAND2_X1   g1715(.A1(new_n1391_), .A2(new_n1382_), .ZN(new_n1765_));
  AOI21_X1   g1716(.A1(new_n1764_), .A2(new_n1765_), .B(new_n1386_), .ZN(new_n1766_));
  NOR3_X1    g1717(.A1(new_n1061_), .A2(new_n1381_), .A3(new_n1380_), .ZN(new_n1767_));
  OAI21_X1   g1718(.A1(new_n939_), .A2(new_n1047_), .B(new_n1767_), .ZN(new_n1768_));
  NOR2_X1    g1719(.A1(new_n1768_), .A2(new_n1391_), .ZN(new_n1769_));
  INV_X1     g1720(.I(new_n1769_), .ZN(new_n1770_));
  NAND2_X1   g1721(.A1(new_n1768_), .A2(new_n1391_), .ZN(new_n1771_));
  AOI21_X1   g1722(.A1(new_n1770_), .A2(new_n1771_), .B(new_n1397_), .ZN(new_n1772_));
  OAI21_X1   g1723(.A1(new_n1772_), .A2(new_n1766_), .B(new_n1762_), .ZN(new_n1773_));
  INV_X1     g1724(.I(new_n1765_), .ZN(new_n1774_));
  OAI21_X1   g1725(.A1(new_n1774_), .A2(new_n1763_), .B(new_n1397_), .ZN(new_n1775_));
  INV_X1     g1726(.I(new_n1771_), .ZN(new_n1776_));
  OAI21_X1   g1727(.A1(new_n1776_), .A2(new_n1769_), .B(new_n1386_), .ZN(new_n1777_));
  NAND3_X1   g1728(.A1(new_n1777_), .A2(new_n1775_), .A3(new_n1761_), .ZN(new_n1778_));
  AOI21_X1   g1729(.A1(new_n1773_), .A2(new_n1778_), .B(new_n1743_), .ZN(new_n1779_));
  OAI21_X1   g1730(.A1(new_n1772_), .A2(new_n1766_), .B(new_n1761_), .ZN(new_n1780_));
  NAND3_X1   g1731(.A1(new_n1777_), .A2(new_n1775_), .A3(new_n1762_), .ZN(new_n1781_));
  AOI21_X1   g1732(.A1(new_n1780_), .A2(new_n1781_), .B(new_n1742_), .ZN(new_n1782_));
  NOR2_X1    g1733(.A1(new_n1779_), .A2(new_n1782_), .ZN(new_n1783_));
  XNOR2_X1   g1734(.A1(new_n1329_), .A2(new_n1335_), .ZN(new_n1784_));
  NOR2_X1    g1735(.A1(new_n1784_), .A2(new_n1343_), .ZN(new_n1785_));
  NOR2_X1    g1736(.A1(new_n1337_), .A2(new_n1344_), .ZN(new_n1786_));
  NOR2_X1    g1737(.A1(new_n1786_), .A2(new_n1342_), .ZN(new_n1787_));
  NOR2_X1    g1738(.A1(new_n1787_), .A2(new_n1785_), .ZN(new_n1788_));
  NOR2_X1    g1739(.A1(new_n1783_), .A2(new_n1788_), .ZN(new_n1789_));
  INV_X1     g1740(.I(new_n1740_), .ZN(new_n1790_));
  INV_X1     g1741(.I(new_n1741_), .ZN(new_n1791_));
  AOI21_X1   g1742(.A1(new_n1791_), .A2(new_n1736_), .B(new_n1790_), .ZN(new_n1792_));
  NAND4_X1   g1743(.A1(new_n1731_), .A2(new_n1728_), .A3(new_n1733_), .A4(new_n1734_), .ZN(new_n1793_));
  INV_X1     g1744(.I(new_n1728_), .ZN(new_n1794_));
  NAND2_X1   g1745(.A1(new_n1735_), .A2(new_n1794_), .ZN(new_n1795_));
  AOI21_X1   g1746(.A1(new_n1795_), .A2(new_n1793_), .B(new_n1740_), .ZN(new_n1796_));
  NOR2_X1    g1747(.A1(new_n651_), .A2(new_n1326_), .ZN(new_n1797_));
  NOR3_X1    g1748(.A1(new_n1792_), .A2(new_n1796_), .A3(new_n1797_), .ZN(new_n1798_));
  NOR2_X1    g1749(.A1(new_n1231_), .A2(new_n1132_), .ZN(new_n1799_));
  AOI21_X1   g1750(.A1(new_n1230_), .A2(new_n1132_), .B(new_n1799_), .ZN(new_n1800_));
  NOR2_X1    g1751(.A1(new_n1110_), .A2(new_n1053_), .ZN(new_n1801_));
  AOI21_X1   g1752(.A1(new_n1053_), .A2(new_n1114_), .B(new_n1801_), .ZN(new_n1802_));
  NAND2_X1   g1753(.A1(new_n1800_), .A2(new_n1802_), .ZN(new_n1803_));
  NOR3_X1    g1754(.A1(new_n1032_), .A2(new_n1034_), .A3(new_n1125_), .ZN(new_n1804_));
  INV_X1     g1755(.I(new_n1804_), .ZN(new_n1805_));
  NAND2_X1   g1756(.A1(new_n1035_), .A2(new_n1153_), .ZN(new_n1806_));
  OAI21_X1   g1757(.A1(new_n1037_), .A2(new_n1153_), .B(new_n1806_), .ZN(new_n1807_));
  OR2_X2     g1758(.A1(new_n1805_), .A2(new_n1807_), .Z(new_n1808_));
  NAND2_X1   g1759(.A1(new_n1803_), .A2(new_n1808_), .ZN(new_n1809_));
  NAND3_X1   g1760(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n1171_), .ZN(new_n1810_));
  NAND2_X1   g1761(.A1(new_n1270_), .A2(new_n943_), .ZN(new_n1811_));
  INV_X1     g1762(.I(new_n1811_), .ZN(new_n1812_));
  NOR2_X1    g1763(.A1(new_n795_), .A2(new_n943_), .ZN(new_n1813_));
  NOR3_X1    g1764(.A1(new_n1812_), .A2(new_n1810_), .A3(new_n1813_), .ZN(new_n1814_));
  INV_X1     g1765(.I(new_n1814_), .ZN(new_n1815_));
  INV_X1     g1766(.I(new_n1808_), .ZN(new_n1816_));
  NAND3_X1   g1767(.A1(new_n1800_), .A2(new_n1816_), .A3(new_n1802_), .ZN(new_n1817_));
  NAND2_X1   g1768(.A1(new_n1815_), .A2(new_n1817_), .ZN(new_n1818_));
  NAND2_X1   g1769(.A1(new_n1818_), .A2(new_n1809_), .ZN(new_n1819_));
  OAI21_X1   g1770(.A1(new_n1792_), .A2(new_n1796_), .B(new_n1797_), .ZN(new_n1820_));
  AOI21_X1   g1771(.A1(new_n1819_), .A2(new_n1820_), .B(new_n1798_), .ZN(new_n1821_));
  AOI21_X1   g1772(.A1(new_n1783_), .A2(new_n1788_), .B(new_n1821_), .ZN(new_n1822_));
  INV_X1     g1773(.I(new_n1312_), .ZN(new_n1823_));
  AOI21_X1   g1774(.A1(new_n1823_), .A2(new_n1313_), .B(new_n1137_), .ZN(new_n1824_));
  NAND2_X1   g1775(.A1(new_n1316_), .A2(new_n1116_), .ZN(new_n1825_));
  AOI21_X1   g1776(.A1(new_n1138_), .A2(new_n1825_), .B(new_n1136_), .ZN(new_n1826_));
  NOR3_X1    g1777(.A1(new_n1824_), .A2(new_n1826_), .A3(new_n1310_), .ZN(new_n1827_));
  OAI21_X1   g1778(.A1(new_n1319_), .A2(new_n1827_), .B(new_n1347_), .ZN(new_n1828_));
  AOI21_X1   g1779(.A1(new_n1318_), .A2(new_n1315_), .B(new_n1310_), .ZN(new_n1829_));
  NOR3_X1    g1780(.A1(new_n1824_), .A2(new_n1826_), .A3(new_n1311_), .ZN(new_n1830_));
  OAI21_X1   g1781(.A1(new_n1829_), .A2(new_n1830_), .B(new_n1346_), .ZN(new_n1831_));
  NAND2_X1   g1782(.A1(new_n1828_), .A2(new_n1831_), .ZN(new_n1832_));
  NAND2_X1   g1783(.A1(new_n1382_), .A2(new_n1397_), .ZN(new_n1833_));
  NOR3_X1    g1784(.A1(new_n1374_), .A2(new_n1833_), .A3(new_n1375_), .ZN(new_n1834_));
  NOR2_X1    g1785(.A1(new_n1768_), .A2(new_n1386_), .ZN(new_n1835_));
  NOR2_X1    g1786(.A1(new_n1376_), .A2(new_n1835_), .ZN(new_n1836_));
  NOR2_X1    g1787(.A1(new_n1768_), .A2(new_n1397_), .ZN(new_n1837_));
  NOR2_X1    g1788(.A1(new_n1382_), .A2(new_n1386_), .ZN(new_n1838_));
  OAI21_X1   g1789(.A1(new_n1837_), .A2(new_n1838_), .B(new_n1398_), .ZN(new_n1839_));
  NOR3_X1    g1790(.A1(new_n1836_), .A2(new_n1839_), .A3(new_n1834_), .ZN(new_n1840_));
  INV_X1     g1791(.I(new_n1375_), .ZN(new_n1841_));
  NAND3_X1   g1792(.A1(new_n1835_), .A2(new_n1841_), .A3(new_n1373_), .ZN(new_n1842_));
  OAI21_X1   g1793(.A1(new_n1374_), .A2(new_n1375_), .B(new_n1833_), .ZN(new_n1843_));
  OR2_X2     g1794(.A1(new_n1837_), .A2(new_n1838_), .Z(new_n1844_));
  AOI22_X1   g1795(.A1(new_n1844_), .A2(new_n1398_), .B1(new_n1842_), .B2(new_n1843_), .ZN(new_n1845_));
  NAND2_X1   g1796(.A1(new_n1762_), .A2(new_n1742_), .ZN(new_n1846_));
  NOR3_X1    g1797(.A1(new_n1845_), .A2(new_n1840_), .A3(new_n1846_), .ZN(new_n1847_));
  NAND4_X1   g1798(.A1(new_n1844_), .A2(new_n1398_), .A3(new_n1842_), .A4(new_n1843_), .ZN(new_n1848_));
  OAI21_X1   g1799(.A1(new_n1836_), .A2(new_n1834_), .B(new_n1839_), .ZN(new_n1849_));
  INV_X1     g1800(.I(new_n1846_), .ZN(new_n1850_));
  AOI21_X1   g1801(.A1(new_n1848_), .A2(new_n1849_), .B(new_n1850_), .ZN(new_n1851_));
  NOR2_X1    g1802(.A1(new_n1742_), .A2(new_n1761_), .ZN(new_n1852_));
  NAND2_X1   g1803(.A1(new_n1742_), .A2(new_n1761_), .ZN(new_n1853_));
  INV_X1     g1804(.I(new_n1853_), .ZN(new_n1854_));
  OAI22_X1   g1805(.A1(new_n1854_), .A2(new_n1852_), .B1(new_n1766_), .B2(new_n1772_), .ZN(new_n1855_));
  NOR3_X1    g1806(.A1(new_n1851_), .A2(new_n1847_), .A3(new_n1855_), .ZN(new_n1856_));
  NAND3_X1   g1807(.A1(new_n1850_), .A2(new_n1849_), .A3(new_n1848_), .ZN(new_n1857_));
  OAI21_X1   g1808(.A1(new_n1845_), .A2(new_n1840_), .B(new_n1846_), .ZN(new_n1858_));
  INV_X1     g1809(.I(new_n1852_), .ZN(new_n1859_));
  AOI22_X1   g1810(.A1(new_n1859_), .A2(new_n1853_), .B1(new_n1775_), .B2(new_n1777_), .ZN(new_n1860_));
  AOI21_X1   g1811(.A1(new_n1857_), .A2(new_n1858_), .B(new_n1860_), .ZN(new_n1861_));
  NOR3_X1    g1812(.A1(new_n1856_), .A2(new_n1861_), .A3(new_n1832_), .ZN(new_n1862_));
  OAI21_X1   g1813(.A1(new_n1824_), .A2(new_n1826_), .B(new_n1310_), .ZN(new_n1863_));
  AOI21_X1   g1814(.A1(new_n1863_), .A2(new_n1348_), .B(new_n1346_), .ZN(new_n1864_));
  OAI21_X1   g1815(.A1(new_n1824_), .A2(new_n1826_), .B(new_n1311_), .ZN(new_n1865_));
  NAND3_X1   g1816(.A1(new_n1318_), .A2(new_n1315_), .A3(new_n1310_), .ZN(new_n1866_));
  AOI21_X1   g1817(.A1(new_n1865_), .A2(new_n1866_), .B(new_n1347_), .ZN(new_n1867_));
  NOR2_X1    g1818(.A1(new_n1864_), .A2(new_n1867_), .ZN(new_n1868_));
  NAND3_X1   g1819(.A1(new_n1857_), .A2(new_n1858_), .A3(new_n1860_), .ZN(new_n1869_));
  OAI21_X1   g1820(.A1(new_n1851_), .A2(new_n1847_), .B(new_n1855_), .ZN(new_n1870_));
  AOI21_X1   g1821(.A1(new_n1870_), .A2(new_n1869_), .B(new_n1868_), .ZN(new_n1871_));
  NOR4_X1    g1822(.A1(new_n1862_), .A2(new_n1871_), .A3(new_n1789_), .A4(new_n1822_), .ZN(new_n1872_));
  AOI21_X1   g1823(.A1(new_n1777_), .A2(new_n1775_), .B(new_n1761_), .ZN(new_n1873_));
  NOR3_X1    g1824(.A1(new_n1772_), .A2(new_n1766_), .A3(new_n1762_), .ZN(new_n1874_));
  OAI21_X1   g1825(.A1(new_n1873_), .A2(new_n1874_), .B(new_n1742_), .ZN(new_n1875_));
  AOI21_X1   g1826(.A1(new_n1777_), .A2(new_n1775_), .B(new_n1762_), .ZN(new_n1876_));
  NOR3_X1    g1827(.A1(new_n1772_), .A2(new_n1766_), .A3(new_n1761_), .ZN(new_n1877_));
  OAI21_X1   g1828(.A1(new_n1876_), .A2(new_n1877_), .B(new_n1743_), .ZN(new_n1878_));
  NAND2_X1   g1829(.A1(new_n1875_), .A2(new_n1878_), .ZN(new_n1879_));
  INV_X1     g1830(.I(new_n1788_), .ZN(new_n1880_));
  NAND2_X1   g1831(.A1(new_n1879_), .A2(new_n1880_), .ZN(new_n1881_));
  INV_X1     g1832(.I(new_n1821_), .ZN(new_n1882_));
  OAI21_X1   g1833(.A1(new_n1879_), .A2(new_n1880_), .B(new_n1882_), .ZN(new_n1883_));
  NAND3_X1   g1834(.A1(new_n1870_), .A2(new_n1869_), .A3(new_n1868_), .ZN(new_n1884_));
  OAI21_X1   g1835(.A1(new_n1856_), .A2(new_n1861_), .B(new_n1832_), .ZN(new_n1885_));
  AOI22_X1   g1836(.A1(new_n1885_), .A2(new_n1884_), .B1(new_n1881_), .B2(new_n1883_), .ZN(new_n1886_));
  NOR2_X1    g1837(.A1(new_n1886_), .A2(new_n1872_), .ZN(new_n1887_));
  NAND2_X1   g1838(.A1(new_n1098_), .A2(new_n1062_), .ZN(new_n1888_));
  NAND2_X1   g1839(.A1(new_n1230_), .A2(new_n1053_), .ZN(new_n1889_));
  NAND2_X1   g1840(.A1(new_n1732_), .A2(new_n1171_), .ZN(new_n1890_));
  NAND2_X1   g1841(.A1(new_n1114_), .A2(new_n939_), .ZN(new_n1891_));
  NAND4_X1   g1842(.A1(new_n1890_), .A2(new_n1888_), .A3(new_n1889_), .A4(new_n1891_), .ZN(new_n1892_));
  NAND3_X1   g1843(.A1(new_n1031_), .A2(new_n1033_), .A3(new_n1134_), .ZN(new_n1893_));
  NAND2_X1   g1844(.A1(new_n1035_), .A2(new_n1126_), .ZN(new_n1894_));
  OAI21_X1   g1845(.A1(new_n1037_), .A2(new_n1126_), .B(new_n1894_), .ZN(new_n1895_));
  NOR2_X1    g1846(.A1(new_n1895_), .A2(new_n1893_), .ZN(new_n1896_));
  NOR2_X1    g1847(.A1(new_n1027_), .A2(new_n576_), .ZN(new_n1897_));
  OAI21_X1   g1848(.A1(new_n1321_), .A2(new_n1153_), .B(new_n937_), .ZN(new_n1898_));
  XOR2_X1    g1849(.A1(new_n1897_), .A2(new_n1898_), .Z(new_n1899_));
  INV_X1     g1850(.I(new_n1899_), .ZN(new_n1900_));
  NAND2_X1   g1851(.A1(new_n1896_), .A2(new_n1900_), .ZN(new_n1901_));
  NOR2_X1    g1852(.A1(new_n1896_), .A2(new_n1900_), .ZN(new_n1902_));
  INV_X1     g1853(.I(new_n1902_), .ZN(new_n1903_));
  AOI21_X1   g1854(.A1(new_n1903_), .A2(new_n1901_), .B(new_n1892_), .ZN(new_n1904_));
  INV_X1     g1855(.I(new_n1892_), .ZN(new_n1905_));
  XOR2_X1    g1856(.A1(new_n1896_), .A2(new_n1899_), .Z(new_n1906_));
  NOR2_X1    g1857(.A1(new_n1906_), .A2(new_n1905_), .ZN(new_n1907_));
  NOR2_X1    g1858(.A1(new_n1907_), .A2(new_n1904_), .ZN(new_n1908_));
  NAND2_X1   g1859(.A1(new_n1098_), .A2(new_n1171_), .ZN(new_n1909_));
  NAND2_X1   g1860(.A1(new_n1230_), .A2(new_n939_), .ZN(new_n1910_));
  NOR2_X1    g1861(.A1(new_n1110_), .A2(new_n62_), .ZN(new_n1911_));
  NOR3_X1    g1862(.A1(new_n1113_), .A2(new_n943_), .A3(new_n1112_), .ZN(new_n1912_));
  NOR2_X1    g1863(.A1(new_n1911_), .A2(new_n1912_), .ZN(new_n1913_));
  NAND3_X1   g1864(.A1(new_n1913_), .A2(new_n1909_), .A3(new_n1910_), .ZN(new_n1914_));
  NAND3_X1   g1865(.A1(new_n1031_), .A2(new_n1033_), .A3(new_n1062_), .ZN(new_n1915_));
  NAND2_X1   g1866(.A1(new_n1035_), .A2(new_n1134_), .ZN(new_n1916_));
  OAI21_X1   g1867(.A1(new_n1037_), .A2(new_n1134_), .B(new_n1916_), .ZN(new_n1917_));
  NOR2_X1    g1868(.A1(new_n1917_), .A2(new_n1915_), .ZN(new_n1918_));
  INV_X1     g1869(.I(new_n1918_), .ZN(new_n1919_));
  NAND2_X1   g1870(.A1(new_n1914_), .A2(new_n1919_), .ZN(new_n1920_));
  XNOR2_X1   g1871(.A1(new_n778_), .A2(new_n494_), .ZN(new_n1921_));
  XOR2_X1    g1872(.A1(new_n752_), .A2(new_n67_), .Z(new_n1922_));
  NOR2_X1    g1873(.A1(new_n1921_), .A2(new_n1922_), .ZN(new_n1923_));
  NOR2_X1    g1874(.A1(new_n1119_), .A2(new_n56_), .ZN(new_n1924_));
  NAND2_X1   g1875(.A1(new_n1498_), .A2(new_n1176_), .ZN(new_n1925_));
  NOR4_X1    g1876(.A1(new_n1924_), .A2(new_n787_), .A3(new_n1923_), .A4(new_n1925_), .ZN(new_n1926_));
  NOR2_X1    g1877(.A1(new_n1914_), .A2(new_n1919_), .ZN(new_n1927_));
  OAI21_X1   g1878(.A1(new_n1926_), .A2(new_n1927_), .B(new_n1920_), .ZN(new_n1928_));
  NAND2_X1   g1879(.A1(new_n1908_), .A2(new_n1928_), .ZN(new_n1929_));
  NAND3_X1   g1880(.A1(new_n1122_), .A2(new_n1119_), .A3(new_n943_), .ZN(new_n1930_));
  NOR2_X1    g1881(.A1(new_n793_), .A2(new_n56_), .ZN(new_n1931_));
  NOR2_X1    g1882(.A1(new_n795_), .A2(new_n1176_), .ZN(new_n1932_));
  NOR3_X1    g1883(.A1(new_n1930_), .A2(new_n1931_), .A3(new_n1932_), .ZN(new_n1933_));
  NOR2_X1    g1884(.A1(new_n1027_), .A2(new_n1153_), .ZN(new_n1934_));
  OAI21_X1   g1885(.A1(new_n1321_), .A2(new_n1126_), .B(new_n937_), .ZN(new_n1935_));
  XOR2_X1    g1886(.A1(new_n1934_), .A2(new_n1935_), .Z(new_n1936_));
  INV_X1     g1887(.I(new_n778_), .ZN(new_n1937_));
  NOR2_X1    g1888(.A1(new_n1937_), .A2(new_n752_), .ZN(new_n1938_));
  NOR2_X1    g1889(.A1(new_n1066_), .A2(new_n778_), .ZN(new_n1939_));
  OAI21_X1   g1890(.A1(new_n1938_), .A2(new_n1939_), .B(new_n67_), .ZN(new_n1940_));
  NOR2_X1    g1891(.A1(new_n1940_), .A2(new_n1120_), .ZN(new_n1941_));
  AOI21_X1   g1892(.A1(new_n1497_), .A2(new_n67_), .B(new_n494_), .ZN(new_n1942_));
  OAI21_X1   g1893(.A1(new_n1941_), .A2(new_n1942_), .B(new_n791_), .ZN(new_n1943_));
  NOR3_X1    g1894(.A1(new_n1943_), .A2(new_n780_), .A3(new_n1936_), .ZN(new_n1944_));
  NOR2_X1    g1895(.A1(new_n1059_), .A2(new_n1326_), .ZN(new_n1945_));
  NOR2_X1    g1896(.A1(new_n1944_), .A2(new_n1945_), .ZN(new_n1946_));
  INV_X1     g1897(.I(new_n1946_), .ZN(new_n1947_));
  NAND2_X1   g1898(.A1(new_n1944_), .A2(new_n1945_), .ZN(new_n1948_));
  AOI21_X1   g1899(.A1(new_n1947_), .A2(new_n1948_), .B(new_n1933_), .ZN(new_n1949_));
  AND3_X2    g1900(.A1(new_n1947_), .A2(new_n1933_), .A3(new_n1948_), .Z(new_n1950_));
  NOR2_X1    g1901(.A1(new_n1950_), .A2(new_n1949_), .ZN(new_n1951_));
  OR2_X2     g1902(.A1(new_n1908_), .A2(new_n1928_), .Z(new_n1952_));
  NAND2_X1   g1903(.A1(new_n1951_), .A2(new_n1952_), .ZN(new_n1953_));
  NAND2_X1   g1904(.A1(new_n1953_), .A2(new_n1929_), .ZN(new_n1954_));
  INV_X1     g1905(.I(new_n1954_), .ZN(new_n1955_));
  NAND2_X1   g1906(.A1(new_n1098_), .A2(new_n943_), .ZN(new_n1956_));
  NAND2_X1   g1907(.A1(new_n1230_), .A2(new_n62_), .ZN(new_n1957_));
  NAND2_X1   g1908(.A1(new_n1732_), .A2(new_n1176_), .ZN(new_n1958_));
  NAND2_X1   g1909(.A1(new_n1114_), .A2(new_n56_), .ZN(new_n1959_));
  AND4_X2    g1910(.A1(new_n1956_), .A2(new_n1958_), .A3(new_n1957_), .A4(new_n1959_), .Z(new_n1960_));
  NAND3_X1   g1911(.A1(new_n1031_), .A2(new_n1033_), .A3(new_n1171_), .ZN(new_n1961_));
  NAND2_X1   g1912(.A1(new_n1035_), .A2(new_n1062_), .ZN(new_n1962_));
  OAI21_X1   g1913(.A1(new_n1037_), .A2(new_n1062_), .B(new_n1962_), .ZN(new_n1963_));
  NOR2_X1    g1914(.A1(new_n1963_), .A2(new_n1961_), .ZN(new_n1964_));
  NOR2_X1    g1915(.A1(new_n1027_), .A2(new_n1126_), .ZN(new_n1965_));
  OAI21_X1   g1916(.A1(new_n1321_), .A2(new_n1134_), .B(new_n937_), .ZN(new_n1966_));
  XOR2_X1    g1917(.A1(new_n1965_), .A2(new_n1966_), .Z(new_n1967_));
  INV_X1     g1918(.I(new_n1967_), .ZN(new_n1968_));
  NAND2_X1   g1919(.A1(new_n1964_), .A2(new_n1968_), .ZN(new_n1969_));
  INV_X1     g1920(.I(new_n1969_), .ZN(new_n1970_));
  NOR2_X1    g1921(.A1(new_n1964_), .A2(new_n1968_), .ZN(new_n1971_));
  OAI21_X1   g1922(.A1(new_n1970_), .A2(new_n1971_), .B(new_n1960_), .ZN(new_n1972_));
  XOR2_X1    g1923(.A1(new_n1964_), .A2(new_n1967_), .Z(new_n1973_));
  OAI21_X1   g1924(.A1(new_n1960_), .A2(new_n1973_), .B(new_n1972_), .ZN(new_n1974_));
  NAND3_X1   g1925(.A1(new_n1497_), .A2(new_n67_), .A3(new_n494_), .ZN(new_n1975_));
  NAND2_X1   g1926(.A1(new_n1940_), .A2(new_n1120_), .ZN(new_n1976_));
  AOI21_X1   g1927(.A1(new_n1976_), .A2(new_n1975_), .B(new_n779_), .ZN(new_n1977_));
  XOR2_X1    g1928(.A1(new_n1977_), .A2(new_n780_), .Z(new_n1978_));
  AOI21_X1   g1929(.A1(new_n1097_), .A2(new_n752_), .B(new_n1176_), .ZN(new_n1979_));
  AOI21_X1   g1930(.A1(new_n1097_), .A2(new_n1066_), .B(new_n56_), .ZN(new_n1980_));
  XOR2_X1    g1931(.A1(new_n830_), .A2(new_n1326_), .Z(new_n1981_));
  NAND2_X1   g1932(.A1(new_n1066_), .A2(new_n1096_), .ZN(new_n1982_));
  NAND2_X1   g1933(.A1(new_n1108_), .A2(new_n752_), .ZN(new_n1983_));
  AOI21_X1   g1934(.A1(new_n1982_), .A2(new_n1983_), .B(new_n1981_), .ZN(new_n1984_));
  NOR4_X1    g1935(.A1(new_n1979_), .A2(new_n1980_), .A3(new_n1984_), .A4(new_n1097_), .ZN(new_n1985_));
  NOR3_X1    g1936(.A1(new_n1096_), .A2(new_n830_), .A3(new_n67_), .ZN(new_n1986_));
  AOI21_X1   g1937(.A1(new_n1096_), .A2(new_n67_), .B(new_n988_), .ZN(new_n1987_));
  OAI21_X1   g1938(.A1(new_n1987_), .A2(new_n1986_), .B(new_n752_), .ZN(new_n1988_));
  INV_X1     g1939(.I(new_n1988_), .ZN(new_n1989_));
  NOR2_X1    g1940(.A1(new_n1027_), .A2(new_n1134_), .ZN(new_n1990_));
  AOI21_X1   g1941(.A1(new_n1027_), .A2(new_n1053_), .B(new_n903_), .ZN(new_n1991_));
  XOR2_X1    g1942(.A1(new_n1991_), .A2(new_n1990_), .Z(new_n1992_));
  NAND2_X1   g1943(.A1(new_n1035_), .A2(new_n1171_), .ZN(new_n1993_));
  OAI21_X1   g1944(.A1(new_n1171_), .A2(new_n1037_), .B(new_n1993_), .ZN(new_n1994_));
  NOR4_X1    g1945(.A1(new_n1994_), .A2(new_n62_), .A3(new_n1032_), .A4(new_n1034_), .ZN(new_n1995_));
  NAND4_X1   g1946(.A1(new_n1985_), .A2(new_n1989_), .A3(new_n1995_), .A4(new_n1992_), .ZN(new_n1996_));
  INV_X1     g1947(.I(new_n1996_), .ZN(new_n1997_));
  INV_X1     g1948(.I(new_n1985_), .ZN(new_n1998_));
  XNOR2_X1   g1949(.A1(new_n1991_), .A2(new_n1990_), .ZN(new_n1999_));
  NOR2_X1    g1950(.A1(new_n1999_), .A2(new_n1989_), .ZN(new_n2000_));
  NOR2_X1    g1951(.A1(new_n1992_), .A2(new_n1988_), .ZN(new_n2001_));
  NOR2_X1    g1952(.A1(new_n2000_), .A2(new_n2001_), .ZN(new_n2002_));
  NAND2_X1   g1953(.A1(new_n1998_), .A2(new_n2002_), .ZN(new_n2003_));
  INV_X1     g1954(.I(new_n1995_), .ZN(new_n2004_));
  NAND2_X1   g1955(.A1(new_n1992_), .A2(new_n1988_), .ZN(new_n2005_));
  NAND2_X1   g1956(.A1(new_n1999_), .A2(new_n1989_), .ZN(new_n2006_));
  NAND2_X1   g1957(.A1(new_n2006_), .A2(new_n2005_), .ZN(new_n2007_));
  NAND2_X1   g1958(.A1(new_n2007_), .A2(new_n1985_), .ZN(new_n2008_));
  NAND2_X1   g1959(.A1(new_n2008_), .A2(new_n2004_), .ZN(new_n2009_));
  NOR2_X1    g1960(.A1(new_n1999_), .A2(new_n1988_), .ZN(new_n2010_));
  AOI21_X1   g1961(.A1(new_n2009_), .A2(new_n2003_), .B(new_n2010_), .ZN(new_n2011_));
  OAI21_X1   g1962(.A1(new_n2011_), .A2(new_n1997_), .B(new_n1978_), .ZN(new_n2012_));
  XOR2_X1    g1963(.A1(new_n1977_), .A2(new_n781_), .Z(new_n2013_));
  NOR2_X1    g1964(.A1(new_n2007_), .A2(new_n1985_), .ZN(new_n2014_));
  AOI21_X1   g1965(.A1(new_n2007_), .A2(new_n1985_), .B(new_n1995_), .ZN(new_n2015_));
  OAI22_X1   g1966(.A1(new_n2015_), .A2(new_n2014_), .B1(new_n1988_), .B2(new_n1999_), .ZN(new_n2016_));
  NAND3_X1   g1967(.A1(new_n2013_), .A2(new_n2016_), .A3(new_n1996_), .ZN(new_n2017_));
  AOI21_X1   g1968(.A1(new_n2012_), .A2(new_n2017_), .B(new_n1974_), .ZN(new_n2018_));
  NOR2_X1    g1969(.A1(new_n2002_), .A2(new_n1985_), .ZN(new_n2019_));
  INV_X1     g1970(.I(new_n2019_), .ZN(new_n2020_));
  NAND2_X1   g1971(.A1(new_n2002_), .A2(new_n1985_), .ZN(new_n2021_));
  AOI21_X1   g1972(.A1(new_n2020_), .A2(new_n2021_), .B(new_n2004_), .ZN(new_n2022_));
  AOI21_X1   g1973(.A1(new_n2003_), .A2(new_n2008_), .B(new_n1995_), .ZN(new_n2023_));
  NAND2_X1   g1974(.A1(new_n1189_), .A2(new_n62_), .ZN(new_n2024_));
  AOI21_X1   g1975(.A1(new_n1188_), .A2(new_n830_), .B(new_n62_), .ZN(new_n2025_));
  NAND2_X1   g1976(.A1(new_n830_), .A2(new_n937_), .ZN(new_n2026_));
  NAND2_X1   g1977(.A1(new_n988_), .A2(new_n903_), .ZN(new_n2027_));
  XOR2_X1    g1978(.A1(new_n978_), .A2(new_n56_), .Z(new_n2028_));
  AOI21_X1   g1979(.A1(new_n2027_), .A2(new_n2026_), .B(new_n2028_), .ZN(new_n2029_));
  NOR3_X1    g1980(.A1(new_n2029_), .A2(new_n2025_), .A3(new_n1188_), .ZN(new_n2030_));
  NAND2_X1   g1981(.A1(new_n1321_), .A2(new_n1053_), .ZN(new_n2031_));
  OAI21_X1   g1982(.A1(new_n1321_), .A2(new_n1171_), .B(new_n937_), .ZN(new_n2032_));
  XOR2_X1    g1983(.A1(new_n2032_), .A2(new_n2031_), .Z(new_n2033_));
  AOI21_X1   g1984(.A1(new_n2030_), .A2(new_n2024_), .B(new_n2033_), .ZN(new_n2034_));
  INV_X1     g1985(.I(new_n904_), .ZN(new_n2035_));
  NAND3_X1   g1986(.A1(new_n1188_), .A2(new_n67_), .A3(new_n988_), .ZN(new_n2036_));
  OAI21_X1   g1987(.A1(new_n980_), .A2(new_n979_), .B(new_n67_), .ZN(new_n2037_));
  NAND2_X1   g1988(.A1(new_n2037_), .A2(new_n830_), .ZN(new_n2038_));
  AOI21_X1   g1989(.A1(new_n2038_), .A2(new_n2036_), .B(new_n2035_), .ZN(new_n2039_));
  AOI21_X1   g1990(.A1(new_n1320_), .A2(new_n1013_), .B(new_n1171_), .ZN(new_n2040_));
  INV_X1     g1991(.I(new_n2040_), .ZN(new_n2041_));
  NAND3_X1   g1992(.A1(new_n1320_), .A2(new_n62_), .A3(new_n1013_), .ZN(new_n2042_));
  NAND2_X1   g1993(.A1(new_n2042_), .A2(new_n937_), .ZN(new_n2043_));
  XOR2_X1    g1994(.A1(new_n2043_), .A2(new_n2041_), .Z(new_n2044_));
  NAND3_X1   g1995(.A1(new_n2039_), .A2(new_n2044_), .A3(new_n905_), .ZN(new_n2045_));
  NAND2_X1   g1996(.A1(new_n1035_), .A2(new_n943_), .ZN(new_n2046_));
  NAND2_X1   g1997(.A1(new_n2027_), .A2(new_n2026_), .ZN(new_n2047_));
  XOR2_X1    g1998(.A1(new_n978_), .A2(new_n1176_), .Z(new_n2048_));
  AOI21_X1   g1999(.A1(new_n2047_), .A2(new_n2048_), .B(new_n1188_), .ZN(new_n2049_));
  NAND4_X1   g2000(.A1(new_n2033_), .A2(new_n2049_), .A3(new_n2024_), .A4(new_n2046_), .ZN(new_n2050_));
  AOI21_X1   g2001(.A1(new_n2045_), .A2(new_n2050_), .B(new_n2034_), .ZN(new_n2051_));
  INV_X1     g2002(.I(new_n2051_), .ZN(new_n2052_));
  OAI21_X1   g2003(.A1(new_n2022_), .A2(new_n2023_), .B(new_n2052_), .ZN(new_n2053_));
  INV_X1     g2004(.I(new_n2024_), .ZN(new_n2054_));
  INV_X1     g2005(.I(new_n2026_), .ZN(new_n2055_));
  NOR2_X1    g2006(.A1(new_n830_), .A2(new_n937_), .ZN(new_n2056_));
  OAI21_X1   g2007(.A1(new_n2055_), .A2(new_n2056_), .B(new_n2048_), .ZN(new_n2057_));
  NAND3_X1   g2008(.A1(new_n2057_), .A2(new_n2046_), .A3(new_n981_), .ZN(new_n2058_));
  XNOR2_X1   g2009(.A1(new_n2032_), .A2(new_n2031_), .ZN(new_n2059_));
  OAI21_X1   g2010(.A1(new_n2058_), .A2(new_n2054_), .B(new_n2059_), .ZN(new_n2060_));
  INV_X1     g2011(.I(new_n905_), .ZN(new_n2061_));
  NOR2_X1    g2012(.A1(new_n2037_), .A2(new_n830_), .ZN(new_n2062_));
  AOI21_X1   g2013(.A1(new_n1188_), .A2(new_n67_), .B(new_n988_), .ZN(new_n2063_));
  OAI21_X1   g2014(.A1(new_n2062_), .A2(new_n2063_), .B(new_n904_), .ZN(new_n2064_));
  AOI21_X1   g2015(.A1(new_n937_), .A2(new_n2042_), .B(new_n2041_), .ZN(new_n2065_));
  NOR2_X1    g2016(.A1(new_n2043_), .A2(new_n2040_), .ZN(new_n2066_));
  NOR2_X1    g2017(.A1(new_n2065_), .A2(new_n2066_), .ZN(new_n2067_));
  NOR3_X1    g2018(.A1(new_n2064_), .A2(new_n2061_), .A3(new_n2067_), .ZN(new_n2068_));
  AOI21_X1   g2019(.A1(new_n2060_), .A2(new_n2050_), .B(new_n2068_), .ZN(new_n2069_));
  NOR3_X1    g2020(.A1(new_n2058_), .A2(new_n2054_), .A3(new_n2059_), .ZN(new_n2070_));
  NOR3_X1    g2021(.A1(new_n2034_), .A2(new_n2070_), .A3(new_n2045_), .ZN(new_n2071_));
  NOR2_X1    g2022(.A1(new_n2071_), .A2(new_n2069_), .ZN(new_n2072_));
  OAI21_X1   g2023(.A1(new_n2064_), .A2(new_n2061_), .B(new_n2044_), .ZN(new_n2073_));
  NAND3_X1   g2024(.A1(new_n2039_), .A2(new_n905_), .A3(new_n2067_), .ZN(new_n2074_));
  NAND2_X1   g2025(.A1(new_n2073_), .A2(new_n2074_), .ZN(new_n2075_));
  AOI21_X1   g2026(.A1(new_n2039_), .A2(new_n905_), .B(new_n2067_), .ZN(new_n2076_));
  NOR3_X1    g2027(.A1(new_n2064_), .A2(new_n2044_), .A3(new_n2061_), .ZN(new_n2077_));
  NAND2_X1   g2028(.A1(new_n1189_), .A2(new_n56_), .ZN(new_n2078_));
  NAND2_X1   g2029(.A1(new_n1035_), .A2(new_n1176_), .ZN(new_n2079_));
  NAND2_X1   g2030(.A1(new_n868_), .A2(new_n67_), .ZN(new_n2080_));
  NAND2_X1   g2031(.A1(new_n978_), .A2(new_n1326_), .ZN(new_n2081_));
  NAND3_X1   g2032(.A1(new_n2047_), .A2(new_n2080_), .A3(new_n2081_), .ZN(new_n2082_));
  NAND4_X1   g2033(.A1(new_n2082_), .A2(new_n2078_), .A3(new_n981_), .A4(new_n2079_), .ZN(new_n2083_));
  OAI21_X1   g2034(.A1(new_n2077_), .A2(new_n2076_), .B(new_n2083_), .ZN(new_n2084_));
  NOR2_X1    g2035(.A1(new_n1037_), .A2(new_n1176_), .ZN(new_n2085_));
  INV_X1     g2036(.I(new_n2079_), .ZN(new_n2086_));
  NAND2_X1   g2037(.A1(new_n2080_), .A2(new_n2081_), .ZN(new_n2087_));
  AOI21_X1   g2038(.A1(new_n2026_), .A2(new_n2027_), .B(new_n2087_), .ZN(new_n2088_));
  NOR4_X1    g2039(.A1(new_n2085_), .A2(new_n2086_), .A3(new_n1188_), .A4(new_n2088_), .ZN(new_n2089_));
  NAND3_X1   g2040(.A1(new_n2073_), .A2(new_n2074_), .A3(new_n2089_), .ZN(new_n2090_));
  NOR2_X1    g2041(.A1(new_n1027_), .A2(new_n943_), .ZN(new_n2091_));
  INV_X1     g2042(.I(new_n2091_), .ZN(new_n2092_));
  AOI21_X1   g2043(.A1(new_n1027_), .A2(new_n56_), .B(new_n903_), .ZN(new_n2093_));
  NOR2_X1    g2044(.A1(new_n2092_), .A2(new_n2093_), .ZN(new_n2094_));
  NAND2_X1   g2045(.A1(new_n2092_), .A2(new_n2093_), .ZN(new_n2095_));
  INV_X1     g2046(.I(new_n2095_), .ZN(new_n2096_));
  NOR2_X1    g2047(.A1(new_n1027_), .A2(new_n1176_), .ZN(new_n2097_));
  NOR3_X1    g2048(.A1(new_n2097_), .A2(new_n67_), .A3(new_n903_), .ZN(new_n2098_));
  OAI21_X1   g2049(.A1(new_n2096_), .A2(new_n2094_), .B(new_n2098_), .ZN(new_n2099_));
  NOR3_X1    g2050(.A1(new_n2096_), .A2(new_n2094_), .A3(new_n2098_), .ZN(new_n2100_));
  NOR2_X1    g2051(.A1(new_n2062_), .A2(new_n2063_), .ZN(new_n2101_));
  MUX2_X1    g2052(.I0(new_n830_), .I1(new_n2101_), .S(new_n904_), .Z(new_n2102_));
  OAI21_X1   g2053(.A1(new_n2102_), .A2(new_n2100_), .B(new_n2099_), .ZN(new_n2103_));
  AOI22_X1   g2054(.A1(new_n2103_), .A2(new_n2075_), .B1(new_n2084_), .B2(new_n2090_), .ZN(new_n2104_));
  NOR2_X1    g2055(.A1(new_n2104_), .A2(new_n2072_), .ZN(new_n2105_));
  OAI21_X1   g2056(.A1(new_n2034_), .A2(new_n2070_), .B(new_n2045_), .ZN(new_n2106_));
  NAND3_X1   g2057(.A1(new_n2060_), .A2(new_n2068_), .A3(new_n2050_), .ZN(new_n2107_));
  NAND2_X1   g2058(.A1(new_n2106_), .A2(new_n2107_), .ZN(new_n2108_));
  NOR2_X1    g2059(.A1(new_n2077_), .A2(new_n2076_), .ZN(new_n2109_));
  AOI21_X1   g2060(.A1(new_n2073_), .A2(new_n2074_), .B(new_n2089_), .ZN(new_n2110_));
  NOR3_X1    g2061(.A1(new_n2077_), .A2(new_n2076_), .A3(new_n2083_), .ZN(new_n2111_));
  INV_X1     g2062(.I(new_n2094_), .ZN(new_n2112_));
  INV_X1     g2063(.I(new_n2098_), .ZN(new_n2113_));
  AOI21_X1   g2064(.A1(new_n2112_), .A2(new_n2095_), .B(new_n2113_), .ZN(new_n2114_));
  NAND3_X1   g2065(.A1(new_n2112_), .A2(new_n2095_), .A3(new_n2113_), .ZN(new_n2115_));
  NAND2_X1   g2066(.A1(new_n2038_), .A2(new_n2036_), .ZN(new_n2116_));
  MUX2_X1    g2067(.I0(new_n988_), .I1(new_n2116_), .S(new_n904_), .Z(new_n2117_));
  AOI21_X1   g2068(.A1(new_n2117_), .A2(new_n2115_), .B(new_n2114_), .ZN(new_n2118_));
  OAI22_X1   g2069(.A1(new_n2118_), .A2(new_n2109_), .B1(new_n2110_), .B2(new_n2111_), .ZN(new_n2119_));
  NOR2_X1    g2070(.A1(new_n2119_), .A2(new_n2108_), .ZN(new_n2120_));
  NAND2_X1   g2071(.A1(new_n1109_), .A2(new_n1107_), .ZN(new_n2121_));
  NOR2_X1    g2072(.A1(new_n2121_), .A2(new_n1326_), .ZN(new_n2122_));
  INV_X1     g2073(.I(new_n2122_), .ZN(new_n2123_));
  OAI22_X1   g2074(.A1(new_n2105_), .A2(new_n2120_), .B1(new_n2072_), .B2(new_n2123_), .ZN(new_n2124_));
  NOR3_X1    g2075(.A1(new_n2022_), .A2(new_n2023_), .A3(new_n2052_), .ZN(new_n2125_));
  OAI21_X1   g2076(.A1(new_n2124_), .A2(new_n2125_), .B(new_n2053_), .ZN(new_n2126_));
  NAND3_X1   g2077(.A1(new_n2012_), .A2(new_n1974_), .A3(new_n2017_), .ZN(new_n2127_));
  AOI21_X1   g2078(.A1(new_n2126_), .A2(new_n2127_), .B(new_n2018_), .ZN(new_n2128_));
  NOR2_X1    g2079(.A1(new_n2015_), .A2(new_n2014_), .ZN(new_n2129_));
  XOR2_X1    g2080(.A1(new_n1978_), .A2(new_n2129_), .Z(new_n2130_));
  OAI21_X1   g2081(.A1(new_n2013_), .A2(new_n2001_), .B(new_n2130_), .ZN(new_n2131_));
  NOR2_X1    g2082(.A1(new_n2128_), .A2(new_n2131_), .ZN(new_n2132_));
  NOR2_X1    g2083(.A1(new_n1231_), .A2(new_n939_), .ZN(new_n2133_));
  NOR2_X1    g2084(.A1(new_n1100_), .A2(new_n1171_), .ZN(new_n2134_));
  NOR4_X1    g2085(.A1(new_n2133_), .A2(new_n2134_), .A3(new_n1911_), .A4(new_n1912_), .ZN(new_n2135_));
  NOR2_X1    g2086(.A1(new_n2135_), .A2(new_n1919_), .ZN(new_n2136_));
  NOR2_X1    g2087(.A1(new_n1914_), .A2(new_n1918_), .ZN(new_n2137_));
  OAI21_X1   g2088(.A1(new_n2136_), .A2(new_n2137_), .B(new_n1926_), .ZN(new_n2138_));
  INV_X1     g2089(.I(new_n1920_), .ZN(new_n2139_));
  INV_X1     g2090(.I(new_n1926_), .ZN(new_n2140_));
  OAI21_X1   g2091(.A1(new_n2139_), .A2(new_n1927_), .B(new_n2140_), .ZN(new_n2141_));
  NAND2_X1   g2092(.A1(new_n2141_), .A2(new_n2138_), .ZN(new_n2142_));
  NOR2_X1    g2093(.A1(new_n1960_), .A2(new_n1970_), .ZN(new_n2143_));
  AOI21_X1   g2094(.A1(new_n1977_), .A2(new_n781_), .B(new_n1936_), .ZN(new_n2144_));
  INV_X1     g2095(.I(new_n1936_), .ZN(new_n2145_));
  NOR3_X1    g2096(.A1(new_n1943_), .A2(new_n780_), .A3(new_n2145_), .ZN(new_n2146_));
  NOR4_X1    g2097(.A1(new_n2143_), .A2(new_n2144_), .A3(new_n2146_), .A4(new_n1971_), .ZN(new_n2147_));
  INV_X1     g2098(.I(new_n1971_), .ZN(new_n2148_));
  NAND4_X1   g2099(.A1(new_n1958_), .A2(new_n1956_), .A3(new_n1957_), .A4(new_n1959_), .ZN(new_n2149_));
  NAND2_X1   g2100(.A1(new_n2149_), .A2(new_n1969_), .ZN(new_n2150_));
  OAI21_X1   g2101(.A1(new_n1943_), .A2(new_n780_), .B(new_n2145_), .ZN(new_n2151_));
  NAND3_X1   g2102(.A1(new_n1977_), .A2(new_n781_), .A3(new_n1936_), .ZN(new_n2152_));
  AOI22_X1   g2103(.A1(new_n2150_), .A2(new_n2148_), .B1(new_n2151_), .B2(new_n2152_), .ZN(new_n2153_));
  NOR2_X1    g2104(.A1(new_n2147_), .A2(new_n2153_), .ZN(new_n2154_));
  NOR2_X1    g2105(.A1(new_n2154_), .A2(new_n2142_), .ZN(new_n2155_));
  XOR2_X1    g2106(.A1(new_n1914_), .A2(new_n1919_), .Z(new_n2156_));
  NAND2_X1   g2107(.A1(new_n2135_), .A2(new_n1918_), .ZN(new_n2157_));
  AOI21_X1   g2108(.A1(new_n2157_), .A2(new_n1920_), .B(new_n1926_), .ZN(new_n2158_));
  AOI21_X1   g2109(.A1(new_n2156_), .A2(new_n1926_), .B(new_n2158_), .ZN(new_n2159_));
  NAND4_X1   g2110(.A1(new_n2150_), .A2(new_n2151_), .A3(new_n2152_), .A4(new_n2148_), .ZN(new_n2160_));
  OAI22_X1   g2111(.A1(new_n2143_), .A2(new_n1971_), .B1(new_n2144_), .B2(new_n2146_), .ZN(new_n2161_));
  NAND2_X1   g2112(.A1(new_n2161_), .A2(new_n2160_), .ZN(new_n2162_));
  NOR2_X1    g2113(.A1(new_n2162_), .A2(new_n2159_), .ZN(new_n2163_));
  NOR2_X1    g2114(.A1(new_n2155_), .A2(new_n2163_), .ZN(new_n2164_));
  AOI21_X1   g2115(.A1(new_n2128_), .A2(new_n2131_), .B(new_n2164_), .ZN(new_n2165_));
  NOR2_X1    g2116(.A1(new_n2143_), .A2(new_n1971_), .ZN(new_n2166_));
  NAND2_X1   g2117(.A1(new_n2151_), .A2(new_n2152_), .ZN(new_n2167_));
  NOR2_X1    g2118(.A1(new_n2166_), .A2(new_n2167_), .ZN(new_n2168_));
  NAND2_X1   g2119(.A1(new_n2166_), .A2(new_n2167_), .ZN(new_n2169_));
  AOI21_X1   g2120(.A1(new_n2142_), .A2(new_n2169_), .B(new_n2168_), .ZN(new_n2170_));
  INV_X1     g2121(.I(new_n2170_), .ZN(new_n2171_));
  OAI21_X1   g2122(.A1(new_n2165_), .A2(new_n2132_), .B(new_n2171_), .ZN(new_n2172_));
  AOI21_X1   g2123(.A1(new_n2148_), .A2(new_n1969_), .B(new_n2149_), .ZN(new_n2173_));
  NOR2_X1    g2124(.A1(new_n1973_), .A2(new_n1960_), .ZN(new_n2174_));
  NOR2_X1    g2125(.A1(new_n2174_), .A2(new_n2173_), .ZN(new_n2175_));
  AOI21_X1   g2126(.A1(new_n1996_), .A2(new_n2016_), .B(new_n2013_), .ZN(new_n2176_));
  NOR3_X1    g2127(.A1(new_n2011_), .A2(new_n1997_), .A3(new_n1978_), .ZN(new_n2177_));
  OAI21_X1   g2128(.A1(new_n2177_), .A2(new_n2176_), .B(new_n2175_), .ZN(new_n2178_));
  INV_X1     g2129(.I(new_n2021_), .ZN(new_n2179_));
  OAI21_X1   g2130(.A1(new_n2179_), .A2(new_n2019_), .B(new_n1995_), .ZN(new_n2180_));
  INV_X1     g2131(.I(new_n2008_), .ZN(new_n2181_));
  OAI21_X1   g2132(.A1(new_n2181_), .A2(new_n2014_), .B(new_n2004_), .ZN(new_n2182_));
  AOI21_X1   g2133(.A1(new_n2180_), .A2(new_n2182_), .B(new_n2051_), .ZN(new_n2183_));
  NAND2_X1   g2134(.A1(new_n2119_), .A2(new_n2108_), .ZN(new_n2184_));
  NAND2_X1   g2135(.A1(new_n2104_), .A2(new_n2072_), .ZN(new_n2185_));
  AOI22_X1   g2136(.A1(new_n2185_), .A2(new_n2184_), .B1(new_n2108_), .B2(new_n2122_), .ZN(new_n2186_));
  NAND3_X1   g2137(.A1(new_n2180_), .A2(new_n2182_), .A3(new_n2051_), .ZN(new_n2187_));
  AOI21_X1   g2138(.A1(new_n2186_), .A2(new_n2187_), .B(new_n2183_), .ZN(new_n2188_));
  NOR3_X1    g2139(.A1(new_n2177_), .A2(new_n2176_), .A3(new_n2175_), .ZN(new_n2189_));
  OAI21_X1   g2140(.A1(new_n2188_), .A2(new_n2189_), .B(new_n2178_), .ZN(new_n2190_));
  XOR2_X1    g2141(.A1(new_n2013_), .A2(new_n2129_), .Z(new_n2191_));
  AOI21_X1   g2142(.A1(new_n1978_), .A2(new_n2006_), .B(new_n2191_), .ZN(new_n2192_));
  NAND2_X1   g2143(.A1(new_n2190_), .A2(new_n2192_), .ZN(new_n2193_));
  NAND2_X1   g2144(.A1(new_n2162_), .A2(new_n2159_), .ZN(new_n2194_));
  NAND2_X1   g2145(.A1(new_n2154_), .A2(new_n2142_), .ZN(new_n2195_));
  NAND2_X1   g2146(.A1(new_n2195_), .A2(new_n2194_), .ZN(new_n2196_));
  OAI21_X1   g2147(.A1(new_n2190_), .A2(new_n2192_), .B(new_n2196_), .ZN(new_n2197_));
  NAND3_X1   g2148(.A1(new_n2197_), .A2(new_n2193_), .A3(new_n2170_), .ZN(new_n2198_));
  NAND2_X1   g2149(.A1(new_n1952_), .A2(new_n1929_), .ZN(new_n2199_));
  XNOR2_X1   g2150(.A1(new_n2199_), .A2(new_n1951_), .ZN(new_n2200_));
  NAND2_X1   g2151(.A1(new_n2198_), .A2(new_n2200_), .ZN(new_n2201_));
  AOI21_X1   g2152(.A1(new_n2201_), .A2(new_n2172_), .B(new_n1955_), .ZN(new_n2202_));
  INV_X1     g2153(.I(new_n2172_), .ZN(new_n2203_));
  NOR2_X1    g2154(.A1(new_n2165_), .A2(new_n2132_), .ZN(new_n2204_));
  XOR2_X1    g2155(.A1(new_n2199_), .A2(new_n1951_), .Z(new_n2205_));
  AOI21_X1   g2156(.A1(new_n2204_), .A2(new_n2170_), .B(new_n2205_), .ZN(new_n2206_));
  INV_X1     g2157(.I(new_n1945_), .ZN(new_n2207_));
  XNOR2_X1   g2158(.A1(new_n1944_), .A2(new_n1933_), .ZN(new_n2208_));
  AOI21_X1   g2159(.A1(new_n1944_), .A2(new_n2207_), .B(new_n2208_), .ZN(new_n2209_));
  AOI21_X1   g2160(.A1(new_n1817_), .A2(new_n1809_), .B(new_n1815_), .ZN(new_n2210_));
  XOR2_X1    g2161(.A1(new_n1803_), .A2(new_n1816_), .Z(new_n2211_));
  NOR2_X1    g2162(.A1(new_n2211_), .A2(new_n1814_), .ZN(new_n2212_));
  NOR3_X1    g2163(.A1(new_n2209_), .A2(new_n2210_), .A3(new_n2212_), .ZN(new_n2213_));
  NOR4_X1    g2164(.A1(new_n1944_), .A2(new_n1930_), .A3(new_n1931_), .A4(new_n1932_), .ZN(new_n2214_));
  NOR2_X1    g2165(.A1(new_n2208_), .A2(new_n2207_), .ZN(new_n2215_));
  NOR2_X1    g2166(.A1(new_n2215_), .A2(new_n2214_), .ZN(new_n2216_));
  NOR2_X1    g2167(.A1(new_n2212_), .A2(new_n2210_), .ZN(new_n2217_));
  NOR2_X1    g2168(.A1(new_n2216_), .A2(new_n2217_), .ZN(new_n2218_));
  NAND3_X1   g2169(.A1(new_n1460_), .A2(new_n1047_), .A3(new_n1176_), .ZN(new_n2219_));
  NOR2_X1    g2170(.A1(new_n1220_), .A2(new_n67_), .ZN(new_n2220_));
  OAI21_X1   g2171(.A1(new_n1046_), .A2(new_n1060_), .B(new_n67_), .ZN(new_n2221_));
  INV_X1     g2172(.I(new_n2221_), .ZN(new_n2222_));
  NOR3_X1    g2173(.A1(new_n2219_), .A2(new_n2220_), .A3(new_n2222_), .ZN(new_n2223_));
  AOI21_X1   g2174(.A1(new_n1892_), .A2(new_n1901_), .B(new_n1902_), .ZN(new_n2224_));
  INV_X1     g2175(.I(new_n2224_), .ZN(new_n2225_));
  NAND2_X1   g2176(.A1(new_n1724_), .A2(new_n416_), .ZN(new_n2226_));
  XNOR2_X1   g2177(.A1(new_n2226_), .A2(new_n1727_), .ZN(new_n2227_));
  INV_X1     g2178(.I(new_n2227_), .ZN(new_n2228_));
  NOR2_X1    g2179(.A1(new_n2228_), .A2(new_n2225_), .ZN(new_n2229_));
  NOR2_X1    g2180(.A1(new_n2227_), .A2(new_n2224_), .ZN(new_n2230_));
  OAI21_X1   g2181(.A1(new_n2229_), .A2(new_n2230_), .B(new_n2223_), .ZN(new_n2231_));
  INV_X1     g2182(.I(new_n2223_), .ZN(new_n2232_));
  XOR2_X1    g2183(.A1(new_n2227_), .A2(new_n2224_), .Z(new_n2233_));
  NAND2_X1   g2184(.A1(new_n2233_), .A2(new_n2232_), .ZN(new_n2234_));
  NAND2_X1   g2185(.A1(new_n2234_), .A2(new_n2231_), .ZN(new_n2235_));
  INV_X1     g2186(.I(new_n2235_), .ZN(new_n2236_));
  NOR3_X1    g2187(.A1(new_n2236_), .A2(new_n2218_), .A3(new_n2213_), .ZN(new_n2237_));
  NAND2_X1   g2188(.A1(new_n2216_), .A2(new_n2217_), .ZN(new_n2238_));
  OAI21_X1   g2189(.A1(new_n2210_), .A2(new_n2212_), .B(new_n2209_), .ZN(new_n2239_));
  AOI21_X1   g2190(.A1(new_n2238_), .A2(new_n2239_), .B(new_n2235_), .ZN(new_n2240_));
  OAI21_X1   g2191(.A1(new_n2237_), .A2(new_n2240_), .B(new_n1955_), .ZN(new_n2241_));
  NOR3_X1    g2192(.A1(new_n2206_), .A2(new_n2241_), .A3(new_n2203_), .ZN(new_n2242_));
  NAND2_X1   g2193(.A1(new_n2217_), .A2(new_n2209_), .ZN(new_n2243_));
  OAI21_X1   g2194(.A1(new_n2209_), .A2(new_n2217_), .B(new_n2236_), .ZN(new_n2244_));
  NAND2_X1   g2195(.A1(new_n2244_), .A2(new_n2243_), .ZN(new_n2245_));
  OAI21_X1   g2196(.A1(new_n2242_), .A2(new_n2202_), .B(new_n2245_), .ZN(new_n2246_));
  OAI21_X1   g2197(.A1(new_n2206_), .A2(new_n2203_), .B(new_n1954_), .ZN(new_n2247_));
  NAND3_X1   g2198(.A1(new_n2238_), .A2(new_n2239_), .A3(new_n2235_), .ZN(new_n2248_));
  OAI21_X1   g2199(.A1(new_n2218_), .A2(new_n2213_), .B(new_n2236_), .ZN(new_n2249_));
  AOI21_X1   g2200(.A1(new_n2249_), .A2(new_n2248_), .B(new_n1954_), .ZN(new_n2250_));
  NAND3_X1   g2201(.A1(new_n2201_), .A2(new_n2172_), .A3(new_n2250_), .ZN(new_n2251_));
  NAND2_X1   g2202(.A1(new_n2228_), .A2(new_n2225_), .ZN(new_n2252_));
  OAI21_X1   g2203(.A1(new_n2223_), .A2(new_n2229_), .B(new_n2252_), .ZN(new_n2253_));
  XOR2_X1    g2204(.A1(new_n1748_), .A2(new_n1752_), .Z(new_n2254_));
  NAND2_X1   g2205(.A1(new_n2254_), .A2(new_n1758_), .ZN(new_n2255_));
  OR2_X2     g2206(.A1(new_n1753_), .A2(new_n1759_), .Z(new_n2256_));
  INV_X1     g2207(.I(new_n2256_), .ZN(new_n2257_));
  OAI21_X1   g2208(.A1(new_n2257_), .A2(new_n1758_), .B(new_n2255_), .ZN(new_n2258_));
  XOR2_X1    g2209(.A1(new_n2253_), .A2(new_n2258_), .Z(new_n2259_));
  INV_X1     g2210(.I(new_n1798_), .ZN(new_n2260_));
  INV_X1     g2211(.I(new_n1819_), .ZN(new_n2261_));
  AOI21_X1   g2212(.A1(new_n2260_), .A2(new_n1820_), .B(new_n2261_), .ZN(new_n2262_));
  INV_X1     g2213(.I(new_n1797_), .ZN(new_n2263_));
  NOR3_X1    g2214(.A1(new_n1792_), .A2(new_n1796_), .A3(new_n2263_), .ZN(new_n2264_));
  INV_X1     g2215(.I(new_n2264_), .ZN(new_n2265_));
  OAI21_X1   g2216(.A1(new_n1792_), .A2(new_n1796_), .B(new_n2263_), .ZN(new_n2266_));
  AOI21_X1   g2217(.A1(new_n2265_), .A2(new_n2266_), .B(new_n1819_), .ZN(new_n2267_));
  OAI21_X1   g2218(.A1(new_n2262_), .A2(new_n2267_), .B(new_n2259_), .ZN(new_n2268_));
  INV_X1     g2219(.I(new_n2259_), .ZN(new_n2269_));
  NOR2_X1    g2220(.A1(new_n2262_), .A2(new_n2267_), .ZN(new_n2270_));
  NAND2_X1   g2221(.A1(new_n2270_), .A2(new_n2269_), .ZN(new_n2271_));
  AOI21_X1   g2222(.A1(new_n2271_), .A2(new_n2268_), .B(new_n2245_), .ZN(new_n2272_));
  NAND3_X1   g2223(.A1(new_n2247_), .A2(new_n2251_), .A3(new_n2272_), .ZN(new_n2273_));
  NAND2_X1   g2224(.A1(new_n1783_), .A2(new_n1880_), .ZN(new_n2274_));
  NAND2_X1   g2225(.A1(new_n1879_), .A2(new_n1788_), .ZN(new_n2275_));
  AOI21_X1   g2226(.A1(new_n2275_), .A2(new_n2274_), .B(new_n1821_), .ZN(new_n2276_));
  NAND2_X1   g2227(.A1(new_n1783_), .A2(new_n1788_), .ZN(new_n2277_));
  NAND2_X1   g2228(.A1(new_n1881_), .A2(new_n2277_), .ZN(new_n2278_));
  AOI21_X1   g2229(.A1(new_n2278_), .A2(new_n1821_), .B(new_n2276_), .ZN(new_n2279_));
  INV_X1     g2230(.I(new_n2279_), .ZN(new_n2280_));
  NAND3_X1   g2231(.A1(new_n2246_), .A2(new_n2273_), .A3(new_n2280_), .ZN(new_n2281_));
  INV_X1     g2232(.I(new_n2258_), .ZN(new_n2282_));
  NOR2_X1    g2233(.A1(new_n2270_), .A2(new_n2282_), .ZN(new_n2283_));
  NAND2_X1   g2234(.A1(new_n2270_), .A2(new_n2282_), .ZN(new_n2284_));
  AOI21_X1   g2235(.A1(new_n2253_), .A2(new_n2284_), .B(new_n2283_), .ZN(new_n2285_));
  INV_X1     g2236(.I(new_n2285_), .ZN(new_n2286_));
  NAND3_X1   g2237(.A1(new_n2281_), .A2(new_n1887_), .A3(new_n2286_), .ZN(new_n2287_));
  AOI21_X1   g2238(.A1(new_n2281_), .A2(new_n2286_), .B(new_n1887_), .ZN(new_n2288_));
  INV_X1     g2239(.I(new_n2288_), .ZN(new_n2289_));
  INV_X1     g2240(.I(new_n1074_), .ZN(new_n2290_));
  NAND2_X1   g2241(.A1(new_n1644_), .A2(new_n915_), .ZN(new_n2291_));
  NOR3_X1    g2242(.A1(new_n2290_), .A2(new_n2291_), .A3(new_n404_), .ZN(new_n2292_));
  NAND2_X1   g2243(.A1(new_n931_), .A2(new_n949_), .ZN(new_n2293_));
  NOR4_X1    g2244(.A1(new_n2293_), .A2(new_n266_), .A3(new_n335_), .A4(new_n393_), .ZN(new_n2294_));
  NOR2_X1    g2245(.A1(new_n454_), .A2(new_n495_), .ZN(new_n2295_));
  NAND4_X1   g2246(.A1(new_n2292_), .A2(new_n728_), .A3(new_n2294_), .A4(new_n2295_), .ZN(new_n2296_));
  NOR4_X1    g2247(.A1(new_n738_), .A2(new_n189_), .A3(new_n384_), .A4(new_n515_), .ZN(new_n2297_));
  NOR4_X1    g2248(.A1(new_n326_), .A2(new_n437_), .A3(new_n747_), .A4(new_n534_), .ZN(new_n2298_));
  NOR4_X1    g2249(.A1(new_n1706_), .A2(new_n483_), .A3(new_n242_), .A4(new_n856_), .ZN(new_n2299_));
  INV_X1     g2250(.I(new_n2299_), .ZN(new_n2300_));
  NAND4_X1   g2251(.A1(new_n2300_), .A2(new_n586_), .A3(new_n2297_), .A4(new_n2298_), .ZN(new_n2301_));
  INV_X1     g2252(.I(new_n718_), .ZN(new_n2302_));
  NAND3_X1   g2253(.A1(new_n2302_), .A2(new_n914_), .A3(new_n742_), .ZN(new_n2303_));
  NOR3_X1    g2254(.A1(new_n642_), .A2(new_n372_), .A3(new_n825_), .ZN(new_n2304_));
  NOR2_X1    g2255(.A1(new_n535_), .A2(new_n593_), .ZN(new_n2305_));
  NAND4_X1   g2256(.A1(new_n800_), .A2(new_n213_), .A3(new_n2304_), .A4(new_n2305_), .ZN(new_n2306_));
  NOR4_X1    g2257(.A1(new_n2296_), .A2(new_n2301_), .A3(new_n2306_), .A4(new_n2303_), .ZN(new_n2307_));
  NAND3_X1   g2258(.A1(new_n2289_), .A2(new_n2287_), .A3(new_n2307_), .ZN(new_n2308_));
  NAND2_X1   g2259(.A1(new_n223_), .A2(new_n458_), .ZN(new_n2309_));
  NOR4_X1    g2260(.A1(new_n2309_), .A2(new_n198_), .A3(new_n327_), .A4(new_n422_), .ZN(new_n2310_));
  INV_X1     g2261(.I(new_n2310_), .ZN(new_n2311_));
  NOR2_X1    g2262(.A1(new_n518_), .A2(new_n278_), .ZN(new_n2312_));
  NOR2_X1    g2263(.A1(new_n594_), .A2(new_n437_), .ZN(new_n2313_));
  NOR2_X1    g2264(.A1(new_n279_), .A2(new_n265_), .ZN(new_n2314_));
  NOR2_X1    g2265(.A1(new_n293_), .A2(new_n2314_), .ZN(new_n2315_));
  INV_X1     g2266(.I(new_n2315_), .ZN(new_n2316_));
  AOI21_X1   g2267(.A1(new_n2312_), .A2(new_n2313_), .B(new_n2316_), .ZN(new_n2317_));
  INV_X1     g2268(.I(new_n2317_), .ZN(new_n2318_));
  NAND2_X1   g2269(.A1(new_n645_), .A2(new_n252_), .ZN(new_n2319_));
  NAND3_X1   g2270(.A1(new_n288_), .A2(new_n539_), .A3(new_n926_), .ZN(new_n2320_));
  NOR4_X1    g2271(.A1(new_n2318_), .A2(new_n2311_), .A3(new_n2319_), .A4(new_n2320_), .ZN(new_n2321_));
  NOR2_X1    g2272(.A1(new_n338_), .A2(new_n473_), .ZN(new_n2322_));
  INV_X1     g2273(.I(new_n2322_), .ZN(new_n2323_));
  NOR3_X1    g2274(.A1(new_n2323_), .A2(new_n1079_), .A3(new_n543_), .ZN(new_n2324_));
  INV_X1     g2275(.I(new_n772_), .ZN(new_n2325_));
  NOR4_X1    g2276(.A1(new_n301_), .A2(new_n378_), .A3(new_n384_), .A4(new_n1091_), .ZN(new_n2326_));
  NOR4_X1    g2277(.A1(new_n825_), .A2(new_n267_), .A3(new_n588_), .A4(new_n266_), .ZN(new_n2327_));
  NOR3_X1    g2278(.A1(new_n2325_), .A2(new_n2326_), .A3(new_n2327_), .ZN(new_n2328_));
  NAND4_X1   g2279(.A1(new_n2321_), .A2(new_n1708_), .A3(new_n2324_), .A4(new_n2328_), .ZN(new_n2329_));
  NOR2_X1    g2280(.A1(new_n2308_), .A2(new_n2329_), .ZN(new_n2330_));
  OAI21_X1   g2281(.A1(new_n1357_), .A2(new_n1539_), .B(new_n1538_), .ZN(new_n2331_));
  XOR2_X1    g2282(.A1(new_n1355_), .A2(new_n1349_), .Z(new_n2332_));
  INV_X1     g2283(.I(new_n2332_), .ZN(new_n2333_));
  NAND2_X1   g2284(.A1(new_n1404_), .A2(new_n2333_), .ZN(new_n2334_));
  NAND2_X1   g2285(.A1(new_n2331_), .A2(new_n2334_), .ZN(new_n2335_));
  INV_X1     g2286(.I(new_n2335_), .ZN(new_n2336_));
  NAND3_X1   g2287(.A1(new_n2246_), .A2(new_n2273_), .A3(new_n2286_), .ZN(new_n2337_));
  INV_X1     g2288(.I(new_n2245_), .ZN(new_n2338_));
  AOI21_X1   g2289(.A1(new_n2247_), .A2(new_n2251_), .B(new_n2338_), .ZN(new_n2339_));
  INV_X1     g2290(.I(new_n2272_), .ZN(new_n2340_));
  NOR3_X1    g2291(.A1(new_n2340_), .A2(new_n2242_), .A3(new_n2202_), .ZN(new_n2341_));
  OAI21_X1   g2292(.A1(new_n2341_), .A2(new_n2339_), .B(new_n2285_), .ZN(new_n2342_));
  NAND2_X1   g2293(.A1(new_n2342_), .A2(new_n2337_), .ZN(new_n2343_));
  NAND2_X1   g2294(.A1(new_n2246_), .A2(new_n2273_), .ZN(new_n2344_));
  NOR3_X1    g2295(.A1(new_n1886_), .A2(new_n1872_), .A3(new_n2285_), .ZN(new_n2345_));
  AOI21_X1   g2296(.A1(new_n2344_), .A2(new_n2345_), .B(new_n2280_), .ZN(new_n2346_));
  NAND2_X1   g2297(.A1(new_n2343_), .A2(new_n2346_), .ZN(new_n2347_));
  NOR2_X1    g2298(.A1(new_n1822_), .A2(new_n1789_), .ZN(new_n2348_));
  OAI21_X1   g2299(.A1(new_n1862_), .A2(new_n1871_), .B(new_n2348_), .ZN(new_n2349_));
  NOR3_X1    g2300(.A1(new_n1868_), .A2(new_n1840_), .A3(new_n1845_), .ZN(new_n2350_));
  AOI21_X1   g2301(.A1(new_n1742_), .A2(new_n1778_), .B(new_n1873_), .ZN(new_n2351_));
  AOI21_X1   g2302(.A1(new_n1848_), .A2(new_n1849_), .B(new_n1832_), .ZN(new_n2352_));
  NOR2_X1    g2303(.A1(new_n2352_), .A2(new_n2351_), .ZN(new_n2353_));
  NOR2_X1    g2304(.A1(new_n2353_), .A2(new_n2350_), .ZN(new_n2354_));
  INV_X1     g2305(.I(new_n2354_), .ZN(new_n2355_));
  AOI21_X1   g2306(.A1(new_n2347_), .A2(new_n2349_), .B(new_n2355_), .ZN(new_n2356_));
  NOR3_X1    g2307(.A1(new_n2341_), .A2(new_n2339_), .A3(new_n2285_), .ZN(new_n2357_));
  AOI21_X1   g2308(.A1(new_n2246_), .A2(new_n2273_), .B(new_n2286_), .ZN(new_n2358_));
  NOR2_X1    g2309(.A1(new_n2357_), .A2(new_n2358_), .ZN(new_n2359_));
  OAI21_X1   g2310(.A1(new_n2341_), .A2(new_n2339_), .B(new_n2345_), .ZN(new_n2360_));
  NAND2_X1   g2311(.A1(new_n2360_), .A2(new_n2279_), .ZN(new_n2361_));
  OAI21_X1   g2312(.A1(new_n2359_), .A2(new_n2361_), .B(new_n2349_), .ZN(new_n2362_));
  NOR2_X1    g2313(.A1(new_n2362_), .A2(new_n2354_), .ZN(new_n2363_));
  OAI21_X1   g2314(.A1(new_n2363_), .A2(new_n2356_), .B(new_n2336_), .ZN(new_n2364_));
  NAND2_X1   g2315(.A1(new_n2362_), .A2(new_n2354_), .ZN(new_n2365_));
  NAND3_X1   g2316(.A1(new_n2347_), .A2(new_n2349_), .A3(new_n2355_), .ZN(new_n2366_));
  NAND3_X1   g2317(.A1(new_n2365_), .A2(new_n2366_), .A3(new_n2335_), .ZN(new_n2367_));
  INV_X1     g2318(.I(new_n2287_), .ZN(new_n2368_));
  INV_X1     g2319(.I(new_n2307_), .ZN(new_n2369_));
  NOR3_X1    g2320(.A1(new_n2368_), .A2(new_n2288_), .A3(new_n2369_), .ZN(new_n2370_));
  INV_X1     g2321(.I(new_n2329_), .ZN(new_n2371_));
  NOR2_X1    g2322(.A1(new_n2370_), .A2(new_n2371_), .ZN(new_n2372_));
  AOI21_X1   g2323(.A1(new_n2364_), .A2(new_n2367_), .B(new_n2372_), .ZN(new_n2373_));
  INV_X1     g2324(.I(new_n432_), .ZN(new_n2374_));
  NOR4_X1    g2325(.A1(new_n642_), .A2(new_n242_), .A3(new_n434_), .A4(new_n399_), .ZN(new_n2375_));
  INV_X1     g2326(.I(new_n449_), .ZN(new_n2376_));
  NOR3_X1    g2327(.A1(new_n2376_), .A2(new_n369_), .A3(new_n478_), .ZN(new_n2377_));
  INV_X1     g2328(.I(new_n2377_), .ZN(new_n2378_));
  NOR3_X1    g2329(.A1(new_n2378_), .A2(new_n817_), .A3(new_n2375_), .ZN(new_n2379_));
  NOR2_X1    g2330(.A1(new_n438_), .A2(new_n535_), .ZN(new_n2380_));
  INV_X1     g2331(.I(new_n2380_), .ZN(new_n2381_));
  NOR4_X1    g2332(.A1(new_n2381_), .A2(new_n865_), .A3(new_n974_), .A4(new_n389_), .ZN(new_n2382_));
  NOR3_X1    g2333(.A1(new_n214_), .A2(new_n2323_), .A3(new_n1085_), .ZN(new_n2383_));
  NAND4_X1   g2334(.A1(new_n2379_), .A2(new_n1704_), .A3(new_n2382_), .A4(new_n2383_), .ZN(new_n2384_));
  INV_X1     g2335(.I(new_n2384_), .ZN(new_n2385_));
  INV_X1     g2336(.I(new_n1067_), .ZN(new_n2386_));
  NOR3_X1    g2337(.A1(new_n801_), .A2(new_n305_), .A3(new_n526_), .ZN(new_n2387_));
  NOR2_X1    g2338(.A1(new_n483_), .A2(new_n263_), .ZN(new_n2388_));
  NAND4_X1   g2339(.A1(new_n2386_), .A2(new_n767_), .A3(new_n2387_), .A4(new_n2388_), .ZN(new_n2389_));
  INV_X1     g2340(.I(new_n614_), .ZN(new_n2390_));
  NOR4_X1    g2341(.A1(new_n204_), .A2(new_n339_), .A3(new_n378_), .A4(new_n488_), .ZN(new_n2391_));
  NOR2_X1    g2342(.A1(new_n306_), .A2(new_n553_), .ZN(new_n2392_));
  INV_X1     g2343(.I(new_n2392_), .ZN(new_n2393_));
  NOR4_X1    g2344(.A1(new_n2393_), .A2(new_n2391_), .A3(new_n307_), .A4(new_n391_), .ZN(new_n2394_));
  NOR2_X1    g2345(.A1(new_n514_), .A2(new_n507_), .ZN(new_n2395_));
  NAND4_X1   g2346(.A1(new_n2394_), .A2(new_n921_), .A3(new_n2390_), .A4(new_n2395_), .ZN(new_n2396_));
  NOR3_X1    g2347(.A1(new_n2396_), .A2(new_n333_), .A3(new_n2389_), .ZN(new_n2397_));
  NAND3_X1   g2348(.A1(new_n2385_), .A2(new_n2397_), .A3(new_n2374_), .ZN(new_n2398_));
  INV_X1     g2349(.I(new_n2398_), .ZN(new_n2399_));
  OAI21_X1   g2350(.A1(new_n2373_), .A2(new_n2330_), .B(new_n2399_), .ZN(new_n2400_));
  AOI21_X1   g2351(.A1(new_n1542_), .A2(new_n1541_), .B(new_n1540_), .ZN(new_n2401_));
  NOR2_X1    g2352(.A1(new_n1428_), .A2(new_n2401_), .ZN(new_n2402_));
  NOR3_X1    g2353(.A1(new_n2373_), .A2(new_n2330_), .A3(new_n2399_), .ZN(new_n2403_));
  OAI21_X1   g2354(.A1(new_n2402_), .A2(new_n2403_), .B(new_n2400_), .ZN(new_n2404_));
  NOR2_X1    g2355(.A1(new_n1546_), .A2(new_n1437_), .ZN(new_n2405_));
  NOR2_X1    g2356(.A1(new_n1433_), .A2(new_n1251_), .ZN(new_n2406_));
  OAI21_X1   g2357(.A1(new_n2406_), .A2(new_n2405_), .B(new_n1435_), .ZN(new_n2407_));
  NOR2_X1    g2358(.A1(new_n1546_), .A2(new_n1251_), .ZN(new_n2408_));
  NOR2_X1    g2359(.A1(new_n1433_), .A2(new_n1437_), .ZN(new_n2409_));
  OAI21_X1   g2360(.A1(new_n2409_), .A2(new_n2408_), .B(new_n1434_), .ZN(new_n2410_));
  NAND3_X1   g2361(.A1(new_n2407_), .A2(new_n2410_), .A3(new_n1428_), .ZN(new_n2411_));
  NAND2_X1   g2362(.A1(new_n1433_), .A2(new_n1251_), .ZN(new_n2412_));
  NAND2_X1   g2363(.A1(new_n1546_), .A2(new_n1437_), .ZN(new_n2413_));
  AOI21_X1   g2364(.A1(new_n2412_), .A2(new_n2413_), .B(new_n1434_), .ZN(new_n2414_));
  NAND2_X1   g2365(.A1(new_n1433_), .A2(new_n1437_), .ZN(new_n2415_));
  NAND2_X1   g2366(.A1(new_n1546_), .A2(new_n1251_), .ZN(new_n2416_));
  AOI21_X1   g2367(.A1(new_n2415_), .A2(new_n2416_), .B(new_n1435_), .ZN(new_n2417_));
  OAI21_X1   g2368(.A1(new_n2414_), .A2(new_n2417_), .B(new_n1543_), .ZN(new_n2418_));
  NAND2_X1   g2369(.A1(new_n2418_), .A2(new_n2411_), .ZN(new_n2419_));
  XNOR2_X1   g2370(.A1(new_n1306_), .A2(new_n1253_), .ZN(new_n2420_));
  INV_X1     g2371(.I(new_n2420_), .ZN(new_n2421_));
  NOR3_X1    g2372(.A1(new_n518_), .A2(new_n306_), .A3(new_n473_), .ZN(new_n2422_));
  NOR4_X1    g2373(.A1(new_n280_), .A2(new_n307_), .A3(new_n878_), .A4(new_n872_), .ZN(new_n2423_));
  NOR2_X1    g2374(.A1(new_n2376_), .A2(new_n832_), .ZN(new_n2424_));
  INV_X1     g2375(.I(new_n2424_), .ZN(new_n2425_));
  NOR4_X1    g2376(.A1(new_n2425_), .A2(new_n500_), .A3(new_n2423_), .A4(new_n402_), .ZN(new_n2426_));
  NAND3_X1   g2377(.A1(new_n2426_), .A2(new_n803_), .A3(new_n2422_), .ZN(new_n2427_));
  INV_X1     g2378(.I(new_n2427_), .ZN(new_n2428_));
  INV_X1     g2379(.I(new_n728_), .ZN(new_n2429_));
  NOR4_X1    g2380(.A1(new_n326_), .A2(new_n438_), .A3(new_n327_), .A4(new_n593_), .ZN(new_n2430_));
  NOR4_X1    g2381(.A1(new_n2430_), .A2(new_n378_), .A3(new_n394_), .A4(new_n517_), .ZN(new_n2431_));
  INV_X1     g2382(.I(new_n2431_), .ZN(new_n2432_));
  NOR4_X1    g2383(.A1(new_n322_), .A2(new_n515_), .A3(new_n278_), .A4(new_n399_), .ZN(new_n2433_));
  NOR4_X1    g2384(.A1(new_n369_), .A2(new_n608_), .A3(new_n372_), .A4(new_n487_), .ZN(new_n2434_));
  NOR4_X1    g2385(.A1(new_n2432_), .A2(new_n2429_), .A3(new_n2433_), .A4(new_n2434_), .ZN(new_n2435_));
  NAND3_X1   g2386(.A1(new_n258_), .A2(new_n2428_), .A3(new_n2435_), .ZN(new_n2436_));
  NAND2_X1   g2387(.A1(new_n1543_), .A2(new_n1548_), .ZN(new_n2437_));
  NAND2_X1   g2388(.A1(new_n2437_), .A2(new_n2436_), .ZN(new_n2438_));
  INV_X1     g2389(.I(new_n2436_), .ZN(new_n2439_));
  NAND3_X1   g2390(.A1(new_n1543_), .A2(new_n1548_), .A3(new_n2439_), .ZN(new_n2440_));
  AOI21_X1   g2391(.A1(new_n2438_), .A2(new_n2440_), .B(new_n2421_), .ZN(new_n2441_));
  AND3_X2    g2392(.A1(new_n2438_), .A2(new_n2421_), .A3(new_n2440_), .Z(new_n2442_));
  NOR2_X1    g2393(.A1(new_n2442_), .A2(new_n2441_), .ZN(new_n2443_));
  NOR4_X1    g2394(.A1(new_n1090_), .A2(new_n435_), .A3(new_n338_), .A4(new_n261_), .ZN(new_n2444_));
  NAND2_X1   g2395(.A1(new_n294_), .A2(new_n146_), .ZN(new_n2445_));
  NOR4_X1    g2396(.A1(new_n2290_), .A2(new_n595_), .A3(new_n2444_), .A4(new_n2445_), .ZN(new_n2446_));
  INV_X1     g2397(.I(new_n2446_), .ZN(new_n2447_));
  NOR4_X1    g2398(.A1(new_n477_), .A2(new_n387_), .A3(new_n417_), .A4(new_n518_), .ZN(new_n2448_));
  NAND2_X1   g2399(.A1(new_n2448_), .A2(new_n2394_), .ZN(new_n2449_));
  NOR4_X1    g2400(.A1(new_n1065_), .A2(new_n2301_), .A3(new_n2447_), .A4(new_n2449_), .ZN(new_n2450_));
  NAND2_X1   g2401(.A1(new_n2443_), .A2(new_n2450_), .ZN(new_n2451_));
  NAND3_X1   g2402(.A1(new_n2404_), .A2(new_n2451_), .A3(new_n2419_), .ZN(new_n2452_));
  NAND2_X1   g2403(.A1(new_n1719_), .A2(new_n1714_), .ZN(new_n2453_));
  NAND2_X1   g2404(.A1(new_n1720_), .A2(new_n1715_), .ZN(new_n2454_));
  XOR2_X1    g2405(.A1(new_n2437_), .A2(new_n2420_), .Z(new_n2455_));
  NOR2_X1    g2406(.A1(new_n2455_), .A2(new_n2439_), .ZN(new_n2456_));
  AOI21_X1   g2407(.A1(new_n2454_), .A2(new_n2453_), .B(new_n2456_), .ZN(new_n2457_));
  AOI22_X1   g2408(.A1(new_n2452_), .A2(new_n2457_), .B1(new_n1715_), .B2(new_n1720_), .ZN(new_n2458_));
  OAI21_X1   g2409(.A1(new_n1678_), .A2(new_n1679_), .B(new_n1696_), .ZN(new_n2459_));
  AOI21_X1   g2410(.A1(new_n2458_), .A2(new_n2459_), .B(new_n1697_), .ZN(new_n2460_));
  AOI21_X1   g2411(.A1(new_n1588_), .A2(new_n1586_), .B(new_n1593_), .ZN(new_n2461_));
  AOI21_X1   g2412(.A1(new_n1490_), .A2(new_n1531_), .B(new_n1587_), .ZN(new_n2462_));
  NOR3_X1    g2413(.A1(new_n1550_), .A2(new_n1553_), .A3(new_n1585_), .ZN(new_n2463_));
  NOR3_X1    g2414(.A1(new_n2462_), .A2(new_n2463_), .A3(new_n1592_), .ZN(new_n2464_));
  NOR2_X1    g2415(.A1(new_n2464_), .A2(new_n2461_), .ZN(new_n2465_));
  NAND4_X1   g2416(.A1(new_n1653_), .A2(new_n211_), .A3(new_n408_), .A4(new_n419_), .ZN(new_n2466_));
  NOR3_X1    g2417(.A1(new_n204_), .A2(new_n434_), .A3(new_n535_), .ZN(new_n2467_));
  NOR4_X1    g2418(.A1(new_n715_), .A2(new_n865_), .A3(new_n500_), .A4(new_n501_), .ZN(new_n2468_));
  NOR2_X1    g2419(.A1(new_n1658_), .A2(new_n2468_), .ZN(new_n2469_));
  NAND4_X1   g2420(.A1(new_n2469_), .A2(new_n972_), .A3(new_n2390_), .A4(new_n2467_), .ZN(new_n2470_));
  NOR4_X1    g2421(.A1(new_n438_), .A2(new_n336_), .A3(new_n1091_), .A4(new_n361_), .ZN(new_n2471_));
  NOR4_X1    g2422(.A1(new_n758_), .A2(new_n2471_), .A3(new_n631_), .A4(new_n2314_), .ZN(new_n2472_));
  INV_X1     g2423(.I(new_n2472_), .ZN(new_n2473_));
  NOR2_X1    g2424(.A1(new_n483_), .A2(new_n471_), .ZN(new_n2474_));
  NOR3_X1    g2425(.A1(new_n271_), .A2(new_n869_), .A3(new_n326_), .ZN(new_n2475_));
  NAND4_X1   g2426(.A1(new_n2475_), .A2(new_n458_), .A3(new_n480_), .A4(new_n2474_), .ZN(new_n2476_));
  NOR4_X1    g2427(.A1(new_n2473_), .A2(new_n2476_), .A3(new_n1011_), .A4(new_n2378_), .ZN(new_n2477_));
  INV_X1     g2428(.I(new_n2477_), .ZN(new_n2478_));
  NOR3_X1    g2429(.A1(new_n2466_), .A2(new_n2470_), .A3(new_n2478_), .ZN(new_n2479_));
  XOR2_X1    g2430(.A1(new_n2465_), .A2(new_n2479_), .Z(new_n2480_));
  INV_X1     g2431(.I(new_n1667_), .ZN(new_n2481_));
  NAND3_X1   g2432(.A1(new_n2481_), .A2(new_n1662_), .A3(new_n1664_), .ZN(new_n2482_));
  OAI21_X1   g2433(.A1(new_n1665_), .A2(new_n1667_), .B(new_n1661_), .ZN(new_n2483_));
  INV_X1     g2434(.I(new_n2465_), .ZN(new_n2484_));
  NOR2_X1    g2435(.A1(new_n2484_), .A2(new_n2479_), .ZN(new_n2485_));
  AOI21_X1   g2436(.A1(new_n2483_), .A2(new_n2482_), .B(new_n2485_), .ZN(new_n2486_));
  OAI21_X1   g2437(.A1(new_n2460_), .A2(new_n2480_), .B(new_n2486_), .ZN(new_n2487_));
  NAND2_X1   g2438(.A1(new_n2487_), .A2(new_n1670_), .ZN(new_n2488_));
  INV_X1     g2439(.I(new_n2488_), .ZN(new_n2489_));
  NAND3_X1   g2440(.A1(new_n1594_), .A2(new_n1596_), .A3(new_n1616_), .ZN(new_n2490_));
  NOR2_X1    g2441(.A1(new_n1550_), .A2(new_n1553_), .ZN(new_n2491_));
  OAI22_X1   g2442(.A1(new_n2462_), .A2(new_n2463_), .B1(new_n2491_), .B2(new_n1592_), .ZN(new_n2492_));
  INV_X1     g2443(.I(new_n1596_), .ZN(new_n2493_));
  INV_X1     g2444(.I(new_n1616_), .ZN(new_n2494_));
  OAI21_X1   g2445(.A1(new_n2492_), .A2(new_n2493_), .B(new_n2494_), .ZN(new_n2495_));
  NAND2_X1   g2446(.A1(new_n2490_), .A2(new_n2495_), .ZN(new_n2496_));
  NAND2_X1   g2447(.A1(new_n2492_), .A2(new_n1596_), .ZN(new_n2497_));
  INV_X1     g2448(.I(new_n2497_), .ZN(new_n2498_));
  NOR2_X1    g2449(.A1(new_n2492_), .A2(new_n1596_), .ZN(new_n2499_));
  OAI21_X1   g2450(.A1(new_n2498_), .A2(new_n2499_), .B(new_n1620_), .ZN(new_n2500_));
  NOR2_X1    g2451(.A1(new_n2500_), .A2(new_n2496_), .ZN(new_n2501_));
  AND2_X2    g2452(.A1(new_n2490_), .A2(new_n2495_), .Z(new_n2502_));
  INV_X1     g2453(.I(new_n2499_), .ZN(new_n2503_));
  AOI22_X1   g2454(.A1(new_n2503_), .A2(new_n2497_), .B1(new_n1617_), .B2(new_n1619_), .ZN(new_n2504_));
  NOR2_X1    g2455(.A1(new_n2504_), .A2(new_n2502_), .ZN(new_n2505_));
  NOR2_X1    g2456(.A1(new_n2505_), .A2(new_n2501_), .ZN(new_n2506_));
  XOR2_X1    g2457(.A1(new_n707_), .A2(new_n670_), .Z(new_n2507_));
  INV_X1     g2458(.I(new_n745_), .ZN(new_n2508_));
  NOR4_X1    g2459(.A1(new_n305_), .A2(new_n435_), .A3(new_n204_), .A4(new_n507_), .ZN(new_n2509_));
  NAND3_X1   g2460(.A1(new_n769_), .A2(new_n310_), .A3(new_n319_), .ZN(new_n2510_));
  INV_X1     g2461(.I(new_n731_), .ZN(new_n2511_));
  OAI21_X1   g2462(.A1(new_n420_), .A2(new_n2511_), .B(new_n1646_), .ZN(new_n2512_));
  NOR4_X1    g2463(.A1(new_n2508_), .A2(new_n2509_), .A3(new_n2510_), .A4(new_n2512_), .ZN(new_n2513_));
  INV_X1     g2464(.I(new_n2513_), .ZN(new_n2514_));
  NAND2_X1   g2465(.A1(new_n284_), .A2(new_n375_), .ZN(new_n2515_));
  NOR4_X1    g2466(.A1(new_n2515_), .A2(new_n307_), .A3(new_n856_), .A4(new_n642_), .ZN(new_n2516_));
  NAND4_X1   g2467(.A1(new_n371_), .A2(new_n480_), .A3(new_n646_), .A4(new_n930_), .ZN(new_n2517_));
  INV_X1     g2468(.I(new_n476_), .ZN(new_n2518_));
  NOR4_X1    g2469(.A1(new_n862_), .A2(new_n620_), .A3(new_n2518_), .A4(new_n717_), .ZN(new_n2519_));
  NAND3_X1   g2470(.A1(new_n2519_), .A2(new_n2516_), .A3(new_n2517_), .ZN(new_n2520_));
  NOR4_X1    g2471(.A1(new_n2514_), .A2(new_n2296_), .A3(new_n2473_), .A4(new_n2520_), .ZN(new_n2521_));
  INV_X1     g2472(.I(new_n2521_), .ZN(new_n2522_));
  NAND2_X1   g2473(.A1(new_n1622_), .A2(new_n1623_), .ZN(new_n2523_));
  NAND2_X1   g2474(.A1(new_n2523_), .A2(new_n2522_), .ZN(new_n2524_));
  NAND3_X1   g2475(.A1(new_n1622_), .A2(new_n1623_), .A3(new_n2521_), .ZN(new_n2525_));
  NAND2_X1   g2476(.A1(new_n2524_), .A2(new_n2525_), .ZN(new_n2526_));
  XNOR2_X1   g2477(.A1(new_n2526_), .A2(new_n2507_), .ZN(new_n2527_));
  INV_X1     g2478(.I(new_n1094_), .ZN(new_n2528_));
  NOR2_X1    g2479(.A1(new_n2376_), .A2(new_n335_), .ZN(new_n2529_));
  NAND4_X1   g2480(.A1(new_n2529_), .A2(new_n395_), .A3(new_n427_), .A4(new_n554_), .ZN(new_n2530_));
  OR4_X2     g2481(.A1(new_n311_), .A2(new_n320_), .A3(new_n361_), .A4(new_n642_), .Z(new_n2531_));
  NOR4_X1    g2482(.A1(new_n2531_), .A2(new_n718_), .A3(new_n759_), .A4(new_n2530_), .ZN(new_n2532_));
  NAND4_X1   g2483(.A1(new_n2532_), .A2(new_n523_), .A3(new_n917_), .A4(new_n2528_), .ZN(new_n2533_));
  NOR2_X1    g2484(.A1(new_n2527_), .A2(new_n2533_), .ZN(new_n2534_));
  NOR3_X1    g2485(.A1(new_n2534_), .A2(new_n2489_), .A3(new_n2506_), .ZN(new_n2535_));
  INV_X1     g2486(.I(new_n2535_), .ZN(new_n2536_));
  XOR2_X1    g2487(.A1(new_n2523_), .A2(new_n2507_), .Z(new_n2537_));
  NOR2_X1    g2488(.A1(new_n2537_), .A2(new_n2521_), .ZN(new_n2538_));
  INV_X1     g2489(.I(new_n2538_), .ZN(new_n2539_));
  NAND3_X1   g2490(.A1(new_n2536_), .A2(new_n1638_), .A3(new_n2539_), .ZN(new_n2540_));
  NAND2_X1   g2491(.A1(new_n2540_), .A2(new_n1637_), .ZN(new_n2541_));
  NAND4_X1   g2492(.A1(new_n390_), .A2(new_n371_), .A3(new_n906_), .A4(new_n440_), .ZN(new_n2542_));
  NOR4_X1    g2493(.A1(new_n518_), .A2(new_n242_), .A3(new_n336_), .A4(new_n478_), .ZN(new_n2543_));
  NOR3_X1    g2494(.A1(new_n2542_), .A2(new_n880_), .A3(new_n2543_), .ZN(new_n2544_));
  INV_X1     g2495(.I(new_n437_), .ZN(new_n2545_));
  NOR3_X1    g2496(.A1(new_n500_), .A2(new_n584_), .A3(new_n246_), .ZN(new_n2546_));
  NAND4_X1   g2497(.A1(new_n2546_), .A2(new_n839_), .A3(new_n757_), .A4(new_n2545_), .ZN(new_n2547_));
  NOR2_X1    g2498(.A1(new_n1709_), .A2(new_n2547_), .ZN(new_n2548_));
  NAND4_X1   g2499(.A1(new_n2548_), .A2(new_n544_), .A3(new_n1013_), .A4(new_n2544_), .ZN(new_n2549_));
  INV_X1     g2500(.I(new_n2549_), .ZN(new_n2550_));
  XOR2_X1    g2501(.A1(new_n2541_), .A2(new_n2550_), .Z(new_n2551_));
  OAI21_X1   g2502(.A1(new_n2535_), .A2(new_n2538_), .B(new_n355_), .ZN(new_n2552_));
  INV_X1     g2503(.I(new_n2552_), .ZN(new_n2553_));
  NOR3_X1    g2504(.A1(new_n2535_), .A2(new_n355_), .A3(new_n2538_), .ZN(new_n2554_));
  OAI21_X1   g2505(.A1(new_n2553_), .A2(new_n2554_), .B(new_n1635_), .ZN(new_n2555_));
  NAND3_X1   g2506(.A1(new_n2536_), .A2(new_n354_), .A3(new_n2539_), .ZN(new_n2556_));
  NAND3_X1   g2507(.A1(new_n2556_), .A2(new_n1636_), .A3(new_n2552_), .ZN(new_n2557_));
  NAND2_X1   g2508(.A1(new_n2555_), .A2(new_n2557_), .ZN(new_n2558_));
  INV_X1     g2509(.I(new_n2558_), .ZN(new_n2559_));
  XOR2_X1    g2510(.A1(new_n2551_), .A2(new_n2559_), .Z(new_n2560_));
  INV_X1     g2511(.I(new_n2506_), .ZN(new_n2561_));
  XOR2_X1    g2512(.A1(new_n2526_), .A2(new_n2507_), .Z(new_n2562_));
  NAND3_X1   g2513(.A1(new_n2488_), .A2(new_n2562_), .A3(new_n2561_), .ZN(new_n2563_));
  INV_X1     g2514(.I(new_n2563_), .ZN(new_n2564_));
  AOI21_X1   g2515(.A1(new_n2488_), .A2(new_n2561_), .B(new_n2562_), .ZN(new_n2565_));
  INV_X1     g2516(.I(new_n2533_), .ZN(new_n2566_));
  NOR2_X1    g2517(.A1(new_n2488_), .A2(new_n2506_), .ZN(new_n2567_));
  AOI21_X1   g2518(.A1(new_n2487_), .A2(new_n1670_), .B(new_n2561_), .ZN(new_n2568_));
  OAI21_X1   g2519(.A1(new_n2567_), .A2(new_n2568_), .B(new_n2566_), .ZN(new_n2569_));
  NOR3_X1    g2520(.A1(new_n2569_), .A2(new_n2564_), .A3(new_n2565_), .ZN(new_n2570_));
  INV_X1     g2521(.I(new_n2565_), .ZN(new_n2571_));
  NAND3_X1   g2522(.A1(new_n2561_), .A2(new_n2487_), .A3(new_n1670_), .ZN(new_n2572_));
  NAND2_X1   g2523(.A1(new_n2488_), .A2(new_n2506_), .ZN(new_n2573_));
  AOI21_X1   g2524(.A1(new_n2573_), .A2(new_n2572_), .B(new_n2533_), .ZN(new_n2574_));
  AOI21_X1   g2525(.A1(new_n2563_), .A2(new_n2571_), .B(new_n2574_), .ZN(new_n2575_));
  NOR2_X1    g2526(.A1(new_n2575_), .A2(new_n2570_), .ZN(new_n2576_));
  INV_X1     g2527(.I(new_n2576_), .ZN(new_n2577_));
  OAI21_X1   g2528(.A1(new_n2505_), .A2(new_n2501_), .B(new_n2566_), .ZN(new_n2578_));
  NAND2_X1   g2529(.A1(new_n2504_), .A2(new_n2502_), .ZN(new_n2579_));
  NAND2_X1   g2530(.A1(new_n2500_), .A2(new_n2496_), .ZN(new_n2580_));
  NAND3_X1   g2531(.A1(new_n2579_), .A2(new_n2580_), .A3(new_n2533_), .ZN(new_n2581_));
  AOI22_X1   g2532(.A1(new_n2487_), .A2(new_n1670_), .B1(new_n2578_), .B2(new_n2581_), .ZN(new_n2582_));
  NAND3_X1   g2533(.A1(new_n2579_), .A2(new_n2580_), .A3(new_n2566_), .ZN(new_n2583_));
  OAI21_X1   g2534(.A1(new_n2505_), .A2(new_n2501_), .B(new_n2533_), .ZN(new_n2584_));
  NAND2_X1   g2535(.A1(new_n2584_), .A2(new_n2583_), .ZN(new_n2585_));
  AOI21_X1   g2536(.A1(new_n2489_), .A2(new_n2585_), .B(new_n2582_), .ZN(new_n2586_));
  OAI21_X1   g2537(.A1(new_n2575_), .A2(new_n2570_), .B(new_n2586_), .ZN(new_n2587_));
  NAND3_X1   g2538(.A1(new_n2574_), .A2(new_n2571_), .A3(new_n2563_), .ZN(new_n2588_));
  OAI21_X1   g2539(.A1(new_n2564_), .A2(new_n2565_), .B(new_n2569_), .ZN(new_n2589_));
  NAND2_X1   g2540(.A1(new_n2578_), .A2(new_n2581_), .ZN(new_n2590_));
  NAND2_X1   g2541(.A1(new_n2488_), .A2(new_n2590_), .ZN(new_n2591_));
  NAND3_X1   g2542(.A1(new_n2585_), .A2(new_n1670_), .A3(new_n2487_), .ZN(new_n2592_));
  NAND2_X1   g2543(.A1(new_n2591_), .A2(new_n2592_), .ZN(new_n2593_));
  NAND3_X1   g2544(.A1(new_n2589_), .A2(new_n2588_), .A3(new_n2593_), .ZN(new_n2594_));
  INV_X1     g2545(.I(new_n1668_), .ZN(new_n2595_));
  NOR2_X1    g2546(.A1(new_n2460_), .A2(new_n2480_), .ZN(new_n2596_));
  OAI21_X1   g2547(.A1(new_n2596_), .A2(new_n2485_), .B(new_n1661_), .ZN(new_n2597_));
  INV_X1     g2548(.I(new_n1679_), .ZN(new_n2598_));
  NAND3_X1   g2549(.A1(new_n2598_), .A2(new_n1677_), .A3(new_n1695_), .ZN(new_n2599_));
  NAND2_X1   g2550(.A1(new_n1720_), .A2(new_n1715_), .ZN(new_n2600_));
  NAND2_X1   g2551(.A1(new_n2452_), .A2(new_n2457_), .ZN(new_n2601_));
  NAND2_X1   g2552(.A1(new_n2601_), .A2(new_n2600_), .ZN(new_n2602_));
  NAND2_X1   g2553(.A1(new_n2459_), .A2(new_n2599_), .ZN(new_n2603_));
  OAI21_X1   g2554(.A1(new_n2603_), .A2(new_n2602_), .B(new_n2599_), .ZN(new_n2604_));
  INV_X1     g2555(.I(new_n2480_), .ZN(new_n2605_));
  NAND2_X1   g2556(.A1(new_n2604_), .A2(new_n2605_), .ZN(new_n2606_));
  INV_X1     g2557(.I(new_n2485_), .ZN(new_n2607_));
  NAND3_X1   g2558(.A1(new_n2606_), .A2(new_n1662_), .A3(new_n2607_), .ZN(new_n2608_));
  AOI21_X1   g2559(.A1(new_n2608_), .A2(new_n2597_), .B(new_n2595_), .ZN(new_n2609_));
  INV_X1     g2560(.I(new_n2597_), .ZN(new_n2610_));
  NOR3_X1    g2561(.A1(new_n2596_), .A2(new_n1661_), .A3(new_n2485_), .ZN(new_n2611_));
  NOR3_X1    g2562(.A1(new_n2610_), .A2(new_n1668_), .A3(new_n2611_), .ZN(new_n2612_));
  NOR3_X1    g2563(.A1(new_n2612_), .A2(new_n2586_), .A3(new_n2609_), .ZN(new_n2613_));
  OAI21_X1   g2564(.A1(new_n2610_), .A2(new_n2611_), .B(new_n1668_), .ZN(new_n2614_));
  NAND3_X1   g2565(.A1(new_n2608_), .A2(new_n2595_), .A3(new_n2597_), .ZN(new_n2615_));
  AOI21_X1   g2566(.A1(new_n2614_), .A2(new_n2615_), .B(new_n2593_), .ZN(new_n2616_));
  NOR2_X1    g2567(.A1(new_n2616_), .A2(new_n2613_), .ZN(new_n2617_));
  NAND3_X1   g2568(.A1(new_n2587_), .A2(new_n2594_), .A3(new_n2617_), .ZN(new_n2618_));
  NOR2_X1    g2569(.A1(new_n2612_), .A2(new_n2609_), .ZN(new_n2619_));
  OAI21_X1   g2570(.A1(new_n2576_), .A2(new_n2619_), .B(new_n2593_), .ZN(new_n2620_));
  NAND2_X1   g2571(.A1(new_n2614_), .A2(new_n2615_), .ZN(new_n2621_));
  NOR2_X1    g2572(.A1(new_n2460_), .A2(new_n2479_), .ZN(new_n2622_));
  INV_X1     g2573(.I(new_n2622_), .ZN(new_n2623_));
  NAND2_X1   g2574(.A1(new_n2460_), .A2(new_n2479_), .ZN(new_n2624_));
  AOI21_X1   g2575(.A1(new_n2623_), .A2(new_n2624_), .B(new_n2484_), .ZN(new_n2625_));
  INV_X1     g2576(.I(new_n2624_), .ZN(new_n2626_));
  NOR3_X1    g2577(.A1(new_n2626_), .A2(new_n2465_), .A3(new_n2622_), .ZN(new_n2627_));
  NOR2_X1    g2578(.A1(new_n2625_), .A2(new_n2627_), .ZN(new_n2628_));
  INV_X1     g2579(.I(new_n2628_), .ZN(new_n2629_));
  INV_X1     g2580(.I(new_n2456_), .ZN(new_n2630_));
  AOI21_X1   g2581(.A1(new_n2452_), .A2(new_n2630_), .B(new_n1714_), .ZN(new_n2631_));
  NAND3_X1   g2582(.A1(new_n2452_), .A2(new_n1714_), .A3(new_n2630_), .ZN(new_n2632_));
  INV_X1     g2583(.I(new_n2632_), .ZN(new_n2633_));
  OAI21_X1   g2584(.A1(new_n2633_), .A2(new_n2631_), .B(new_n1719_), .ZN(new_n2634_));
  INV_X1     g2585(.I(new_n2631_), .ZN(new_n2635_));
  NAND3_X1   g2586(.A1(new_n2635_), .A2(new_n1720_), .A3(new_n2632_), .ZN(new_n2636_));
  NAND2_X1   g2587(.A1(new_n2636_), .A2(new_n2634_), .ZN(new_n2637_));
  NAND3_X1   g2588(.A1(new_n2404_), .A2(new_n2419_), .A3(new_n2443_), .ZN(new_n2638_));
  INV_X1     g2589(.I(new_n2330_), .ZN(new_n2639_));
  AOI21_X1   g2590(.A1(new_n2365_), .A2(new_n2366_), .B(new_n2335_), .ZN(new_n2640_));
  NOR3_X1    g2591(.A1(new_n2363_), .A2(new_n2356_), .A3(new_n2336_), .ZN(new_n2641_));
  NAND2_X1   g2592(.A1(new_n2308_), .A2(new_n2329_), .ZN(new_n2642_));
  OAI21_X1   g2593(.A1(new_n2641_), .A2(new_n2640_), .B(new_n2642_), .ZN(new_n2643_));
  AOI21_X1   g2594(.A1(new_n2643_), .A2(new_n2639_), .B(new_n2398_), .ZN(new_n2644_));
  INV_X1     g2595(.I(new_n2402_), .ZN(new_n2645_));
  NAND3_X1   g2596(.A1(new_n2643_), .A2(new_n2639_), .A3(new_n2398_), .ZN(new_n2646_));
  AOI21_X1   g2597(.A1(new_n2645_), .A2(new_n2646_), .B(new_n2644_), .ZN(new_n2647_));
  INV_X1     g2598(.I(new_n2419_), .ZN(new_n2648_));
  OAI22_X1   g2599(.A1(new_n2647_), .A2(new_n2648_), .B1(new_n2441_), .B2(new_n2442_), .ZN(new_n2649_));
  NAND2_X1   g2600(.A1(new_n2649_), .A2(new_n2638_), .ZN(new_n2650_));
  NAND2_X1   g2601(.A1(new_n2364_), .A2(new_n2367_), .ZN(new_n2651_));
  AOI21_X1   g2602(.A1(new_n2651_), .A2(new_n2642_), .B(new_n2330_), .ZN(new_n2652_));
  AOI21_X1   g2603(.A1(new_n2652_), .A2(new_n2398_), .B(new_n2402_), .ZN(new_n2653_));
  NOR3_X1    g2604(.A1(new_n2653_), .A2(new_n2644_), .A3(new_n2648_), .ZN(new_n2654_));
  NOR2_X1    g2605(.A1(new_n2647_), .A2(new_n2419_), .ZN(new_n2655_));
  OAI21_X1   g2606(.A1(new_n2655_), .A2(new_n2654_), .B(new_n2450_), .ZN(new_n2656_));
  NOR2_X1    g2607(.A1(new_n2650_), .A2(new_n2656_), .ZN(new_n2657_));
  NAND2_X1   g2608(.A1(new_n2646_), .A2(new_n2645_), .ZN(new_n2658_));
  NAND3_X1   g2609(.A1(new_n2658_), .A2(new_n2400_), .A3(new_n2419_), .ZN(new_n2659_));
  NAND2_X1   g2610(.A1(new_n2404_), .A2(new_n2648_), .ZN(new_n2660_));
  NAND2_X1   g2611(.A1(new_n2660_), .A2(new_n2659_), .ZN(new_n2661_));
  AOI22_X1   g2612(.A1(new_n2661_), .A2(new_n2450_), .B1(new_n2638_), .B2(new_n2649_), .ZN(new_n2662_));
  NOR2_X1    g2613(.A1(new_n2657_), .A2(new_n2662_), .ZN(new_n2663_));
  AOI21_X1   g2614(.A1(new_n2646_), .A2(new_n2400_), .B(new_n2402_), .ZN(new_n2664_));
  NAND3_X1   g2615(.A1(new_n2643_), .A2(new_n2639_), .A3(new_n2399_), .ZN(new_n2665_));
  OAI21_X1   g2616(.A1(new_n2373_), .A2(new_n2330_), .B(new_n2398_), .ZN(new_n2666_));
  AOI21_X1   g2617(.A1(new_n2665_), .A2(new_n2666_), .B(new_n2645_), .ZN(new_n2667_));
  NOR2_X1    g2618(.A1(new_n2664_), .A2(new_n2667_), .ZN(new_n2668_));
  AOI22_X1   g2619(.A1(new_n2639_), .A2(new_n2642_), .B1(new_n2364_), .B2(new_n2367_), .ZN(new_n2669_));
  XOR2_X1    g2620(.A1(new_n2308_), .A2(new_n2371_), .Z(new_n2670_));
  NOR2_X1    g2621(.A1(new_n2670_), .A2(new_n2651_), .ZN(new_n2671_));
  NOR2_X1    g2622(.A1(new_n2671_), .A2(new_n2669_), .ZN(new_n2672_));
  INV_X1     g2623(.I(new_n2672_), .ZN(new_n2673_));
  OAI21_X1   g2624(.A1(new_n2644_), .A2(new_n2403_), .B(new_n2645_), .ZN(new_n2674_));
  NOR3_X1    g2625(.A1(new_n2373_), .A2(new_n2330_), .A3(new_n2398_), .ZN(new_n2675_));
  AOI21_X1   g2626(.A1(new_n2643_), .A2(new_n2639_), .B(new_n2399_), .ZN(new_n2676_));
  OAI21_X1   g2627(.A1(new_n2676_), .A2(new_n2675_), .B(new_n2402_), .ZN(new_n2677_));
  NOR3_X1    g2628(.A1(new_n2288_), .A2(new_n2368_), .A3(new_n2307_), .ZN(new_n2678_));
  AOI21_X1   g2629(.A1(new_n2289_), .A2(new_n2287_), .B(new_n2369_), .ZN(new_n2679_));
  NOR2_X1    g2630(.A1(new_n2678_), .A2(new_n2679_), .ZN(new_n2680_));
  AOI21_X1   g2631(.A1(new_n2674_), .A2(new_n2677_), .B(new_n2680_), .ZN(new_n2681_));
  NOR2_X1    g2632(.A1(new_n2681_), .A2(new_n2673_), .ZN(new_n2682_));
  NAND3_X1   g2633(.A1(new_n2418_), .A2(new_n2411_), .A3(new_n2450_), .ZN(new_n2683_));
  AOI21_X1   g2634(.A1(new_n2418_), .A2(new_n2411_), .B(new_n2450_), .ZN(new_n2684_));
  INV_X1     g2635(.I(new_n2684_), .ZN(new_n2685_));
  NAND2_X1   g2636(.A1(new_n2685_), .A2(new_n2683_), .ZN(new_n2686_));
  NOR3_X1    g2637(.A1(new_n2653_), .A2(new_n2644_), .A3(new_n2686_), .ZN(new_n2687_));
  INV_X1     g2638(.I(new_n2683_), .ZN(new_n2688_));
  NOR2_X1    g2639(.A1(new_n2688_), .A2(new_n2684_), .ZN(new_n2689_));
  AOI21_X1   g2640(.A1(new_n2658_), .A2(new_n2400_), .B(new_n2689_), .ZN(new_n2690_));
  NOR2_X1    g2641(.A1(new_n2690_), .A2(new_n2687_), .ZN(new_n2691_));
  NAND2_X1   g2642(.A1(new_n2637_), .A2(new_n2663_), .ZN(new_n2692_));
  INV_X1     g2643(.I(new_n2692_), .ZN(new_n2693_));
  NAND3_X1   g2644(.A1(new_n2458_), .A2(new_n2599_), .A3(new_n2459_), .ZN(new_n2694_));
  NAND2_X1   g2645(.A1(new_n2603_), .A2(new_n2602_), .ZN(new_n2695_));
  NAND2_X1   g2646(.A1(new_n2695_), .A2(new_n2694_), .ZN(new_n2696_));
  AND2_X2    g2647(.A1(new_n2636_), .A2(new_n2634_), .Z(new_n2697_));
  NAND4_X1   g2648(.A1(new_n2661_), .A2(new_n2450_), .A3(new_n2638_), .A4(new_n2649_), .ZN(new_n2698_));
  NAND2_X1   g2649(.A1(new_n2650_), .A2(new_n2656_), .ZN(new_n2699_));
  NAND2_X1   g2650(.A1(new_n2699_), .A2(new_n2698_), .ZN(new_n2700_));
  NAND2_X1   g2651(.A1(new_n2674_), .A2(new_n2677_), .ZN(new_n2701_));
  OAI21_X1   g2652(.A1(new_n2668_), .A2(new_n2680_), .B(new_n2672_), .ZN(new_n2702_));
  OAI21_X1   g2653(.A1(new_n2701_), .A2(new_n2702_), .B(new_n2663_), .ZN(new_n2703_));
  OAI21_X1   g2654(.A1(new_n2700_), .A2(new_n2703_), .B(new_n2697_), .ZN(new_n2704_));
  AOI21_X1   g2655(.A1(new_n2704_), .A2(new_n2696_), .B(new_n2693_), .ZN(new_n2705_));
  OAI21_X1   g2656(.A1(new_n2621_), .A2(new_n2705_), .B(new_n2629_), .ZN(new_n2706_));
  INV_X1     g2657(.I(new_n2706_), .ZN(new_n2707_));
  INV_X1     g2658(.I(new_n2696_), .ZN(new_n2708_));
  AOI21_X1   g2659(.A1(new_n2668_), .A2(new_n2682_), .B(new_n2700_), .ZN(new_n2709_));
  AOI21_X1   g2660(.A1(new_n2709_), .A2(new_n2663_), .B(new_n2637_), .ZN(new_n2710_));
  OAI21_X1   g2661(.A1(new_n2710_), .A2(new_n2708_), .B(new_n2692_), .ZN(new_n2711_));
  NAND3_X1   g2662(.A1(new_n2619_), .A2(new_n2628_), .A3(new_n2711_), .ZN(new_n2712_));
  NAND2_X1   g2663(.A1(new_n2712_), .A2(new_n2708_), .ZN(new_n2713_));
  OAI21_X1   g2664(.A1(new_n2621_), .A2(new_n2705_), .B(new_n2628_), .ZN(new_n2714_));
  OAI21_X1   g2665(.A1(new_n2713_), .A2(new_n2707_), .B(new_n2714_), .ZN(new_n2715_));
  NAND3_X1   g2666(.A1(new_n2715_), .A2(new_n2618_), .A3(new_n2620_), .ZN(new_n2716_));
  NAND3_X1   g2667(.A1(new_n2706_), .A2(new_n2712_), .A3(new_n2708_), .ZN(new_n2717_));
  NAND4_X1   g2668(.A1(new_n2618_), .A2(new_n2593_), .A3(new_n2717_), .A4(new_n2714_), .ZN(new_n2718_));
  AOI21_X1   g2669(.A1(new_n2716_), .A2(new_n2718_), .B(new_n2577_), .ZN(new_n2719_));
  NAND3_X1   g2670(.A1(new_n2716_), .A2(new_n2718_), .A3(new_n2577_), .ZN(new_n2720_));
  AOI21_X1   g2671(.A1(new_n2558_), .A2(new_n2720_), .B(new_n2719_), .ZN(new_n2721_));
  NAND2_X1   g2672(.A1(new_n2721_), .A2(new_n2560_), .ZN(new_n2722_));
  XOR2_X1    g2673(.A1(new_n2551_), .A2(new_n2558_), .Z(new_n2723_));
  AOI21_X1   g2674(.A1(new_n2589_), .A2(new_n2588_), .B(new_n2593_), .ZN(new_n2724_));
  NOR3_X1    g2675(.A1(new_n2575_), .A2(new_n2570_), .A3(new_n2586_), .ZN(new_n2725_));
  NOR4_X1    g2676(.A1(new_n2725_), .A2(new_n2724_), .A3(new_n2613_), .A4(new_n2616_), .ZN(new_n2726_));
  NOR2_X1    g2677(.A1(new_n2621_), .A2(new_n2705_), .ZN(new_n2727_));
  AOI21_X1   g2678(.A1(new_n2727_), .A2(new_n2628_), .B(new_n2696_), .ZN(new_n2728_));
  INV_X1     g2679(.I(new_n2714_), .ZN(new_n2729_));
  AOI21_X1   g2680(.A1(new_n2728_), .A2(new_n2706_), .B(new_n2729_), .ZN(new_n2730_));
  NOR3_X1    g2681(.A1(new_n2730_), .A2(new_n2726_), .A3(new_n2593_), .ZN(new_n2731_));
  AOI21_X1   g2682(.A1(new_n2715_), .A2(new_n2618_), .B(new_n2620_), .ZN(new_n2732_));
  OAI21_X1   g2683(.A1(new_n2731_), .A2(new_n2732_), .B(new_n2576_), .ZN(new_n2733_));
  NOR3_X1    g2684(.A1(new_n2731_), .A2(new_n2732_), .A3(new_n2576_), .ZN(new_n2734_));
  OAI21_X1   g2685(.A1(new_n2559_), .A2(new_n2734_), .B(new_n2733_), .ZN(new_n2735_));
  NAND2_X1   g2686(.A1(new_n2735_), .A2(new_n2723_), .ZN(new_n2736_));
  AOI21_X1   g2687(.A1(new_n2736_), .A2(new_n2722_), .B(new_n72_), .ZN(new_n2737_));
  XOR2_X1    g2688(.A1(new_n62_), .A2(new_n1326_), .Z(new_n2738_));
  INV_X1     g2689(.I(new_n69_), .ZN(new_n2739_));
  XOR2_X1    g2690(.A1(new_n62_), .A2(new_n2739_), .Z(new_n2740_));
  NOR3_X1    g2691(.A1(new_n63_), .A2(new_n2738_), .A3(new_n2740_), .ZN(new_n2741_));
  INV_X1     g2692(.I(new_n2741_), .ZN(new_n2742_));
  NOR2_X1    g2693(.A1(new_n2576_), .A2(new_n2742_), .ZN(new_n2743_));
  INV_X1     g2694(.I(new_n2743_), .ZN(new_n2744_));
  INV_X1     g2695(.I(new_n2551_), .ZN(new_n2745_));
  INV_X1     g2696(.I(new_n70_), .ZN(new_n2746_));
  NAND2_X1   g2697(.A1(new_n63_), .A2(new_n2746_), .ZN(new_n2747_));
  INV_X1     g2698(.I(new_n2747_), .ZN(new_n2748_));
  NAND2_X1   g2699(.A1(new_n2745_), .A2(new_n2748_), .ZN(new_n2749_));
  NOR3_X1    g2700(.A1(new_n1326_), .A2(new_n56_), .A3(new_n2739_), .ZN(new_n2750_));
  NOR3_X1    g2701(.A1(new_n1176_), .A2(new_n67_), .A3(new_n69_), .ZN(new_n2751_));
  NOR2_X1    g2702(.A1(new_n2751_), .A2(new_n2750_), .ZN(new_n2752_));
  INV_X1     g2703(.I(new_n2752_), .ZN(new_n2753_));
  AOI22_X1   g2704(.A1(new_n2749_), .A2(new_n2744_), .B1(new_n2559_), .B2(new_n2753_), .ZN(new_n2754_));
  INV_X1     g2705(.I(new_n2754_), .ZN(new_n2755_));
  NOR2_X1    g2706(.A1(new_n2737_), .A2(new_n2755_), .ZN(new_n2756_));
  NOR2_X1    g2707(.A1(new_n2619_), .A2(new_n2628_), .ZN(new_n2757_));
  AOI21_X1   g2708(.A1(new_n2717_), .A2(new_n2714_), .B(new_n2621_), .ZN(new_n2758_));
  OAI21_X1   g2709(.A1(new_n2758_), .A2(new_n2757_), .B(new_n2593_), .ZN(new_n2759_));
  NAND2_X1   g2710(.A1(new_n2621_), .A2(new_n2628_), .ZN(new_n2760_));
  NAND3_X1   g2711(.A1(new_n2717_), .A2(new_n2619_), .A3(new_n2714_), .ZN(new_n2761_));
  NAND2_X1   g2712(.A1(new_n2761_), .A2(new_n2760_), .ZN(new_n2762_));
  INV_X1     g2713(.I(new_n2762_), .ZN(new_n2763_));
  OAI21_X1   g2714(.A1(new_n2763_), .A2(new_n2593_), .B(new_n2759_), .ZN(new_n2764_));
  NOR3_X1    g2715(.A1(new_n1171_), .A2(new_n943_), .A3(new_n1053_), .ZN(new_n2765_));
  NOR2_X1    g2716(.A1(new_n1062_), .A2(new_n62_), .ZN(new_n2766_));
  AOI21_X1   g2717(.A1(new_n1171_), .A2(new_n2766_), .B(new_n2765_), .ZN(new_n2767_));
  NOR2_X1    g2718(.A1(new_n943_), .A2(new_n1053_), .ZN(new_n2768_));
  XOR2_X1    g2719(.A1(new_n939_), .A2(new_n943_), .Z(new_n2769_));
  INV_X1     g2720(.I(new_n2769_), .ZN(new_n2770_));
  OR3_X2     g2721(.A1(new_n2770_), .A2(new_n2768_), .A3(new_n2766_), .Z(new_n2771_));
  XOR2_X1    g2722(.A1(new_n1132_), .A2(new_n943_), .Z(new_n2772_));
  AND2_X2    g2723(.A1(new_n2771_), .A2(new_n2772_), .Z(new_n2773_));
  INV_X1     g2724(.I(new_n2773_), .ZN(new_n2774_));
  OAI22_X1   g2725(.A1(new_n2619_), .A2(new_n2767_), .B1(new_n2629_), .B2(new_n2774_), .ZN(new_n2775_));
  NOR2_X1    g2726(.A1(new_n1451_), .A2(new_n2770_), .ZN(new_n2776_));
  NAND2_X1   g2727(.A1(new_n2586_), .A2(new_n2776_), .ZN(new_n2777_));
  NOR2_X1    g2728(.A1(new_n1451_), .A2(new_n2769_), .ZN(new_n2778_));
  INV_X1     g2729(.I(new_n2778_), .ZN(new_n2779_));
  AOI21_X1   g2730(.A1(new_n2775_), .A2(new_n2777_), .B(new_n2779_), .ZN(new_n2780_));
  NAND3_X1   g2731(.A1(new_n2764_), .A2(new_n1132_), .A3(new_n2780_), .ZN(new_n2781_));
  INV_X1     g2732(.I(new_n2757_), .ZN(new_n2782_));
  NAND2_X1   g2733(.A1(new_n2715_), .A2(new_n2619_), .ZN(new_n2783_));
  AOI21_X1   g2734(.A1(new_n2783_), .A2(new_n2782_), .B(new_n2586_), .ZN(new_n2784_));
  AOI21_X1   g2735(.A1(new_n2761_), .A2(new_n2760_), .B(new_n2593_), .ZN(new_n2785_));
  OAI21_X1   g2736(.A1(new_n2784_), .A2(new_n2785_), .B(new_n2780_), .ZN(new_n2786_));
  NAND2_X1   g2737(.A1(new_n2786_), .A2(new_n1134_), .ZN(new_n2787_));
  INV_X1     g2738(.I(new_n2680_), .ZN(new_n2788_));
  XOR2_X1    g2739(.A1(new_n2672_), .A2(new_n2788_), .Z(new_n2789_));
  NOR2_X1    g2740(.A1(new_n685_), .A2(new_n1628_), .ZN(new_n2790_));
  INV_X1     g2741(.I(new_n2790_), .ZN(new_n2791_));
  NOR3_X1    g2742(.A1(new_n582_), .A2(new_n576_), .A3(new_n667_), .ZN(new_n2792_));
  NOR2_X1    g2743(.A1(new_n790_), .A2(new_n678_), .ZN(new_n2793_));
  AOI21_X1   g2744(.A1(new_n582_), .A2(new_n2793_), .B(new_n2792_), .ZN(new_n2794_));
  INV_X1     g2745(.I(new_n2794_), .ZN(new_n2795_));
  NAND2_X1   g2746(.A1(new_n686_), .A2(new_n1628_), .ZN(new_n2796_));
  AOI21_X1   g2747(.A1(new_n2680_), .A2(new_n2795_), .B(new_n2796_), .ZN(new_n2797_));
  OAI21_X1   g2748(.A1(new_n2673_), .A2(new_n2791_), .B(new_n2797_), .ZN(new_n2798_));
  NOR3_X1    g2749(.A1(new_n2789_), .A2(new_n2798_), .A3(new_n659_), .ZN(new_n2799_));
  NOR2_X1    g2750(.A1(new_n2789_), .A2(new_n2798_), .ZN(new_n2800_));
  NOR2_X1    g2751(.A1(new_n2800_), .A2(new_n658_), .ZN(new_n2801_));
  NOR2_X1    g2752(.A1(new_n2801_), .A2(new_n2799_), .ZN(new_n2802_));
  NOR2_X1    g2753(.A1(new_n2788_), .A2(new_n685_), .ZN(new_n2803_));
  NOR2_X1    g2754(.A1(new_n2803_), .A2(new_n659_), .ZN(new_n2804_));
  NAND2_X1   g2755(.A1(new_n2802_), .A2(new_n2804_), .ZN(new_n2805_));
  NAND3_X1   g2756(.A1(new_n2364_), .A2(new_n2367_), .A3(new_n2370_), .ZN(new_n2806_));
  INV_X1     g2757(.I(new_n2806_), .ZN(new_n2807_));
  AOI21_X1   g2758(.A1(new_n2364_), .A2(new_n2367_), .B(new_n2370_), .ZN(new_n2808_));
  OAI21_X1   g2759(.A1(new_n2807_), .A2(new_n2808_), .B(new_n2329_), .ZN(new_n2809_));
  INV_X1     g2760(.I(new_n2808_), .ZN(new_n2810_));
  NAND3_X1   g2761(.A1(new_n2810_), .A2(new_n2371_), .A3(new_n2806_), .ZN(new_n2811_));
  AOI21_X1   g2762(.A1(new_n2811_), .A2(new_n2809_), .B(new_n2788_), .ZN(new_n2812_));
  OAI21_X1   g2763(.A1(new_n2373_), .A2(new_n2330_), .B(new_n2402_), .ZN(new_n2813_));
  NOR3_X1    g2764(.A1(new_n2373_), .A2(new_n2330_), .A3(new_n2402_), .ZN(new_n2814_));
  INV_X1     g2765(.I(new_n2814_), .ZN(new_n2815_));
  AOI21_X1   g2766(.A1(new_n2815_), .A2(new_n2813_), .B(new_n2399_), .ZN(new_n2816_));
  INV_X1     g2767(.I(new_n2816_), .ZN(new_n2817_));
  NAND3_X1   g2768(.A1(new_n2815_), .A2(new_n2399_), .A3(new_n2813_), .ZN(new_n2818_));
  AOI21_X1   g2769(.A1(new_n2817_), .A2(new_n2818_), .B(new_n2812_), .ZN(new_n2819_));
  INV_X1     g2770(.I(new_n2812_), .ZN(new_n2820_));
  INV_X1     g2771(.I(new_n2818_), .ZN(new_n2821_));
  NOR3_X1    g2772(.A1(new_n2820_), .A2(new_n2821_), .A3(new_n2816_), .ZN(new_n2822_));
  NOR2_X1    g2773(.A1(new_n2822_), .A2(new_n2819_), .ZN(new_n2823_));
  INV_X1     g2774(.I(new_n2796_), .ZN(new_n2824_));
  NOR2_X1    g2775(.A1(new_n576_), .A2(new_n667_), .ZN(new_n2825_));
  NOR3_X1    g2776(.A1(new_n686_), .A2(new_n2825_), .A3(new_n2793_), .ZN(new_n2826_));
  XOR2_X1    g2777(.A1(new_n576_), .A2(new_n658_), .Z(new_n2827_));
  INV_X1     g2778(.I(new_n2827_), .ZN(new_n2828_));
  NOR2_X1    g2779(.A1(new_n2826_), .A2(new_n2828_), .ZN(new_n2829_));
  INV_X1     g2780(.I(new_n2829_), .ZN(new_n2830_));
  OAI22_X1   g2781(.A1(new_n2673_), .A2(new_n2794_), .B1(new_n2788_), .B2(new_n2830_), .ZN(new_n2831_));
  OAI21_X1   g2782(.A1(new_n2701_), .A2(new_n2791_), .B(new_n2831_), .ZN(new_n2832_));
  NAND2_X1   g2783(.A1(new_n2832_), .A2(new_n2824_), .ZN(new_n2833_));
  NOR2_X1    g2784(.A1(new_n2833_), .A2(new_n2823_), .ZN(new_n2834_));
  XOR2_X1    g2785(.A1(new_n2834_), .A2(new_n658_), .Z(new_n2835_));
  XOR2_X1    g2786(.A1(new_n2835_), .A2(new_n2805_), .Z(new_n2836_));
  INV_X1     g2787(.I(new_n2836_), .ZN(new_n2837_));
  NAND4_X1   g2788(.A1(new_n2637_), .A2(new_n2663_), .A3(new_n2668_), .A4(new_n2682_), .ZN(new_n2838_));
  NOR3_X1    g2789(.A1(new_n2700_), .A2(new_n2701_), .A3(new_n2702_), .ZN(new_n2839_));
  OR2_X2     g2790(.A1(new_n2839_), .A2(new_n2637_), .Z(new_n2840_));
  NAND2_X1   g2791(.A1(new_n2840_), .A2(new_n2838_), .ZN(new_n2841_));
  NAND3_X1   g2792(.A1(new_n2658_), .A2(new_n2400_), .A3(new_n2689_), .ZN(new_n2842_));
  OAI21_X1   g2793(.A1(new_n2653_), .A2(new_n2644_), .B(new_n2686_), .ZN(new_n2843_));
  NAND2_X1   g2794(.A1(new_n2843_), .A2(new_n2842_), .ZN(new_n2844_));
  XOR2_X1    g2795(.A1(new_n576_), .A2(new_n1125_), .Z(new_n2845_));
  XOR2_X1    g2796(.A1(new_n576_), .A2(new_n1132_), .Z(new_n2846_));
  XOR2_X1    g2797(.A1(new_n576_), .A2(new_n1106_), .Z(new_n2847_));
  NOR3_X1    g2798(.A1(new_n2845_), .A2(new_n2846_), .A3(new_n2847_), .ZN(new_n2848_));
  NOR3_X1    g2799(.A1(new_n1153_), .A2(new_n1132_), .A3(new_n1125_), .ZN(new_n2849_));
  AOI21_X1   g2800(.A1(new_n1576_), .A2(new_n1132_), .B(new_n2849_), .ZN(new_n2850_));
  INV_X1     g2801(.I(new_n2850_), .ZN(new_n2851_));
  AOI22_X1   g2802(.A1(new_n2700_), .A2(new_n2851_), .B1(new_n2844_), .B2(new_n2848_), .ZN(new_n2852_));
  INV_X1     g2803(.I(new_n2847_), .ZN(new_n2853_));
  XNOR2_X1   g2804(.A1(new_n1132_), .A2(new_n1125_), .ZN(new_n2854_));
  NOR2_X1    g2805(.A1(new_n2853_), .A2(new_n2854_), .ZN(new_n2855_));
  INV_X1     g2806(.I(new_n2855_), .ZN(new_n2856_));
  NOR2_X1    g2807(.A1(new_n2637_), .A2(new_n2856_), .ZN(new_n2857_));
  NOR2_X1    g2808(.A1(new_n2847_), .A2(new_n2854_), .ZN(new_n2858_));
  OAI21_X1   g2809(.A1(new_n2857_), .A2(new_n2852_), .B(new_n2858_), .ZN(new_n2859_));
  INV_X1     g2810(.I(new_n2859_), .ZN(new_n2860_));
  NAND3_X1   g2811(.A1(new_n2860_), .A2(new_n2841_), .A3(new_n790_), .ZN(new_n2861_));
  INV_X1     g2812(.I(new_n2838_), .ZN(new_n2862_));
  NOR2_X1    g2813(.A1(new_n2839_), .A2(new_n2637_), .ZN(new_n2863_));
  NOR2_X1    g2814(.A1(new_n2862_), .A2(new_n2863_), .ZN(new_n2864_));
  OAI21_X1   g2815(.A1(new_n2864_), .A2(new_n2859_), .B(new_n576_), .ZN(new_n2865_));
  NAND2_X1   g2816(.A1(new_n2865_), .A2(new_n2861_), .ZN(new_n2866_));
  NOR2_X1    g2817(.A1(new_n2866_), .A2(new_n2837_), .ZN(new_n2867_));
  AOI21_X1   g2818(.A1(new_n2861_), .A2(new_n2865_), .B(new_n2836_), .ZN(new_n2868_));
  NOR2_X1    g2819(.A1(new_n2682_), .A2(new_n2844_), .ZN(new_n2869_));
  NOR3_X1    g2820(.A1(new_n2691_), .A2(new_n2673_), .A3(new_n2681_), .ZN(new_n2870_));
  NAND3_X1   g2821(.A1(new_n2701_), .A2(new_n2672_), .A3(new_n2680_), .ZN(new_n2871_));
  NAND2_X1   g2822(.A1(new_n2668_), .A2(new_n2673_), .ZN(new_n2872_));
  NAND2_X1   g2823(.A1(new_n2871_), .A2(new_n2872_), .ZN(new_n2873_));
  NOR3_X1    g2824(.A1(new_n2869_), .A2(new_n2873_), .A3(new_n2870_), .ZN(new_n2874_));
  NOR2_X1    g2825(.A1(new_n2874_), .A2(new_n2700_), .ZN(new_n2875_));
  NAND2_X1   g2826(.A1(new_n2702_), .A2(new_n2691_), .ZN(new_n2876_));
  NAND2_X1   g2827(.A1(new_n2682_), .A2(new_n2844_), .ZN(new_n2877_));
  NAND4_X1   g2828(.A1(new_n2877_), .A2(new_n2876_), .A3(new_n2871_), .A4(new_n2872_), .ZN(new_n2878_));
  NOR2_X1    g2829(.A1(new_n2878_), .A2(new_n2663_), .ZN(new_n2879_));
  NOR2_X1    g2830(.A1(new_n2879_), .A2(new_n2875_), .ZN(new_n2880_));
  INV_X1     g2831(.I(new_n2858_), .ZN(new_n2881_));
  INV_X1     g2832(.I(new_n2848_), .ZN(new_n2882_));
  OAI22_X1   g2833(.A1(new_n2691_), .A2(new_n2850_), .B1(new_n2701_), .B2(new_n2882_), .ZN(new_n2883_));
  NAND2_X1   g2834(.A1(new_n2700_), .A2(new_n2855_), .ZN(new_n2884_));
  AOI21_X1   g2835(.A1(new_n2884_), .A2(new_n2883_), .B(new_n2881_), .ZN(new_n2885_));
  NAND3_X1   g2836(.A1(new_n2880_), .A2(new_n2885_), .A3(new_n790_), .ZN(new_n2886_));
  AOI21_X1   g2837(.A1(new_n2880_), .A2(new_n2885_), .B(new_n790_), .ZN(new_n2887_));
  INV_X1     g2838(.I(new_n2887_), .ZN(new_n2888_));
  NAND2_X1   g2839(.A1(new_n2888_), .A2(new_n2886_), .ZN(new_n2889_));
  INV_X1     g2840(.I(new_n2889_), .ZN(new_n2890_));
  XNOR2_X1   g2841(.A1(new_n2802_), .A2(new_n2804_), .ZN(new_n2891_));
  NAND2_X1   g2842(.A1(new_n2890_), .A2(new_n2891_), .ZN(new_n2892_));
  INV_X1     g2843(.I(new_n2891_), .ZN(new_n2893_));
  NAND2_X1   g2844(.A1(new_n2889_), .A2(new_n2893_), .ZN(new_n2894_));
  AOI21_X1   g2845(.A1(new_n2871_), .A2(new_n2872_), .B(new_n2691_), .ZN(new_n2895_));
  NAND2_X1   g2846(.A1(new_n2668_), .A2(new_n2672_), .ZN(new_n2896_));
  OAI22_X1   g2847(.A1(new_n2673_), .A2(new_n2788_), .B1(new_n2664_), .B2(new_n2667_), .ZN(new_n2897_));
  AOI21_X1   g2848(.A1(new_n2896_), .A2(new_n2897_), .B(new_n2844_), .ZN(new_n2898_));
  NOR2_X1    g2849(.A1(new_n2895_), .A2(new_n2898_), .ZN(new_n2899_));
  OAI22_X1   g2850(.A1(new_n2701_), .A2(new_n2850_), .B1(new_n2673_), .B2(new_n2882_), .ZN(new_n2900_));
  OAI21_X1   g2851(.A1(new_n2691_), .A2(new_n2856_), .B(new_n2900_), .ZN(new_n2901_));
  NAND3_X1   g2852(.A1(new_n2899_), .A2(new_n2858_), .A3(new_n2901_), .ZN(new_n2902_));
  XOR2_X1    g2853(.A1(new_n2902_), .A2(new_n576_), .Z(new_n2903_));
  INV_X1     g2854(.I(new_n2803_), .ZN(new_n2904_));
  AOI21_X1   g2855(.A1(new_n2680_), .A2(new_n2851_), .B(new_n2881_), .ZN(new_n2905_));
  OAI21_X1   g2856(.A1(new_n2673_), .A2(new_n2856_), .B(new_n2905_), .ZN(new_n2906_));
  NOR3_X1    g2857(.A1(new_n2789_), .A2(new_n2906_), .A3(new_n576_), .ZN(new_n2907_));
  NOR2_X1    g2858(.A1(new_n2789_), .A2(new_n2906_), .ZN(new_n2908_));
  NOR2_X1    g2859(.A1(new_n2908_), .A2(new_n790_), .ZN(new_n2909_));
  NOR2_X1    g2860(.A1(new_n2909_), .A2(new_n2907_), .ZN(new_n2910_));
  NOR2_X1    g2861(.A1(new_n2788_), .A2(new_n2854_), .ZN(new_n2911_));
  OAI21_X1   g2862(.A1(new_n2816_), .A2(new_n2821_), .B(new_n2820_), .ZN(new_n2912_));
  NAND3_X1   g2863(.A1(new_n2817_), .A2(new_n2812_), .A3(new_n2818_), .ZN(new_n2913_));
  NAND2_X1   g2864(.A1(new_n2912_), .A2(new_n2913_), .ZN(new_n2914_));
  OAI22_X1   g2865(.A1(new_n2673_), .A2(new_n2850_), .B1(new_n2788_), .B2(new_n2882_), .ZN(new_n2915_));
  NAND2_X1   g2866(.A1(new_n2668_), .A2(new_n2855_), .ZN(new_n2916_));
  NAND2_X1   g2867(.A1(new_n2916_), .A2(new_n2915_), .ZN(new_n2917_));
  NAND3_X1   g2868(.A1(new_n2914_), .A2(new_n2858_), .A3(new_n2917_), .ZN(new_n2918_));
  NOR4_X1    g2869(.A1(new_n2918_), .A2(new_n2910_), .A3(new_n576_), .A4(new_n2911_), .ZN(new_n2919_));
  NOR2_X1    g2870(.A1(new_n2919_), .A2(new_n2904_), .ZN(new_n2920_));
  INV_X1     g2871(.I(new_n2911_), .ZN(new_n2921_));
  INV_X1     g2872(.I(new_n2917_), .ZN(new_n2922_));
  NOR3_X1    g2873(.A1(new_n2922_), .A2(new_n2823_), .A3(new_n2881_), .ZN(new_n2923_));
  NAND4_X1   g2874(.A1(new_n2923_), .A2(new_n790_), .A3(new_n2908_), .A4(new_n2921_), .ZN(new_n2924_));
  NOR2_X1    g2875(.A1(new_n2924_), .A2(new_n2803_), .ZN(new_n2925_));
  NOR2_X1    g2876(.A1(new_n2920_), .A2(new_n2925_), .ZN(new_n2926_));
  NOR2_X1    g2877(.A1(new_n2924_), .A2(new_n2904_), .ZN(new_n2927_));
  INV_X1     g2878(.I(new_n2927_), .ZN(new_n2928_));
  OAI21_X1   g2879(.A1(new_n2926_), .A2(new_n2903_), .B(new_n2928_), .ZN(new_n2929_));
  INV_X1     g2880(.I(new_n2929_), .ZN(new_n2930_));
  NAND2_X1   g2881(.A1(new_n2894_), .A2(new_n2930_), .ZN(new_n2931_));
  NAND2_X1   g2882(.A1(new_n2931_), .A2(new_n2892_), .ZN(new_n2932_));
  OAI22_X1   g2883(.A1(new_n2932_), .A2(new_n2837_), .B1(new_n2867_), .B2(new_n2868_), .ZN(new_n2933_));
  NAND2_X1   g2884(.A1(new_n2637_), .A2(new_n2700_), .ZN(new_n2934_));
  NAND3_X1   g2885(.A1(new_n2697_), .A2(new_n2709_), .A3(new_n2663_), .ZN(new_n2935_));
  AOI21_X1   g2886(.A1(new_n2935_), .A2(new_n2934_), .B(new_n2708_), .ZN(new_n2936_));
  AOI21_X1   g2887(.A1(new_n2704_), .A2(new_n2692_), .B(new_n2696_), .ZN(new_n2937_));
  OAI22_X1   g2888(.A1(new_n2637_), .A2(new_n2850_), .B1(new_n2663_), .B2(new_n2882_), .ZN(new_n2938_));
  NAND2_X1   g2889(.A1(new_n2708_), .A2(new_n2855_), .ZN(new_n2939_));
  AOI21_X1   g2890(.A1(new_n2939_), .A2(new_n2938_), .B(new_n2881_), .ZN(new_n2940_));
  OAI21_X1   g2891(.A1(new_n2937_), .A2(new_n2936_), .B(new_n2940_), .ZN(new_n2941_));
  NOR2_X1    g2892(.A1(new_n2941_), .A2(new_n576_), .ZN(new_n2942_));
  NAND2_X1   g2893(.A1(new_n2941_), .A2(new_n576_), .ZN(new_n2943_));
  INV_X1     g2894(.I(new_n2943_), .ZN(new_n2944_));
  NAND3_X1   g2895(.A1(new_n2914_), .A2(new_n2824_), .A3(new_n2832_), .ZN(new_n2945_));
  NOR4_X1    g2896(.A1(new_n2945_), .A2(new_n659_), .A3(new_n2800_), .A4(new_n2803_), .ZN(new_n2946_));
  NOR3_X1    g2897(.A1(new_n2668_), .A2(new_n2673_), .A3(new_n2788_), .ZN(new_n2947_));
  NOR2_X1    g2898(.A1(new_n2701_), .A2(new_n2672_), .ZN(new_n2948_));
  OAI21_X1   g2899(.A1(new_n2947_), .A2(new_n2948_), .B(new_n2844_), .ZN(new_n2949_));
  NOR2_X1    g2900(.A1(new_n2701_), .A2(new_n2673_), .ZN(new_n2950_));
  AOI22_X1   g2901(.A1(new_n2674_), .A2(new_n2677_), .B1(new_n2672_), .B2(new_n2680_), .ZN(new_n2951_));
  OAI21_X1   g2902(.A1(new_n2950_), .A2(new_n2951_), .B(new_n2691_), .ZN(new_n2952_));
  OAI22_X1   g2903(.A1(new_n2701_), .A2(new_n2794_), .B1(new_n2673_), .B2(new_n2830_), .ZN(new_n2953_));
  AOI21_X1   g2904(.A1(new_n2843_), .A2(new_n2842_), .B(new_n2791_), .ZN(new_n2954_));
  INV_X1     g2905(.I(new_n2954_), .ZN(new_n2955_));
  AOI21_X1   g2906(.A1(new_n2955_), .A2(new_n2953_), .B(new_n2796_), .ZN(new_n2956_));
  NAND4_X1   g2907(.A1(new_n2956_), .A2(new_n2949_), .A3(new_n2952_), .A4(new_n658_), .ZN(new_n2957_));
  NAND2_X1   g2908(.A1(new_n2949_), .A2(new_n2952_), .ZN(new_n2958_));
  AOI22_X1   g2909(.A1(new_n2668_), .A2(new_n2795_), .B1(new_n2672_), .B2(new_n2829_), .ZN(new_n2959_));
  OAI21_X1   g2910(.A1(new_n2959_), .A2(new_n2954_), .B(new_n2824_), .ZN(new_n2960_));
  OAI21_X1   g2911(.A1(new_n2958_), .A2(new_n2960_), .B(new_n659_), .ZN(new_n2961_));
  NOR2_X1    g2912(.A1(new_n2788_), .A2(new_n659_), .ZN(new_n2962_));
  INV_X1     g2913(.I(new_n2962_), .ZN(new_n2963_));
  NAND3_X1   g2914(.A1(new_n2961_), .A2(new_n2957_), .A3(new_n2963_), .ZN(new_n2964_));
  NAND4_X1   g2915(.A1(new_n2899_), .A2(new_n658_), .A3(new_n2680_), .A4(new_n2956_), .ZN(new_n2965_));
  AOI21_X1   g2916(.A1(new_n2964_), .A2(new_n2965_), .B(new_n2946_), .ZN(new_n2966_));
  NAND4_X1   g2917(.A1(new_n2834_), .A2(new_n2802_), .A3(new_n658_), .A4(new_n2904_), .ZN(new_n2967_));
  NOR4_X1    g2918(.A1(new_n2960_), .A2(new_n2895_), .A3(new_n2898_), .A4(new_n659_), .ZN(new_n2968_));
  AOI21_X1   g2919(.A1(new_n2899_), .A2(new_n2956_), .B(new_n658_), .ZN(new_n2969_));
  NOR3_X1    g2920(.A1(new_n2969_), .A2(new_n2968_), .A3(new_n2962_), .ZN(new_n2970_));
  INV_X1     g2921(.I(new_n2965_), .ZN(new_n2971_));
  NOR3_X1    g2922(.A1(new_n2970_), .A2(new_n2971_), .A3(new_n2967_), .ZN(new_n2972_));
  NOR2_X1    g2923(.A1(new_n2972_), .A2(new_n2966_), .ZN(new_n2973_));
  INV_X1     g2924(.I(new_n2973_), .ZN(new_n2974_));
  OAI21_X1   g2925(.A1(new_n2944_), .A2(new_n2942_), .B(new_n2974_), .ZN(new_n2975_));
  INV_X1     g2926(.I(new_n2942_), .ZN(new_n2976_));
  NAND3_X1   g2927(.A1(new_n2976_), .A2(new_n2943_), .A3(new_n2973_), .ZN(new_n2977_));
  AOI21_X1   g2928(.A1(new_n2975_), .A2(new_n2977_), .B(new_n2933_), .ZN(new_n2978_));
  NOR2_X1    g2929(.A1(new_n2867_), .A2(new_n2868_), .ZN(new_n2979_));
  NOR2_X1    g2930(.A1(new_n2889_), .A2(new_n2893_), .ZN(new_n2980_));
  AOI21_X1   g2931(.A1(new_n2889_), .A2(new_n2893_), .B(new_n2929_), .ZN(new_n2981_));
  NOR2_X1    g2932(.A1(new_n2981_), .A2(new_n2980_), .ZN(new_n2982_));
  AOI21_X1   g2933(.A1(new_n2836_), .A2(new_n2982_), .B(new_n2979_), .ZN(new_n2983_));
  NOR3_X1    g2934(.A1(new_n2944_), .A2(new_n2942_), .A3(new_n2973_), .ZN(new_n2984_));
  INV_X1     g2935(.I(new_n2984_), .ZN(new_n2985_));
  AOI21_X1   g2936(.A1(new_n2976_), .A2(new_n2943_), .B(new_n2974_), .ZN(new_n2986_));
  INV_X1     g2937(.I(new_n2986_), .ZN(new_n2987_));
  AOI21_X1   g2938(.A1(new_n2985_), .A2(new_n2987_), .B(new_n2983_), .ZN(new_n2988_));
  NOR2_X1    g2939(.A1(new_n2988_), .A2(new_n2978_), .ZN(new_n2989_));
  NAND3_X1   g2940(.A1(new_n2781_), .A2(new_n2989_), .A3(new_n2787_), .ZN(new_n2990_));
  NOR2_X1    g2941(.A1(new_n2786_), .A2(new_n1134_), .ZN(new_n2991_));
  AOI21_X1   g2942(.A1(new_n2764_), .A2(new_n2780_), .B(new_n1132_), .ZN(new_n2992_));
  NAND2_X1   g2943(.A1(new_n2975_), .A2(new_n2977_), .ZN(new_n2993_));
  NAND2_X1   g2944(.A1(new_n2983_), .A2(new_n2993_), .ZN(new_n2994_));
  OAI21_X1   g2945(.A1(new_n2984_), .A2(new_n2986_), .B(new_n2933_), .ZN(new_n2995_));
  NAND2_X1   g2946(.A1(new_n2995_), .A2(new_n2994_), .ZN(new_n2996_));
  OAI21_X1   g2947(.A1(new_n2992_), .A2(new_n2991_), .B(new_n2996_), .ZN(new_n2997_));
  NAND3_X1   g2948(.A1(new_n2710_), .A2(new_n2692_), .A3(new_n2696_), .ZN(new_n2998_));
  NAND2_X1   g2949(.A1(new_n2693_), .A2(new_n2708_), .ZN(new_n2999_));
  NAND2_X1   g2950(.A1(new_n2998_), .A2(new_n2999_), .ZN(new_n3000_));
  INV_X1     g2951(.I(new_n3000_), .ZN(new_n3001_));
  NOR2_X1    g2952(.A1(new_n2629_), .A2(new_n2705_), .ZN(new_n3002_));
  NOR2_X1    g2953(.A1(new_n2711_), .A2(new_n2628_), .ZN(new_n3003_));
  NOR4_X1    g2954(.A1(new_n3001_), .A2(new_n3002_), .A3(new_n2621_), .A4(new_n3003_), .ZN(new_n3004_));
  NOR3_X1    g2955(.A1(new_n3001_), .A2(new_n3002_), .A3(new_n3003_), .ZN(new_n3005_));
  NOR2_X1    g2956(.A1(new_n3005_), .A2(new_n2619_), .ZN(new_n3006_));
  INV_X1     g2957(.I(new_n2776_), .ZN(new_n3007_));
  OAI22_X1   g2958(.A1(new_n2619_), .A2(new_n3007_), .B1(new_n2696_), .B2(new_n2774_), .ZN(new_n3008_));
  INV_X1     g2959(.I(new_n2767_), .ZN(new_n3009_));
  NAND2_X1   g2960(.A1(new_n2628_), .A2(new_n3009_), .ZN(new_n3010_));
  AOI21_X1   g2961(.A1(new_n3008_), .A2(new_n3010_), .B(new_n2779_), .ZN(new_n3011_));
  OAI21_X1   g2962(.A1(new_n3006_), .A2(new_n3004_), .B(new_n3011_), .ZN(new_n3012_));
  NOR2_X1    g2963(.A1(new_n3012_), .A2(new_n1134_), .ZN(new_n3013_));
  XOR2_X1    g2964(.A1(new_n3005_), .A2(new_n2621_), .Z(new_n3014_));
  AOI21_X1   g2965(.A1(new_n3014_), .A2(new_n3011_), .B(new_n1132_), .ZN(new_n3015_));
  INV_X1     g2966(.I(new_n2805_), .ZN(new_n3016_));
  INV_X1     g2967(.I(new_n2866_), .ZN(new_n3017_));
  AOI21_X1   g2968(.A1(new_n2931_), .A2(new_n2892_), .B(new_n3017_), .ZN(new_n3018_));
  NOR3_X1    g2969(.A1(new_n2981_), .A2(new_n2980_), .A3(new_n2866_), .ZN(new_n3019_));
  OAI21_X1   g2970(.A1(new_n3018_), .A2(new_n3019_), .B(new_n2835_), .ZN(new_n3020_));
  INV_X1     g2971(.I(new_n2835_), .ZN(new_n3021_));
  OAI21_X1   g2972(.A1(new_n2981_), .A2(new_n2980_), .B(new_n2866_), .ZN(new_n3022_));
  NAND3_X1   g2973(.A1(new_n2931_), .A2(new_n3017_), .A3(new_n2892_), .ZN(new_n3023_));
  NAND3_X1   g2974(.A1(new_n3023_), .A2(new_n3022_), .A3(new_n3021_), .ZN(new_n3024_));
  AOI21_X1   g2975(.A1(new_n3020_), .A2(new_n3024_), .B(new_n3016_), .ZN(new_n3025_));
  AOI21_X1   g2976(.A1(new_n3023_), .A2(new_n3022_), .B(new_n3021_), .ZN(new_n3026_));
  NOR3_X1    g2977(.A1(new_n3018_), .A2(new_n3019_), .A3(new_n2835_), .ZN(new_n3027_));
  NOR3_X1    g2978(.A1(new_n3027_), .A2(new_n3026_), .A3(new_n2805_), .ZN(new_n3028_));
  OAI22_X1   g2979(.A1(new_n3028_), .A2(new_n3025_), .B1(new_n3013_), .B2(new_n3015_), .ZN(new_n3029_));
  NAND2_X1   g2980(.A1(new_n2929_), .A2(new_n2891_), .ZN(new_n3030_));
  INV_X1     g2981(.I(new_n3030_), .ZN(new_n3031_));
  NOR2_X1    g2982(.A1(new_n2929_), .A2(new_n2891_), .ZN(new_n3032_));
  OAI21_X1   g2983(.A1(new_n3031_), .A2(new_n3032_), .B(new_n2890_), .ZN(new_n3033_));
  XOR2_X1    g2984(.A1(new_n2902_), .A2(new_n790_), .Z(new_n3034_));
  OAI21_X1   g2985(.A1(new_n2920_), .A2(new_n2925_), .B(new_n3034_), .ZN(new_n3035_));
  NAND3_X1   g2986(.A1(new_n3035_), .A2(new_n2893_), .A3(new_n2928_), .ZN(new_n3036_));
  NAND3_X1   g2987(.A1(new_n3036_), .A2(new_n3030_), .A3(new_n2889_), .ZN(new_n3037_));
  NAND2_X1   g2988(.A1(new_n3033_), .A2(new_n3037_), .ZN(new_n3038_));
  NAND2_X1   g2989(.A1(new_n3000_), .A2(new_n2629_), .ZN(new_n3039_));
  XOR2_X1    g2990(.A1(new_n2711_), .A2(new_n2696_), .Z(new_n3040_));
  OAI21_X1   g2991(.A1(new_n3040_), .A2(new_n2629_), .B(new_n3039_), .ZN(new_n3041_));
  AOI22_X1   g2992(.A1(new_n2708_), .A2(new_n3009_), .B1(new_n2697_), .B2(new_n2773_), .ZN(new_n3042_));
  INV_X1     g2993(.I(new_n3042_), .ZN(new_n3043_));
  NAND2_X1   g2994(.A1(new_n2628_), .A2(new_n2776_), .ZN(new_n3044_));
  AOI21_X1   g2995(.A1(new_n3044_), .A2(new_n3043_), .B(new_n2779_), .ZN(new_n3045_));
  NAND3_X1   g2996(.A1(new_n3041_), .A2(new_n1132_), .A3(new_n3045_), .ZN(new_n3046_));
  INV_X1     g2997(.I(new_n3039_), .ZN(new_n3047_));
  XOR2_X1    g2998(.A1(new_n2711_), .A2(new_n2708_), .Z(new_n3048_));
  AOI21_X1   g2999(.A1(new_n3048_), .A2(new_n2628_), .B(new_n3047_), .ZN(new_n3049_));
  INV_X1     g3000(.I(new_n3045_), .ZN(new_n3050_));
  OAI21_X1   g3001(.A1(new_n3049_), .A2(new_n3050_), .B(new_n1134_), .ZN(new_n3051_));
  AOI21_X1   g3002(.A1(new_n3051_), .A2(new_n3046_), .B(new_n3038_), .ZN(new_n3052_));
  OR2_X2     g3003(.A1(new_n2937_), .A2(new_n2936_), .Z(new_n3053_));
  OAI22_X1   g3004(.A1(new_n2637_), .A2(new_n2767_), .B1(new_n2663_), .B2(new_n2774_), .ZN(new_n3054_));
  NAND2_X1   g3005(.A1(new_n2708_), .A2(new_n2776_), .ZN(new_n3055_));
  AOI21_X1   g3006(.A1(new_n3055_), .A2(new_n3054_), .B(new_n2779_), .ZN(new_n3056_));
  NAND3_X1   g3007(.A1(new_n3053_), .A2(new_n1132_), .A3(new_n3056_), .ZN(new_n3057_));
  AOI21_X1   g3008(.A1(new_n3053_), .A2(new_n3056_), .B(new_n1132_), .ZN(new_n3058_));
  INV_X1     g3009(.I(new_n3058_), .ZN(new_n3059_));
  XOR2_X1    g3010(.A1(new_n2903_), .A2(new_n2904_), .Z(new_n3060_));
  XOR2_X1    g3011(.A1(new_n3034_), .A2(new_n2904_), .Z(new_n3061_));
  MUX2_X1    g3012(.I0(new_n3061_), .I1(new_n3060_), .S(new_n2919_), .Z(new_n3062_));
  NAND3_X1   g3013(.A1(new_n3062_), .A2(new_n3059_), .A3(new_n3057_), .ZN(new_n3063_));
  NAND3_X1   g3014(.A1(new_n2908_), .A2(new_n790_), .A3(new_n2921_), .ZN(new_n3064_));
  XOR2_X1    g3015(.A1(new_n2918_), .A2(new_n790_), .Z(new_n3065_));
  XOR2_X1    g3016(.A1(new_n3065_), .A2(new_n3064_), .Z(new_n3066_));
  OAI22_X1   g3017(.A1(new_n2663_), .A2(new_n2767_), .B1(new_n2691_), .B2(new_n2774_), .ZN(new_n3067_));
  NAND2_X1   g3018(.A1(new_n2697_), .A2(new_n2776_), .ZN(new_n3068_));
  AOI21_X1   g3019(.A1(new_n3068_), .A2(new_n3067_), .B(new_n2779_), .ZN(new_n3069_));
  AND3_X2    g3020(.A1(new_n2841_), .A2(new_n3069_), .A3(new_n1132_), .Z(new_n3070_));
  AOI21_X1   g3021(.A1(new_n2841_), .A2(new_n3069_), .B(new_n1132_), .ZN(new_n3071_));
  OAI21_X1   g3022(.A1(new_n3070_), .A2(new_n3071_), .B(new_n3066_), .ZN(new_n3072_));
  INV_X1     g3023(.I(new_n3072_), .ZN(new_n3073_));
  OAI22_X1   g3024(.A1(new_n2691_), .A2(new_n2767_), .B1(new_n2701_), .B2(new_n2774_), .ZN(new_n3074_));
  NAND2_X1   g3025(.A1(new_n2700_), .A2(new_n2776_), .ZN(new_n3075_));
  AOI21_X1   g3026(.A1(new_n3075_), .A2(new_n3074_), .B(new_n2779_), .ZN(new_n3076_));
  NAND2_X1   g3027(.A1(new_n2880_), .A2(new_n3076_), .ZN(new_n3077_));
  NOR2_X1    g3028(.A1(new_n3077_), .A2(new_n1134_), .ZN(new_n3078_));
  INV_X1     g3029(.I(new_n3078_), .ZN(new_n3079_));
  NAND2_X1   g3030(.A1(new_n3077_), .A2(new_n1134_), .ZN(new_n3080_));
  NOR2_X1    g3031(.A1(new_n2911_), .A2(new_n576_), .ZN(new_n3081_));
  XOR2_X1    g3032(.A1(new_n2910_), .A2(new_n3081_), .Z(new_n3082_));
  NAND3_X1   g3033(.A1(new_n3079_), .A2(new_n3080_), .A3(new_n3082_), .ZN(new_n3083_));
  OAI22_X1   g3034(.A1(new_n2701_), .A2(new_n2767_), .B1(new_n2673_), .B2(new_n2774_), .ZN(new_n3084_));
  OAI21_X1   g3035(.A1(new_n2691_), .A2(new_n3007_), .B(new_n3084_), .ZN(new_n3085_));
  NAND3_X1   g3036(.A1(new_n2899_), .A2(new_n2778_), .A3(new_n3085_), .ZN(new_n3086_));
  XOR2_X1    g3037(.A1(new_n3086_), .A2(new_n1134_), .Z(new_n3087_));
  XOR2_X1    g3038(.A1(new_n2672_), .A2(new_n2680_), .Z(new_n3088_));
  NAND2_X1   g3039(.A1(new_n2672_), .A2(new_n2776_), .ZN(new_n3089_));
  NAND2_X1   g3040(.A1(new_n2680_), .A2(new_n3009_), .ZN(new_n3090_));
  NAND4_X1   g3041(.A1(new_n3088_), .A2(new_n2778_), .A3(new_n3089_), .A4(new_n3090_), .ZN(new_n3091_));
  XOR2_X1    g3042(.A1(new_n3091_), .A2(new_n1134_), .Z(new_n3092_));
  NOR2_X1    g3043(.A1(new_n2788_), .A2(new_n2769_), .ZN(new_n3093_));
  INV_X1     g3044(.I(new_n3093_), .ZN(new_n3094_));
  AOI22_X1   g3045(.A1(new_n2672_), .A2(new_n3009_), .B1(new_n2680_), .B2(new_n2773_), .ZN(new_n3095_));
  AOI21_X1   g3046(.A1(new_n2668_), .A2(new_n2776_), .B(new_n3095_), .ZN(new_n3096_));
  NAND2_X1   g3047(.A1(new_n2914_), .A2(new_n2778_), .ZN(new_n3097_));
  NOR2_X1    g3048(.A1(new_n3097_), .A2(new_n3096_), .ZN(new_n3098_));
  NAND4_X1   g3049(.A1(new_n3098_), .A2(new_n3092_), .A3(new_n1132_), .A4(new_n3094_), .ZN(new_n3099_));
  XOR2_X1    g3050(.A1(new_n3099_), .A2(new_n2921_), .Z(new_n3100_));
  NOR2_X1    g3051(.A1(new_n3099_), .A2(new_n2921_), .ZN(new_n3101_));
  AOI21_X1   g3052(.A1(new_n3100_), .A2(new_n3087_), .B(new_n3101_), .ZN(new_n3102_));
  INV_X1     g3053(.I(new_n3102_), .ZN(new_n3103_));
  AOI21_X1   g3054(.A1(new_n3079_), .A2(new_n3080_), .B(new_n3082_), .ZN(new_n3104_));
  OAI21_X1   g3055(.A1(new_n3103_), .A2(new_n3104_), .B(new_n3083_), .ZN(new_n3105_));
  INV_X1     g3056(.I(new_n3066_), .ZN(new_n3106_));
  NOR2_X1    g3057(.A1(new_n3070_), .A2(new_n3071_), .ZN(new_n3107_));
  NAND2_X1   g3058(.A1(new_n3107_), .A2(new_n3106_), .ZN(new_n3108_));
  AOI21_X1   g3059(.A1(new_n3105_), .A2(new_n3108_), .B(new_n3073_), .ZN(new_n3109_));
  AOI21_X1   g3060(.A1(new_n3059_), .A2(new_n3057_), .B(new_n3062_), .ZN(new_n3110_));
  OAI21_X1   g3061(.A1(new_n3110_), .A2(new_n3109_), .B(new_n3063_), .ZN(new_n3111_));
  NAND3_X1   g3062(.A1(new_n3051_), .A2(new_n3038_), .A3(new_n3046_), .ZN(new_n3112_));
  AOI21_X1   g3063(.A1(new_n3111_), .A2(new_n3112_), .B(new_n3052_), .ZN(new_n3113_));
  NAND3_X1   g3064(.A1(new_n3014_), .A2(new_n1132_), .A3(new_n3011_), .ZN(new_n3114_));
  NAND2_X1   g3065(.A1(new_n3012_), .A2(new_n1134_), .ZN(new_n3115_));
  OAI21_X1   g3066(.A1(new_n3027_), .A2(new_n3026_), .B(new_n2805_), .ZN(new_n3116_));
  NAND3_X1   g3067(.A1(new_n3020_), .A2(new_n3024_), .A3(new_n3016_), .ZN(new_n3117_));
  NAND4_X1   g3068(.A1(new_n3116_), .A2(new_n3117_), .A3(new_n3114_), .A4(new_n3115_), .ZN(new_n3118_));
  NAND3_X1   g3069(.A1(new_n3029_), .A2(new_n3118_), .A3(new_n3113_), .ZN(new_n3119_));
  NAND4_X1   g3070(.A1(new_n2990_), .A2(new_n3119_), .A3(new_n2997_), .A4(new_n3029_), .ZN(new_n3120_));
  NOR3_X1    g3071(.A1(new_n2992_), .A2(new_n2991_), .A3(new_n2996_), .ZN(new_n3121_));
  AOI21_X1   g3072(.A1(new_n2781_), .A2(new_n2787_), .B(new_n2989_), .ZN(new_n3122_));
  INV_X1     g3073(.I(new_n3052_), .ZN(new_n3123_));
  NAND2_X1   g3074(.A1(new_n3111_), .A2(new_n3112_), .ZN(new_n3124_));
  NAND2_X1   g3075(.A1(new_n3124_), .A2(new_n3123_), .ZN(new_n3125_));
  NOR4_X1    g3076(.A1(new_n3028_), .A2(new_n3025_), .A3(new_n3013_), .A4(new_n3015_), .ZN(new_n3126_));
  OAI21_X1   g3077(.A1(new_n3125_), .A2(new_n3126_), .B(new_n3029_), .ZN(new_n3127_));
  OAI21_X1   g3078(.A1(new_n3121_), .A2(new_n3122_), .B(new_n3127_), .ZN(new_n3128_));
  NAND3_X1   g3079(.A1(new_n3128_), .A2(new_n3120_), .A3(new_n943_), .ZN(new_n3129_));
  NOR3_X1    g3080(.A1(new_n3127_), .A2(new_n3122_), .A3(new_n3121_), .ZN(new_n3130_));
  AOI22_X1   g3081(.A1(new_n2990_), .A2(new_n2997_), .B1(new_n3119_), .B2(new_n3029_), .ZN(new_n3131_));
  OAI21_X1   g3082(.A1(new_n3131_), .A2(new_n3130_), .B(new_n62_), .ZN(new_n3132_));
  AOI21_X1   g3083(.A1(new_n3129_), .A2(new_n3132_), .B(new_n2756_), .ZN(new_n3133_));
  NAND3_X1   g3084(.A1(new_n3129_), .A2(new_n3132_), .A3(new_n2756_), .ZN(new_n3134_));
  INV_X1     g3085(.I(new_n3134_), .ZN(new_n3135_));
  AOI22_X1   g3086(.A1(new_n3116_), .A2(new_n3117_), .B1(new_n3114_), .B2(new_n3115_), .ZN(new_n3136_));
  OAI21_X1   g3087(.A1(new_n3136_), .A2(new_n3126_), .B(new_n3125_), .ZN(new_n3137_));
  NAND2_X1   g3088(.A1(new_n2716_), .A2(new_n2718_), .ZN(new_n3138_));
  NAND3_X1   g3089(.A1(new_n2555_), .A2(new_n2557_), .A3(new_n2576_), .ZN(new_n3139_));
  AOI21_X1   g3090(.A1(new_n2555_), .A2(new_n2557_), .B(new_n2576_), .ZN(new_n3140_));
  INV_X1     g3091(.I(new_n3140_), .ZN(new_n3141_));
  NAND2_X1   g3092(.A1(new_n3141_), .A2(new_n3139_), .ZN(new_n3142_));
  NOR2_X1    g3093(.A1(new_n3138_), .A2(new_n3142_), .ZN(new_n3143_));
  INV_X1     g3094(.I(new_n3139_), .ZN(new_n3144_));
  NOR2_X1    g3095(.A1(new_n3144_), .A2(new_n3140_), .ZN(new_n3145_));
  AOI21_X1   g3096(.A1(new_n2716_), .A2(new_n2718_), .B(new_n3145_), .ZN(new_n3146_));
  OAI22_X1   g3097(.A1(new_n2576_), .A2(new_n2752_), .B1(new_n2593_), .B2(new_n2742_), .ZN(new_n3147_));
  NAND2_X1   g3098(.A1(new_n2559_), .A2(new_n2748_), .ZN(new_n3148_));
  AOI21_X1   g3099(.A1(new_n3148_), .A2(new_n3147_), .B(new_n72_), .ZN(new_n3149_));
  OAI21_X1   g3100(.A1(new_n3146_), .A2(new_n3143_), .B(new_n3149_), .ZN(new_n3150_));
  XOR2_X1    g3101(.A1(new_n3150_), .A2(new_n62_), .Z(new_n3151_));
  NAND3_X1   g3102(.A1(new_n3151_), .A2(new_n3119_), .A3(new_n3137_), .ZN(new_n3152_));
  NAND2_X1   g3103(.A1(new_n3137_), .A2(new_n3119_), .ZN(new_n3153_));
  XOR2_X1    g3104(.A1(new_n3150_), .A2(new_n943_), .Z(new_n3154_));
  NAND2_X1   g3105(.A1(new_n3153_), .A2(new_n3154_), .ZN(new_n3155_));
  NAND2_X1   g3106(.A1(new_n3155_), .A2(new_n3152_), .ZN(new_n3156_));
  INV_X1     g3107(.I(new_n3057_), .ZN(new_n3157_));
  XOR2_X1    g3108(.A1(new_n3034_), .A2(new_n2904_), .Z(new_n3158_));
  NOR2_X1    g3109(.A1(new_n3158_), .A2(new_n2924_), .ZN(new_n3159_));
  XOR2_X1    g3110(.A1(new_n2903_), .A2(new_n2904_), .Z(new_n3160_));
  NOR2_X1    g3111(.A1(new_n3160_), .A2(new_n2919_), .ZN(new_n3161_));
  NOR2_X1    g3112(.A1(new_n3159_), .A2(new_n3161_), .ZN(new_n3162_));
  OAI21_X1   g3113(.A1(new_n3157_), .A2(new_n3058_), .B(new_n3162_), .ZN(new_n3163_));
  AOI21_X1   g3114(.A1(new_n3163_), .A2(new_n3063_), .B(new_n3109_), .ZN(new_n3164_));
  INV_X1     g3115(.I(new_n3083_), .ZN(new_n3165_));
  INV_X1     g3116(.I(new_n3104_), .ZN(new_n3166_));
  AOI21_X1   g3117(.A1(new_n3102_), .A2(new_n3166_), .B(new_n3165_), .ZN(new_n3167_));
  INV_X1     g3118(.I(new_n3108_), .ZN(new_n3168_));
  OAI21_X1   g3119(.A1(new_n3168_), .A2(new_n3167_), .B(new_n3072_), .ZN(new_n3169_));
  OAI21_X1   g3120(.A1(new_n3157_), .A2(new_n3058_), .B(new_n3062_), .ZN(new_n3170_));
  NAND3_X1   g3121(.A1(new_n3162_), .A2(new_n3057_), .A3(new_n3059_), .ZN(new_n3171_));
  AOI21_X1   g3122(.A1(new_n3170_), .A2(new_n3171_), .B(new_n3169_), .ZN(new_n3172_));
  NOR2_X1    g3123(.A1(new_n3172_), .A2(new_n3164_), .ZN(new_n3173_));
  OAI22_X1   g3124(.A1(new_n2619_), .A2(new_n2752_), .B1(new_n2629_), .B2(new_n2742_), .ZN(new_n3174_));
  NAND2_X1   g3125(.A1(new_n2586_), .A2(new_n2748_), .ZN(new_n3175_));
  AOI21_X1   g3126(.A1(new_n3174_), .A2(new_n3175_), .B(new_n72_), .ZN(new_n3176_));
  OAI21_X1   g3127(.A1(new_n2784_), .A2(new_n2785_), .B(new_n3176_), .ZN(new_n3177_));
  NOR2_X1    g3128(.A1(new_n3177_), .A2(new_n943_), .ZN(new_n3178_));
  AOI21_X1   g3129(.A1(new_n2764_), .A2(new_n3176_), .B(new_n62_), .ZN(new_n3179_));
  OAI21_X1   g3130(.A1(new_n3179_), .A2(new_n3178_), .B(new_n3173_), .ZN(new_n3180_));
  INV_X1     g3131(.I(new_n3063_), .ZN(new_n3181_));
  OAI21_X1   g3132(.A1(new_n3181_), .A2(new_n3110_), .B(new_n3169_), .ZN(new_n3182_));
  AOI21_X1   g3133(.A1(new_n3059_), .A2(new_n3057_), .B(new_n3162_), .ZN(new_n3183_));
  NOR3_X1    g3134(.A1(new_n3062_), .A2(new_n3157_), .A3(new_n3058_), .ZN(new_n3184_));
  OAI21_X1   g3135(.A1(new_n3183_), .A2(new_n3184_), .B(new_n3109_), .ZN(new_n3185_));
  NAND2_X1   g3136(.A1(new_n3182_), .A2(new_n3185_), .ZN(new_n3186_));
  NAND3_X1   g3137(.A1(new_n2764_), .A2(new_n62_), .A3(new_n3176_), .ZN(new_n3187_));
  NAND2_X1   g3138(.A1(new_n3177_), .A2(new_n943_), .ZN(new_n3188_));
  NAND3_X1   g3139(.A1(new_n3186_), .A2(new_n3187_), .A3(new_n3188_), .ZN(new_n3189_));
  NAND2_X1   g3140(.A1(new_n3108_), .A2(new_n3072_), .ZN(new_n3190_));
  OAI21_X1   g3141(.A1(new_n3070_), .A2(new_n3071_), .B(new_n3106_), .ZN(new_n3191_));
  NAND2_X1   g3142(.A1(new_n3107_), .A2(new_n3066_), .ZN(new_n3192_));
  AOI21_X1   g3143(.A1(new_n3191_), .A2(new_n3192_), .B(new_n3105_), .ZN(new_n3193_));
  AOI21_X1   g3144(.A1(new_n3190_), .A2(new_n3105_), .B(new_n3193_), .ZN(new_n3194_));
  OAI22_X1   g3145(.A1(new_n2619_), .A2(new_n2747_), .B1(new_n2696_), .B2(new_n2742_), .ZN(new_n3195_));
  NAND2_X1   g3146(.A1(new_n2628_), .A2(new_n2753_), .ZN(new_n3196_));
  AOI21_X1   g3147(.A1(new_n3195_), .A2(new_n3196_), .B(new_n72_), .ZN(new_n3197_));
  NAND3_X1   g3148(.A1(new_n3014_), .A2(new_n62_), .A3(new_n3197_), .ZN(new_n3198_));
  INV_X1     g3149(.I(new_n3198_), .ZN(new_n3199_));
  AOI21_X1   g3150(.A1(new_n3014_), .A2(new_n3197_), .B(new_n62_), .ZN(new_n3200_));
  OAI21_X1   g3151(.A1(new_n3199_), .A2(new_n3200_), .B(new_n3194_), .ZN(new_n3201_));
  NOR3_X1    g3152(.A1(new_n3199_), .A2(new_n3194_), .A3(new_n3200_), .ZN(new_n3202_));
  NAND2_X1   g3153(.A1(new_n3079_), .A2(new_n3080_), .ZN(new_n3203_));
  NOR2_X1    g3154(.A1(new_n3203_), .A2(new_n3082_), .ZN(new_n3204_));
  INV_X1     g3155(.I(new_n3080_), .ZN(new_n3205_));
  NOR2_X1    g3156(.A1(new_n3205_), .A2(new_n3078_), .ZN(new_n3206_));
  INV_X1     g3157(.I(new_n3082_), .ZN(new_n3207_));
  NOR2_X1    g3158(.A1(new_n3206_), .A2(new_n3207_), .ZN(new_n3208_));
  OAI21_X1   g3159(.A1(new_n3204_), .A2(new_n3208_), .B(new_n3103_), .ZN(new_n3209_));
  NAND2_X1   g3160(.A1(new_n3206_), .A2(new_n3207_), .ZN(new_n3210_));
  NAND2_X1   g3161(.A1(new_n3203_), .A2(new_n3082_), .ZN(new_n3211_));
  NAND3_X1   g3162(.A1(new_n3210_), .A2(new_n3211_), .A3(new_n3102_), .ZN(new_n3212_));
  NAND2_X1   g3163(.A1(new_n3209_), .A2(new_n3212_), .ZN(new_n3213_));
  OAI22_X1   g3164(.A1(new_n2637_), .A2(new_n2752_), .B1(new_n2663_), .B2(new_n2742_), .ZN(new_n3214_));
  NAND2_X1   g3165(.A1(new_n2708_), .A2(new_n2748_), .ZN(new_n3215_));
  AOI21_X1   g3166(.A1(new_n3215_), .A2(new_n3214_), .B(new_n72_), .ZN(new_n3216_));
  OAI21_X1   g3167(.A1(new_n2937_), .A2(new_n2936_), .B(new_n3216_), .ZN(new_n3217_));
  NOR2_X1    g3168(.A1(new_n3217_), .A2(new_n943_), .ZN(new_n3218_));
  INV_X1     g3169(.I(new_n3218_), .ZN(new_n3219_));
  NAND2_X1   g3170(.A1(new_n3217_), .A2(new_n943_), .ZN(new_n3220_));
  XOR2_X1    g3171(.A1(new_n3086_), .A2(new_n1132_), .Z(new_n3221_));
  NAND2_X1   g3172(.A1(new_n3221_), .A2(new_n2911_), .ZN(new_n3222_));
  NAND2_X1   g3173(.A1(new_n3087_), .A2(new_n2921_), .ZN(new_n3223_));
  AND2_X2    g3174(.A1(new_n3222_), .A2(new_n3223_), .Z(new_n3224_));
  NOR2_X1    g3175(.A1(new_n3221_), .A2(new_n2921_), .ZN(new_n3225_));
  NOR2_X1    g3176(.A1(new_n3087_), .A2(new_n2911_), .ZN(new_n3226_));
  OAI21_X1   g3177(.A1(new_n3226_), .A2(new_n3225_), .B(new_n3099_), .ZN(new_n3227_));
  OAI21_X1   g3178(.A1(new_n3224_), .A2(new_n3099_), .B(new_n3227_), .ZN(new_n3228_));
  NAND3_X1   g3179(.A1(new_n3228_), .A2(new_n3219_), .A3(new_n3220_), .ZN(new_n3229_));
  NOR2_X1    g3180(.A1(new_n3093_), .A2(new_n1134_), .ZN(new_n3230_));
  NAND2_X1   g3181(.A1(new_n3092_), .A2(new_n3230_), .ZN(new_n3231_));
  NAND2_X1   g3182(.A1(new_n3098_), .A2(new_n1132_), .ZN(new_n3232_));
  INV_X1     g3183(.I(new_n3232_), .ZN(new_n3233_));
  NOR2_X1    g3184(.A1(new_n3098_), .A2(new_n1132_), .ZN(new_n3234_));
  OAI21_X1   g3185(.A1(new_n3233_), .A2(new_n3234_), .B(new_n3231_), .ZN(new_n3235_));
  INV_X1     g3186(.I(new_n3231_), .ZN(new_n3236_));
  INV_X1     g3187(.I(new_n3234_), .ZN(new_n3237_));
  NAND3_X1   g3188(.A1(new_n3237_), .A2(new_n3236_), .A3(new_n3232_), .ZN(new_n3238_));
  NAND2_X1   g3189(.A1(new_n3235_), .A2(new_n3238_), .ZN(new_n3239_));
  AOI22_X1   g3190(.A1(new_n2700_), .A2(new_n2753_), .B1(new_n2844_), .B2(new_n2741_), .ZN(new_n3240_));
  NOR2_X1    g3191(.A1(new_n2637_), .A2(new_n2747_), .ZN(new_n3241_));
  OAI21_X1   g3192(.A1(new_n3241_), .A2(new_n3240_), .B(new_n71_), .ZN(new_n3242_));
  INV_X1     g3193(.I(new_n3242_), .ZN(new_n3243_));
  NAND3_X1   g3194(.A1(new_n3243_), .A2(new_n2841_), .A3(new_n62_), .ZN(new_n3244_));
  OAI21_X1   g3195(.A1(new_n2864_), .A2(new_n3242_), .B(new_n943_), .ZN(new_n3245_));
  NAND3_X1   g3196(.A1(new_n3239_), .A2(new_n3245_), .A3(new_n3244_), .ZN(new_n3246_));
  AOI21_X1   g3197(.A1(new_n3237_), .A2(new_n3232_), .B(new_n3236_), .ZN(new_n3247_));
  NOR3_X1    g3198(.A1(new_n3233_), .A2(new_n3231_), .A3(new_n3234_), .ZN(new_n3248_));
  NOR2_X1    g3199(.A1(new_n3247_), .A2(new_n3248_), .ZN(new_n3249_));
  INV_X1     g3200(.I(new_n3244_), .ZN(new_n3250_));
  AOI21_X1   g3201(.A1(new_n3243_), .A2(new_n2841_), .B(new_n62_), .ZN(new_n3251_));
  OAI21_X1   g3202(.A1(new_n3250_), .A2(new_n3251_), .B(new_n3249_), .ZN(new_n3252_));
  XNOR2_X1   g3203(.A1(new_n3092_), .A2(new_n3230_), .ZN(new_n3253_));
  NOR2_X1    g3204(.A1(new_n2673_), .A2(new_n2747_), .ZN(new_n3254_));
  NOR2_X1    g3205(.A1(new_n2788_), .A2(new_n2752_), .ZN(new_n3255_));
  NOR4_X1    g3206(.A1(new_n2789_), .A2(new_n72_), .A3(new_n3254_), .A4(new_n3255_), .ZN(new_n3256_));
  XOR2_X1    g3207(.A1(new_n3256_), .A2(new_n943_), .Z(new_n3257_));
  NOR2_X1    g3208(.A1(new_n2788_), .A2(new_n70_), .ZN(new_n3258_));
  NOR2_X1    g3209(.A1(new_n3258_), .A2(new_n943_), .ZN(new_n3259_));
  AOI22_X1   g3210(.A1(new_n2672_), .A2(new_n2753_), .B1(new_n2680_), .B2(new_n2741_), .ZN(new_n3260_));
  NOR2_X1    g3211(.A1(new_n2701_), .A2(new_n2747_), .ZN(new_n3261_));
  NOR2_X1    g3212(.A1(new_n3261_), .A2(new_n3260_), .ZN(new_n3262_));
  INV_X1     g3213(.I(new_n3262_), .ZN(new_n3263_));
  NAND4_X1   g3214(.A1(new_n3263_), .A2(new_n2914_), .A3(new_n62_), .A4(new_n71_), .ZN(new_n3264_));
  OAI21_X1   g3215(.A1(new_n2822_), .A2(new_n2819_), .B(new_n71_), .ZN(new_n3265_));
  OAI21_X1   g3216(.A1(new_n3265_), .A2(new_n3262_), .B(new_n943_), .ZN(new_n3266_));
  NAND2_X1   g3217(.A1(new_n3264_), .A2(new_n3266_), .ZN(new_n3267_));
  NAND4_X1   g3218(.A1(new_n3267_), .A2(new_n3093_), .A3(new_n3257_), .A4(new_n3259_), .ZN(new_n3268_));
  AOI22_X1   g3219(.A1(new_n2668_), .A2(new_n2753_), .B1(new_n2672_), .B2(new_n2741_), .ZN(new_n3269_));
  NOR2_X1    g3220(.A1(new_n2691_), .A2(new_n2747_), .ZN(new_n3270_));
  OAI21_X1   g3221(.A1(new_n3270_), .A2(new_n3269_), .B(new_n71_), .ZN(new_n3271_));
  NOR2_X1    g3222(.A1(new_n2958_), .A2(new_n3271_), .ZN(new_n3272_));
  XOR2_X1    g3223(.A1(new_n3272_), .A2(new_n943_), .Z(new_n3273_));
  INV_X1     g3224(.I(new_n3258_), .ZN(new_n3274_));
  NOR2_X1    g3225(.A1(new_n3265_), .A2(new_n3262_), .ZN(new_n3275_));
  NAND4_X1   g3226(.A1(new_n3275_), .A2(new_n62_), .A3(new_n3256_), .A4(new_n3274_), .ZN(new_n3276_));
  AND4_X2    g3227(.A1(new_n62_), .A2(new_n3256_), .A3(new_n3093_), .A4(new_n3274_), .Z(new_n3277_));
  AOI22_X1   g3228(.A1(new_n3267_), .A2(new_n3277_), .B1(new_n3276_), .B2(new_n3094_), .ZN(new_n3278_));
  NAND2_X1   g3229(.A1(new_n3273_), .A2(new_n3278_), .ZN(new_n3279_));
  NAND3_X1   g3230(.A1(new_n3279_), .A2(new_n3253_), .A3(new_n3268_), .ZN(new_n3280_));
  OAI22_X1   g3231(.A1(new_n2691_), .A2(new_n2752_), .B1(new_n2701_), .B2(new_n2742_), .ZN(new_n3281_));
  NAND2_X1   g3232(.A1(new_n2700_), .A2(new_n2748_), .ZN(new_n3282_));
  AOI21_X1   g3233(.A1(new_n3282_), .A2(new_n3281_), .B(new_n72_), .ZN(new_n3283_));
  NAND2_X1   g3234(.A1(new_n2880_), .A2(new_n3283_), .ZN(new_n3284_));
  XOR2_X1    g3235(.A1(new_n3284_), .A2(new_n62_), .Z(new_n3285_));
  AOI21_X1   g3236(.A1(new_n3279_), .A2(new_n3268_), .B(new_n3253_), .ZN(new_n3286_));
  OAI21_X1   g3237(.A1(new_n3285_), .A2(new_n3286_), .B(new_n3280_), .ZN(new_n3287_));
  AOI22_X1   g3238(.A1(new_n3239_), .A2(new_n3287_), .B1(new_n3252_), .B2(new_n3246_), .ZN(new_n3288_));
  NAND2_X1   g3239(.A1(new_n3219_), .A2(new_n3220_), .ZN(new_n3289_));
  AOI21_X1   g3240(.A1(new_n3223_), .A2(new_n3222_), .B(new_n3099_), .ZN(new_n3290_));
  OR2_X2     g3241(.A1(new_n3225_), .A2(new_n3226_), .Z(new_n3291_));
  AOI21_X1   g3242(.A1(new_n3291_), .A2(new_n3099_), .B(new_n3290_), .ZN(new_n3292_));
  NAND2_X1   g3243(.A1(new_n3289_), .A2(new_n3292_), .ZN(new_n3293_));
  NAND2_X1   g3244(.A1(new_n3293_), .A2(new_n3288_), .ZN(new_n3294_));
  NAND3_X1   g3245(.A1(new_n3294_), .A2(new_n3213_), .A3(new_n3229_), .ZN(new_n3295_));
  INV_X1     g3246(.I(new_n3213_), .ZN(new_n3296_));
  NAND2_X1   g3247(.A1(new_n3252_), .A2(new_n3246_), .ZN(new_n3297_));
  AOI21_X1   g3248(.A1(new_n3245_), .A2(new_n3244_), .B(new_n3239_), .ZN(new_n3298_));
  INV_X1     g3249(.I(new_n3287_), .ZN(new_n3299_));
  AOI21_X1   g3250(.A1(new_n3297_), .A2(new_n3299_), .B(new_n3298_), .ZN(new_n3300_));
  AOI21_X1   g3251(.A1(new_n3219_), .A2(new_n3220_), .B(new_n3228_), .ZN(new_n3301_));
  OAI21_X1   g3252(.A1(new_n3300_), .A2(new_n3301_), .B(new_n3229_), .ZN(new_n3302_));
  NAND2_X1   g3253(.A1(new_n3302_), .A2(new_n3296_), .ZN(new_n3303_));
  AOI22_X1   g3254(.A1(new_n2708_), .A2(new_n2753_), .B1(new_n2697_), .B2(new_n2741_), .ZN(new_n3304_));
  INV_X1     g3255(.I(new_n3304_), .ZN(new_n3305_));
  NAND2_X1   g3256(.A1(new_n2628_), .A2(new_n2748_), .ZN(new_n3306_));
  AOI21_X1   g3257(.A1(new_n3306_), .A2(new_n3305_), .B(new_n72_), .ZN(new_n3307_));
  NAND3_X1   g3258(.A1(new_n3041_), .A2(new_n62_), .A3(new_n3307_), .ZN(new_n3308_));
  NAND2_X1   g3259(.A1(new_n3041_), .A2(new_n3307_), .ZN(new_n3309_));
  NAND2_X1   g3260(.A1(new_n3309_), .A2(new_n943_), .ZN(new_n3310_));
  NAND2_X1   g3261(.A1(new_n3310_), .A2(new_n3308_), .ZN(new_n3311_));
  AOI22_X1   g3262(.A1(new_n3303_), .A2(new_n3295_), .B1(new_n3213_), .B2(new_n3311_), .ZN(new_n3312_));
  OAI21_X1   g3263(.A1(new_n3312_), .A2(new_n3202_), .B(new_n3201_), .ZN(new_n3313_));
  NAND3_X1   g3264(.A1(new_n3313_), .A2(new_n3180_), .A3(new_n3189_), .ZN(new_n3314_));
  NOR2_X1    g3265(.A1(new_n2715_), .A2(new_n2593_), .ZN(new_n3315_));
  NOR2_X1    g3266(.A1(new_n2730_), .A2(new_n2586_), .ZN(new_n3316_));
  NOR2_X1    g3267(.A1(new_n3316_), .A2(new_n3315_), .ZN(new_n3317_));
  NOR3_X1    g3268(.A1(new_n3317_), .A2(new_n2763_), .A3(new_n2577_), .ZN(new_n3318_));
  NAND2_X1   g3269(.A1(new_n2730_), .A2(new_n2586_), .ZN(new_n3319_));
  NAND2_X1   g3270(.A1(new_n2715_), .A2(new_n2593_), .ZN(new_n3320_));
  NAND2_X1   g3271(.A1(new_n3319_), .A2(new_n3320_), .ZN(new_n3321_));
  AOI21_X1   g3272(.A1(new_n3321_), .A2(new_n2762_), .B(new_n2576_), .ZN(new_n3322_));
  OAI22_X1   g3273(.A1(new_n2576_), .A2(new_n2747_), .B1(new_n2619_), .B2(new_n2742_), .ZN(new_n3323_));
  NAND2_X1   g3274(.A1(new_n2586_), .A2(new_n2753_), .ZN(new_n3324_));
  AOI21_X1   g3275(.A1(new_n3323_), .A2(new_n3324_), .B(new_n72_), .ZN(new_n3325_));
  OAI21_X1   g3276(.A1(new_n3318_), .A2(new_n3322_), .B(new_n3325_), .ZN(new_n3326_));
  NOR2_X1    g3277(.A1(new_n3326_), .A2(new_n943_), .ZN(new_n3327_));
  NAND3_X1   g3278(.A1(new_n3321_), .A2(new_n2576_), .A3(new_n2762_), .ZN(new_n3328_));
  OAI21_X1   g3279(.A1(new_n3317_), .A2(new_n2763_), .B(new_n2577_), .ZN(new_n3329_));
  NAND2_X1   g3280(.A1(new_n3329_), .A2(new_n3328_), .ZN(new_n3330_));
  AOI21_X1   g3281(.A1(new_n3330_), .A2(new_n3325_), .B(new_n62_), .ZN(new_n3331_));
  NOR2_X1    g3282(.A1(new_n3327_), .A2(new_n3331_), .ZN(new_n3332_));
  NAND2_X1   g3283(.A1(new_n3314_), .A2(new_n3332_), .ZN(new_n3333_));
  AOI21_X1   g3284(.A1(new_n3187_), .A2(new_n3188_), .B(new_n3186_), .ZN(new_n3334_));
  NOR3_X1    g3285(.A1(new_n3173_), .A2(new_n3179_), .A3(new_n3178_), .ZN(new_n3335_));
  NAND2_X1   g3286(.A1(new_n3190_), .A2(new_n3105_), .ZN(new_n3336_));
  NAND2_X1   g3287(.A1(new_n3191_), .A2(new_n3192_), .ZN(new_n3337_));
  NAND2_X1   g3288(.A1(new_n3337_), .A2(new_n3167_), .ZN(new_n3338_));
  NAND2_X1   g3289(.A1(new_n3338_), .A2(new_n3336_), .ZN(new_n3339_));
  INV_X1     g3290(.I(new_n3200_), .ZN(new_n3340_));
  AOI21_X1   g3291(.A1(new_n3340_), .A2(new_n3198_), .B(new_n3339_), .ZN(new_n3341_));
  NAND3_X1   g3292(.A1(new_n3340_), .A2(new_n3339_), .A3(new_n3198_), .ZN(new_n3342_));
  NOR2_X1    g3293(.A1(new_n3302_), .A2(new_n3296_), .ZN(new_n3343_));
  AOI21_X1   g3294(.A1(new_n3294_), .A2(new_n3229_), .B(new_n3213_), .ZN(new_n3344_));
  INV_X1     g3295(.I(new_n3311_), .ZN(new_n3345_));
  OAI22_X1   g3296(.A1(new_n3343_), .A2(new_n3344_), .B1(new_n3345_), .B2(new_n3296_), .ZN(new_n3346_));
  AOI21_X1   g3297(.A1(new_n3346_), .A2(new_n3342_), .B(new_n3341_), .ZN(new_n3347_));
  NOR3_X1    g3298(.A1(new_n3347_), .A2(new_n3334_), .A3(new_n3335_), .ZN(new_n3348_));
  XOR2_X1    g3299(.A1(new_n3326_), .A2(new_n62_), .Z(new_n3349_));
  NAND2_X1   g3300(.A1(new_n3348_), .A2(new_n3349_), .ZN(new_n3350_));
  NAND2_X1   g3301(.A1(new_n3123_), .A2(new_n3112_), .ZN(new_n3351_));
  NAND2_X1   g3302(.A1(new_n3051_), .A2(new_n3046_), .ZN(new_n3352_));
  XOR2_X1    g3303(.A1(new_n3352_), .A2(new_n3038_), .Z(new_n3353_));
  NOR2_X1    g3304(.A1(new_n3353_), .A2(new_n3111_), .ZN(new_n3354_));
  AOI21_X1   g3305(.A1(new_n3111_), .A2(new_n3351_), .B(new_n3354_), .ZN(new_n3355_));
  INV_X1     g3306(.I(new_n3355_), .ZN(new_n3356_));
  AOI22_X1   g3307(.A1(new_n3350_), .A2(new_n3333_), .B1(new_n3314_), .B2(new_n3356_), .ZN(new_n3357_));
  OAI21_X1   g3308(.A1(new_n3357_), .A2(new_n3156_), .B(new_n3152_), .ZN(new_n3358_));
  NOR3_X1    g3309(.A1(new_n3358_), .A2(new_n3133_), .A3(new_n3135_), .ZN(new_n3359_));
  NOR2_X1    g3310(.A1(new_n3135_), .A2(new_n3133_), .ZN(new_n3360_));
  NOR2_X1    g3311(.A1(new_n3153_), .A2(new_n3154_), .ZN(new_n3361_));
  AOI21_X1   g3312(.A1(new_n3119_), .A2(new_n3137_), .B(new_n3151_), .ZN(new_n3362_));
  NOR2_X1    g3313(.A1(new_n3362_), .A2(new_n3361_), .ZN(new_n3363_));
  NOR2_X1    g3314(.A1(new_n3348_), .A2(new_n3349_), .ZN(new_n3364_));
  NOR4_X1    g3315(.A1(new_n3332_), .A2(new_n3334_), .A3(new_n3335_), .A4(new_n3347_), .ZN(new_n3365_));
  OAI22_X1   g3316(.A1(new_n3364_), .A2(new_n3365_), .B1(new_n3355_), .B2(new_n3348_), .ZN(new_n3366_));
  AOI21_X1   g3317(.A1(new_n3366_), .A2(new_n3363_), .B(new_n3361_), .ZN(new_n3367_));
  NOR2_X1    g3318(.A1(new_n3360_), .A2(new_n3367_), .ZN(new_n3368_));
  NOR2_X1    g3319(.A1(new_n3368_), .A2(new_n3359_), .ZN(new_n3369_));
  INV_X1     g3320(.I(new_n3369_), .ZN(new_n3370_));
  NOR4_X1    g3321(.A1(new_n563_), .A2(new_n387_), .A3(new_n620_), .A4(new_n865_), .ZN(new_n3371_));
  NOR2_X1    g3322(.A1(new_n198_), .A2(new_n553_), .ZN(new_n3372_));
  INV_X1     g3323(.I(new_n3372_), .ZN(new_n3373_));
  NOR3_X1    g3324(.A1(new_n3373_), .A2(new_n369_), .A3(new_n642_), .ZN(new_n3374_));
  NAND3_X1   g3325(.A1(new_n769_), .A2(new_n309_), .A3(new_n549_), .ZN(new_n3375_));
  NOR3_X1    g3326(.A1(new_n3374_), .A2(new_n3371_), .A3(new_n3375_), .ZN(new_n3376_));
  NOR2_X1    g3327(.A1(new_n825_), .A2(new_n402_), .ZN(new_n3377_));
  NAND4_X1   g3328(.A1(new_n3377_), .A2(new_n371_), .A3(new_n550_), .A4(new_n950_), .ZN(new_n3378_));
  NOR4_X1    g3329(.A1(new_n3378_), .A2(new_n209_), .A3(new_n1647_), .A4(new_n1706_), .ZN(new_n3379_));
  AND2_X2    g3330(.A1(new_n3376_), .A2(new_n3379_), .Z(new_n3380_));
  INV_X1     g3331(.I(new_n2422_), .ZN(new_n3381_));
  INV_X1     g3332(.I(new_n319_), .ZN(new_n3382_));
  NOR3_X1    g3333(.A1(new_n3382_), .A2(new_n266_), .A3(new_n890_), .ZN(new_n3383_));
  NAND4_X1   g3334(.A1(new_n418_), .A2(new_n475_), .A3(new_n481_), .A4(new_n458_), .ZN(new_n3384_));
  NAND4_X1   g3335(.A1(new_n2545_), .A2(new_n223_), .A3(new_n363_), .A4(new_n556_), .ZN(new_n3385_));
  NAND3_X1   g3336(.A1(new_n3385_), .A2(new_n3383_), .A3(new_n3384_), .ZN(new_n3386_));
  NOR4_X1    g3337(.A1(new_n3386_), .A2(new_n257_), .A3(new_n713_), .A4(new_n3381_), .ZN(new_n3387_));
  NAND3_X1   g3338(.A1(new_n3380_), .A2(new_n737_), .A3(new_n3387_), .ZN(new_n3388_));
  NOR2_X1    g3339(.A1(new_n3388_), .A2(new_n2549_), .ZN(new_n3389_));
  INV_X1     g3340(.I(new_n3389_), .ZN(new_n3390_));
  INV_X1     g3341(.I(new_n405_), .ZN(new_n3391_));
  NAND4_X1   g3342(.A1(new_n719_), .A2(new_n720_), .A3(new_n837_), .A4(new_n1019_), .ZN(new_n3392_));
  INV_X1     g3343(.I(new_n764_), .ZN(new_n3393_));
  NOR2_X1    g3344(.A1(new_n2376_), .A2(new_n324_), .ZN(new_n3394_));
  NAND4_X1   g3345(.A1(new_n1077_), .A2(new_n3394_), .A3(new_n3393_), .A4(new_n2380_), .ZN(new_n3395_));
  INV_X1     g3346(.I(new_n3395_), .ZN(new_n3396_));
  NAND4_X1   g3347(.A1(new_n3396_), .A2(new_n1640_), .A3(new_n1704_), .A4(new_n3392_), .ZN(new_n3397_));
  NOR3_X1    g3348(.A1(new_n3397_), .A2(new_n606_), .A3(new_n3391_), .ZN(new_n3398_));
  INV_X1     g3349(.I(new_n3398_), .ZN(new_n3399_));
  NOR2_X1    g3350(.A1(new_n3390_), .A2(new_n3399_), .ZN(new_n3400_));
  NAND2_X1   g3351(.A1(new_n2541_), .A2(new_n3400_), .ZN(new_n3401_));
  INV_X1     g3352(.I(new_n649_), .ZN(new_n3402_));
  INV_X1     g3353(.I(new_n624_), .ZN(new_n3403_));
  NOR2_X1    g3354(.A1(new_n589_), .A2(new_n267_), .ZN(new_n3404_));
  INV_X1     g3355(.I(new_n3404_), .ZN(new_n3405_));
  NOR3_X1    g3356(.A1(new_n3405_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n3406_));
  NOR3_X1    g3357(.A1(new_n282_), .A2(new_n975_), .A3(new_n2314_), .ZN(new_n3407_));
  NAND4_X1   g3358(.A1(new_n3403_), .A2(new_n373_), .A3(new_n3406_), .A4(new_n3407_), .ZN(new_n3408_));
  INV_X1     g3359(.I(new_n3408_), .ZN(new_n3409_));
  NAND4_X1   g3360(.A1(new_n3409_), .A2(new_n600_), .A3(new_n405_), .A4(new_n3402_), .ZN(new_n3410_));
  NAND2_X1   g3361(.A1(new_n3401_), .A2(new_n3410_), .ZN(new_n3411_));
  NOR2_X1    g3362(.A1(new_n3401_), .A2(new_n3410_), .ZN(new_n3412_));
  INV_X1     g3363(.I(new_n3412_), .ZN(new_n3413_));
  NAND2_X1   g3364(.A1(new_n3413_), .A2(new_n3411_), .ZN(new_n3414_));
  INV_X1     g3365(.I(new_n2541_), .ZN(new_n3415_));
  INV_X1     g3366(.I(new_n3388_), .ZN(new_n3416_));
  NOR2_X1    g3367(.A1(new_n3415_), .A2(new_n2549_), .ZN(new_n3417_));
  OAI22_X1   g3368(.A1(new_n3417_), .A2(new_n3416_), .B1(new_n3415_), .B2(new_n3390_), .ZN(new_n3418_));
  INV_X1     g3369(.I(new_n3418_), .ZN(new_n3419_));
  OAI21_X1   g3370(.A1(new_n2721_), .A2(new_n3418_), .B(new_n2551_), .ZN(new_n3420_));
  NAND2_X1   g3371(.A1(new_n2720_), .A2(new_n2558_), .ZN(new_n3421_));
  AOI21_X1   g3372(.A1(new_n3421_), .A2(new_n2733_), .B(new_n3418_), .ZN(new_n3422_));
  AOI21_X1   g3373(.A1(new_n3422_), .A2(new_n2745_), .B(new_n2558_), .ZN(new_n3423_));
  AOI21_X1   g3374(.A1(new_n2735_), .A2(new_n3419_), .B(new_n2551_), .ZN(new_n3424_));
  AOI21_X1   g3375(.A1(new_n3423_), .A2(new_n3420_), .B(new_n3424_), .ZN(new_n3425_));
  NAND2_X1   g3376(.A1(new_n3425_), .A2(new_n3419_), .ZN(new_n3426_));
  AOI21_X1   g3377(.A1(new_n2735_), .A2(new_n3419_), .B(new_n2745_), .ZN(new_n3427_));
  NOR2_X1    g3378(.A1(new_n2734_), .A2(new_n2559_), .ZN(new_n3428_));
  OAI21_X1   g3379(.A1(new_n3428_), .A2(new_n2719_), .B(new_n3419_), .ZN(new_n3429_));
  OAI21_X1   g3380(.A1(new_n3429_), .A2(new_n2551_), .B(new_n2559_), .ZN(new_n3430_));
  NAND2_X1   g3381(.A1(new_n3429_), .A2(new_n2745_), .ZN(new_n3431_));
  OAI21_X1   g3382(.A1(new_n3430_), .A2(new_n3427_), .B(new_n3431_), .ZN(new_n3432_));
  NAND2_X1   g3383(.A1(new_n3432_), .A2(new_n3418_), .ZN(new_n3433_));
  NAND3_X1   g3384(.A1(new_n3417_), .A2(new_n3416_), .A3(new_n3399_), .ZN(new_n3434_));
  NAND2_X1   g3385(.A1(new_n3417_), .A2(new_n3416_), .ZN(new_n3435_));
  NAND2_X1   g3386(.A1(new_n3435_), .A2(new_n3398_), .ZN(new_n3436_));
  AOI21_X1   g3387(.A1(new_n3436_), .A2(new_n3434_), .B(new_n3418_), .ZN(new_n3437_));
  NAND3_X1   g3388(.A1(new_n3436_), .A2(new_n3418_), .A3(new_n3434_), .ZN(new_n3438_));
  INV_X1     g3389(.I(new_n3438_), .ZN(new_n3439_));
  NOR2_X1    g3390(.A1(new_n3439_), .A2(new_n3437_), .ZN(new_n3440_));
  INV_X1     g3391(.I(new_n3440_), .ZN(new_n3441_));
  NAND3_X1   g3392(.A1(new_n3433_), .A2(new_n3426_), .A3(new_n3441_), .ZN(new_n3442_));
  NOR2_X1    g3393(.A1(new_n3442_), .A2(new_n3414_), .ZN(new_n3443_));
  INV_X1     g3394(.I(new_n3414_), .ZN(new_n3444_));
  OAI21_X1   g3395(.A1(new_n3425_), .A2(new_n3419_), .B(new_n3441_), .ZN(new_n3445_));
  AOI21_X1   g3396(.A1(new_n3419_), .A2(new_n3425_), .B(new_n3445_), .ZN(new_n3446_));
  NOR2_X1    g3397(.A1(new_n3446_), .A2(new_n3444_), .ZN(new_n3447_));
  NOR2_X1    g3398(.A1(new_n3447_), .A2(new_n3443_), .ZN(new_n3448_));
  NAND2_X1   g3399(.A1(new_n3436_), .A2(new_n3434_), .ZN(new_n3449_));
  NOR2_X1    g3400(.A1(new_n65_), .A2(\a[2] ), .ZN(new_n3450_));
  INV_X1     g3401(.I(new_n3450_), .ZN(new_n3451_));
  INV_X1     g3402(.I(\a[0] ), .ZN(new_n3452_));
  NAND2_X1   g3403(.A1(new_n3452_), .A2(\a[1] ), .ZN(new_n3453_));
  OAI22_X1   g3404(.A1(new_n3449_), .A2(new_n3453_), .B1(new_n3419_), .B2(new_n3451_), .ZN(new_n3454_));
  XNOR2_X1   g3405(.A1(\a[1] ), .A2(\a[2] ), .ZN(new_n3455_));
  NOR2_X1    g3406(.A1(new_n3455_), .A2(\a[0] ), .ZN(new_n3456_));
  INV_X1     g3407(.I(new_n3456_), .ZN(new_n3457_));
  OAI21_X1   g3408(.A1(new_n3444_), .A2(new_n3457_), .B(new_n3454_), .ZN(new_n3458_));
  NOR2_X1    g3409(.A1(new_n3455_), .A2(new_n3452_), .ZN(new_n3459_));
  NAND2_X1   g3410(.A1(new_n3458_), .A2(new_n3459_), .ZN(new_n3460_));
  NOR3_X1    g3411(.A1(new_n3448_), .A2(new_n2739_), .A3(new_n3460_), .ZN(new_n3461_));
  NAND2_X1   g3412(.A1(new_n3446_), .A2(new_n3444_), .ZN(new_n3462_));
  NAND2_X1   g3413(.A1(new_n3442_), .A2(new_n3414_), .ZN(new_n3463_));
  NAND2_X1   g3414(.A1(new_n3462_), .A2(new_n3463_), .ZN(new_n3464_));
  INV_X1     g3415(.I(new_n3460_), .ZN(new_n3465_));
  AOI21_X1   g3416(.A1(new_n3464_), .A2(new_n3465_), .B(new_n69_), .ZN(new_n3466_));
  NOR2_X1    g3417(.A1(new_n3461_), .A2(new_n3466_), .ZN(new_n3467_));
  INV_X1     g3418(.I(new_n3467_), .ZN(new_n3468_));
  NOR2_X1    g3419(.A1(new_n2735_), .A2(new_n2745_), .ZN(new_n3469_));
  NOR2_X1    g3420(.A1(new_n2721_), .A2(new_n2551_), .ZN(new_n3470_));
  OAI21_X1   g3421(.A1(new_n3469_), .A2(new_n3470_), .B(new_n2723_), .ZN(new_n3471_));
  XOR2_X1    g3422(.A1(new_n3471_), .A2(new_n3419_), .Z(new_n3472_));
  INV_X1     g3423(.I(new_n3459_), .ZN(new_n3473_));
  OAI22_X1   g3424(.A1(new_n2551_), .A2(new_n3453_), .B1(new_n2558_), .B2(new_n3451_), .ZN(new_n3474_));
  NAND2_X1   g3425(.A1(new_n3418_), .A2(new_n3456_), .ZN(new_n3475_));
  AOI21_X1   g3426(.A1(new_n3475_), .A2(new_n3474_), .B(new_n3473_), .ZN(new_n3476_));
  NAND3_X1   g3427(.A1(new_n3472_), .A2(new_n69_), .A3(new_n3476_), .ZN(new_n3477_));
  AOI21_X1   g3428(.A1(new_n3472_), .A2(new_n3476_), .B(new_n69_), .ZN(new_n3478_));
  INV_X1     g3429(.I(new_n3478_), .ZN(new_n3479_));
  OAI21_X1   g3430(.A1(new_n3364_), .A2(new_n3365_), .B(new_n3355_), .ZN(new_n3480_));
  NAND3_X1   g3431(.A1(new_n3350_), .A2(new_n3333_), .A3(new_n3356_), .ZN(new_n3481_));
  NAND2_X1   g3432(.A1(new_n3481_), .A2(new_n3480_), .ZN(new_n3482_));
  NAND3_X1   g3433(.A1(new_n3482_), .A2(new_n3479_), .A3(new_n3477_), .ZN(new_n3483_));
  NAND3_X1   g3434(.A1(new_n3145_), .A2(new_n2716_), .A3(new_n2718_), .ZN(new_n3484_));
  NAND2_X1   g3435(.A1(new_n3138_), .A2(new_n3142_), .ZN(new_n3485_));
  AOI21_X1   g3436(.A1(new_n3485_), .A2(new_n3484_), .B(new_n3473_), .ZN(new_n3486_));
  INV_X1     g3437(.I(new_n3453_), .ZN(new_n3487_));
  AOI22_X1   g3438(.A1(new_n2577_), .A2(new_n3487_), .B1(new_n2586_), .B2(new_n3450_), .ZN(new_n3488_));
  AOI21_X1   g3439(.A1(new_n2559_), .A2(new_n3456_), .B(new_n3488_), .ZN(new_n3489_));
  INV_X1     g3440(.I(new_n3489_), .ZN(new_n3490_));
  OAI21_X1   g3441(.A1(new_n3486_), .A2(new_n3490_), .B(new_n2739_), .ZN(new_n3491_));
  OAI21_X1   g3442(.A1(new_n3146_), .A2(new_n3143_), .B(new_n3459_), .ZN(new_n3492_));
  NAND3_X1   g3443(.A1(new_n3492_), .A2(new_n69_), .A3(new_n3489_), .ZN(new_n3493_));
  NAND2_X1   g3444(.A1(new_n3493_), .A2(new_n3491_), .ZN(new_n3494_));
  NAND3_X1   g3445(.A1(new_n3312_), .A2(new_n3201_), .A3(new_n3342_), .ZN(new_n3495_));
  INV_X1     g3446(.I(new_n3495_), .ZN(new_n3496_));
  AOI21_X1   g3447(.A1(new_n3201_), .A2(new_n3342_), .B(new_n3312_), .ZN(new_n3497_));
  NOR2_X1    g3448(.A1(new_n3496_), .A2(new_n3497_), .ZN(new_n3498_));
  NOR2_X1    g3449(.A1(new_n3498_), .A2(new_n3494_), .ZN(new_n3499_));
  AOI21_X1   g3450(.A1(new_n3293_), .A2(new_n3229_), .B(new_n3288_), .ZN(new_n3500_));
  AND3_X2    g3451(.A1(new_n3293_), .A2(new_n3229_), .A3(new_n3288_), .Z(new_n3501_));
  NOR2_X1    g3452(.A1(new_n3501_), .A2(new_n3500_), .ZN(new_n3502_));
  INV_X1     g3453(.I(new_n3502_), .ZN(new_n3503_));
  OAI22_X1   g3454(.A1(new_n2619_), .A2(new_n3453_), .B1(new_n2629_), .B2(new_n3451_), .ZN(new_n3504_));
  NAND2_X1   g3455(.A1(new_n2586_), .A2(new_n3456_), .ZN(new_n3505_));
  AOI21_X1   g3456(.A1(new_n3504_), .A2(new_n3505_), .B(new_n3473_), .ZN(new_n3506_));
  NAND3_X1   g3457(.A1(new_n2764_), .A2(new_n69_), .A3(new_n3506_), .ZN(new_n3507_));
  AOI21_X1   g3458(.A1(new_n2764_), .A2(new_n3506_), .B(new_n69_), .ZN(new_n3508_));
  INV_X1     g3459(.I(new_n3508_), .ZN(new_n3509_));
  NAND3_X1   g3460(.A1(new_n3509_), .A2(new_n3503_), .A3(new_n3507_), .ZN(new_n3510_));
  INV_X1     g3461(.I(new_n3507_), .ZN(new_n3511_));
  OAI21_X1   g3462(.A1(new_n3511_), .A2(new_n3508_), .B(new_n3502_), .ZN(new_n3512_));
  AOI21_X1   g3463(.A1(new_n2708_), .A2(new_n3450_), .B(new_n3473_), .ZN(new_n3513_));
  OAI21_X1   g3464(.A1(new_n2629_), .A2(new_n3453_), .B(new_n3513_), .ZN(new_n3514_));
  AOI21_X1   g3465(.A1(new_n2621_), .A2(new_n3456_), .B(new_n3514_), .ZN(new_n3515_));
  AND3_X2    g3466(.A1(new_n3014_), .A2(new_n69_), .A3(new_n3515_), .Z(new_n3516_));
  AOI21_X1   g3467(.A1(new_n3014_), .A2(new_n3515_), .B(new_n69_), .ZN(new_n3517_));
  NOR2_X1    g3468(.A1(new_n3516_), .A2(new_n3517_), .ZN(new_n3518_));
  NOR2_X1    g3469(.A1(new_n3233_), .A2(new_n3234_), .ZN(new_n3519_));
  INV_X1     g3470(.I(new_n3519_), .ZN(new_n3520_));
  NOR2_X1    g3471(.A1(new_n3250_), .A2(new_n3251_), .ZN(new_n3521_));
  NOR2_X1    g3472(.A1(new_n3287_), .A2(new_n3521_), .ZN(new_n3522_));
  INV_X1     g3473(.I(new_n3522_), .ZN(new_n3523_));
  NAND2_X1   g3474(.A1(new_n3287_), .A2(new_n3521_), .ZN(new_n3524_));
  AOI21_X1   g3475(.A1(new_n3523_), .A2(new_n3524_), .B(new_n3520_), .ZN(new_n3525_));
  INV_X1     g3476(.I(new_n3525_), .ZN(new_n3526_));
  NAND3_X1   g3477(.A1(new_n3523_), .A2(new_n3520_), .A3(new_n3524_), .ZN(new_n3527_));
  AOI21_X1   g3478(.A1(new_n3526_), .A2(new_n3527_), .B(new_n3236_), .ZN(new_n3528_));
  INV_X1     g3479(.I(new_n3528_), .ZN(new_n3529_));
  NAND3_X1   g3480(.A1(new_n3526_), .A2(new_n3236_), .A3(new_n3527_), .ZN(new_n3530_));
  NAND3_X1   g3481(.A1(new_n3529_), .A2(new_n3518_), .A3(new_n3530_), .ZN(new_n3531_));
  XOR2_X1    g3482(.A1(new_n3273_), .A2(new_n3278_), .Z(new_n3532_));
  NAND2_X1   g3483(.A1(new_n2878_), .A2(new_n2663_), .ZN(new_n3533_));
  NAND2_X1   g3484(.A1(new_n2874_), .A2(new_n2700_), .ZN(new_n3534_));
  NAND2_X1   g3485(.A1(new_n3533_), .A2(new_n3534_), .ZN(new_n3535_));
  NAND2_X1   g3486(.A1(new_n2817_), .A2(new_n2818_), .ZN(new_n3536_));
  XOR2_X1    g3487(.A1(new_n2404_), .A2(new_n2686_), .Z(new_n3537_));
  AOI22_X1   g3488(.A1(new_n3537_), .A2(new_n3453_), .B1(new_n3536_), .B2(new_n3451_), .ZN(new_n3538_));
  NOR2_X1    g3489(.A1(new_n2663_), .A2(new_n3457_), .ZN(new_n3539_));
  OAI21_X1   g3490(.A1(new_n3539_), .A2(new_n3538_), .B(new_n3459_), .ZN(new_n3540_));
  OR2_X2     g3491(.A1(new_n3535_), .A2(new_n3540_), .Z(new_n3541_));
  NOR2_X1    g3492(.A1(new_n3541_), .A2(new_n2739_), .ZN(new_n3542_));
  NOR2_X1    g3493(.A1(new_n3535_), .A2(new_n3540_), .ZN(new_n3543_));
  NOR2_X1    g3494(.A1(new_n3543_), .A2(new_n69_), .ZN(new_n3544_));
  XNOR2_X1   g3495(.A1(new_n3257_), .A2(new_n3259_), .ZN(new_n3545_));
  INV_X1     g3496(.I(new_n3545_), .ZN(new_n3546_));
  NOR3_X1    g3497(.A1(new_n3542_), .A2(new_n3544_), .A3(new_n3546_), .ZN(new_n3547_));
  NAND2_X1   g3498(.A1(new_n2672_), .A2(new_n3487_), .ZN(new_n3548_));
  NAND2_X1   g3499(.A1(new_n2680_), .A2(new_n3450_), .ZN(new_n3549_));
  NAND4_X1   g3500(.A1(new_n2668_), .A2(new_n3456_), .A3(new_n3548_), .A4(new_n3549_), .ZN(new_n3550_));
  OAI21_X1   g3501(.A1(\a[0] ), .A2(\a[1] ), .B(new_n2680_), .ZN(new_n3551_));
  AOI22_X1   g3502(.A1(new_n2672_), .A2(new_n3456_), .B1(new_n69_), .B2(new_n3551_), .ZN(new_n3552_));
  NOR4_X1    g3503(.A1(new_n3088_), .A2(new_n2739_), .A3(new_n3459_), .A4(new_n3552_), .ZN(new_n3553_));
  NAND3_X1   g3504(.A1(new_n2823_), .A2(new_n3550_), .A3(new_n3553_), .ZN(new_n3554_));
  NOR2_X1    g3505(.A1(new_n2869_), .A2(new_n2870_), .ZN(new_n3555_));
  XOR2_X1    g3506(.A1(new_n3555_), .A2(new_n2701_), .Z(new_n3556_));
  NOR2_X1    g3507(.A1(new_n3556_), .A2(new_n3473_), .ZN(new_n3557_));
  AOI22_X1   g3508(.A1(new_n2668_), .A2(new_n3487_), .B1(new_n2672_), .B2(new_n3450_), .ZN(new_n3558_));
  NOR2_X1    g3509(.A1(new_n2691_), .A2(new_n3457_), .ZN(new_n3559_));
  NOR2_X1    g3510(.A1(new_n3559_), .A2(new_n3558_), .ZN(new_n3560_));
  INV_X1     g3511(.I(new_n3560_), .ZN(new_n3561_));
  NOR3_X1    g3512(.A1(new_n3557_), .A2(new_n2739_), .A3(new_n3561_), .ZN(new_n3562_));
  INV_X1     g3513(.I(new_n3562_), .ZN(new_n3563_));
  OAI21_X1   g3514(.A1(new_n3557_), .A2(new_n3561_), .B(new_n2739_), .ZN(new_n3564_));
  AOI22_X1   g3515(.A1(new_n3563_), .A2(new_n3564_), .B1(new_n3274_), .B2(new_n3554_), .ZN(new_n3565_));
  OAI21_X1   g3516(.A1(new_n3542_), .A2(new_n3544_), .B(new_n3546_), .ZN(new_n3566_));
  NOR2_X1    g3517(.A1(new_n3554_), .A2(new_n3274_), .ZN(new_n3567_));
  INV_X1     g3518(.I(new_n3567_), .ZN(new_n3568_));
  NAND2_X1   g3519(.A1(new_n3566_), .A2(new_n3568_), .ZN(new_n3569_));
  NOR2_X1    g3520(.A1(new_n3569_), .A2(new_n3565_), .ZN(new_n3570_));
  OAI22_X1   g3521(.A1(new_n2663_), .A2(new_n3453_), .B1(new_n2691_), .B2(new_n3451_), .ZN(new_n3571_));
  NAND2_X1   g3522(.A1(new_n2697_), .A2(new_n3456_), .ZN(new_n3572_));
  AOI21_X1   g3523(.A1(new_n3572_), .A2(new_n3571_), .B(new_n3473_), .ZN(new_n3573_));
  NAND3_X1   g3524(.A1(new_n2841_), .A2(new_n3573_), .A3(new_n69_), .ZN(new_n3574_));
  AOI21_X1   g3525(.A1(new_n2841_), .A2(new_n3573_), .B(new_n69_), .ZN(new_n3575_));
  INV_X1     g3526(.I(new_n3575_), .ZN(new_n3576_));
  NAND2_X1   g3527(.A1(new_n3576_), .A2(new_n3574_), .ZN(new_n3577_));
  INV_X1     g3528(.I(new_n3577_), .ZN(new_n3578_));
  NOR3_X1    g3529(.A1(new_n3570_), .A2(new_n3547_), .A3(new_n3578_), .ZN(new_n3579_));
  INV_X1     g3530(.I(new_n3547_), .ZN(new_n3580_));
  INV_X1     g3531(.I(new_n3554_), .ZN(new_n3581_));
  INV_X1     g3532(.I(new_n3564_), .ZN(new_n3582_));
  OAI22_X1   g3533(.A1(new_n3582_), .A2(new_n3562_), .B1(new_n3258_), .B2(new_n3581_), .ZN(new_n3583_));
  NAND3_X1   g3534(.A1(new_n3583_), .A2(new_n3566_), .A3(new_n3568_), .ZN(new_n3584_));
  INV_X1     g3535(.I(new_n3574_), .ZN(new_n3585_));
  NAND2_X1   g3536(.A1(new_n3257_), .A2(new_n3259_), .ZN(new_n3586_));
  XOR2_X1    g3537(.A1(new_n3586_), .A2(new_n3267_), .Z(new_n3587_));
  OR3_X2     g3538(.A1(new_n3585_), .A2(new_n3575_), .A3(new_n3587_), .Z(new_n3588_));
  AOI21_X1   g3539(.A1(new_n3584_), .A2(new_n3580_), .B(new_n3588_), .ZN(new_n3589_));
  NOR3_X1    g3540(.A1(new_n3579_), .A2(new_n3589_), .A3(new_n3532_), .ZN(new_n3590_));
  INV_X1     g3541(.I(new_n3532_), .ZN(new_n3591_));
  NAND3_X1   g3542(.A1(new_n3584_), .A2(new_n3580_), .A3(new_n3577_), .ZN(new_n3592_));
  NOR2_X1    g3543(.A1(new_n3577_), .A2(new_n3587_), .ZN(new_n3593_));
  OAI21_X1   g3544(.A1(new_n3570_), .A2(new_n3547_), .B(new_n3593_), .ZN(new_n3594_));
  AOI21_X1   g3545(.A1(new_n3594_), .A2(new_n3592_), .B(new_n3591_), .ZN(new_n3595_));
  OAI22_X1   g3546(.A1(new_n2637_), .A2(new_n3453_), .B1(new_n2663_), .B2(new_n3451_), .ZN(new_n3596_));
  NAND2_X1   g3547(.A1(new_n2708_), .A2(new_n3456_), .ZN(new_n3597_));
  AOI21_X1   g3548(.A1(new_n3597_), .A2(new_n3596_), .B(new_n3473_), .ZN(new_n3598_));
  NAND2_X1   g3549(.A1(new_n3053_), .A2(new_n3598_), .ZN(new_n3599_));
  XOR2_X1    g3550(.A1(new_n3599_), .A2(new_n2739_), .Z(new_n3600_));
  OAI22_X1   g3551(.A1(new_n3590_), .A2(new_n3595_), .B1(new_n3532_), .B2(new_n3600_), .ZN(new_n3601_));
  OAI22_X1   g3552(.A1(new_n2637_), .A2(new_n3451_), .B1(new_n2696_), .B2(new_n3453_), .ZN(new_n3602_));
  NAND2_X1   g3553(.A1(new_n2628_), .A2(new_n3456_), .ZN(new_n3603_));
  AOI21_X1   g3554(.A1(new_n3603_), .A2(new_n3602_), .B(new_n3473_), .ZN(new_n3604_));
  NAND2_X1   g3555(.A1(new_n3041_), .A2(new_n3604_), .ZN(new_n3605_));
  XOR2_X1    g3556(.A1(new_n3605_), .A2(new_n2739_), .Z(new_n3606_));
  NOR2_X1    g3557(.A1(new_n3601_), .A2(new_n3606_), .ZN(new_n3607_));
  NAND2_X1   g3558(.A1(new_n3279_), .A2(new_n3268_), .ZN(new_n3608_));
  XOR2_X1    g3559(.A1(new_n3285_), .A2(new_n3253_), .Z(new_n3609_));
  XNOR2_X1   g3560(.A1(new_n3609_), .A2(new_n3608_), .ZN(new_n3610_));
  AOI21_X1   g3561(.A1(new_n3601_), .A2(new_n3606_), .B(new_n3610_), .ZN(new_n3611_));
  NOR2_X1    g3562(.A1(new_n3611_), .A2(new_n3607_), .ZN(new_n3612_));
  AOI21_X1   g3563(.A1(new_n3529_), .A2(new_n3530_), .B(new_n3518_), .ZN(new_n3613_));
  OAI21_X1   g3564(.A1(new_n3612_), .A2(new_n3613_), .B(new_n3531_), .ZN(new_n3614_));
  AOI22_X1   g3565(.A1(new_n3614_), .A2(new_n3503_), .B1(new_n3510_), .B2(new_n3512_), .ZN(new_n3615_));
  OAI22_X1   g3566(.A1(new_n2576_), .A2(new_n3457_), .B1(new_n2619_), .B2(new_n3451_), .ZN(new_n3616_));
  NAND2_X1   g3567(.A1(new_n2586_), .A2(new_n3487_), .ZN(new_n3617_));
  AOI21_X1   g3568(.A1(new_n3616_), .A2(new_n3617_), .B(new_n3473_), .ZN(new_n3618_));
  NAND3_X1   g3569(.A1(new_n3330_), .A2(new_n69_), .A3(new_n3618_), .ZN(new_n3619_));
  AOI21_X1   g3570(.A1(new_n3330_), .A2(new_n3618_), .B(new_n69_), .ZN(new_n3620_));
  INV_X1     g3571(.I(new_n3620_), .ZN(new_n3621_));
  NOR2_X1    g3572(.A1(new_n3208_), .A2(new_n3204_), .ZN(new_n3622_));
  INV_X1     g3573(.I(new_n3622_), .ZN(new_n3623_));
  NAND3_X1   g3574(.A1(new_n3311_), .A2(new_n3294_), .A3(new_n3229_), .ZN(new_n3624_));
  NAND2_X1   g3575(.A1(new_n3345_), .A2(new_n3302_), .ZN(new_n3625_));
  AOI21_X1   g3576(.A1(new_n3625_), .A2(new_n3624_), .B(new_n3623_), .ZN(new_n3626_));
  INV_X1     g3577(.I(new_n3624_), .ZN(new_n3627_));
  AOI21_X1   g3578(.A1(new_n3229_), .A2(new_n3294_), .B(new_n3311_), .ZN(new_n3628_));
  NOR3_X1    g3579(.A1(new_n3627_), .A2(new_n3628_), .A3(new_n3622_), .ZN(new_n3629_));
  OAI21_X1   g3580(.A1(new_n3629_), .A2(new_n3626_), .B(new_n3103_), .ZN(new_n3630_));
  OAI21_X1   g3581(.A1(new_n3627_), .A2(new_n3628_), .B(new_n3622_), .ZN(new_n3631_));
  NAND3_X1   g3582(.A1(new_n3625_), .A2(new_n3623_), .A3(new_n3624_), .ZN(new_n3632_));
  NAND3_X1   g3583(.A1(new_n3631_), .A2(new_n3632_), .A3(new_n3102_), .ZN(new_n3633_));
  AOI22_X1   g3584(.A1(new_n3630_), .A2(new_n3633_), .B1(new_n3621_), .B2(new_n3619_), .ZN(new_n3634_));
  INV_X1     g3585(.I(new_n3634_), .ZN(new_n3635_));
  NAND2_X1   g3586(.A1(new_n3635_), .A2(new_n3615_), .ZN(new_n3636_));
  OAI21_X1   g3587(.A1(new_n3341_), .A2(new_n3202_), .B(new_n3346_), .ZN(new_n3637_));
  NAND3_X1   g3588(.A1(new_n3494_), .A2(new_n3637_), .A3(new_n3495_), .ZN(new_n3638_));
  AND2_X2    g3589(.A1(new_n3493_), .A2(new_n3491_), .Z(new_n3639_));
  NAND2_X1   g3590(.A1(new_n3637_), .A2(new_n3495_), .ZN(new_n3640_));
  NAND2_X1   g3591(.A1(new_n3639_), .A2(new_n3640_), .ZN(new_n3641_));
  INV_X1     g3592(.I(new_n3619_), .ZN(new_n3642_));
  AOI21_X1   g3593(.A1(new_n3631_), .A2(new_n3632_), .B(new_n3102_), .ZN(new_n3643_));
  NOR3_X1    g3594(.A1(new_n3629_), .A2(new_n3626_), .A3(new_n3103_), .ZN(new_n3644_));
  NOR4_X1    g3595(.A1(new_n3644_), .A2(new_n3643_), .A3(new_n3642_), .A4(new_n3620_), .ZN(new_n3645_));
  AOI21_X1   g3596(.A1(new_n3641_), .A2(new_n3638_), .B(new_n3645_), .ZN(new_n3646_));
  AOI21_X1   g3597(.A1(new_n3636_), .A2(new_n3646_), .B(new_n3499_), .ZN(new_n3647_));
  NAND3_X1   g3598(.A1(new_n3347_), .A2(new_n3180_), .A3(new_n3189_), .ZN(new_n3648_));
  OAI21_X1   g3599(.A1(new_n3334_), .A2(new_n3335_), .B(new_n3313_), .ZN(new_n3649_));
  NAND2_X1   g3600(.A1(new_n3649_), .A2(new_n3648_), .ZN(new_n3650_));
  INV_X1     g3601(.I(new_n3650_), .ZN(new_n3651_));
  NOR2_X1    g3602(.A1(new_n3647_), .A2(new_n3651_), .ZN(new_n3652_));
  NAND2_X1   g3603(.A1(new_n2736_), .A2(new_n2722_), .ZN(new_n3653_));
  NAND2_X1   g3604(.A1(new_n2559_), .A2(new_n3487_), .ZN(new_n3654_));
  NAND2_X1   g3605(.A1(new_n2745_), .A2(new_n3456_), .ZN(new_n3655_));
  AOI21_X1   g3606(.A1(new_n2577_), .A2(new_n3450_), .B(new_n3473_), .ZN(new_n3656_));
  NAND4_X1   g3607(.A1(new_n3653_), .A2(new_n3654_), .A3(new_n3655_), .A4(new_n3656_), .ZN(new_n3657_));
  XOR2_X1    g3608(.A1(new_n3657_), .A2(new_n2739_), .Z(new_n3658_));
  AOI21_X1   g3609(.A1(new_n3647_), .A2(new_n3651_), .B(new_n3658_), .ZN(new_n3659_));
  NOR3_X1    g3610(.A1(new_n3659_), .A2(new_n3652_), .A3(new_n3483_), .ZN(new_n3660_));
  NOR2_X1    g3611(.A1(new_n3366_), .A2(new_n3156_), .ZN(new_n3661_));
  NOR2_X1    g3612(.A1(new_n3357_), .A2(new_n3363_), .ZN(new_n3662_));
  NOR2_X1    g3613(.A1(new_n3662_), .A2(new_n3661_), .ZN(new_n3663_));
  XOR2_X1    g3614(.A1(new_n3449_), .A2(new_n3418_), .Z(new_n3664_));
  NOR2_X1    g3615(.A1(new_n3432_), .A2(new_n3664_), .ZN(new_n3665_));
  NOR2_X1    g3616(.A1(new_n3425_), .A2(new_n3440_), .ZN(new_n3666_));
  OAI21_X1   g3617(.A1(new_n3665_), .A2(new_n3666_), .B(new_n3459_), .ZN(new_n3667_));
  INV_X1     g3618(.I(new_n3449_), .ZN(new_n3668_));
  NAND2_X1   g3619(.A1(new_n3418_), .A2(new_n3487_), .ZN(new_n3669_));
  NAND2_X1   g3620(.A1(new_n2745_), .A2(new_n3450_), .ZN(new_n3670_));
  AOI22_X1   g3621(.A1(new_n3668_), .A2(new_n3456_), .B1(new_n3669_), .B2(new_n3670_), .ZN(new_n3671_));
  NAND2_X1   g3622(.A1(new_n3667_), .A2(new_n3671_), .ZN(new_n3672_));
  NOR2_X1    g3623(.A1(new_n3672_), .A2(new_n2739_), .ZN(new_n3673_));
  AOI21_X1   g3624(.A1(new_n3667_), .A2(new_n3671_), .B(new_n69_), .ZN(new_n3674_));
  NOR2_X1    g3625(.A1(new_n3673_), .A2(new_n3674_), .ZN(new_n3675_));
  OAI21_X1   g3626(.A1(new_n3675_), .A2(new_n3663_), .B(new_n3483_), .ZN(new_n3676_));
  NOR2_X1    g3627(.A1(new_n3660_), .A2(new_n3676_), .ZN(new_n3677_));
  INV_X1     g3628(.I(new_n3672_), .ZN(new_n3678_));
  NAND2_X1   g3629(.A1(new_n3357_), .A2(new_n3363_), .ZN(new_n3679_));
  NAND2_X1   g3630(.A1(new_n3366_), .A2(new_n3156_), .ZN(new_n3680_));
  AOI21_X1   g3631(.A1(new_n3679_), .A2(new_n3680_), .B(new_n2739_), .ZN(new_n3681_));
  NOR3_X1    g3632(.A1(new_n3662_), .A2(new_n3661_), .A3(new_n69_), .ZN(new_n3682_));
  OAI21_X1   g3633(.A1(new_n3682_), .A2(new_n3681_), .B(new_n3678_), .ZN(new_n3683_));
  OAI21_X1   g3634(.A1(new_n3662_), .A2(new_n3661_), .B(new_n69_), .ZN(new_n3684_));
  NAND3_X1   g3635(.A1(new_n3679_), .A2(new_n3680_), .A3(new_n2739_), .ZN(new_n3685_));
  NAND3_X1   g3636(.A1(new_n3684_), .A2(new_n3685_), .A3(new_n3672_), .ZN(new_n3686_));
  NAND2_X1   g3637(.A1(new_n3683_), .A2(new_n3686_), .ZN(new_n3687_));
  INV_X1     g3638(.I(new_n3687_), .ZN(new_n3688_));
  AOI21_X1   g3639(.A1(new_n3688_), .A2(new_n3677_), .B(new_n3468_), .ZN(new_n3689_));
  INV_X1     g3640(.I(new_n3477_), .ZN(new_n3690_));
  AND2_X2    g3641(.A1(new_n3481_), .A2(new_n3480_), .Z(new_n3691_));
  NOR3_X1    g3642(.A1(new_n3691_), .A2(new_n3690_), .A3(new_n3478_), .ZN(new_n3692_));
  INV_X1     g3643(.I(new_n3499_), .ZN(new_n3693_));
  NAND2_X1   g3644(.A1(new_n3510_), .A2(new_n3512_), .ZN(new_n3694_));
  NAND2_X1   g3645(.A1(new_n3694_), .A2(new_n3502_), .ZN(new_n3695_));
  NAND3_X1   g3646(.A1(new_n3594_), .A2(new_n3592_), .A3(new_n3591_), .ZN(new_n3696_));
  OAI21_X1   g3647(.A1(new_n3579_), .A2(new_n3589_), .B(new_n3532_), .ZN(new_n3697_));
  INV_X1     g3648(.I(new_n3600_), .ZN(new_n3698_));
  AOI22_X1   g3649(.A1(new_n3697_), .A2(new_n3696_), .B1(new_n3591_), .B2(new_n3698_), .ZN(new_n3699_));
  INV_X1     g3650(.I(new_n3606_), .ZN(new_n3700_));
  NAND2_X1   g3651(.A1(new_n3699_), .A2(new_n3700_), .ZN(new_n3701_));
  INV_X1     g3652(.I(new_n3610_), .ZN(new_n3702_));
  OAI21_X1   g3653(.A1(new_n3699_), .A2(new_n3700_), .B(new_n3702_), .ZN(new_n3703_));
  NAND2_X1   g3654(.A1(new_n3703_), .A2(new_n3701_), .ZN(new_n3704_));
  AND3_X2    g3655(.A1(new_n3526_), .A2(new_n3236_), .A3(new_n3527_), .Z(new_n3705_));
  OAI22_X1   g3656(.A1(new_n3705_), .A2(new_n3528_), .B1(new_n3516_), .B2(new_n3517_), .ZN(new_n3706_));
  NAND2_X1   g3657(.A1(new_n3704_), .A2(new_n3706_), .ZN(new_n3707_));
  NAND3_X1   g3658(.A1(new_n3694_), .A2(new_n3707_), .A3(new_n3531_), .ZN(new_n3708_));
  AOI21_X1   g3659(.A1(new_n3708_), .A2(new_n3695_), .B(new_n3634_), .ZN(new_n3709_));
  INV_X1     g3660(.I(new_n3638_), .ZN(new_n3710_));
  NOR2_X1    g3661(.A1(new_n3498_), .A2(new_n3494_), .ZN(new_n3711_));
  NAND4_X1   g3662(.A1(new_n3630_), .A2(new_n3633_), .A3(new_n3621_), .A4(new_n3619_), .ZN(new_n3712_));
  OAI21_X1   g3663(.A1(new_n3711_), .A2(new_n3710_), .B(new_n3712_), .ZN(new_n3713_));
  OAI21_X1   g3664(.A1(new_n3713_), .A2(new_n3709_), .B(new_n3693_), .ZN(new_n3714_));
  NAND2_X1   g3665(.A1(new_n3714_), .A2(new_n3650_), .ZN(new_n3715_));
  INV_X1     g3666(.I(new_n3658_), .ZN(new_n3716_));
  OAI21_X1   g3667(.A1(new_n3714_), .A2(new_n3650_), .B(new_n3716_), .ZN(new_n3717_));
  NAND3_X1   g3668(.A1(new_n3692_), .A2(new_n3717_), .A3(new_n3715_), .ZN(new_n3718_));
  NAND2_X1   g3669(.A1(new_n3679_), .A2(new_n3680_), .ZN(new_n3719_));
  OAI21_X1   g3670(.A1(new_n3673_), .A2(new_n3674_), .B(new_n3719_), .ZN(new_n3720_));
  NAND3_X1   g3671(.A1(new_n3718_), .A2(new_n3483_), .A3(new_n3720_), .ZN(new_n3721_));
  NOR3_X1    g3672(.A1(new_n3721_), .A2(new_n3467_), .A3(new_n3687_), .ZN(new_n3722_));
  NOR2_X1    g3673(.A1(new_n3689_), .A2(new_n3722_), .ZN(new_n3723_));
  NOR2_X1    g3674(.A1(new_n3723_), .A2(new_n3370_), .ZN(new_n3724_));
  NOR3_X1    g3675(.A1(new_n3689_), .A2(new_n3369_), .A3(new_n3722_), .ZN(new_n3725_));
  NAND2_X1   g3676(.A1(new_n3717_), .A2(new_n3715_), .ZN(new_n3726_));
  NOR2_X1    g3677(.A1(new_n3690_), .A2(new_n3478_), .ZN(new_n3727_));
  NOR2_X1    g3678(.A1(new_n3727_), .A2(new_n3482_), .ZN(new_n3728_));
  AOI21_X1   g3679(.A1(new_n3726_), .A2(new_n3483_), .B(new_n3728_), .ZN(new_n3729_));
  INV_X1     g3680(.I(new_n3729_), .ZN(new_n3730_));
  XOR2_X1    g3681(.A1(new_n3675_), .A2(new_n3719_), .Z(new_n3731_));
  NOR4_X1    g3682(.A1(new_n393_), .A2(new_n389_), .A3(new_n878_), .A4(new_n426_), .ZN(new_n3732_));
  NOR4_X1    g3683(.A1(new_n1688_), .A2(new_n615_), .A3(new_n2378_), .A4(new_n3732_), .ZN(new_n3733_));
  INV_X1     g3684(.I(new_n3733_), .ZN(new_n3734_));
  INV_X1     g3685(.I(new_n303_), .ZN(new_n3735_));
  NAND4_X1   g3686(.A1(new_n3735_), .A2(new_n256_), .A3(new_n765_), .A4(new_n341_), .ZN(new_n3736_));
  NOR2_X1    g3687(.A1(new_n3373_), .A2(new_n289_), .ZN(new_n3737_));
  INV_X1     g3688(.I(new_n317_), .ZN(new_n3738_));
  NOR4_X1    g3689(.A1(new_n595_), .A2(new_n272_), .A3(new_n246_), .A4(new_n472_), .ZN(new_n3739_));
  NOR4_X1    g3690(.A1(new_n3739_), .A2(new_n483_), .A3(new_n3738_), .A4(new_n738_), .ZN(new_n3740_));
  NAND4_X1   g3691(.A1(new_n3740_), .A2(new_n2322_), .A3(new_n3737_), .A4(new_n2395_), .ZN(new_n3741_));
  OR3_X2     g3692(.A1(new_n3736_), .A2(new_n2432_), .A3(new_n3741_), .Z(new_n3742_));
  OAI22_X1   g3693(.A1(new_n3730_), .A2(new_n3731_), .B1(new_n3734_), .B2(new_n3742_), .ZN(new_n3743_));
  AOI21_X1   g3694(.A1(new_n3730_), .A2(new_n3731_), .B(new_n3743_), .ZN(new_n3744_));
  NOR4_X1    g3695(.A1(new_n398_), .A2(new_n632_), .A3(new_n438_), .A4(new_n643_), .ZN(new_n3745_));
  NOR4_X1    g3696(.A1(new_n212_), .A2(new_n181_), .A3(new_n306_), .A4(new_n384_), .ZN(new_n3746_));
  NOR4_X1    g3697(.A1(new_n194_), .A2(new_n198_), .A3(new_n3746_), .A4(new_n204_), .ZN(new_n3747_));
  NAND3_X1   g3698(.A1(new_n3747_), .A2(new_n855_), .A3(new_n3745_), .ZN(new_n3748_));
  NOR4_X1    g3699(.A1(new_n3748_), .A2(new_n339_), .A3(new_n593_), .A4(new_n2325_), .ZN(new_n3749_));
  INV_X1     g3700(.I(new_n767_), .ZN(new_n3750_));
  NAND2_X1   g3701(.A1(new_n252_), .A2(new_n774_), .ZN(new_n3751_));
  NOR4_X1    g3702(.A1(new_n1706_), .A2(new_n3751_), .A3(new_n338_), .A4(new_n520_), .ZN(new_n3752_));
  INV_X1     g3703(.I(new_n3752_), .ZN(new_n3753_));
  NOR4_X1    g3704(.A1(new_n326_), .A2(new_n597_), .A3(new_n272_), .A4(new_n434_), .ZN(new_n3754_));
  NOR4_X1    g3705(.A1(new_n715_), .A2(new_n209_), .A3(new_n239_), .A4(new_n377_), .ZN(new_n3755_));
  NOR4_X1    g3706(.A1(new_n3753_), .A2(new_n3750_), .A3(new_n3754_), .A4(new_n3755_), .ZN(new_n3756_));
  NOR4_X1    g3707(.A1(new_n376_), .A2(new_n872_), .A3(new_n335_), .A4(new_n534_), .ZN(new_n3757_));
  NOR4_X1    g3708(.A1(new_n869_), .A2(new_n387_), .A3(new_n238_), .A4(new_n524_), .ZN(new_n3758_));
  NAND3_X1   g3709(.A1(new_n3758_), .A2(new_n291_), .A3(new_n411_), .ZN(new_n3759_));
  NOR3_X1    g3710(.A1(new_n2318_), .A2(new_n3759_), .A3(new_n3757_), .ZN(new_n3760_));
  NAND2_X1   g3711(.A1(new_n3760_), .A2(new_n3756_), .ZN(new_n3761_));
  NOR3_X1    g3712(.A1(new_n3744_), .A2(new_n3749_), .A3(new_n3761_), .ZN(new_n3762_));
  OAI21_X1   g3713(.A1(new_n3724_), .A2(new_n3725_), .B(new_n3762_), .ZN(new_n3763_));
  NOR2_X1    g3714(.A1(new_n3724_), .A2(new_n3725_), .ZN(new_n3764_));
  NAND2_X1   g3715(.A1(new_n3764_), .A2(new_n3744_), .ZN(new_n3765_));
  NAND2_X1   g3716(.A1(new_n3763_), .A2(new_n3765_), .ZN(new_n3766_));
  NOR2_X1    g3717(.A1(new_n741_), .A2(new_n435_), .ZN(new_n3767_));
  NOR2_X1    g3718(.A1(new_n242_), .A2(new_n378_), .ZN(new_n3768_));
  INV_X1     g3719(.I(new_n3768_), .ZN(new_n3769_));
  AOI21_X1   g3720(.A1(new_n3767_), .A2(new_n621_), .B(new_n3769_), .ZN(new_n3770_));
  NAND4_X1   g3721(.A1(new_n530_), .A2(new_n321_), .A3(new_n481_), .A4(new_n545_), .ZN(new_n3771_));
  NAND4_X1   g3722(.A1(new_n809_), .A2(new_n503_), .A3(new_n211_), .A4(new_n930_), .ZN(new_n3772_));
  INV_X1     g3723(.I(new_n1651_), .ZN(new_n3773_));
  NOR2_X1    g3724(.A1(new_n801_), .A2(new_n2376_), .ZN(new_n3774_));
  INV_X1     g3725(.I(new_n3774_), .ZN(new_n3775_));
  NOR2_X1    g3726(.A1(new_n3775_), .A2(new_n3773_), .ZN(new_n3776_));
  NAND4_X1   g3727(.A1(new_n3776_), .A2(new_n3770_), .A3(new_n3771_), .A4(new_n3772_), .ZN(new_n3777_));
  NOR4_X1    g3728(.A1(new_n533_), .A2(new_n324_), .A3(new_n563_), .A4(new_n526_), .ZN(new_n3778_));
  INV_X1     g3729(.I(new_n3778_), .ZN(new_n3779_));
  NOR2_X1    g3730(.A1(new_n3777_), .A2(new_n3779_), .ZN(new_n3780_));
  NOR4_X1    g3731(.A1(new_n597_), .A2(new_n608_), .A3(new_n500_), .A4(new_n747_), .ZN(new_n3781_));
  NAND2_X1   g3732(.A1(new_n465_), .A2(new_n3781_), .ZN(new_n3782_));
  NOR2_X1    g3733(.A1(new_n3782_), .A2(new_n3378_), .ZN(new_n3783_));
  INV_X1     g3734(.I(new_n3383_), .ZN(new_n3784_));
  INV_X1     g3735(.I(new_n264_), .ZN(new_n3785_));
  NOR2_X1    g3736(.A1(new_n189_), .A2(new_n588_), .ZN(new_n3786_));
  INV_X1     g3737(.I(new_n3786_), .ZN(new_n3787_));
  NOR4_X1    g3738(.A1(new_n3787_), .A2(new_n3785_), .A3(new_n501_), .A4(new_n543_), .ZN(new_n3788_));
  INV_X1     g3739(.I(new_n3788_), .ZN(new_n3789_));
  NOR4_X1    g3740(.A1(new_n1706_), .A2(new_n974_), .A3(new_n209_), .A4(new_n488_), .ZN(new_n3790_));
  NOR4_X1    g3741(.A1(new_n432_), .A2(new_n3784_), .A3(new_n3789_), .A4(new_n3790_), .ZN(new_n3791_));
  NAND3_X1   g3742(.A1(new_n3780_), .A2(new_n3791_), .A3(new_n3783_), .ZN(new_n3792_));
  NOR2_X1    g3743(.A1(new_n3766_), .A2(new_n3792_), .ZN(new_n3793_));
  NAND2_X1   g3744(.A1(new_n3467_), .A2(new_n3369_), .ZN(new_n3794_));
  INV_X1     g3745(.I(new_n3794_), .ZN(new_n3795_));
  INV_X1     g3746(.I(new_n3359_), .ZN(new_n3796_));
  OAI21_X1   g3747(.A1(new_n3133_), .A2(new_n3135_), .B(new_n3358_), .ZN(new_n3797_));
  NAND3_X1   g3748(.A1(new_n3464_), .A2(new_n69_), .A3(new_n3465_), .ZN(new_n3798_));
  OAI21_X1   g3749(.A1(new_n3448_), .A2(new_n3460_), .B(new_n2739_), .ZN(new_n3799_));
  AOI22_X1   g3750(.A1(new_n3796_), .A2(new_n3797_), .B1(new_n3799_), .B2(new_n3798_), .ZN(new_n3800_));
  NOR3_X1    g3751(.A1(new_n3721_), .A2(new_n3687_), .A3(new_n3800_), .ZN(new_n3801_));
  NOR2_X1    g3752(.A1(new_n3801_), .A2(new_n3795_), .ZN(new_n3802_));
  OAI22_X1   g3753(.A1(new_n2551_), .A2(new_n2752_), .B1(new_n2558_), .B2(new_n2742_), .ZN(new_n3803_));
  NAND2_X1   g3754(.A1(new_n3418_), .A2(new_n2748_), .ZN(new_n3804_));
  AOI21_X1   g3755(.A1(new_n3804_), .A2(new_n3803_), .B(new_n72_), .ZN(new_n3805_));
  NAND3_X1   g3756(.A1(new_n3472_), .A2(new_n62_), .A3(new_n3805_), .ZN(new_n3806_));
  NOR2_X1    g3757(.A1(new_n3471_), .A2(new_n3418_), .ZN(new_n3807_));
  OR2_X2     g3758(.A1(new_n3469_), .A2(new_n3470_), .Z(new_n3808_));
  AOI21_X1   g3759(.A1(new_n3808_), .A2(new_n2723_), .B(new_n3419_), .ZN(new_n3809_));
  OAI21_X1   g3760(.A1(new_n3809_), .A2(new_n3807_), .B(new_n3805_), .ZN(new_n3810_));
  NAND2_X1   g3761(.A1(new_n3810_), .A2(new_n943_), .ZN(new_n3811_));
  NAND2_X1   g3762(.A1(new_n3811_), .A2(new_n3806_), .ZN(new_n3812_));
  OAI22_X1   g3763(.A1(new_n2576_), .A2(new_n3007_), .B1(new_n2619_), .B2(new_n2774_), .ZN(new_n3813_));
  NAND2_X1   g3764(.A1(new_n2586_), .A2(new_n3009_), .ZN(new_n3814_));
  AOI21_X1   g3765(.A1(new_n3813_), .A2(new_n3814_), .B(new_n2779_), .ZN(new_n3815_));
  NAND3_X1   g3766(.A1(new_n3330_), .A2(new_n1132_), .A3(new_n3815_), .ZN(new_n3816_));
  INV_X1     g3767(.I(new_n3816_), .ZN(new_n3817_));
  AOI21_X1   g3768(.A1(new_n3330_), .A2(new_n3815_), .B(new_n1132_), .ZN(new_n3818_));
  NAND2_X1   g3769(.A1(new_n2983_), .A2(new_n2987_), .ZN(new_n3819_));
  OAI22_X1   g3770(.A1(new_n2637_), .A2(new_n2882_), .B1(new_n2696_), .B2(new_n2850_), .ZN(new_n3820_));
  NAND2_X1   g3771(.A1(new_n2628_), .A2(new_n2855_), .ZN(new_n3821_));
  AOI21_X1   g3772(.A1(new_n3821_), .A2(new_n3820_), .B(new_n2881_), .ZN(new_n3822_));
  NAND3_X1   g3773(.A1(new_n3041_), .A2(new_n790_), .A3(new_n3822_), .ZN(new_n3823_));
  AOI21_X1   g3774(.A1(new_n3041_), .A2(new_n3822_), .B(new_n790_), .ZN(new_n3824_));
  INV_X1     g3775(.I(new_n3824_), .ZN(new_n3825_));
  NAND2_X1   g3776(.A1(new_n2673_), .A2(new_n658_), .ZN(new_n3826_));
  AOI21_X1   g3777(.A1(new_n2961_), .A2(new_n2957_), .B(new_n2963_), .ZN(new_n3827_));
  NAND3_X1   g3778(.A1(new_n3533_), .A2(new_n3534_), .A3(new_n2824_), .ZN(new_n3828_));
  NAND2_X1   g3779(.A1(new_n2844_), .A2(new_n2795_), .ZN(new_n3829_));
  NAND2_X1   g3780(.A1(new_n2668_), .A2(new_n2829_), .ZN(new_n3830_));
  AOI22_X1   g3781(.A1(new_n2700_), .A2(new_n2790_), .B1(new_n3829_), .B2(new_n3830_), .ZN(new_n3831_));
  NAND2_X1   g3782(.A1(new_n3828_), .A2(new_n3831_), .ZN(new_n3832_));
  NOR3_X1    g3783(.A1(new_n2966_), .A2(new_n3832_), .A3(new_n3827_), .ZN(new_n3833_));
  OAI22_X1   g3784(.A1(new_n2970_), .A2(new_n2971_), .B1(new_n2967_), .B2(new_n2962_), .ZN(new_n3834_));
  INV_X1     g3785(.I(new_n3831_), .ZN(new_n3835_));
  AOI21_X1   g3786(.A1(new_n2880_), .A2(new_n2824_), .B(new_n3835_), .ZN(new_n3836_));
  NOR2_X1    g3787(.A1(new_n3834_), .A2(new_n3836_), .ZN(new_n3837_));
  NOR2_X1    g3788(.A1(new_n3837_), .A2(new_n3833_), .ZN(new_n3838_));
  XNOR2_X1   g3789(.A1(new_n3838_), .A2(new_n3826_), .ZN(new_n3839_));
  INV_X1     g3790(.I(new_n3839_), .ZN(new_n3840_));
  NAND3_X1   g3791(.A1(new_n3825_), .A2(new_n3840_), .A3(new_n3823_), .ZN(new_n3841_));
  INV_X1     g3792(.I(new_n3823_), .ZN(new_n3842_));
  OAI21_X1   g3793(.A1(new_n3842_), .A2(new_n3824_), .B(new_n3839_), .ZN(new_n3843_));
  AOI22_X1   g3794(.A1(new_n3819_), .A2(new_n2985_), .B1(new_n3843_), .B2(new_n3841_), .ZN(new_n3844_));
  OAI21_X1   g3795(.A1(new_n2933_), .A2(new_n2986_), .B(new_n2985_), .ZN(new_n3845_));
  OAI21_X1   g3796(.A1(new_n3842_), .A2(new_n3824_), .B(new_n3840_), .ZN(new_n3846_));
  NAND3_X1   g3797(.A1(new_n3825_), .A2(new_n3823_), .A3(new_n3839_), .ZN(new_n3847_));
  AOI21_X1   g3798(.A1(new_n3846_), .A2(new_n3847_), .B(new_n3845_), .ZN(new_n3848_));
  NOR2_X1    g3799(.A1(new_n3844_), .A2(new_n3848_), .ZN(new_n3849_));
  INV_X1     g3800(.I(new_n3849_), .ZN(new_n3850_));
  NOR3_X1    g3801(.A1(new_n3817_), .A2(new_n3850_), .A3(new_n3818_), .ZN(new_n3851_));
  INV_X1     g3802(.I(new_n3818_), .ZN(new_n3852_));
  AOI21_X1   g3803(.A1(new_n3852_), .A2(new_n3816_), .B(new_n3849_), .ZN(new_n3853_));
  NAND3_X1   g3804(.A1(new_n3127_), .A2(new_n2990_), .A3(new_n2997_), .ZN(new_n3854_));
  INV_X1     g3805(.I(new_n3854_), .ZN(new_n3855_));
  NOR3_X1    g3806(.A1(new_n3855_), .A2(new_n3851_), .A3(new_n3853_), .ZN(new_n3856_));
  NAND3_X1   g3807(.A1(new_n3852_), .A2(new_n3816_), .A3(new_n3849_), .ZN(new_n3857_));
  OAI21_X1   g3808(.A1(new_n3817_), .A2(new_n3818_), .B(new_n3850_), .ZN(new_n3858_));
  AOI21_X1   g3809(.A1(new_n3858_), .A2(new_n3857_), .B(new_n3854_), .ZN(new_n3859_));
  NOR2_X1    g3810(.A1(new_n3856_), .A2(new_n3859_), .ZN(new_n3860_));
  INV_X1     g3811(.I(new_n2756_), .ZN(new_n3861_));
  NOR3_X1    g3812(.A1(new_n3131_), .A2(new_n3130_), .A3(new_n62_), .ZN(new_n3862_));
  AOI21_X1   g3813(.A1(new_n3128_), .A2(new_n3120_), .B(new_n943_), .ZN(new_n3863_));
  OAI21_X1   g3814(.A1(new_n3863_), .A2(new_n3862_), .B(new_n3861_), .ZN(new_n3864_));
  NOR2_X1    g3815(.A1(new_n2735_), .A2(new_n2723_), .ZN(new_n3865_));
  NOR2_X1    g3816(.A1(new_n2721_), .A2(new_n2560_), .ZN(new_n3866_));
  OAI21_X1   g3817(.A1(new_n3865_), .A2(new_n3866_), .B(new_n71_), .ZN(new_n3867_));
  NAND3_X1   g3818(.A1(new_n3867_), .A2(new_n62_), .A3(new_n2754_), .ZN(new_n3868_));
  OAI21_X1   g3819(.A1(new_n2737_), .A2(new_n2755_), .B(new_n943_), .ZN(new_n3869_));
  NAND2_X1   g3820(.A1(new_n3869_), .A2(new_n3868_), .ZN(new_n3870_));
  NAND3_X1   g3821(.A1(new_n3870_), .A2(new_n3120_), .A3(new_n3128_), .ZN(new_n3871_));
  NAND3_X1   g3822(.A1(new_n3864_), .A2(new_n3134_), .A3(new_n3871_), .ZN(new_n3872_));
  OAI21_X1   g3823(.A1(new_n3872_), .A2(new_n3367_), .B(new_n3860_), .ZN(new_n3873_));
  NAND3_X1   g3824(.A1(new_n3858_), .A2(new_n3857_), .A3(new_n3854_), .ZN(new_n3874_));
  INV_X1     g3825(.I(new_n3859_), .ZN(new_n3875_));
  NAND2_X1   g3826(.A1(new_n3875_), .A2(new_n3874_), .ZN(new_n3876_));
  NAND4_X1   g3827(.A1(new_n3360_), .A2(new_n3358_), .A3(new_n3876_), .A4(new_n3871_), .ZN(new_n3877_));
  AOI21_X1   g3828(.A1(new_n3877_), .A2(new_n3873_), .B(new_n3812_), .ZN(new_n3878_));
  NOR2_X1    g3829(.A1(new_n3810_), .A2(new_n943_), .ZN(new_n3879_));
  AOI21_X1   g3830(.A1(new_n3472_), .A2(new_n3805_), .B(new_n62_), .ZN(new_n3880_));
  NOR2_X1    g3831(.A1(new_n3879_), .A2(new_n3880_), .ZN(new_n3881_));
  INV_X1     g3832(.I(new_n3873_), .ZN(new_n3882_));
  NOR3_X1    g3833(.A1(new_n3872_), .A2(new_n3367_), .A3(new_n3860_), .ZN(new_n3883_));
  NOR3_X1    g3834(.A1(new_n3882_), .A2(new_n3881_), .A3(new_n3883_), .ZN(new_n3884_));
  NOR2_X1    g3835(.A1(new_n3884_), .A2(new_n3878_), .ZN(new_n3885_));
  INV_X1     g3836(.I(new_n3885_), .ZN(new_n3886_));
  NOR2_X1    g3837(.A1(new_n3391_), .A2(new_n591_), .ZN(new_n3887_));
  NOR3_X1    g3838(.A1(new_n649_), .A2(new_n280_), .A3(new_n631_), .ZN(new_n3888_));
  NOR4_X1    g3839(.A1(new_n617_), .A2(new_n500_), .A3(new_n378_), .A4(new_n595_), .ZN(new_n3889_));
  NAND4_X1   g3840(.A1(new_n3889_), .A2(new_n3887_), .A3(new_n636_), .A4(new_n3888_), .ZN(new_n3890_));
  INV_X1     g3841(.I(new_n3890_), .ZN(new_n3891_));
  NAND2_X1   g3842(.A1(new_n3413_), .A2(new_n3891_), .ZN(new_n3892_));
  NAND2_X1   g3843(.A1(new_n3412_), .A2(new_n3890_), .ZN(new_n3893_));
  NAND2_X1   g3844(.A1(new_n3892_), .A2(new_n3893_), .ZN(new_n3894_));
  INV_X1     g3845(.I(new_n3894_), .ZN(new_n3895_));
  INV_X1     g3846(.I(new_n3437_), .ZN(new_n3896_));
  AOI21_X1   g3847(.A1(new_n3434_), .A2(new_n3436_), .B(new_n3414_), .ZN(new_n3897_));
  INV_X1     g3848(.I(new_n3897_), .ZN(new_n3898_));
  NAND3_X1   g3849(.A1(new_n3414_), .A2(new_n3436_), .A3(new_n3434_), .ZN(new_n3899_));
  NAND4_X1   g3850(.A1(new_n3898_), .A2(new_n3896_), .A3(new_n3438_), .A4(new_n3899_), .ZN(new_n3900_));
  NAND3_X1   g3851(.A1(new_n3432_), .A2(new_n3668_), .A3(new_n3900_), .ZN(new_n3901_));
  NAND3_X1   g3852(.A1(new_n3425_), .A2(new_n3449_), .A3(new_n3900_), .ZN(new_n3902_));
  NAND2_X1   g3853(.A1(new_n3901_), .A2(new_n3902_), .ZN(new_n3903_));
  NAND2_X1   g3854(.A1(new_n3903_), .A2(new_n3414_), .ZN(new_n3904_));
  INV_X1     g3855(.I(new_n3899_), .ZN(new_n3905_));
  NOR4_X1    g3856(.A1(new_n3905_), .A2(new_n3439_), .A3(new_n3437_), .A4(new_n3897_), .ZN(new_n3906_));
  NOR3_X1    g3857(.A1(new_n3425_), .A2(new_n3449_), .A3(new_n3906_), .ZN(new_n3907_));
  NOR3_X1    g3858(.A1(new_n2721_), .A2(new_n2551_), .A3(new_n3418_), .ZN(new_n3908_));
  NOR3_X1    g3859(.A1(new_n3427_), .A2(new_n3908_), .A3(new_n2558_), .ZN(new_n3909_));
  NOR4_X1    g3860(.A1(new_n3909_), .A2(new_n3424_), .A3(new_n3668_), .A4(new_n3906_), .ZN(new_n3910_));
  NOR2_X1    g3861(.A1(new_n3907_), .A2(new_n3910_), .ZN(new_n3911_));
  NAND2_X1   g3862(.A1(new_n3911_), .A2(new_n3444_), .ZN(new_n3912_));
  AOI21_X1   g3863(.A1(new_n3904_), .A2(new_n3912_), .B(new_n3895_), .ZN(new_n3913_));
  NOR3_X1    g3864(.A1(new_n3907_), .A2(new_n3910_), .A3(new_n3444_), .ZN(new_n3914_));
  AOI21_X1   g3865(.A1(new_n3901_), .A2(new_n3902_), .B(new_n3414_), .ZN(new_n3915_));
  NOR2_X1    g3866(.A1(new_n3915_), .A2(new_n3914_), .ZN(new_n3916_));
  NOR2_X1    g3867(.A1(new_n3916_), .A2(new_n3894_), .ZN(new_n3917_));
  AOI22_X1   g3868(.A1(new_n3668_), .A2(new_n3450_), .B1(new_n3414_), .B2(new_n3487_), .ZN(new_n3918_));
  AOI21_X1   g3869(.A1(new_n3456_), .A2(new_n3895_), .B(new_n3918_), .ZN(new_n3919_));
  NOR2_X1    g3870(.A1(new_n3919_), .A2(new_n3473_), .ZN(new_n3920_));
  OAI21_X1   g3871(.A1(new_n3917_), .A2(new_n3913_), .B(new_n3920_), .ZN(new_n3921_));
  NOR2_X1    g3872(.A1(new_n3921_), .A2(new_n2739_), .ZN(new_n3922_));
  NOR2_X1    g3873(.A1(new_n3911_), .A2(new_n3444_), .ZN(new_n3923_));
  NOR2_X1    g3874(.A1(new_n3903_), .A2(new_n3414_), .ZN(new_n3924_));
  OAI21_X1   g3875(.A1(new_n3924_), .A2(new_n3923_), .B(new_n3894_), .ZN(new_n3925_));
  OAI21_X1   g3876(.A1(new_n3894_), .A2(new_n3916_), .B(new_n3925_), .ZN(new_n3926_));
  AOI21_X1   g3877(.A1(new_n3926_), .A2(new_n3920_), .B(new_n69_), .ZN(new_n3927_));
  NOR2_X1    g3878(.A1(new_n3927_), .A2(new_n3922_), .ZN(new_n3928_));
  NOR2_X1    g3879(.A1(new_n3886_), .A2(new_n3928_), .ZN(new_n3929_));
  INV_X1     g3880(.I(new_n3928_), .ZN(new_n3930_));
  NOR2_X1    g3881(.A1(new_n3930_), .A2(new_n3885_), .ZN(new_n3931_));
  NOR2_X1    g3882(.A1(new_n3929_), .A2(new_n3931_), .ZN(new_n3932_));
  NOR2_X1    g3883(.A1(new_n3932_), .A2(new_n3802_), .ZN(new_n3933_));
  INV_X1     g3884(.I(new_n3802_), .ZN(new_n3934_));
  INV_X1     g3885(.I(new_n3932_), .ZN(new_n3935_));
  NOR2_X1    g3886(.A1(new_n3935_), .A2(new_n3934_), .ZN(new_n3936_));
  NOR2_X1    g3887(.A1(new_n3936_), .A2(new_n3933_), .ZN(new_n3937_));
  AOI21_X1   g3888(.A1(new_n3766_), .A2(new_n3792_), .B(new_n3937_), .ZN(new_n3938_));
  NOR2_X1    g3889(.A1(new_n3938_), .A2(new_n3793_), .ZN(new_n3939_));
  NOR2_X1    g3890(.A1(new_n3146_), .A2(new_n3143_), .ZN(new_n3940_));
  AOI22_X1   g3891(.A1(new_n2577_), .A2(new_n3009_), .B1(new_n2586_), .B2(new_n2773_), .ZN(new_n3941_));
  AOI21_X1   g3892(.A1(new_n2559_), .A2(new_n2776_), .B(new_n3941_), .ZN(new_n3942_));
  NOR3_X1    g3893(.A1(new_n3940_), .A2(new_n2779_), .A3(new_n3942_), .ZN(new_n3943_));
  NAND2_X1   g3894(.A1(new_n3943_), .A2(new_n1132_), .ZN(new_n3944_));
  OR2_X2     g3895(.A1(new_n3943_), .A2(new_n1132_), .Z(new_n3945_));
  NAND2_X1   g3896(.A1(new_n3945_), .A2(new_n3944_), .ZN(new_n3946_));
  OAI22_X1   g3897(.A1(new_n2619_), .A2(new_n2856_), .B1(new_n2696_), .B2(new_n2882_), .ZN(new_n3947_));
  NAND2_X1   g3898(.A1(new_n2628_), .A2(new_n2851_), .ZN(new_n3948_));
  AOI21_X1   g3899(.A1(new_n3947_), .A2(new_n3948_), .B(new_n2881_), .ZN(new_n3949_));
  OAI21_X1   g3900(.A1(new_n3006_), .A2(new_n3004_), .B(new_n3949_), .ZN(new_n3950_));
  XOR2_X1    g3901(.A1(new_n3950_), .A2(new_n790_), .Z(new_n3951_));
  NAND2_X1   g3902(.A1(new_n3834_), .A2(new_n3836_), .ZN(new_n3952_));
  AOI22_X1   g3903(.A1(new_n2964_), .A2(new_n2965_), .B1(new_n2946_), .B2(new_n2963_), .ZN(new_n3953_));
  NAND2_X1   g3904(.A1(new_n3953_), .A2(new_n3832_), .ZN(new_n3954_));
  AOI22_X1   g3905(.A1(new_n3952_), .A2(new_n3954_), .B1(new_n658_), .B2(new_n3836_), .ZN(new_n3955_));
  INV_X1     g3906(.I(new_n3955_), .ZN(new_n3956_));
  NOR3_X1    g3907(.A1(new_n3834_), .A2(new_n658_), .A3(new_n3832_), .ZN(new_n3957_));
  INV_X1     g3908(.I(new_n3957_), .ZN(new_n3958_));
  AOI21_X1   g3909(.A1(new_n3952_), .A2(new_n3954_), .B(new_n659_), .ZN(new_n3959_));
  NOR3_X1    g3910(.A1(new_n3837_), .A2(new_n3833_), .A3(new_n658_), .ZN(new_n3960_));
  OAI21_X1   g3911(.A1(new_n3959_), .A2(new_n3960_), .B(new_n2672_), .ZN(new_n3961_));
  NAND3_X1   g3912(.A1(new_n3961_), .A2(new_n3956_), .A3(new_n3958_), .ZN(new_n3962_));
  AOI21_X1   g3913(.A1(new_n2840_), .A2(new_n2838_), .B(new_n2796_), .ZN(new_n3963_));
  OAI22_X1   g3914(.A1(new_n2663_), .A2(new_n2794_), .B1(new_n2691_), .B2(new_n2830_), .ZN(new_n3964_));
  OAI21_X1   g3915(.A1(new_n2637_), .A2(new_n2791_), .B(new_n3964_), .ZN(new_n3965_));
  NOR2_X1    g3916(.A1(new_n2668_), .A2(new_n659_), .ZN(new_n3966_));
  INV_X1     g3917(.I(new_n3966_), .ZN(new_n3967_));
  OAI21_X1   g3918(.A1(new_n3963_), .A2(new_n3965_), .B(new_n3967_), .ZN(new_n3968_));
  NOR3_X1    g3919(.A1(new_n3963_), .A2(new_n3965_), .A3(new_n3967_), .ZN(new_n3969_));
  INV_X1     g3920(.I(new_n3969_), .ZN(new_n3970_));
  NAND2_X1   g3921(.A1(new_n3970_), .A2(new_n3968_), .ZN(new_n3971_));
  AND2_X2    g3922(.A1(new_n3962_), .A2(new_n3971_), .Z(new_n3972_));
  NOR2_X1    g3923(.A1(new_n3962_), .A2(new_n3971_), .ZN(new_n3973_));
  OAI21_X1   g3924(.A1(new_n3972_), .A2(new_n3973_), .B(new_n3951_), .ZN(new_n3974_));
  XOR2_X1    g3925(.A1(new_n3950_), .A2(new_n576_), .Z(new_n3975_));
  NAND4_X1   g3926(.A1(new_n3961_), .A2(new_n3956_), .A3(new_n3958_), .A4(new_n3971_), .ZN(new_n3976_));
  INV_X1     g3927(.I(new_n3968_), .ZN(new_n3977_));
  NOR2_X1    g3928(.A1(new_n3977_), .A2(new_n3969_), .ZN(new_n3978_));
  NAND2_X1   g3929(.A1(new_n3962_), .A2(new_n3978_), .ZN(new_n3979_));
  NAND2_X1   g3930(.A1(new_n3979_), .A2(new_n3976_), .ZN(new_n3980_));
  NAND2_X1   g3931(.A1(new_n3975_), .A2(new_n3980_), .ZN(new_n3981_));
  INV_X1     g3932(.I(new_n3841_), .ZN(new_n3982_));
  AOI21_X1   g3933(.A1(new_n3845_), .A2(new_n3843_), .B(new_n3982_), .ZN(new_n3983_));
  NAND3_X1   g3934(.A1(new_n3974_), .A2(new_n3983_), .A3(new_n3981_), .ZN(new_n3984_));
  INV_X1     g3935(.I(new_n3984_), .ZN(new_n3985_));
  AOI21_X1   g3936(.A1(new_n3974_), .A2(new_n3981_), .B(new_n3983_), .ZN(new_n3986_));
  NOR3_X1    g3937(.A1(new_n3946_), .A2(new_n3985_), .A3(new_n3986_), .ZN(new_n3987_));
  INV_X1     g3938(.I(new_n3946_), .ZN(new_n3988_));
  INV_X1     g3939(.I(new_n3986_), .ZN(new_n3989_));
  AOI21_X1   g3940(.A1(new_n3984_), .A2(new_n3989_), .B(new_n3988_), .ZN(new_n3990_));
  NOR2_X1    g3941(.A1(new_n3990_), .A2(new_n3987_), .ZN(new_n3991_));
  INV_X1     g3942(.I(new_n3991_), .ZN(new_n3992_));
  NOR2_X1    g3943(.A1(new_n3665_), .A2(new_n3666_), .ZN(new_n3993_));
  INV_X1     g3944(.I(new_n3993_), .ZN(new_n3994_));
  OAI22_X1   g3945(.A1(new_n3419_), .A2(new_n2752_), .B1(new_n2551_), .B2(new_n2742_), .ZN(new_n3995_));
  NAND2_X1   g3946(.A1(new_n3668_), .A2(new_n2748_), .ZN(new_n3996_));
  AOI21_X1   g3947(.A1(new_n3996_), .A2(new_n3995_), .B(new_n72_), .ZN(new_n3997_));
  NAND3_X1   g3948(.A1(new_n3994_), .A2(new_n62_), .A3(new_n3997_), .ZN(new_n3998_));
  AOI21_X1   g3949(.A1(new_n3994_), .A2(new_n3997_), .B(new_n62_), .ZN(new_n3999_));
  INV_X1     g3950(.I(new_n3999_), .ZN(new_n4000_));
  NAND2_X1   g3951(.A1(new_n4000_), .A2(new_n3998_), .ZN(new_n4001_));
  NOR2_X1    g3952(.A1(new_n4001_), .A2(new_n3992_), .ZN(new_n4002_));
  INV_X1     g3953(.I(new_n3998_), .ZN(new_n4003_));
  NOR2_X1    g3954(.A1(new_n4003_), .A2(new_n3999_), .ZN(new_n4004_));
  NOR2_X1    g3955(.A1(new_n4004_), .A2(new_n3991_), .ZN(new_n4005_));
  NOR2_X1    g3956(.A1(new_n4002_), .A2(new_n4005_), .ZN(new_n4006_));
  NAND3_X1   g3957(.A1(new_n3901_), .A2(new_n3902_), .A3(new_n3414_), .ZN(new_n4007_));
  OAI21_X1   g3958(.A1(new_n3907_), .A2(new_n3910_), .B(new_n3444_), .ZN(new_n4008_));
  NAND2_X1   g3959(.A1(new_n4007_), .A2(new_n4008_), .ZN(new_n4009_));
  NAND2_X1   g3960(.A1(new_n3412_), .A2(new_n3891_), .ZN(new_n4010_));
  NOR3_X1    g3961(.A1(new_n3775_), .A2(new_n588_), .A3(new_n3382_), .ZN(new_n4011_));
  NOR4_X1    g3962(.A1(new_n326_), .A2(new_n250_), .A3(new_n873_), .A4(new_n384_), .ZN(new_n4012_));
  NOR3_X1    g3963(.A1(new_n4011_), .A2(new_n477_), .A3(new_n4012_), .ZN(new_n4013_));
  INV_X1     g3964(.I(new_n422_), .ZN(new_n4014_));
  NOR2_X1    g3965(.A1(new_n385_), .A2(new_n391_), .ZN(new_n4015_));
  NOR2_X1    g3966(.A1(new_n3738_), .A2(new_n518_), .ZN(new_n4016_));
  NAND4_X1   g3967(.A1(new_n4016_), .A2(new_n4014_), .A3(new_n2380_), .A4(new_n4015_), .ZN(new_n4017_));
  NOR4_X1    g3968(.A1(new_n533_), .A2(new_n242_), .A3(new_n472_), .A4(new_n529_), .ZN(new_n4018_));
  NOR4_X1    g3969(.A1(new_n313_), .A2(new_n4017_), .A3(new_n154_), .A4(new_n4018_), .ZN(new_n4019_));
  NAND3_X1   g3970(.A1(new_n4013_), .A2(new_n4019_), .A3(new_n958_), .ZN(new_n4020_));
  AND2_X2    g3971(.A1(new_n4010_), .A2(new_n4020_), .Z(new_n4021_));
  NOR2_X1    g3972(.A1(new_n4010_), .A2(new_n4020_), .ZN(new_n4022_));
  NOR2_X1    g3973(.A1(new_n4021_), .A2(new_n4022_), .ZN(new_n4023_));
  OAI21_X1   g3974(.A1(new_n3907_), .A2(new_n3910_), .B(new_n3895_), .ZN(new_n4024_));
  NAND3_X1   g3975(.A1(new_n3901_), .A2(new_n3902_), .A3(new_n3894_), .ZN(new_n4025_));
  NAND2_X1   g3976(.A1(new_n4025_), .A2(new_n4024_), .ZN(new_n4026_));
  NAND3_X1   g3977(.A1(new_n4009_), .A2(new_n4026_), .A3(new_n4023_), .ZN(new_n4027_));
  INV_X1     g3978(.I(new_n4023_), .ZN(new_n4028_));
  AOI21_X1   g3979(.A1(new_n3901_), .A2(new_n3902_), .B(new_n3894_), .ZN(new_n4029_));
  NOR3_X1    g3980(.A1(new_n3907_), .A2(new_n3910_), .A3(new_n3895_), .ZN(new_n4030_));
  NOR2_X1    g3981(.A1(new_n4029_), .A2(new_n4030_), .ZN(new_n4031_));
  OAI21_X1   g3982(.A1(new_n3916_), .A2(new_n4031_), .B(new_n4028_), .ZN(new_n4032_));
  AOI21_X1   g3983(.A1(new_n4032_), .A2(new_n4027_), .B(new_n3473_), .ZN(new_n4033_));
  NOR2_X1    g3984(.A1(new_n3444_), .A2(new_n3451_), .ZN(new_n4034_));
  NOR2_X1    g3985(.A1(new_n3894_), .A2(new_n3453_), .ZN(new_n4035_));
  OAI22_X1   g3986(.A1(new_n4035_), .A2(new_n4034_), .B1(new_n4023_), .B2(new_n3457_), .ZN(new_n4036_));
  NOR2_X1    g3987(.A1(new_n3872_), .A2(new_n3367_), .ZN(new_n4037_));
  NOR3_X1    g3988(.A1(new_n3876_), .A2(new_n3879_), .A3(new_n3880_), .ZN(new_n4038_));
  NAND2_X1   g3989(.A1(new_n3812_), .A2(new_n3876_), .ZN(new_n4039_));
  AOI21_X1   g3990(.A1(new_n4037_), .A2(new_n4039_), .B(new_n4038_), .ZN(new_n4040_));
  OAI21_X1   g3991(.A1(new_n4033_), .A2(new_n4036_), .B(new_n4040_), .ZN(new_n4041_));
  INV_X1     g3992(.I(new_n4033_), .ZN(new_n4042_));
  INV_X1     g3993(.I(new_n4036_), .ZN(new_n4043_));
  NAND4_X1   g3994(.A1(new_n3358_), .A2(new_n3864_), .A3(new_n3134_), .A4(new_n3871_), .ZN(new_n4044_));
  NAND2_X1   g3995(.A1(new_n3881_), .A2(new_n3860_), .ZN(new_n4045_));
  AOI21_X1   g3996(.A1(new_n3806_), .A2(new_n3811_), .B(new_n3860_), .ZN(new_n4046_));
  OAI21_X1   g3997(.A1(new_n4044_), .A2(new_n4046_), .B(new_n4045_), .ZN(new_n4047_));
  NAND3_X1   g3998(.A1(new_n4042_), .A2(new_n4047_), .A3(new_n4043_), .ZN(new_n4048_));
  AOI21_X1   g3999(.A1(new_n4048_), .A2(new_n4041_), .B(new_n2739_), .ZN(new_n4049_));
  NOR2_X1    g4000(.A1(new_n4033_), .A2(new_n4036_), .ZN(new_n4050_));
  NOR2_X1    g4001(.A1(new_n4050_), .A2(new_n4047_), .ZN(new_n4051_));
  NOR3_X1    g4002(.A1(new_n4040_), .A2(new_n4033_), .A3(new_n4036_), .ZN(new_n4052_));
  NOR3_X1    g4003(.A1(new_n4051_), .A2(new_n69_), .A3(new_n4052_), .ZN(new_n4053_));
  OAI21_X1   g4004(.A1(new_n4053_), .A2(new_n4049_), .B(new_n4006_), .ZN(new_n4054_));
  NAND2_X1   g4005(.A1(new_n4004_), .A2(new_n3991_), .ZN(new_n4055_));
  NAND2_X1   g4006(.A1(new_n4001_), .A2(new_n3992_), .ZN(new_n4056_));
  NAND2_X1   g4007(.A1(new_n4056_), .A2(new_n4055_), .ZN(new_n4057_));
  OAI21_X1   g4008(.A1(new_n4051_), .A2(new_n4052_), .B(new_n69_), .ZN(new_n4058_));
  NAND3_X1   g4009(.A1(new_n4048_), .A2(new_n4041_), .A3(new_n2739_), .ZN(new_n4059_));
  NAND3_X1   g4010(.A1(new_n4058_), .A2(new_n4059_), .A3(new_n4057_), .ZN(new_n4060_));
  NAND4_X1   g4011(.A1(new_n3934_), .A2(new_n3886_), .A3(new_n4054_), .A4(new_n4060_), .ZN(new_n4061_));
  AOI21_X1   g4012(.A1(new_n4058_), .A2(new_n4059_), .B(new_n4057_), .ZN(new_n4062_));
  NOR3_X1    g4013(.A1(new_n4053_), .A2(new_n4049_), .A3(new_n4006_), .ZN(new_n4063_));
  NAND2_X1   g4014(.A1(new_n3934_), .A2(new_n3886_), .ZN(new_n4064_));
  OAI21_X1   g4015(.A1(new_n4062_), .A2(new_n4063_), .B(new_n4064_), .ZN(new_n4065_));
  NAND2_X1   g4016(.A1(new_n3802_), .A2(new_n3885_), .ZN(new_n4066_));
  NAND3_X1   g4017(.A1(new_n4064_), .A2(new_n3928_), .A3(new_n4066_), .ZN(new_n4067_));
  AND3_X2    g4018(.A1(new_n4065_), .A2(new_n4061_), .A3(new_n4067_), .Z(new_n4068_));
  AOI21_X1   g4019(.A1(new_n4065_), .A2(new_n4061_), .B(new_n4067_), .ZN(new_n4069_));
  NOR2_X1    g4020(.A1(new_n4068_), .A2(new_n4069_), .ZN(new_n4070_));
  NOR3_X1    g4021(.A1(new_n3784_), .A2(new_n1011_), .A3(new_n876_), .ZN(new_n4071_));
  NAND3_X1   g4022(.A1(new_n813_), .A2(new_n542_), .A3(new_n929_), .ZN(new_n4072_));
  NOR4_X1    g4023(.A1(new_n3775_), .A2(new_n555_), .A3(new_n3750_), .A4(new_n4072_), .ZN(new_n4073_));
  NAND4_X1   g4024(.A1(new_n1684_), .A2(new_n513_), .A3(new_n4071_), .A4(new_n4073_), .ZN(new_n4074_));
  NAND2_X1   g4025(.A1(new_n4070_), .A2(new_n4074_), .ZN(new_n4075_));
  NOR2_X1    g4026(.A1(new_n4070_), .A2(new_n4074_), .ZN(new_n4076_));
  INV_X1     g4027(.I(new_n4076_), .ZN(new_n4077_));
  NAND2_X1   g4028(.A1(new_n4077_), .A2(new_n4075_), .ZN(new_n4078_));
  INV_X1     g4029(.I(new_n3792_), .ZN(new_n4079_));
  AOI21_X1   g4030(.A1(new_n3763_), .A2(new_n3765_), .B(new_n3934_), .ZN(new_n4080_));
  INV_X1     g4031(.I(new_n4080_), .ZN(new_n4081_));
  NAND3_X1   g4032(.A1(new_n3763_), .A2(new_n3765_), .A3(new_n3934_), .ZN(new_n4082_));
  AOI21_X1   g4033(.A1(new_n4081_), .A2(new_n4082_), .B(new_n4079_), .ZN(new_n4083_));
  NAND3_X1   g4034(.A1(new_n4081_), .A2(new_n4079_), .A3(new_n4082_), .ZN(new_n4084_));
  INV_X1     g4035(.I(new_n4084_), .ZN(new_n4085_));
  OAI21_X1   g4036(.A1(new_n4085_), .A2(new_n4083_), .B(new_n3932_), .ZN(new_n4086_));
  INV_X1     g4037(.I(new_n4082_), .ZN(new_n4087_));
  OAI21_X1   g4038(.A1(new_n4087_), .A2(new_n4080_), .B(new_n3792_), .ZN(new_n4088_));
  NAND3_X1   g4039(.A1(new_n4084_), .A2(new_n4088_), .A3(new_n3935_), .ZN(new_n4089_));
  NAND2_X1   g4040(.A1(new_n4086_), .A2(new_n4089_), .ZN(new_n4090_));
  NAND2_X1   g4041(.A1(new_n4090_), .A2(new_n4078_), .ZN(new_n4091_));
  INV_X1     g4042(.I(new_n4078_), .ZN(new_n4092_));
  AND2_X2    g4043(.A1(new_n4086_), .A2(new_n4089_), .Z(new_n4093_));
  NAND2_X1   g4044(.A1(new_n4093_), .A2(new_n4092_), .ZN(new_n4094_));
  AOI21_X1   g4045(.A1(new_n4094_), .A2(new_n4091_), .B(new_n3939_), .ZN(new_n4095_));
  INV_X1     g4046(.I(new_n3939_), .ZN(new_n4096_));
  NAND2_X1   g4047(.A1(new_n4090_), .A2(new_n4092_), .ZN(new_n4097_));
  NAND2_X1   g4048(.A1(new_n4093_), .A2(new_n4078_), .ZN(new_n4098_));
  AOI21_X1   g4049(.A1(new_n4098_), .A2(new_n4097_), .B(new_n4096_), .ZN(new_n4099_));
  NOR2_X1    g4050(.A1(new_n4099_), .A2(new_n4095_), .ZN(new_n4100_));
  INV_X1     g4051(.I(new_n4100_), .ZN(\sin[0] ));
  XOR2_X1    g4052(.A1(\a[22] ), .A2(\a[23] ), .Z(new_n4102_));
  NAND2_X1   g4053(.A1(\sin[0] ), .A2(new_n4102_), .ZN(new_n4103_));
  NAND2_X1   g4054(.A1(new_n4078_), .A2(new_n4096_), .ZN(new_n4104_));
  NAND2_X1   g4055(.A1(new_n4092_), .A2(new_n3939_), .ZN(new_n4105_));
  AOI21_X1   g4056(.A1(new_n4105_), .A2(new_n4104_), .B(new_n4090_), .ZN(new_n4106_));
  INV_X1     g4057(.I(new_n4106_), .ZN(new_n4107_));
  INV_X1     g4058(.I(new_n4074_), .ZN(new_n4108_));
  XOR2_X1    g4059(.A1(new_n4023_), .A2(new_n3895_), .Z(new_n4109_));
  NOR2_X1    g4060(.A1(new_n3895_), .A2(new_n3414_), .ZN(new_n4110_));
  NOR2_X1    g4061(.A1(new_n3894_), .A2(new_n3444_), .ZN(new_n4111_));
  OR3_X2     g4062(.A1(new_n4109_), .A2(new_n4110_), .A3(new_n4111_), .Z(new_n4112_));
  NAND3_X1   g4063(.A1(new_n3911_), .A2(new_n4112_), .A3(new_n3895_), .ZN(new_n4113_));
  NAND3_X1   g4064(.A1(new_n3903_), .A2(new_n3894_), .A3(new_n4112_), .ZN(new_n4114_));
  NAND2_X1   g4065(.A1(new_n4114_), .A2(new_n4113_), .ZN(new_n4115_));
  INV_X1     g4066(.I(new_n4115_), .ZN(new_n4116_));
  NOR4_X1    g4067(.A1(new_n311_), .A2(new_n525_), .A3(new_n747_), .A4(new_n488_), .ZN(new_n4117_));
  INV_X1     g4068(.I(new_n4117_), .ZN(new_n4118_));
  NOR2_X1    g4069(.A1(new_n2429_), .A2(new_n3773_), .ZN(new_n4119_));
  NAND4_X1   g4070(.A1(new_n4119_), .A2(new_n382_), .A3(new_n2395_), .A4(new_n4118_), .ZN(new_n4120_));
  INV_X1     g4071(.I(new_n4120_), .ZN(new_n4121_));
  NOR4_X1    g4072(.A1(new_n204_), .A2(new_n856_), .A3(new_n484_), .A4(new_n643_), .ZN(new_n4122_));
  NAND4_X1   g4073(.A1(new_n1077_), .A2(new_n329_), .A3(new_n330_), .A4(new_n918_), .ZN(new_n4123_));
  NOR4_X1    g4074(.A1(new_n766_), .A2(new_n1023_), .A3(new_n4122_), .A4(new_n4123_), .ZN(new_n4124_));
  NAND3_X1   g4075(.A1(new_n2385_), .A2(new_n4121_), .A3(new_n4124_), .ZN(new_n4125_));
  NOR2_X1    g4076(.A1(new_n4022_), .A2(new_n4125_), .ZN(new_n4126_));
  NAND2_X1   g4077(.A1(new_n4022_), .A2(new_n4125_), .ZN(new_n4127_));
  INV_X1     g4078(.I(new_n4127_), .ZN(new_n4128_));
  NOR2_X1    g4079(.A1(new_n4128_), .A2(new_n4126_), .ZN(new_n4129_));
  NOR2_X1    g4080(.A1(new_n4129_), .A2(new_n4028_), .ZN(new_n4130_));
  INV_X1     g4081(.I(new_n4129_), .ZN(new_n4131_));
  NOR2_X1    g4082(.A1(new_n4131_), .A2(new_n4023_), .ZN(new_n4132_));
  NOR2_X1    g4083(.A1(new_n4132_), .A2(new_n4130_), .ZN(new_n4133_));
  NOR2_X1    g4084(.A1(new_n4116_), .A2(new_n4133_), .ZN(new_n4134_));
  XOR2_X1    g4085(.A1(new_n4129_), .A2(new_n4023_), .Z(new_n4135_));
  NOR2_X1    g4086(.A1(new_n4115_), .A2(new_n4135_), .ZN(new_n4136_));
  OAI22_X1   g4087(.A1(new_n4023_), .A2(new_n3453_), .B1(new_n3451_), .B2(new_n3894_), .ZN(new_n4137_));
  NAND2_X1   g4088(.A1(new_n4131_), .A2(new_n3456_), .ZN(new_n4138_));
  AOI21_X1   g4089(.A1(new_n4138_), .A2(new_n4137_), .B(new_n3473_), .ZN(new_n4139_));
  OAI21_X1   g4090(.A1(new_n4134_), .A2(new_n4136_), .B(new_n4139_), .ZN(new_n4140_));
  XOR2_X1    g4091(.A1(new_n4140_), .A2(new_n2739_), .Z(new_n4141_));
  AOI21_X1   g4092(.A1(new_n2736_), .A2(new_n2722_), .B(new_n2779_), .ZN(new_n4142_));
  OAI22_X1   g4093(.A1(new_n2551_), .A2(new_n3007_), .B1(new_n2576_), .B2(new_n2774_), .ZN(new_n4143_));
  OAI21_X1   g4094(.A1(new_n2558_), .A2(new_n2767_), .B(new_n4143_), .ZN(new_n4144_));
  NOR2_X1    g4095(.A1(new_n4142_), .A2(new_n4144_), .ZN(new_n4145_));
  OAI22_X1   g4096(.A1(new_n2619_), .A2(new_n2850_), .B1(new_n2629_), .B2(new_n2882_), .ZN(new_n4146_));
  NAND2_X1   g4097(.A1(new_n2586_), .A2(new_n2855_), .ZN(new_n4147_));
  AOI21_X1   g4098(.A1(new_n4146_), .A2(new_n4147_), .B(new_n2881_), .ZN(new_n4148_));
  NAND3_X1   g4099(.A1(new_n2764_), .A2(new_n790_), .A3(new_n4148_), .ZN(new_n4149_));
  INV_X1     g4100(.I(new_n4149_), .ZN(new_n4150_));
  AOI21_X1   g4101(.A1(new_n2764_), .A2(new_n4148_), .B(new_n790_), .ZN(new_n4151_));
  NOR4_X1    g4102(.A1(new_n3963_), .A2(new_n659_), .A3(new_n2701_), .A4(new_n3965_), .ZN(new_n4152_));
  INV_X1     g4103(.I(new_n4152_), .ZN(new_n4153_));
  NAND2_X1   g4104(.A1(new_n3976_), .A2(new_n4153_), .ZN(new_n4154_));
  NAND2_X1   g4105(.A1(new_n3053_), .A2(new_n2824_), .ZN(new_n4155_));
  AOI22_X1   g4106(.A1(new_n2697_), .A2(new_n2795_), .B1(new_n2700_), .B2(new_n2829_), .ZN(new_n4156_));
  AOI21_X1   g4107(.A1(new_n2708_), .A2(new_n2790_), .B(new_n4156_), .ZN(new_n4157_));
  NAND2_X1   g4108(.A1(new_n4155_), .A2(new_n4157_), .ZN(new_n4158_));
  NOR2_X1    g4109(.A1(new_n2844_), .A2(new_n659_), .ZN(new_n4159_));
  XOR2_X1    g4110(.A1(new_n4158_), .A2(new_n4159_), .Z(new_n4160_));
  XOR2_X1    g4111(.A1(new_n4160_), .A2(new_n4154_), .Z(new_n4161_));
  NOR3_X1    g4112(.A1(new_n4150_), .A2(new_n4161_), .A3(new_n4151_), .ZN(new_n4162_));
  INV_X1     g4113(.I(new_n4162_), .ZN(new_n4163_));
  INV_X1     g4114(.I(new_n4151_), .ZN(new_n4164_));
  NAND2_X1   g4115(.A1(new_n4164_), .A2(new_n4149_), .ZN(new_n4165_));
  NAND2_X1   g4116(.A1(new_n4165_), .A2(new_n4161_), .ZN(new_n4166_));
  OR2_X2     g4117(.A1(new_n3972_), .A2(new_n3973_), .Z(new_n4167_));
  AOI22_X1   g4118(.A1(new_n3983_), .A2(new_n3981_), .B1(new_n3951_), .B2(new_n4167_), .ZN(new_n4168_));
  NAND3_X1   g4119(.A1(new_n4163_), .A2(new_n4166_), .A3(new_n4168_), .ZN(new_n4169_));
  XNOR2_X1   g4120(.A1(new_n4160_), .A2(new_n4154_), .ZN(new_n4170_));
  AOI21_X1   g4121(.A1(new_n4149_), .A2(new_n4164_), .B(new_n4170_), .ZN(new_n4171_));
  INV_X1     g4122(.I(new_n3981_), .ZN(new_n4172_));
  NAND2_X1   g4123(.A1(new_n3845_), .A2(new_n3843_), .ZN(new_n4173_));
  NAND2_X1   g4124(.A1(new_n4173_), .A2(new_n3841_), .ZN(new_n4174_));
  OAI21_X1   g4125(.A1(new_n4172_), .A2(new_n4174_), .B(new_n3974_), .ZN(new_n4175_));
  OAI21_X1   g4126(.A1(new_n4171_), .A2(new_n4162_), .B(new_n4175_), .ZN(new_n4176_));
  NAND3_X1   g4127(.A1(new_n4169_), .A2(new_n4176_), .A3(new_n1134_), .ZN(new_n4177_));
  NOR3_X1    g4128(.A1(new_n4171_), .A2(new_n4175_), .A3(new_n4162_), .ZN(new_n4178_));
  AOI21_X1   g4129(.A1(new_n4163_), .A2(new_n4166_), .B(new_n4168_), .ZN(new_n4179_));
  OAI21_X1   g4130(.A1(new_n4179_), .A2(new_n4178_), .B(new_n1132_), .ZN(new_n4180_));
  AOI21_X1   g4131(.A1(new_n4180_), .A2(new_n4177_), .B(new_n4145_), .ZN(new_n4181_));
  INV_X1     g4132(.I(new_n4145_), .ZN(new_n4182_));
  NOR3_X1    g4133(.A1(new_n4179_), .A2(new_n4178_), .A3(new_n1132_), .ZN(new_n4183_));
  AOI21_X1   g4134(.A1(new_n4169_), .A2(new_n4176_), .B(new_n1134_), .ZN(new_n4184_));
  NOR3_X1    g4135(.A1(new_n4183_), .A2(new_n4184_), .A3(new_n4182_), .ZN(new_n4185_));
  OAI21_X1   g4136(.A1(new_n3985_), .A2(new_n3986_), .B(new_n3946_), .ZN(new_n4186_));
  NOR3_X1    g4137(.A1(new_n4185_), .A2(new_n4181_), .A3(new_n4186_), .ZN(new_n4187_));
  OAI21_X1   g4138(.A1(new_n4183_), .A2(new_n4184_), .B(new_n4182_), .ZN(new_n4188_));
  NAND3_X1   g4139(.A1(new_n4180_), .A2(new_n4177_), .A3(new_n4145_), .ZN(new_n4189_));
  INV_X1     g4140(.I(new_n4186_), .ZN(new_n4190_));
  AOI21_X1   g4141(.A1(new_n4188_), .A2(new_n4189_), .B(new_n4190_), .ZN(new_n4191_));
  OAI22_X1   g4142(.A1(new_n3449_), .A2(new_n2752_), .B1(new_n2742_), .B2(new_n3419_), .ZN(new_n4192_));
  OAI21_X1   g4143(.A1(new_n2747_), .A2(new_n3444_), .B(new_n4192_), .ZN(new_n4193_));
  NAND2_X1   g4144(.A1(new_n4193_), .A2(new_n71_), .ZN(new_n4194_));
  NOR3_X1    g4145(.A1(new_n3448_), .A2(new_n943_), .A3(new_n4194_), .ZN(new_n4195_));
  INV_X1     g4146(.I(new_n4194_), .ZN(new_n4196_));
  AOI21_X1   g4147(.A1(new_n3464_), .A2(new_n4196_), .B(new_n62_), .ZN(new_n4197_));
  NOR4_X1    g4148(.A1(new_n4195_), .A2(new_n4197_), .A3(new_n4187_), .A4(new_n4191_), .ZN(new_n4198_));
  NAND3_X1   g4149(.A1(new_n4188_), .A2(new_n4189_), .A3(new_n4190_), .ZN(new_n4199_));
  OAI21_X1   g4150(.A1(new_n4185_), .A2(new_n4181_), .B(new_n4186_), .ZN(new_n4200_));
  NAND3_X1   g4151(.A1(new_n3464_), .A2(new_n62_), .A3(new_n4196_), .ZN(new_n4201_));
  OAI21_X1   g4152(.A1(new_n3448_), .A2(new_n4194_), .B(new_n943_), .ZN(new_n4202_));
  AOI22_X1   g4153(.A1(new_n4202_), .A2(new_n4201_), .B1(new_n4199_), .B2(new_n4200_), .ZN(new_n4203_));
  NOR3_X1    g4154(.A1(new_n4046_), .A2(new_n3367_), .A3(new_n3872_), .ZN(new_n4204_));
  OAI21_X1   g4155(.A1(new_n4204_), .A2(new_n4038_), .B(new_n3992_), .ZN(new_n4205_));
  NOR3_X1    g4156(.A1(new_n4198_), .A2(new_n4203_), .A3(new_n4205_), .ZN(new_n4206_));
  NAND4_X1   g4157(.A1(new_n4202_), .A2(new_n4201_), .A3(new_n4199_), .A4(new_n4200_), .ZN(new_n4207_));
  OAI22_X1   g4158(.A1(new_n4195_), .A2(new_n4197_), .B1(new_n4187_), .B2(new_n4191_), .ZN(new_n4208_));
  NOR2_X1    g4159(.A1(new_n4040_), .A2(new_n3991_), .ZN(new_n4209_));
  AOI21_X1   g4160(.A1(new_n4207_), .A2(new_n4208_), .B(new_n4209_), .ZN(new_n4210_));
  NOR3_X1    g4161(.A1(new_n4204_), .A2(new_n3992_), .A3(new_n4038_), .ZN(new_n4211_));
  NOR3_X1    g4162(.A1(new_n4209_), .A2(new_n4001_), .A3(new_n4211_), .ZN(new_n4212_));
  NOR3_X1    g4163(.A1(new_n4210_), .A2(new_n4212_), .A3(new_n4206_), .ZN(new_n4213_));
  NAND3_X1   g4164(.A1(new_n4209_), .A2(new_n4208_), .A3(new_n4207_), .ZN(new_n4214_));
  OAI21_X1   g4165(.A1(new_n4203_), .A2(new_n4198_), .B(new_n4205_), .ZN(new_n4215_));
  NAND2_X1   g4166(.A1(new_n4040_), .A2(new_n3991_), .ZN(new_n4216_));
  NAND3_X1   g4167(.A1(new_n4216_), .A2(new_n4004_), .A3(new_n4205_), .ZN(new_n4217_));
  AOI21_X1   g4168(.A1(new_n4214_), .A2(new_n4215_), .B(new_n4217_), .ZN(new_n4218_));
  NOR2_X1    g4169(.A1(new_n4213_), .A2(new_n4218_), .ZN(new_n4219_));
  XOR2_X1    g4170(.A1(new_n4219_), .A2(new_n4141_), .Z(new_n4220_));
  INV_X1     g4171(.I(new_n4220_), .ZN(new_n4221_));
  NOR2_X1    g4172(.A1(new_n1089_), .A2(new_n488_), .ZN(new_n4222_));
  NAND4_X1   g4173(.A1(new_n728_), .A2(new_n1698_), .A3(new_n4222_), .A4(new_n554_), .ZN(new_n4223_));
  INV_X1     g4174(.I(new_n3375_), .ZN(new_n4224_));
  INV_X1     g4175(.I(new_n2314_), .ZN(new_n4225_));
  NAND4_X1   g4176(.A1(new_n4225_), .A2(new_n223_), .A3(new_n837_), .A4(new_n820_), .ZN(new_n4226_));
  NAND4_X1   g4177(.A1(new_n727_), .A2(new_n310_), .A3(new_n547_), .A4(new_n343_), .ZN(new_n4227_));
  NAND4_X1   g4178(.A1(new_n4224_), .A2(new_n3383_), .A3(new_n4226_), .A4(new_n4227_), .ZN(new_n4228_));
  OR4_X2     g4179(.A1(new_n2470_), .A2(new_n3777_), .A3(new_n4223_), .A4(new_n4228_), .Z(new_n4229_));
  OAI21_X1   g4180(.A1(new_n3882_), .A2(new_n3883_), .B(new_n3881_), .ZN(new_n4230_));
  NAND3_X1   g4181(.A1(new_n3877_), .A2(new_n3812_), .A3(new_n3873_), .ZN(new_n4231_));
  NAND3_X1   g4182(.A1(new_n3926_), .A2(new_n69_), .A3(new_n3920_), .ZN(new_n4232_));
  NAND2_X1   g4183(.A1(new_n3921_), .A2(new_n2739_), .ZN(new_n4233_));
  AOI22_X1   g4184(.A1(new_n4230_), .A2(new_n4231_), .B1(new_n4232_), .B2(new_n4233_), .ZN(new_n4234_));
  OAI21_X1   g4185(.A1(new_n3801_), .A2(new_n3795_), .B(new_n4234_), .ZN(new_n4235_));
  NAND3_X1   g4186(.A1(new_n4054_), .A2(new_n4060_), .A3(new_n4235_), .ZN(new_n4236_));
  NOR2_X1    g4187(.A1(new_n3886_), .A2(new_n3930_), .ZN(new_n4237_));
  NAND2_X1   g4188(.A1(new_n4236_), .A2(new_n4237_), .ZN(new_n4238_));
  OAI21_X1   g4189(.A1(new_n4033_), .A2(new_n4036_), .B(new_n2739_), .ZN(new_n4239_));
  NAND2_X1   g4190(.A1(new_n4050_), .A2(new_n69_), .ZN(new_n4240_));
  NAND2_X1   g4191(.A1(new_n4240_), .A2(new_n4239_), .ZN(new_n4241_));
  NAND2_X1   g4192(.A1(new_n4057_), .A2(new_n4047_), .ZN(new_n4242_));
  NAND2_X1   g4193(.A1(new_n4006_), .A2(new_n4040_), .ZN(new_n4243_));
  NAND2_X1   g4194(.A1(new_n4243_), .A2(new_n4242_), .ZN(new_n4244_));
  NAND2_X1   g4195(.A1(new_n4244_), .A2(new_n4241_), .ZN(new_n4245_));
  NAND2_X1   g4196(.A1(new_n4238_), .A2(new_n4245_), .ZN(new_n4246_));
  XOR2_X1    g4197(.A1(new_n4246_), .A2(new_n4229_), .Z(new_n4247_));
  NOR2_X1    g4198(.A1(new_n4247_), .A2(new_n4221_), .ZN(new_n4248_));
  AND2_X2    g4199(.A1(new_n4247_), .A2(new_n4221_), .Z(new_n4249_));
  OR2_X2     g4200(.A1(new_n4249_), .A2(new_n4248_), .Z(new_n4250_));
  NOR3_X1    g4201(.A1(new_n3938_), .A2(new_n3793_), .A3(new_n4074_), .ZN(new_n4251_));
  NOR2_X1    g4202(.A1(new_n3939_), .A2(new_n4108_), .ZN(new_n4252_));
  OAI21_X1   g4203(.A1(new_n4252_), .A2(new_n4251_), .B(new_n4070_), .ZN(new_n4253_));
  NOR2_X1    g4204(.A1(new_n4250_), .A2(new_n4253_), .ZN(new_n4254_));
  INV_X1     g4205(.I(new_n4254_), .ZN(new_n4255_));
  NAND2_X1   g4206(.A1(new_n4250_), .A2(new_n4253_), .ZN(new_n4256_));
  NAND4_X1   g4207(.A1(new_n4255_), .A2(new_n4256_), .A3(new_n4096_), .A4(new_n4108_), .ZN(new_n4257_));
  INV_X1     g4208(.I(new_n4256_), .ZN(new_n4258_));
  NAND2_X1   g4209(.A1(new_n4096_), .A2(new_n4108_), .ZN(new_n4259_));
  OAI21_X1   g4210(.A1(new_n4258_), .A2(new_n4254_), .B(new_n4259_), .ZN(new_n4260_));
  NAND2_X1   g4211(.A1(new_n4257_), .A2(new_n4260_), .ZN(new_n4261_));
  XOR2_X1    g4212(.A1(new_n4261_), .A2(new_n4107_), .Z(new_n4262_));
  XOR2_X1    g4213(.A1(new_n4262_), .A2(new_n4103_), .Z(\sin[1] ));
  AOI21_X1   g4214(.A1(new_n4257_), .A2(new_n4260_), .B(new_n4107_), .ZN(new_n4264_));
  NOR3_X1    g4215(.A1(new_n4213_), .A2(new_n4218_), .A3(new_n4141_), .ZN(new_n4265_));
  AOI22_X1   g4216(.A1(new_n4243_), .A2(new_n4242_), .B1(new_n4239_), .B2(new_n4240_), .ZN(new_n4266_));
  OAI21_X1   g4217(.A1(new_n4213_), .A2(new_n4218_), .B(new_n4141_), .ZN(new_n4267_));
  XOR2_X1    g4218(.A1(new_n4140_), .A2(new_n69_), .Z(new_n4268_));
  NAND3_X1   g4219(.A1(new_n4214_), .A2(new_n4215_), .A3(new_n4217_), .ZN(new_n4269_));
  NAND2_X1   g4220(.A1(new_n4208_), .A2(new_n4207_), .ZN(new_n4270_));
  NAND4_X1   g4221(.A1(new_n4270_), .A2(new_n4004_), .A3(new_n4205_), .A4(new_n4216_), .ZN(new_n4271_));
  NAND3_X1   g4222(.A1(new_n4269_), .A2(new_n4268_), .A3(new_n4271_), .ZN(new_n4272_));
  AOI21_X1   g4223(.A1(new_n4267_), .A2(new_n4272_), .B(new_n4266_), .ZN(new_n4273_));
  AOI21_X1   g4224(.A1(new_n4238_), .A2(new_n4273_), .B(new_n4265_), .ZN(new_n4274_));
  OAI22_X1   g4225(.A1(new_n2551_), .A2(new_n2767_), .B1(new_n2558_), .B2(new_n2774_), .ZN(new_n4275_));
  NAND2_X1   g4226(.A1(new_n3418_), .A2(new_n2776_), .ZN(new_n4276_));
  AOI21_X1   g4227(.A1(new_n4276_), .A2(new_n4275_), .B(new_n2779_), .ZN(new_n4277_));
  OAI21_X1   g4228(.A1(new_n3809_), .A2(new_n3807_), .B(new_n4277_), .ZN(new_n4278_));
  XOR2_X1    g4229(.A1(new_n4278_), .A2(new_n1134_), .Z(new_n4279_));
  OAI22_X1   g4230(.A1(new_n2576_), .A2(new_n2856_), .B1(new_n2619_), .B2(new_n2882_), .ZN(new_n4280_));
  NAND2_X1   g4231(.A1(new_n2586_), .A2(new_n2851_), .ZN(new_n4281_));
  AOI21_X1   g4232(.A1(new_n4280_), .A2(new_n4281_), .B(new_n2881_), .ZN(new_n4282_));
  NAND3_X1   g4233(.A1(new_n3330_), .A2(new_n790_), .A3(new_n4282_), .ZN(new_n4283_));
  INV_X1     g4234(.I(new_n4283_), .ZN(new_n4284_));
  AOI21_X1   g4235(.A1(new_n3330_), .A2(new_n4282_), .B(new_n790_), .ZN(new_n4285_));
  NOR2_X1    g4236(.A1(new_n4284_), .A2(new_n4285_), .ZN(new_n4286_));
  INV_X1     g4237(.I(new_n4159_), .ZN(new_n4287_));
  NAND2_X1   g4238(.A1(new_n4154_), .A2(new_n4287_), .ZN(new_n4288_));
  INV_X1     g4239(.I(new_n4288_), .ZN(new_n4289_));
  OAI21_X1   g4240(.A1(new_n3837_), .A2(new_n3833_), .B(new_n658_), .ZN(new_n4290_));
  NAND3_X1   g4241(.A1(new_n3952_), .A2(new_n3954_), .A3(new_n659_), .ZN(new_n4291_));
  AOI21_X1   g4242(.A1(new_n4290_), .A2(new_n4291_), .B(new_n2673_), .ZN(new_n4292_));
  NOR4_X1    g4243(.A1(new_n4292_), .A2(new_n3955_), .A3(new_n3978_), .A4(new_n3957_), .ZN(new_n4293_));
  OAI21_X1   g4244(.A1(new_n4293_), .A2(new_n4152_), .B(new_n4287_), .ZN(new_n4294_));
  NAND3_X1   g4245(.A1(new_n3976_), .A2(new_n4153_), .A3(new_n4159_), .ZN(new_n4295_));
  AOI21_X1   g4246(.A1(new_n4294_), .A2(new_n4295_), .B(new_n659_), .ZN(new_n4296_));
  AOI21_X1   g4247(.A1(new_n3976_), .A2(new_n4153_), .B(new_n4159_), .ZN(new_n4297_));
  NOR3_X1    g4248(.A1(new_n4293_), .A2(new_n4152_), .A3(new_n4287_), .ZN(new_n4298_));
  NOR3_X1    g4249(.A1(new_n4298_), .A2(new_n4297_), .A3(new_n658_), .ZN(new_n4299_));
  OAI21_X1   g4250(.A1(new_n4299_), .A2(new_n4296_), .B(new_n4158_), .ZN(new_n4300_));
  NOR2_X1    g4251(.A1(new_n4300_), .A2(new_n4289_), .ZN(new_n4301_));
  OAI21_X1   g4252(.A1(new_n4298_), .A2(new_n4297_), .B(new_n658_), .ZN(new_n4302_));
  NAND3_X1   g4253(.A1(new_n4294_), .A2(new_n4295_), .A3(new_n659_), .ZN(new_n4303_));
  NAND2_X1   g4254(.A1(new_n4302_), .A2(new_n4303_), .ZN(new_n4304_));
  AOI21_X1   g4255(.A1(new_n4304_), .A2(new_n4158_), .B(new_n4288_), .ZN(new_n4305_));
  AOI22_X1   g4256(.A1(new_n2708_), .A2(new_n2795_), .B1(new_n2697_), .B2(new_n2829_), .ZN(new_n4306_));
  AOI21_X1   g4257(.A1(new_n2628_), .A2(new_n2790_), .B(new_n4306_), .ZN(new_n4307_));
  OAI21_X1   g4258(.A1(new_n3049_), .A2(new_n2796_), .B(new_n4307_), .ZN(new_n4308_));
  NOR2_X1    g4259(.A1(new_n2700_), .A2(new_n659_), .ZN(new_n4309_));
  INV_X1     g4260(.I(new_n4309_), .ZN(new_n4310_));
  XOR2_X1    g4261(.A1(new_n4308_), .A2(new_n4310_), .Z(new_n4311_));
  NOR3_X1    g4262(.A1(new_n4301_), .A2(new_n4305_), .A3(new_n4311_), .ZN(new_n4312_));
  NAND3_X1   g4263(.A1(new_n4304_), .A2(new_n4158_), .A3(new_n4288_), .ZN(new_n4313_));
  NAND2_X1   g4264(.A1(new_n4300_), .A2(new_n4289_), .ZN(new_n4314_));
  INV_X1     g4265(.I(new_n4311_), .ZN(new_n4315_));
  AOI21_X1   g4266(.A1(new_n4314_), .A2(new_n4313_), .B(new_n4315_), .ZN(new_n4316_));
  OAI21_X1   g4267(.A1(new_n4312_), .A2(new_n4316_), .B(new_n4286_), .ZN(new_n4317_));
  INV_X1     g4268(.I(new_n4285_), .ZN(new_n4318_));
  NAND2_X1   g4269(.A1(new_n4318_), .A2(new_n4283_), .ZN(new_n4319_));
  NAND3_X1   g4270(.A1(new_n4314_), .A2(new_n4313_), .A3(new_n4315_), .ZN(new_n4320_));
  OAI21_X1   g4271(.A1(new_n4301_), .A2(new_n4305_), .B(new_n4311_), .ZN(new_n4321_));
  NAND3_X1   g4272(.A1(new_n4319_), .A2(new_n4321_), .A3(new_n4320_), .ZN(new_n4322_));
  NAND2_X1   g4273(.A1(new_n4175_), .A2(new_n4170_), .ZN(new_n4323_));
  NAND2_X1   g4274(.A1(new_n4168_), .A2(new_n4161_), .ZN(new_n4324_));
  AOI21_X1   g4275(.A1(new_n4323_), .A2(new_n4324_), .B(new_n4165_), .ZN(new_n4325_));
  NAND3_X1   g4276(.A1(new_n4317_), .A2(new_n4325_), .A3(new_n4322_), .ZN(new_n4326_));
  AOI21_X1   g4277(.A1(new_n4320_), .A2(new_n4321_), .B(new_n4319_), .ZN(new_n4327_));
  NOR3_X1    g4278(.A1(new_n4286_), .A2(new_n4312_), .A3(new_n4316_), .ZN(new_n4328_));
  INV_X1     g4279(.I(new_n4165_), .ZN(new_n4329_));
  NOR2_X1    g4280(.A1(new_n4168_), .A2(new_n4161_), .ZN(new_n4330_));
  NOR2_X1    g4281(.A1(new_n4175_), .A2(new_n4170_), .ZN(new_n4331_));
  OAI21_X1   g4282(.A1(new_n4331_), .A2(new_n4330_), .B(new_n4329_), .ZN(new_n4332_));
  OAI21_X1   g4283(.A1(new_n4327_), .A2(new_n4328_), .B(new_n4332_), .ZN(new_n4333_));
  NOR2_X1    g4284(.A1(new_n4175_), .A2(new_n4161_), .ZN(new_n4334_));
  NAND3_X1   g4285(.A1(new_n4333_), .A2(new_n4326_), .A3(new_n4334_), .ZN(new_n4335_));
  NOR3_X1    g4286(.A1(new_n4327_), .A2(new_n4332_), .A3(new_n4328_), .ZN(new_n4336_));
  AOI21_X1   g4287(.A1(new_n4317_), .A2(new_n4322_), .B(new_n4325_), .ZN(new_n4337_));
  INV_X1     g4288(.I(new_n4334_), .ZN(new_n4338_));
  OAI21_X1   g4289(.A1(new_n4337_), .A2(new_n4336_), .B(new_n4338_), .ZN(new_n4339_));
  NAND2_X1   g4290(.A1(new_n4339_), .A2(new_n4335_), .ZN(new_n4340_));
  NAND2_X1   g4291(.A1(new_n4145_), .A2(new_n1132_), .ZN(new_n4341_));
  NAND2_X1   g4292(.A1(new_n4182_), .A2(new_n1134_), .ZN(new_n4342_));
  NAND2_X1   g4293(.A1(new_n4342_), .A2(new_n4341_), .ZN(new_n4343_));
  NAND3_X1   g4294(.A1(new_n4343_), .A2(new_n4169_), .A3(new_n4176_), .ZN(new_n4344_));
  NAND4_X1   g4295(.A1(new_n4344_), .A2(new_n4188_), .A3(new_n4189_), .A4(new_n4186_), .ZN(new_n4345_));
  XOR2_X1    g4296(.A1(new_n4340_), .A2(new_n4345_), .Z(new_n4346_));
  NAND2_X1   g4297(.A1(new_n4346_), .A2(new_n4279_), .ZN(new_n4347_));
  NAND3_X1   g4298(.A1(new_n3472_), .A2(new_n1132_), .A3(new_n4277_), .ZN(new_n4348_));
  NAND2_X1   g4299(.A1(new_n4278_), .A2(new_n1134_), .ZN(new_n4349_));
  NAND2_X1   g4300(.A1(new_n4349_), .A2(new_n4348_), .ZN(new_n4350_));
  NOR3_X1    g4301(.A1(new_n4337_), .A2(new_n4336_), .A3(new_n4338_), .ZN(new_n4351_));
  AOI21_X1   g4302(.A1(new_n4333_), .A2(new_n4326_), .B(new_n4334_), .ZN(new_n4352_));
  NOR2_X1    g4303(.A1(new_n4351_), .A2(new_n4352_), .ZN(new_n4353_));
  XOR2_X1    g4304(.A1(new_n4353_), .A2(new_n4345_), .Z(new_n4354_));
  NAND2_X1   g4305(.A1(new_n4354_), .A2(new_n4350_), .ZN(new_n4355_));
  OAI22_X1   g4306(.A1(new_n3449_), .A2(new_n2742_), .B1(new_n3444_), .B2(new_n2752_), .ZN(new_n4356_));
  NAND2_X1   g4307(.A1(new_n3895_), .A2(new_n2748_), .ZN(new_n4357_));
  AOI21_X1   g4308(.A1(new_n4357_), .A2(new_n4356_), .B(new_n72_), .ZN(new_n4358_));
  NAND2_X1   g4309(.A1(new_n3926_), .A2(new_n4358_), .ZN(new_n4359_));
  XOR2_X1    g4310(.A1(new_n4359_), .A2(new_n943_), .Z(new_n4360_));
  NAND3_X1   g4311(.A1(new_n4360_), .A2(new_n4347_), .A3(new_n4355_), .ZN(new_n4361_));
  NAND2_X1   g4312(.A1(new_n4347_), .A2(new_n4355_), .ZN(new_n4362_));
  INV_X1     g4313(.I(new_n4360_), .ZN(new_n4363_));
  NAND2_X1   g4314(.A1(new_n4362_), .A2(new_n4363_), .ZN(new_n4364_));
  NOR2_X1    g4315(.A1(new_n4056_), .A2(new_n4040_), .ZN(new_n4365_));
  NOR2_X1    g4316(.A1(new_n4270_), .A2(new_n4365_), .ZN(new_n4366_));
  OAI21_X1   g4317(.A1(new_n4366_), .A2(new_n4055_), .B(new_n4208_), .ZN(new_n4367_));
  NAND3_X1   g4318(.A1(new_n4364_), .A2(new_n4361_), .A3(new_n4367_), .ZN(new_n4368_));
  INV_X1     g4319(.I(new_n4361_), .ZN(new_n4369_));
  AOI21_X1   g4320(.A1(new_n4347_), .A2(new_n4355_), .B(new_n4360_), .ZN(new_n4370_));
  INV_X1     g4321(.I(new_n4367_), .ZN(new_n4371_));
  OAI21_X1   g4322(.A1(new_n4369_), .A2(new_n4370_), .B(new_n4371_), .ZN(new_n4372_));
  NAND2_X1   g4323(.A1(new_n4372_), .A2(new_n4368_), .ZN(new_n4373_));
  NAND2_X1   g4324(.A1(new_n4116_), .A2(new_n4132_), .ZN(new_n4374_));
  NAND2_X1   g4325(.A1(new_n4115_), .A2(new_n4130_), .ZN(new_n4375_));
  NAND2_X1   g4326(.A1(new_n4374_), .A2(new_n4375_), .ZN(new_n4376_));
  OAI21_X1   g4327(.A1(new_n4023_), .A2(new_n3451_), .B(new_n3459_), .ZN(new_n4377_));
  AOI21_X1   g4328(.A1(new_n4131_), .A2(new_n3487_), .B(new_n4377_), .ZN(new_n4378_));
  AND3_X2    g4329(.A1(new_n4376_), .A2(new_n69_), .A3(new_n4378_), .Z(new_n4379_));
  AOI21_X1   g4330(.A1(new_n4376_), .A2(new_n4378_), .B(new_n69_), .ZN(new_n4380_));
  NOR2_X1    g4331(.A1(new_n4379_), .A2(new_n4380_), .ZN(new_n4381_));
  INV_X1     g4332(.I(new_n4381_), .ZN(new_n4382_));
  XOR2_X1    g4333(.A1(new_n4373_), .A2(new_n4382_), .Z(new_n4383_));
  NOR2_X1    g4334(.A1(new_n4383_), .A2(new_n4274_), .ZN(new_n4384_));
  OAI22_X1   g4335(.A1(new_n3461_), .A2(new_n3466_), .B1(new_n3368_), .B2(new_n3359_), .ZN(new_n4385_));
  NAND4_X1   g4336(.A1(new_n3677_), .A2(new_n3683_), .A3(new_n4385_), .A4(new_n3686_), .ZN(new_n4386_));
  OAI22_X1   g4337(.A1(new_n3884_), .A2(new_n3878_), .B1(new_n3927_), .B2(new_n3922_), .ZN(new_n4387_));
  AOI21_X1   g4338(.A1(new_n4386_), .A2(new_n3794_), .B(new_n4387_), .ZN(new_n4388_));
  NOR3_X1    g4339(.A1(new_n4063_), .A2(new_n4062_), .A3(new_n4388_), .ZN(new_n4389_));
  INV_X1     g4340(.I(new_n4237_), .ZN(new_n4390_));
  NOR2_X1    g4341(.A1(new_n4389_), .A2(new_n4390_), .ZN(new_n4391_));
  INV_X1     g4342(.I(new_n4265_), .ZN(new_n4392_));
  AOI21_X1   g4343(.A1(new_n4269_), .A2(new_n4271_), .B(new_n4268_), .ZN(new_n4393_));
  NOR3_X1    g4344(.A1(new_n4213_), .A2(new_n4218_), .A3(new_n4141_), .ZN(new_n4394_));
  OAI21_X1   g4345(.A1(new_n4394_), .A2(new_n4393_), .B(new_n4245_), .ZN(new_n4395_));
  OAI21_X1   g4346(.A1(new_n4391_), .A2(new_n4395_), .B(new_n4392_), .ZN(new_n4396_));
  XOR2_X1    g4347(.A1(new_n4373_), .A2(new_n4381_), .Z(new_n4397_));
  NOR2_X1    g4348(.A1(new_n4397_), .A2(new_n4396_), .ZN(new_n4398_));
  NOR2_X1    g4349(.A1(new_n4384_), .A2(new_n4398_), .ZN(new_n4399_));
  INV_X1     g4350(.I(new_n4399_), .ZN(new_n4400_));
  NOR2_X1    g4351(.A1(new_n435_), .A2(new_n584_), .ZN(new_n4401_));
  NOR2_X1    g4352(.A1(new_n377_), .A2(new_n501_), .ZN(new_n4402_));
  NAND4_X1   g4353(.A1(new_n4401_), .A2(new_n4402_), .A3(new_n275_), .A4(new_n4014_), .ZN(new_n4403_));
  NOR4_X1    g4354(.A1(new_n2393_), .A2(new_n361_), .A3(new_n507_), .A4(new_n520_), .ZN(new_n4404_));
  INV_X1     g4355(.I(new_n4404_), .ZN(new_n4405_));
  NOR4_X1    g4356(.A1(new_n326_), .A2(new_n339_), .A3(new_n238_), .A4(new_n856_), .ZN(new_n4406_));
  NOR4_X1    g4357(.A1(new_n4405_), .A2(new_n531_), .A3(new_n4403_), .A4(new_n4406_), .ZN(new_n4407_));
  INV_X1     g4358(.I(new_n4407_), .ZN(new_n4408_));
  NOR3_X1    g4359(.A1(new_n4408_), .A2(new_n761_), .A3(new_n3734_), .ZN(new_n4409_));
  INV_X1     g4360(.I(new_n4409_), .ZN(new_n4410_));
  NOR4_X1    g4361(.A1(new_n4249_), .A2(new_n4248_), .A3(new_n3939_), .A4(new_n4074_), .ZN(new_n4411_));
  NOR2_X1    g4362(.A1(new_n4246_), .A2(new_n4220_), .ZN(new_n4412_));
  NAND2_X1   g4363(.A1(new_n4246_), .A2(new_n4220_), .ZN(new_n4413_));
  NAND2_X1   g4364(.A1(new_n4413_), .A2(new_n4229_), .ZN(new_n4414_));
  NOR2_X1    g4365(.A1(new_n4414_), .A2(new_n4412_), .ZN(new_n4415_));
  OAI21_X1   g4366(.A1(new_n4411_), .A2(new_n4253_), .B(new_n4415_), .ZN(new_n4416_));
  NAND2_X1   g4367(.A1(new_n4416_), .A2(new_n4410_), .ZN(new_n4417_));
  NOR2_X1    g4368(.A1(new_n4416_), .A2(new_n4410_), .ZN(new_n4418_));
  INV_X1     g4369(.I(new_n4418_), .ZN(new_n4419_));
  AOI21_X1   g4370(.A1(new_n4419_), .A2(new_n4417_), .B(new_n4400_), .ZN(new_n4420_));
  INV_X1     g4371(.I(new_n4420_), .ZN(new_n4421_));
  NAND3_X1   g4372(.A1(new_n4419_), .A2(new_n4400_), .A3(new_n4417_), .ZN(new_n4422_));
  NAND2_X1   g4373(.A1(new_n4421_), .A2(new_n4422_), .ZN(new_n4423_));
  NOR3_X1    g4374(.A1(new_n4258_), .A2(new_n4254_), .A3(new_n4259_), .ZN(new_n4424_));
  AOI22_X1   g4375(.A1(new_n4255_), .A2(new_n4256_), .B1(new_n4096_), .B2(new_n4108_), .ZN(new_n4425_));
  NOR3_X1    g4376(.A1(new_n4425_), .A2(new_n4424_), .A3(new_n4106_), .ZN(new_n4426_));
  OAI21_X1   g4377(.A1(new_n4426_), .A2(new_n4264_), .B(new_n4100_), .ZN(new_n4427_));
  NAND2_X1   g4378(.A1(new_n4427_), .A2(new_n4102_), .ZN(new_n4428_));
  XOR2_X1    g4379(.A1(new_n4428_), .A2(new_n4423_), .Z(new_n4429_));
  XOR2_X1    g4380(.A1(new_n4429_), .A2(new_n4264_), .Z(\sin[2] ));
  OAI21_X1   g4381(.A1(new_n4425_), .A2(new_n4424_), .B(new_n4106_), .ZN(new_n4431_));
  INV_X1     g4382(.I(new_n4417_), .ZN(new_n4432_));
  NOR3_X1    g4383(.A1(new_n4432_), .A2(new_n4399_), .A3(new_n4418_), .ZN(new_n4433_));
  NOR3_X1    g4384(.A1(new_n4431_), .A2(new_n4433_), .A3(new_n4420_), .ZN(new_n4434_));
  NOR2_X1    g4385(.A1(new_n4411_), .A2(new_n4253_), .ZN(new_n4435_));
  XOR2_X1    g4386(.A1(new_n4399_), .A2(new_n4410_), .Z(new_n4436_));
  NAND2_X1   g4387(.A1(new_n4436_), .A2(new_n4415_), .ZN(new_n4437_));
  OAI22_X1   g4388(.A1(new_n4437_), .A2(new_n4435_), .B1(new_n4399_), .B2(new_n4409_), .ZN(new_n4438_));
  AOI21_X1   g4389(.A1(new_n4115_), .A2(new_n4023_), .B(new_n4129_), .ZN(new_n4439_));
  AOI22_X1   g4390(.A1(new_n4439_), .A2(new_n3459_), .B1(new_n3450_), .B2(new_n4131_), .ZN(new_n4440_));
  AOI22_X1   g4391(.A1(new_n2577_), .A2(new_n2851_), .B1(new_n2586_), .B2(new_n2848_), .ZN(new_n4441_));
  AOI21_X1   g4392(.A1(new_n2559_), .A2(new_n2855_), .B(new_n4441_), .ZN(new_n4442_));
  OR3_X2     g4393(.A1(new_n3940_), .A2(new_n2881_), .A3(new_n4442_), .Z(new_n4443_));
  XOR2_X1    g4394(.A1(new_n4443_), .A2(new_n576_), .Z(new_n4444_));
  NOR2_X1    g4395(.A1(new_n2697_), .A2(new_n659_), .ZN(new_n4445_));
  NOR3_X1    g4396(.A1(new_n4301_), .A2(new_n4305_), .A3(new_n4309_), .ZN(new_n4446_));
  INV_X1     g4397(.I(new_n4446_), .ZN(new_n4447_));
  NOR3_X1    g4398(.A1(new_n4301_), .A2(new_n4305_), .A3(new_n4309_), .ZN(new_n4448_));
  AOI21_X1   g4399(.A1(new_n4314_), .A2(new_n4313_), .B(new_n4310_), .ZN(new_n4449_));
  OAI21_X1   g4400(.A1(new_n4448_), .A2(new_n4449_), .B(new_n658_), .ZN(new_n4450_));
  NAND3_X1   g4401(.A1(new_n4314_), .A2(new_n4313_), .A3(new_n4310_), .ZN(new_n4451_));
  OAI21_X1   g4402(.A1(new_n4301_), .A2(new_n4305_), .B(new_n4309_), .ZN(new_n4452_));
  NAND3_X1   g4403(.A1(new_n4452_), .A2(new_n4451_), .A3(new_n659_), .ZN(new_n4453_));
  NAND2_X1   g4404(.A1(new_n4450_), .A2(new_n4453_), .ZN(new_n4454_));
  NAND3_X1   g4405(.A1(new_n4454_), .A2(new_n4308_), .A3(new_n4447_), .ZN(new_n4455_));
  AOI21_X1   g4406(.A1(new_n4452_), .A2(new_n4451_), .B(new_n659_), .ZN(new_n4456_));
  NOR3_X1    g4407(.A1(new_n4448_), .A2(new_n4449_), .A3(new_n658_), .ZN(new_n4457_));
  OAI21_X1   g4408(.A1(new_n4457_), .A2(new_n4456_), .B(new_n4308_), .ZN(new_n4458_));
  NAND2_X1   g4409(.A1(new_n4458_), .A2(new_n4446_), .ZN(new_n4459_));
  AND2_X2    g4410(.A1(new_n3014_), .A2(new_n2824_), .Z(new_n4460_));
  OAI22_X1   g4411(.A1(new_n2619_), .A2(new_n2791_), .B1(new_n2696_), .B2(new_n2830_), .ZN(new_n4461_));
  OAI21_X1   g4412(.A1(new_n2629_), .A2(new_n2794_), .B(new_n4461_), .ZN(new_n4462_));
  NOR2_X1    g4413(.A1(new_n4460_), .A2(new_n4462_), .ZN(new_n4463_));
  NAND3_X1   g4414(.A1(new_n4459_), .A2(new_n4455_), .A3(new_n4463_), .ZN(new_n4464_));
  NOR2_X1    g4415(.A1(new_n4458_), .A2(new_n4446_), .ZN(new_n4465_));
  AOI21_X1   g4416(.A1(new_n4454_), .A2(new_n4308_), .B(new_n4447_), .ZN(new_n4466_));
  INV_X1     g4417(.I(new_n4463_), .ZN(new_n4467_));
  OAI21_X1   g4418(.A1(new_n4465_), .A2(new_n4466_), .B(new_n4467_), .ZN(new_n4468_));
  AOI21_X1   g4419(.A1(new_n4468_), .A2(new_n4464_), .B(new_n4445_), .ZN(new_n4469_));
  INV_X1     g4420(.I(new_n4445_), .ZN(new_n4470_));
  NOR3_X1    g4421(.A1(new_n4465_), .A2(new_n4466_), .A3(new_n4467_), .ZN(new_n4471_));
  AOI21_X1   g4422(.A1(new_n4459_), .A2(new_n4455_), .B(new_n4463_), .ZN(new_n4472_));
  NOR3_X1    g4423(.A1(new_n4471_), .A2(new_n4472_), .A3(new_n4470_), .ZN(new_n4473_));
  NAND2_X1   g4424(.A1(new_n4165_), .A2(new_n4161_), .ZN(new_n4474_));
  NAND3_X1   g4425(.A1(new_n4317_), .A2(new_n4322_), .A3(new_n4474_), .ZN(new_n4475_));
  INV_X1     g4426(.I(new_n4475_), .ZN(new_n4476_));
  NOR3_X1    g4427(.A1(new_n4473_), .A2(new_n4469_), .A3(new_n4476_), .ZN(new_n4477_));
  OAI21_X1   g4428(.A1(new_n4471_), .A2(new_n4472_), .B(new_n4470_), .ZN(new_n4478_));
  NAND3_X1   g4429(.A1(new_n4468_), .A2(new_n4464_), .A3(new_n4445_), .ZN(new_n4479_));
  AOI21_X1   g4430(.A1(new_n4478_), .A2(new_n4479_), .B(new_n4475_), .ZN(new_n4480_));
  OAI21_X1   g4431(.A1(new_n4477_), .A2(new_n4480_), .B(new_n4444_), .ZN(new_n4481_));
  INV_X1     g4432(.I(new_n4444_), .ZN(new_n4482_));
  NAND3_X1   g4433(.A1(new_n4478_), .A2(new_n4479_), .A3(new_n4475_), .ZN(new_n4483_));
  OAI21_X1   g4434(.A1(new_n4473_), .A2(new_n4469_), .B(new_n4476_), .ZN(new_n4484_));
  NAND3_X1   g4435(.A1(new_n4484_), .A2(new_n4483_), .A3(new_n4482_), .ZN(new_n4485_));
  OAI22_X1   g4436(.A1(new_n3419_), .A2(new_n2767_), .B1(new_n2551_), .B2(new_n2774_), .ZN(new_n4486_));
  NAND2_X1   g4437(.A1(new_n3668_), .A2(new_n2776_), .ZN(new_n4487_));
  AOI21_X1   g4438(.A1(new_n4487_), .A2(new_n4486_), .B(new_n2779_), .ZN(new_n4488_));
  NAND2_X1   g4439(.A1(new_n3994_), .A2(new_n4488_), .ZN(new_n4489_));
  XOR2_X1    g4440(.A1(new_n4489_), .A2(new_n1134_), .Z(new_n4490_));
  INV_X1     g4441(.I(new_n4490_), .ZN(new_n4491_));
  NAND3_X1   g4442(.A1(new_n4481_), .A2(new_n4485_), .A3(new_n4491_), .ZN(new_n4492_));
  AOI21_X1   g4443(.A1(new_n4484_), .A2(new_n4483_), .B(new_n4482_), .ZN(new_n4493_));
  NOR3_X1    g4444(.A1(new_n4477_), .A2(new_n4480_), .A3(new_n4444_), .ZN(new_n4494_));
  OAI21_X1   g4445(.A1(new_n4494_), .A2(new_n4493_), .B(new_n4490_), .ZN(new_n4495_));
  NAND2_X1   g4446(.A1(new_n4169_), .A2(new_n4176_), .ZN(new_n4496_));
  AOI21_X1   g4447(.A1(new_n4341_), .A2(new_n4342_), .B(new_n4496_), .ZN(new_n4497_));
  NOR4_X1    g4448(.A1(new_n4181_), .A2(new_n4185_), .A3(new_n4497_), .A4(new_n4190_), .ZN(new_n4498_));
  AOI21_X1   g4449(.A1(new_n4339_), .A2(new_n4335_), .B(new_n4350_), .ZN(new_n4499_));
  NOR3_X1    g4450(.A1(new_n4279_), .A2(new_n4351_), .A3(new_n4352_), .ZN(new_n4500_));
  OAI22_X1   g4451(.A1(new_n4500_), .A2(new_n4499_), .B1(new_n4353_), .B2(new_n4498_), .ZN(new_n4501_));
  NAND2_X1   g4452(.A1(new_n4032_), .A2(new_n4027_), .ZN(new_n4502_));
  AOI22_X1   g4453(.A1(new_n3895_), .A2(new_n2753_), .B1(new_n2741_), .B2(new_n3414_), .ZN(new_n4503_));
  AOI21_X1   g4454(.A1(new_n2748_), .A2(new_n4028_), .B(new_n4503_), .ZN(new_n4504_));
  NOR2_X1    g4455(.A1(new_n4504_), .A2(new_n72_), .ZN(new_n4505_));
  NAND3_X1   g4456(.A1(new_n4502_), .A2(new_n62_), .A3(new_n4505_), .ZN(new_n4506_));
  NOR3_X1    g4457(.A1(new_n3916_), .A2(new_n4031_), .A3(new_n4028_), .ZN(new_n4507_));
  AOI21_X1   g4458(.A1(new_n4009_), .A2(new_n4026_), .B(new_n4023_), .ZN(new_n4508_));
  OAI21_X1   g4459(.A1(new_n4507_), .A2(new_n4508_), .B(new_n4505_), .ZN(new_n4509_));
  NAND2_X1   g4460(.A1(new_n4509_), .A2(new_n943_), .ZN(new_n4510_));
  AOI21_X1   g4461(.A1(new_n4506_), .A2(new_n4510_), .B(new_n4501_), .ZN(new_n4511_));
  OAI21_X1   g4462(.A1(new_n4351_), .A2(new_n4352_), .B(new_n4279_), .ZN(new_n4512_));
  NAND3_X1   g4463(.A1(new_n4339_), .A2(new_n4335_), .A3(new_n4350_), .ZN(new_n4513_));
  AOI22_X1   g4464(.A1(new_n4512_), .A2(new_n4513_), .B1(new_n4340_), .B2(new_n4345_), .ZN(new_n4514_));
  NOR2_X1    g4465(.A1(new_n4509_), .A2(new_n943_), .ZN(new_n4515_));
  AOI21_X1   g4466(.A1(new_n4502_), .A2(new_n4505_), .B(new_n62_), .ZN(new_n4516_));
  NOR3_X1    g4467(.A1(new_n4514_), .A2(new_n4515_), .A3(new_n4516_), .ZN(new_n4517_));
  NOR2_X1    g4468(.A1(new_n4511_), .A2(new_n4517_), .ZN(new_n4518_));
  AOI21_X1   g4469(.A1(new_n4495_), .A2(new_n4492_), .B(new_n4518_), .ZN(new_n4519_));
  NOR3_X1    g4470(.A1(new_n4494_), .A2(new_n4493_), .A3(new_n4490_), .ZN(new_n4520_));
  AOI21_X1   g4471(.A1(new_n4481_), .A2(new_n4485_), .B(new_n4491_), .ZN(new_n4521_));
  AOI21_X1   g4472(.A1(new_n4506_), .A2(new_n4510_), .B(new_n4514_), .ZN(new_n4522_));
  NOR3_X1    g4473(.A1(new_n4501_), .A2(new_n4515_), .A3(new_n4516_), .ZN(new_n4523_));
  NOR2_X1    g4474(.A1(new_n4522_), .A2(new_n4523_), .ZN(new_n4524_));
  NOR3_X1    g4475(.A1(new_n4520_), .A2(new_n4521_), .A3(new_n4524_), .ZN(new_n4525_));
  OAI21_X1   g4476(.A1(new_n4525_), .A2(new_n4519_), .B(new_n2739_), .ZN(new_n4526_));
  OAI21_X1   g4477(.A1(new_n4515_), .A2(new_n4516_), .B(new_n4514_), .ZN(new_n4527_));
  NAND3_X1   g4478(.A1(new_n4501_), .A2(new_n4510_), .A3(new_n4506_), .ZN(new_n4528_));
  NAND2_X1   g4479(.A1(new_n4527_), .A2(new_n4528_), .ZN(new_n4529_));
  OAI21_X1   g4480(.A1(new_n4520_), .A2(new_n4521_), .B(new_n4529_), .ZN(new_n4530_));
  OAI21_X1   g4481(.A1(new_n4515_), .A2(new_n4516_), .B(new_n4501_), .ZN(new_n4531_));
  NAND3_X1   g4482(.A1(new_n4514_), .A2(new_n4510_), .A3(new_n4506_), .ZN(new_n4532_));
  NAND2_X1   g4483(.A1(new_n4531_), .A2(new_n4532_), .ZN(new_n4533_));
  NAND3_X1   g4484(.A1(new_n4495_), .A2(new_n4492_), .A3(new_n4533_), .ZN(new_n4534_));
  NAND3_X1   g4485(.A1(new_n4530_), .A2(new_n4534_), .A3(new_n69_), .ZN(new_n4535_));
  AOI21_X1   g4486(.A1(new_n4526_), .A2(new_n4535_), .B(new_n4440_), .ZN(new_n4536_));
  INV_X1     g4487(.I(new_n4440_), .ZN(new_n4537_));
  NAND3_X1   g4488(.A1(new_n4530_), .A2(new_n4534_), .A3(new_n2739_), .ZN(new_n4538_));
  OAI21_X1   g4489(.A1(new_n4525_), .A2(new_n4519_), .B(new_n69_), .ZN(new_n4539_));
  AOI21_X1   g4490(.A1(new_n4539_), .A2(new_n4538_), .B(new_n4537_), .ZN(new_n4540_));
  NOR3_X1    g4491(.A1(new_n4369_), .A2(new_n4371_), .A3(new_n4370_), .ZN(new_n4541_));
  NOR2_X1    g4492(.A1(new_n4541_), .A2(new_n4370_), .ZN(new_n4542_));
  NOR3_X1    g4493(.A1(new_n4536_), .A2(new_n4540_), .A3(new_n4542_), .ZN(new_n4543_));
  AOI21_X1   g4494(.A1(new_n4530_), .A2(new_n4534_), .B(new_n69_), .ZN(new_n4544_));
  NOR3_X1    g4495(.A1(new_n4525_), .A2(new_n4519_), .A3(new_n2739_), .ZN(new_n4545_));
  OAI21_X1   g4496(.A1(new_n4545_), .A2(new_n4544_), .B(new_n4537_), .ZN(new_n4546_));
  NOR3_X1    g4497(.A1(new_n4525_), .A2(new_n4519_), .A3(new_n69_), .ZN(new_n4547_));
  AOI21_X1   g4498(.A1(new_n4530_), .A2(new_n4534_), .B(new_n2739_), .ZN(new_n4548_));
  OAI21_X1   g4499(.A1(new_n4547_), .A2(new_n4548_), .B(new_n4440_), .ZN(new_n4549_));
  NAND2_X1   g4500(.A1(new_n4368_), .A2(new_n4364_), .ZN(new_n4550_));
  AOI21_X1   g4501(.A1(new_n4546_), .A2(new_n4549_), .B(new_n4550_), .ZN(new_n4551_));
  AOI21_X1   g4502(.A1(new_n4364_), .A2(new_n4361_), .B(new_n4367_), .ZN(new_n4552_));
  NOR2_X1    g4503(.A1(new_n4541_), .A2(new_n4552_), .ZN(new_n4553_));
  NOR2_X1    g4504(.A1(new_n4274_), .A2(new_n4553_), .ZN(new_n4554_));
  INV_X1     g4505(.I(new_n4554_), .ZN(new_n4555_));
  NOR3_X1    g4506(.A1(new_n4551_), .A2(new_n4543_), .A3(new_n4555_), .ZN(new_n4556_));
  NAND3_X1   g4507(.A1(new_n4546_), .A2(new_n4549_), .A3(new_n4550_), .ZN(new_n4557_));
  OAI21_X1   g4508(.A1(new_n4536_), .A2(new_n4540_), .B(new_n4542_), .ZN(new_n4558_));
  AOI21_X1   g4509(.A1(new_n4557_), .A2(new_n4558_), .B(new_n4554_), .ZN(new_n4559_));
  XOR2_X1    g4510(.A1(new_n4274_), .A2(new_n4553_), .Z(new_n4560_));
  NAND2_X1   g4511(.A1(new_n4560_), .A2(new_n4382_), .ZN(new_n4561_));
  NOR3_X1    g4512(.A1(new_n4561_), .A2(new_n4556_), .A3(new_n4559_), .ZN(new_n4562_));
  NOR2_X1    g4513(.A1(new_n4556_), .A2(new_n4559_), .ZN(new_n4563_));
  AOI21_X1   g4514(.A1(new_n4382_), .A2(new_n4560_), .B(new_n4563_), .ZN(new_n4564_));
  NAND3_X1   g4515(.A1(new_n749_), .A2(new_n182_), .A3(new_n3752_), .ZN(new_n4565_));
  NOR3_X1    g4516(.A1(new_n615_), .A2(new_n300_), .A3(new_n974_), .ZN(new_n4566_));
  INV_X1     g4517(.I(new_n4566_), .ZN(new_n4567_));
  NOR4_X1    g4518(.A1(new_n3738_), .A2(new_n801_), .A3(new_n198_), .A4(new_n261_), .ZN(new_n4568_));
  NOR4_X1    g4519(.A1(new_n4567_), .A2(new_n823_), .A3(new_n1699_), .A4(new_n4568_), .ZN(new_n4569_));
  INV_X1     g4520(.I(new_n4569_), .ZN(new_n4570_));
  NOR4_X1    g4521(.A1(new_n4570_), .A2(new_n1014_), .A3(new_n2473_), .A4(new_n4565_), .ZN(new_n4571_));
  INV_X1     g4522(.I(new_n4571_), .ZN(new_n4572_));
  NOR3_X1    g4523(.A1(new_n4564_), .A2(new_n4562_), .A3(new_n4572_), .ZN(new_n4573_));
  OAI21_X1   g4524(.A1(new_n4564_), .A2(new_n4562_), .B(new_n4572_), .ZN(new_n4574_));
  INV_X1     g4525(.I(new_n4574_), .ZN(new_n4575_));
  NOR2_X1    g4526(.A1(new_n4575_), .A2(new_n4573_), .ZN(new_n4576_));
  NOR2_X1    g4527(.A1(new_n4438_), .A2(new_n4576_), .ZN(new_n4577_));
  INV_X1     g4528(.I(new_n4577_), .ZN(new_n4578_));
  NAND2_X1   g4529(.A1(new_n4438_), .A2(new_n4576_), .ZN(new_n4579_));
  AOI21_X1   g4530(.A1(new_n4579_), .A2(new_n4578_), .B(new_n4434_), .ZN(new_n4580_));
  NAND3_X1   g4531(.A1(new_n4421_), .A2(new_n4264_), .A3(new_n4422_), .ZN(new_n4581_));
  INV_X1     g4532(.I(new_n4579_), .ZN(new_n4582_));
  NOR3_X1    g4533(.A1(new_n4581_), .A2(new_n4577_), .A3(new_n4582_), .ZN(new_n4583_));
  NOR2_X1    g4534(.A1(new_n4583_), .A2(new_n4580_), .ZN(new_n4584_));
  INV_X1     g4535(.I(new_n4102_), .ZN(new_n4585_));
  OAI21_X1   g4536(.A1(new_n4420_), .A2(new_n4433_), .B(new_n4431_), .ZN(new_n4586_));
  AOI21_X1   g4537(.A1(new_n4581_), .A2(new_n4586_), .B(new_n4427_), .ZN(new_n4587_));
  NOR2_X1    g4538(.A1(new_n4587_), .A2(new_n4585_), .ZN(new_n4588_));
  XOR2_X1    g4539(.A1(new_n4588_), .A2(new_n4584_), .Z(\sin[3] ));
  OAI21_X1   g4540(.A1(new_n4577_), .A2(new_n4582_), .B(new_n4434_), .ZN(new_n4590_));
  OAI21_X1   g4541(.A1(new_n4520_), .A2(new_n4521_), .B(new_n4501_), .ZN(new_n4591_));
  NAND3_X1   g4542(.A1(new_n4495_), .A2(new_n4492_), .A3(new_n4514_), .ZN(new_n4592_));
  NAND2_X1   g4543(.A1(new_n4591_), .A2(new_n4592_), .ZN(new_n4593_));
  INV_X1     g4544(.I(new_n4593_), .ZN(new_n4594_));
  NOR2_X1    g4545(.A1(new_n4515_), .A2(new_n4516_), .ZN(new_n4595_));
  XNOR2_X1   g4546(.A1(new_n4593_), .A2(new_n4595_), .ZN(new_n4596_));
  XOR2_X1    g4547(.A1(new_n4440_), .A2(new_n69_), .Z(new_n4597_));
  OAI21_X1   g4548(.A1(new_n4594_), .A2(new_n4597_), .B(new_n4596_), .ZN(new_n4598_));
  AOI21_X1   g4549(.A1(new_n4495_), .A2(new_n4514_), .B(new_n4520_), .ZN(new_n4599_));
  INV_X1     g4550(.I(new_n4599_), .ZN(new_n4600_));
  OAI22_X1   g4551(.A1(new_n4023_), .A2(new_n2752_), .B1(new_n2742_), .B2(new_n3894_), .ZN(new_n4601_));
  NAND2_X1   g4552(.A1(new_n4131_), .A2(new_n2748_), .ZN(new_n4602_));
  AOI21_X1   g4553(.A1(new_n4602_), .A2(new_n4601_), .B(new_n72_), .ZN(new_n4603_));
  OAI21_X1   g4554(.A1(new_n4134_), .A2(new_n4136_), .B(new_n4603_), .ZN(new_n4604_));
  XOR2_X1    g4555(.A1(new_n4604_), .A2(new_n943_), .Z(new_n4605_));
  INV_X1     g4556(.I(new_n4605_), .ZN(new_n4606_));
  OAI22_X1   g4557(.A1(new_n2551_), .A2(new_n2856_), .B1(new_n2576_), .B2(new_n2882_), .ZN(new_n4607_));
  NAND2_X1   g4558(.A1(new_n2559_), .A2(new_n2851_), .ZN(new_n4608_));
  AOI21_X1   g4559(.A1(new_n4607_), .A2(new_n4608_), .B(new_n2881_), .ZN(new_n4609_));
  NAND2_X1   g4560(.A1(new_n3653_), .A2(new_n4609_), .ZN(new_n4610_));
  XOR2_X1    g4561(.A1(new_n4610_), .A2(new_n576_), .Z(new_n4611_));
  OAI22_X1   g4562(.A1(new_n2619_), .A2(new_n2794_), .B1(new_n2629_), .B2(new_n2830_), .ZN(new_n4612_));
  NAND2_X1   g4563(.A1(new_n2586_), .A2(new_n2790_), .ZN(new_n4613_));
  AOI21_X1   g4564(.A1(new_n4612_), .A2(new_n4613_), .B(new_n2796_), .ZN(new_n4614_));
  NAND2_X1   g4565(.A1(new_n2764_), .A2(new_n4614_), .ZN(new_n4615_));
  XOR2_X1    g4566(.A1(new_n4615_), .A2(new_n658_), .Z(new_n4616_));
  NOR2_X1    g4567(.A1(new_n2696_), .A2(new_n659_), .ZN(new_n4617_));
  XOR2_X1    g4568(.A1(new_n4617_), .A2(new_n2739_), .Z(new_n4618_));
  XOR2_X1    g4569(.A1(new_n4616_), .A2(new_n4618_), .Z(new_n4619_));
  OAI22_X1   g4570(.A1(new_n4471_), .A2(new_n4472_), .B1(new_n659_), .B2(new_n4467_), .ZN(new_n4620_));
  OAI21_X1   g4571(.A1(new_n4471_), .A2(new_n4472_), .B(new_n658_), .ZN(new_n4621_));
  NAND3_X1   g4572(.A1(new_n4468_), .A2(new_n4464_), .A3(new_n659_), .ZN(new_n4622_));
  NAND2_X1   g4573(.A1(new_n4621_), .A2(new_n4622_), .ZN(new_n4623_));
  NOR4_X1    g4574(.A1(new_n4471_), .A2(new_n4472_), .A3(new_n658_), .A4(new_n4467_), .ZN(new_n4624_));
  AOI21_X1   g4575(.A1(new_n4623_), .A2(new_n2697_), .B(new_n4624_), .ZN(new_n4625_));
  NAND2_X1   g4576(.A1(new_n4625_), .A2(new_n4620_), .ZN(new_n4626_));
  NAND2_X1   g4577(.A1(new_n4626_), .A2(new_n4619_), .ZN(new_n4627_));
  INV_X1     g4578(.I(new_n4619_), .ZN(new_n4628_));
  NAND3_X1   g4579(.A1(new_n4625_), .A2(new_n4628_), .A3(new_n4620_), .ZN(new_n4629_));
  AOI21_X1   g4580(.A1(new_n4627_), .A2(new_n4629_), .B(new_n4611_), .ZN(new_n4630_));
  INV_X1     g4581(.I(new_n4611_), .ZN(new_n4631_));
  NAND2_X1   g4582(.A1(new_n4626_), .A2(new_n4628_), .ZN(new_n4632_));
  NAND3_X1   g4583(.A1(new_n4625_), .A2(new_n4619_), .A3(new_n4620_), .ZN(new_n4633_));
  AOI21_X1   g4584(.A1(new_n4632_), .A2(new_n4633_), .B(new_n4631_), .ZN(new_n4634_));
  OAI22_X1   g4585(.A1(new_n3449_), .A2(new_n2767_), .B1(new_n2774_), .B2(new_n3419_), .ZN(new_n4635_));
  NAND2_X1   g4586(.A1(new_n3414_), .A2(new_n2776_), .ZN(new_n4636_));
  AOI21_X1   g4587(.A1(new_n4635_), .A2(new_n4636_), .B(new_n2779_), .ZN(new_n4637_));
  NAND2_X1   g4588(.A1(new_n3464_), .A2(new_n4637_), .ZN(new_n4638_));
  XOR2_X1    g4589(.A1(new_n4638_), .A2(new_n1134_), .Z(new_n4639_));
  INV_X1     g4590(.I(new_n4639_), .ZN(new_n4640_));
  OAI21_X1   g4591(.A1(new_n4630_), .A2(new_n4634_), .B(new_n4640_), .ZN(new_n4641_));
  NOR3_X1    g4592(.A1(new_n4630_), .A2(new_n4634_), .A3(new_n4640_), .ZN(new_n4642_));
  INV_X1     g4593(.I(new_n4642_), .ZN(new_n4643_));
  AOI21_X1   g4594(.A1(new_n4643_), .A2(new_n4641_), .B(new_n4606_), .ZN(new_n4644_));
  INV_X1     g4595(.I(new_n4641_), .ZN(new_n4645_));
  NOR3_X1    g4596(.A1(new_n4645_), .A2(new_n4605_), .A3(new_n4642_), .ZN(new_n4646_));
  OAI21_X1   g4597(.A1(new_n4646_), .A2(new_n4644_), .B(new_n4600_), .ZN(new_n4647_));
  AOI21_X1   g4598(.A1(new_n4643_), .A2(new_n4641_), .B(new_n4605_), .ZN(new_n4648_));
  NOR3_X1    g4599(.A1(new_n4645_), .A2(new_n4606_), .A3(new_n4642_), .ZN(new_n4649_));
  OAI21_X1   g4600(.A1(new_n4649_), .A2(new_n4648_), .B(new_n4599_), .ZN(new_n4650_));
  NAND2_X1   g4601(.A1(new_n4647_), .A2(new_n4650_), .ZN(new_n4651_));
  XOR2_X1    g4602(.A1(new_n4651_), .A2(new_n4598_), .Z(new_n4652_));
  NAND4_X1   g4603(.A1(new_n564_), .A2(new_n2380_), .A3(new_n291_), .A4(new_n639_), .ZN(new_n4653_));
  NOR2_X1    g4604(.A1(new_n2518_), .A2(new_n461_), .ZN(new_n4654_));
  NAND4_X1   g4605(.A1(new_n4654_), .A2(new_n275_), .A3(new_n350_), .A4(new_n950_), .ZN(new_n4655_));
  NOR3_X1    g4606(.A1(new_n1087_), .A2(new_n4655_), .A3(new_n4653_), .ZN(new_n4656_));
  NAND3_X1   g4607(.A1(new_n2321_), .A2(new_n723_), .A3(new_n4656_), .ZN(new_n4657_));
  INV_X1     g4608(.I(new_n4657_), .ZN(new_n4658_));
  OAI21_X1   g4609(.A1(new_n4396_), .A2(new_n4373_), .B(new_n4382_), .ZN(new_n4659_));
  NOR3_X1    g4610(.A1(new_n4551_), .A2(new_n4543_), .A3(new_n4659_), .ZN(new_n4660_));
  OAI21_X1   g4611(.A1(new_n4536_), .A2(new_n4540_), .B(new_n4550_), .ZN(new_n4661_));
  OAI21_X1   g4612(.A1(new_n4660_), .A2(new_n4555_), .B(new_n4661_), .ZN(new_n4662_));
  XOR2_X1    g4613(.A1(new_n4662_), .A2(new_n4658_), .Z(new_n4663_));
  XOR2_X1    g4614(.A1(new_n4663_), .A2(new_n4652_), .Z(new_n4664_));
  OAI21_X1   g4615(.A1(new_n4438_), .A2(new_n4573_), .B(new_n4574_), .ZN(new_n4665_));
  XOR2_X1    g4616(.A1(new_n4665_), .A2(new_n4664_), .Z(new_n4666_));
  XOR2_X1    g4617(.A1(new_n4666_), .A2(new_n4590_), .Z(new_n4667_));
  OAI21_X1   g4618(.A1(new_n4580_), .A2(new_n4583_), .B(new_n4587_), .ZN(new_n4668_));
  NAND2_X1   g4619(.A1(new_n4668_), .A2(new_n4102_), .ZN(new_n4669_));
  XNOR2_X1   g4620(.A1(new_n4669_), .A2(new_n4667_), .ZN(\sin[4] ));
  NOR2_X1    g4621(.A1(new_n4666_), .A2(new_n4590_), .ZN(new_n4671_));
  INV_X1     g4622(.I(new_n4671_), .ZN(new_n4672_));
  INV_X1     g4623(.I(new_n4598_), .ZN(new_n4673_));
  OAI21_X1   g4624(.A1(new_n4645_), .A2(new_n4642_), .B(new_n4605_), .ZN(new_n4674_));
  NAND3_X1   g4625(.A1(new_n4643_), .A2(new_n4606_), .A3(new_n4641_), .ZN(new_n4675_));
  AOI21_X1   g4626(.A1(new_n4674_), .A2(new_n4675_), .B(new_n4599_), .ZN(new_n4676_));
  OAI21_X1   g4627(.A1(new_n4645_), .A2(new_n4642_), .B(new_n4606_), .ZN(new_n4677_));
  NAND3_X1   g4628(.A1(new_n4643_), .A2(new_n4605_), .A3(new_n4641_), .ZN(new_n4678_));
  AOI21_X1   g4629(.A1(new_n4677_), .A2(new_n4678_), .B(new_n4600_), .ZN(new_n4679_));
  NOR2_X1    g4630(.A1(new_n4676_), .A2(new_n4679_), .ZN(new_n4680_));
  NAND2_X1   g4631(.A1(new_n4662_), .A2(new_n4680_), .ZN(new_n4681_));
  AOI21_X1   g4632(.A1(new_n4274_), .A2(new_n4553_), .B(new_n4381_), .ZN(new_n4682_));
  NAND3_X1   g4633(.A1(new_n4557_), .A2(new_n4558_), .A3(new_n4682_), .ZN(new_n4683_));
  NAND2_X1   g4634(.A1(new_n4683_), .A2(new_n4554_), .ZN(new_n4684_));
  NAND3_X1   g4635(.A1(new_n4684_), .A2(new_n4651_), .A3(new_n4661_), .ZN(new_n4685_));
  AOI22_X1   g4636(.A1(new_n4681_), .A2(new_n4685_), .B1(new_n4673_), .B2(new_n4662_), .ZN(new_n4686_));
  AOI21_X1   g4637(.A1(new_n4600_), .A2(new_n4677_), .B(new_n4649_), .ZN(new_n4687_));
  NAND2_X1   g4638(.A1(new_n4131_), .A2(new_n2753_), .ZN(new_n4688_));
  NAND2_X1   g4639(.A1(new_n4028_), .A2(new_n2741_), .ZN(new_n4689_));
  NAND4_X1   g4640(.A1(new_n4376_), .A2(new_n71_), .A3(new_n4688_), .A4(new_n4689_), .ZN(new_n4690_));
  XOR2_X1    g4641(.A1(new_n4690_), .A2(new_n943_), .Z(new_n4691_));
  OAI22_X1   g4642(.A1(new_n2576_), .A2(new_n2791_), .B1(new_n2619_), .B2(new_n2830_), .ZN(new_n4692_));
  NAND2_X1   g4643(.A1(new_n2586_), .A2(new_n2795_), .ZN(new_n4693_));
  AOI21_X1   g4644(.A1(new_n4692_), .A2(new_n4693_), .B(new_n2796_), .ZN(new_n4694_));
  NAND2_X1   g4645(.A1(new_n3330_), .A2(new_n4694_), .ZN(new_n4695_));
  XOR2_X1    g4646(.A1(new_n4695_), .A2(new_n659_), .Z(new_n4696_));
  INV_X1     g4647(.I(new_n4696_), .ZN(new_n4697_));
  NOR2_X1    g4648(.A1(new_n2629_), .A2(new_n659_), .ZN(new_n4698_));
  NAND2_X1   g4649(.A1(new_n658_), .A2(new_n69_), .ZN(new_n4699_));
  OAI22_X1   g4650(.A1(new_n4698_), .A2(new_n69_), .B1(new_n2629_), .B2(new_n4699_), .ZN(new_n4700_));
  OAI22_X1   g4651(.A1(new_n2551_), .A2(new_n2850_), .B1(new_n2558_), .B2(new_n2882_), .ZN(new_n4701_));
  NAND2_X1   g4652(.A1(new_n3418_), .A2(new_n2855_), .ZN(new_n4702_));
  AOI21_X1   g4653(.A1(new_n4702_), .A2(new_n4701_), .B(new_n2881_), .ZN(new_n4703_));
  NAND2_X1   g4654(.A1(new_n3472_), .A2(new_n4703_), .ZN(new_n4704_));
  XOR2_X1    g4655(.A1(new_n4704_), .A2(new_n576_), .Z(new_n4705_));
  NOR2_X1    g4656(.A1(new_n4616_), .A2(new_n2739_), .ZN(new_n4706_));
  INV_X1     g4657(.I(new_n4617_), .ZN(new_n4707_));
  AOI21_X1   g4658(.A1(new_n4616_), .A2(new_n2739_), .B(new_n4707_), .ZN(new_n4708_));
  NOR2_X1    g4659(.A1(new_n4708_), .A2(new_n4706_), .ZN(new_n4709_));
  XOR2_X1    g4660(.A1(new_n4705_), .A2(new_n4709_), .Z(new_n4710_));
  NOR2_X1    g4661(.A1(new_n4710_), .A2(new_n4700_), .ZN(new_n4711_));
  INV_X1     g4662(.I(new_n4711_), .ZN(new_n4712_));
  NAND2_X1   g4663(.A1(new_n4710_), .A2(new_n4700_), .ZN(new_n4713_));
  AOI21_X1   g4664(.A1(new_n4712_), .A2(new_n4713_), .B(new_n4697_), .ZN(new_n4714_));
  INV_X1     g4665(.I(new_n4713_), .ZN(new_n4715_));
  NOR3_X1    g4666(.A1(new_n4715_), .A2(new_n4696_), .A3(new_n4711_), .ZN(new_n4716_));
  NOR2_X1    g4667(.A1(new_n4714_), .A2(new_n4716_), .ZN(new_n4717_));
  INV_X1     g4668(.I(new_n3926_), .ZN(new_n4718_));
  NOR2_X1    g4669(.A1(new_n4718_), .A2(new_n2779_), .ZN(new_n4719_));
  OAI22_X1   g4670(.A1(new_n2774_), .A2(new_n3449_), .B1(new_n3444_), .B2(new_n2767_), .ZN(new_n4720_));
  OAI21_X1   g4671(.A1(new_n3007_), .A2(new_n3894_), .B(new_n4720_), .ZN(new_n4721_));
  NOR2_X1    g4672(.A1(new_n4719_), .A2(new_n4721_), .ZN(new_n4722_));
  INV_X1     g4673(.I(new_n4722_), .ZN(new_n4723_));
  NAND2_X1   g4674(.A1(new_n4633_), .A2(new_n4611_), .ZN(new_n4724_));
  NAND2_X1   g4675(.A1(new_n4724_), .A2(new_n4632_), .ZN(new_n4725_));
  NAND2_X1   g4676(.A1(new_n4725_), .A2(new_n4723_), .ZN(new_n4726_));
  NOR2_X1    g4677(.A1(new_n4725_), .A2(new_n4723_), .ZN(new_n4727_));
  INV_X1     g4678(.I(new_n4727_), .ZN(new_n4728_));
  AOI21_X1   g4679(.A1(new_n4728_), .A2(new_n4726_), .B(new_n1134_), .ZN(new_n4729_));
  INV_X1     g4680(.I(new_n4726_), .ZN(new_n4730_));
  NOR3_X1    g4681(.A1(new_n4730_), .A2(new_n1132_), .A3(new_n4727_), .ZN(new_n4731_));
  OAI21_X1   g4682(.A1(new_n4729_), .A2(new_n4731_), .B(new_n4717_), .ZN(new_n4732_));
  INV_X1     g4683(.I(new_n4717_), .ZN(new_n4733_));
  OAI21_X1   g4684(.A1(new_n4730_), .A2(new_n4727_), .B(new_n1132_), .ZN(new_n4734_));
  NAND3_X1   g4685(.A1(new_n4728_), .A2(new_n1134_), .A3(new_n4726_), .ZN(new_n4735_));
  NAND3_X1   g4686(.A1(new_n4734_), .A2(new_n4735_), .A3(new_n4733_), .ZN(new_n4736_));
  NAND2_X1   g4687(.A1(new_n4732_), .A2(new_n4736_), .ZN(new_n4737_));
  NAND2_X1   g4688(.A1(new_n4737_), .A2(new_n4641_), .ZN(new_n4738_));
  NAND3_X1   g4689(.A1(new_n4732_), .A2(new_n4736_), .A3(new_n4645_), .ZN(new_n4739_));
  AOI21_X1   g4690(.A1(new_n4738_), .A2(new_n4739_), .B(new_n4691_), .ZN(new_n4740_));
  INV_X1     g4691(.I(new_n4691_), .ZN(new_n4741_));
  NAND2_X1   g4692(.A1(new_n4737_), .A2(new_n4645_), .ZN(new_n4742_));
  NAND3_X1   g4693(.A1(new_n4732_), .A2(new_n4736_), .A3(new_n4641_), .ZN(new_n4743_));
  AOI21_X1   g4694(.A1(new_n4742_), .A2(new_n4743_), .B(new_n4741_), .ZN(new_n4744_));
  NOR2_X1    g4695(.A1(new_n4740_), .A2(new_n4744_), .ZN(new_n4745_));
  NAND2_X1   g4696(.A1(new_n4745_), .A2(new_n4687_), .ZN(new_n4746_));
  INV_X1     g4697(.I(new_n4746_), .ZN(new_n4747_));
  NOR2_X1    g4698(.A1(new_n4745_), .A2(new_n4687_), .ZN(new_n4748_));
  NOR3_X1    g4699(.A1(new_n3738_), .A2(new_n399_), .A3(new_n434_), .ZN(new_n4749_));
  NAND4_X1   g4700(.A1(new_n449_), .A2(new_n893_), .A3(new_n445_), .A4(new_n344_), .ZN(new_n4750_));
  NAND3_X1   g4701(.A1(new_n4749_), .A2(new_n4226_), .A3(new_n4750_), .ZN(new_n4751_));
  NAND4_X1   g4702(.A1(new_n193_), .A2(new_n598_), .A3(new_n768_), .A4(new_n968_), .ZN(new_n4752_));
  NOR3_X1    g4703(.A1(new_n4751_), .A2(new_n1691_), .A3(new_n4752_), .ZN(new_n4753_));
  NAND3_X1   g4704(.A1(new_n3380_), .A2(new_n4121_), .A3(new_n4753_), .ZN(new_n4754_));
  INV_X1     g4705(.I(new_n4754_), .ZN(new_n4755_));
  OAI21_X1   g4706(.A1(new_n4747_), .A2(new_n4748_), .B(new_n4755_), .ZN(new_n4756_));
  INV_X1     g4707(.I(new_n4748_), .ZN(new_n4757_));
  NAND3_X1   g4708(.A1(new_n4757_), .A2(new_n4746_), .A3(new_n4754_), .ZN(new_n4758_));
  NAND2_X1   g4709(.A1(new_n4756_), .A2(new_n4758_), .ZN(new_n4759_));
  NOR3_X1    g4710(.A1(new_n4747_), .A2(new_n4748_), .A3(new_n4754_), .ZN(new_n4760_));
  AOI21_X1   g4711(.A1(new_n4757_), .A2(new_n4746_), .B(new_n4755_), .ZN(new_n4761_));
  NOR2_X1    g4712(.A1(new_n4761_), .A2(new_n4760_), .ZN(new_n4762_));
  NOR2_X1    g4713(.A1(new_n4762_), .A2(new_n4686_), .ZN(new_n4763_));
  AOI21_X1   g4714(.A1(new_n4686_), .A2(new_n4759_), .B(new_n4763_), .ZN(new_n4764_));
  XNOR2_X1   g4715(.A1(new_n4652_), .A2(new_n4662_), .ZN(new_n4765_));
  OAI22_X1   g4716(.A1(new_n4665_), .A2(new_n4664_), .B1(new_n4658_), .B2(new_n4765_), .ZN(new_n4766_));
  NAND2_X1   g4717(.A1(new_n4764_), .A2(new_n4766_), .ZN(new_n4767_));
  NAND2_X1   g4718(.A1(new_n4759_), .A2(new_n4686_), .ZN(new_n4768_));
  OAI21_X1   g4719(.A1(new_n4686_), .A2(new_n4762_), .B(new_n4768_), .ZN(new_n4769_));
  INV_X1     g4720(.I(new_n4766_), .ZN(new_n4770_));
  NAND2_X1   g4721(.A1(new_n4769_), .A2(new_n4770_), .ZN(new_n4771_));
  NAND2_X1   g4722(.A1(new_n4767_), .A2(new_n4771_), .ZN(new_n4772_));
  AOI21_X1   g4723(.A1(new_n4578_), .A2(new_n4579_), .B(new_n4581_), .ZN(new_n4773_));
  NOR2_X1    g4724(.A1(new_n4773_), .A2(new_n4666_), .ZN(new_n4774_));
  INV_X1     g4725(.I(new_n4666_), .ZN(new_n4775_));
  NOR2_X1    g4726(.A1(new_n4775_), .A2(new_n4590_), .ZN(new_n4776_));
  NOR3_X1    g4727(.A1(new_n4776_), .A2(new_n4668_), .A3(new_n4774_), .ZN(new_n4777_));
  NOR2_X1    g4728(.A1(new_n4777_), .A2(new_n4585_), .ZN(new_n4778_));
  XOR2_X1    g4729(.A1(new_n4778_), .A2(new_n4772_), .Z(new_n4779_));
  XOR2_X1    g4730(.A1(new_n4779_), .A2(new_n4672_), .Z(\sin[5] ));
  NOR2_X1    g4731(.A1(new_n4769_), .A2(new_n4770_), .ZN(new_n4781_));
  NOR2_X1    g4732(.A1(new_n4764_), .A2(new_n4766_), .ZN(new_n4782_));
  OAI21_X1   g4733(.A1(new_n4781_), .A2(new_n4782_), .B(new_n4671_), .ZN(new_n4783_));
  INV_X1     g4734(.I(new_n4783_), .ZN(new_n4784_));
  INV_X1     g4735(.I(new_n4739_), .ZN(new_n4785_));
  AOI21_X1   g4736(.A1(new_n4737_), .A2(new_n4641_), .B(new_n4741_), .ZN(new_n4786_));
  XOR2_X1    g4737(.A1(new_n4722_), .A2(new_n1132_), .Z(new_n4787_));
  INV_X1     g4738(.I(new_n4787_), .ZN(new_n4788_));
  NAND2_X1   g4739(.A1(new_n4788_), .A2(new_n4717_), .ZN(new_n4789_));
  NAND2_X1   g4740(.A1(new_n4733_), .A2(new_n4787_), .ZN(new_n4790_));
  AOI22_X1   g4741(.A1(new_n4790_), .A2(new_n4789_), .B1(new_n4725_), .B2(new_n4788_), .ZN(new_n4791_));
  AOI22_X1   g4742(.A1(new_n4439_), .A2(new_n71_), .B1(new_n2741_), .B2(new_n4131_), .ZN(new_n4792_));
  INV_X1     g4743(.I(new_n4792_), .ZN(new_n4793_));
  NOR2_X1    g4744(.A1(new_n4507_), .A2(new_n4508_), .ZN(new_n4794_));
  AOI22_X1   g4745(.A1(new_n3895_), .A2(new_n3009_), .B1(new_n2773_), .B2(new_n3414_), .ZN(new_n4795_));
  AOI21_X1   g4746(.A1(new_n2776_), .A2(new_n4028_), .B(new_n4795_), .ZN(new_n4796_));
  OR3_X2     g4747(.A1(new_n4794_), .A2(new_n2779_), .A3(new_n4796_), .Z(new_n4797_));
  NOR2_X1    g4748(.A1(new_n4797_), .A2(new_n1134_), .ZN(new_n4798_));
  INV_X1     g4749(.I(new_n4798_), .ZN(new_n4799_));
  NAND2_X1   g4750(.A1(new_n4797_), .A2(new_n1134_), .ZN(new_n4800_));
  NAND2_X1   g4751(.A1(new_n4799_), .A2(new_n4800_), .ZN(new_n4801_));
  NAND2_X1   g4752(.A1(new_n3668_), .A2(new_n2855_), .ZN(new_n4802_));
  NAND2_X1   g4753(.A1(new_n3418_), .A2(new_n2851_), .ZN(new_n4803_));
  AOI21_X1   g4754(.A1(new_n2745_), .A2(new_n2848_), .B(new_n2881_), .ZN(new_n4804_));
  NAND4_X1   g4755(.A1(new_n3994_), .A2(new_n4802_), .A3(new_n4803_), .A4(new_n4804_), .ZN(new_n4805_));
  XOR2_X1    g4756(.A1(new_n4805_), .A2(new_n790_), .Z(new_n4806_));
  NOR2_X1    g4757(.A1(new_n2619_), .A2(new_n659_), .ZN(new_n4807_));
  INV_X1     g4758(.I(new_n4807_), .ZN(new_n4808_));
  INV_X1     g4759(.I(new_n4698_), .ZN(new_n4809_));
  NOR3_X1    g4760(.A1(new_n4709_), .A2(new_n69_), .A3(new_n4809_), .ZN(new_n4810_));
  NAND3_X1   g4761(.A1(new_n4709_), .A2(new_n69_), .A3(new_n4809_), .ZN(new_n4811_));
  INV_X1     g4762(.I(new_n4811_), .ZN(new_n4812_));
  OAI21_X1   g4763(.A1(new_n4812_), .A2(new_n4810_), .B(new_n4808_), .ZN(new_n4813_));
  INV_X1     g4764(.I(new_n4813_), .ZN(new_n4814_));
  INV_X1     g4765(.I(new_n4810_), .ZN(new_n4815_));
  NAND3_X1   g4766(.A1(new_n4815_), .A2(new_n4811_), .A3(new_n4807_), .ZN(new_n4816_));
  INV_X1     g4767(.I(new_n4816_), .ZN(new_n4817_));
  AOI22_X1   g4768(.A1(new_n2577_), .A2(new_n2795_), .B1(new_n2586_), .B2(new_n2829_), .ZN(new_n4818_));
  AOI21_X1   g4769(.A1(new_n2559_), .A2(new_n2790_), .B(new_n4818_), .ZN(new_n4819_));
  OR3_X2     g4770(.A1(new_n3940_), .A2(new_n2796_), .A3(new_n4819_), .Z(new_n4820_));
  XOR2_X1    g4771(.A1(new_n4820_), .A2(new_n659_), .Z(new_n4821_));
  NOR3_X1    g4772(.A1(new_n4817_), .A2(new_n4814_), .A3(new_n4821_), .ZN(new_n4822_));
  INV_X1     g4773(.I(new_n4821_), .ZN(new_n4823_));
  AOI21_X1   g4774(.A1(new_n4816_), .A2(new_n4813_), .B(new_n4823_), .ZN(new_n4824_));
  OAI21_X1   g4775(.A1(new_n4822_), .A2(new_n4824_), .B(new_n4806_), .ZN(new_n4825_));
  XOR2_X1    g4776(.A1(new_n4805_), .A2(new_n576_), .Z(new_n4826_));
  AOI21_X1   g4777(.A1(new_n4816_), .A2(new_n4813_), .B(new_n4821_), .ZN(new_n4827_));
  NOR3_X1    g4778(.A1(new_n4817_), .A2(new_n4814_), .A3(new_n4823_), .ZN(new_n4828_));
  OAI21_X1   g4779(.A1(new_n4828_), .A2(new_n4827_), .B(new_n4826_), .ZN(new_n4829_));
  NAND2_X1   g4780(.A1(new_n4825_), .A2(new_n4829_), .ZN(new_n4830_));
  NOR2_X1    g4781(.A1(new_n4705_), .A2(new_n4696_), .ZN(new_n4831_));
  NAND2_X1   g4782(.A1(new_n4705_), .A2(new_n4696_), .ZN(new_n4832_));
  XOR2_X1    g4783(.A1(new_n4709_), .A2(new_n4700_), .Z(new_n4833_));
  AOI21_X1   g4784(.A1(new_n4832_), .A2(new_n4833_), .B(new_n4831_), .ZN(new_n4834_));
  INV_X1     g4785(.I(new_n4834_), .ZN(new_n4835_));
  NAND2_X1   g4786(.A1(new_n4830_), .A2(new_n4835_), .ZN(new_n4836_));
  NAND3_X1   g4787(.A1(new_n4825_), .A2(new_n4829_), .A3(new_n4834_), .ZN(new_n4837_));
  NAND2_X1   g4788(.A1(new_n4836_), .A2(new_n4837_), .ZN(new_n4838_));
  NAND2_X1   g4789(.A1(new_n4838_), .A2(new_n4801_), .ZN(new_n4839_));
  INV_X1     g4790(.I(new_n4800_), .ZN(new_n4840_));
  NOR2_X1    g4791(.A1(new_n4840_), .A2(new_n4798_), .ZN(new_n4841_));
  NOR2_X1    g4792(.A1(new_n4830_), .A2(new_n4834_), .ZN(new_n4842_));
  AOI21_X1   g4793(.A1(new_n4825_), .A2(new_n4829_), .B(new_n4835_), .ZN(new_n4843_));
  OAI21_X1   g4794(.A1(new_n4842_), .A2(new_n4843_), .B(new_n4841_), .ZN(new_n4844_));
  AOI21_X1   g4795(.A1(new_n4839_), .A2(new_n4844_), .B(new_n4793_), .ZN(new_n4845_));
  AOI21_X1   g4796(.A1(new_n4836_), .A2(new_n4837_), .B(new_n4841_), .ZN(new_n4846_));
  NOR2_X1    g4797(.A1(new_n4842_), .A2(new_n4843_), .ZN(new_n4847_));
  NOR2_X1    g4798(.A1(new_n4847_), .A2(new_n4801_), .ZN(new_n4848_));
  NOR3_X1    g4799(.A1(new_n4848_), .A2(new_n4846_), .A3(new_n4792_), .ZN(new_n4849_));
  OAI21_X1   g4800(.A1(new_n4849_), .A2(new_n4845_), .B(new_n62_), .ZN(new_n4850_));
  OAI21_X1   g4801(.A1(new_n4848_), .A2(new_n4846_), .B(new_n4792_), .ZN(new_n4851_));
  NAND3_X1   g4802(.A1(new_n4839_), .A2(new_n4844_), .A3(new_n4793_), .ZN(new_n4852_));
  NAND3_X1   g4803(.A1(new_n4851_), .A2(new_n4852_), .A3(new_n943_), .ZN(new_n4853_));
  NAND2_X1   g4804(.A1(new_n4850_), .A2(new_n4853_), .ZN(new_n4854_));
  XOR2_X1    g4805(.A1(new_n4854_), .A2(new_n4791_), .Z(new_n4855_));
  NOR3_X1    g4806(.A1(new_n4855_), .A2(new_n4786_), .A3(new_n4785_), .ZN(new_n4856_));
  INV_X1     g4807(.I(new_n4786_), .ZN(new_n4857_));
  INV_X1     g4808(.I(new_n4791_), .ZN(new_n4858_));
  XOR2_X1    g4809(.A1(new_n4854_), .A2(new_n4858_), .Z(new_n4859_));
  AOI21_X1   g4810(.A1(new_n4857_), .A2(new_n4739_), .B(new_n4859_), .ZN(new_n4860_));
  NOR2_X1    g4811(.A1(new_n4860_), .A2(new_n4856_), .ZN(new_n4861_));
  NOR2_X1    g4812(.A1(new_n4662_), .A2(new_n4680_), .ZN(new_n4862_));
  AOI21_X1   g4813(.A1(new_n4681_), .A2(new_n4685_), .B(new_n4673_), .ZN(new_n4863_));
  NOR3_X1    g4814(.A1(new_n4863_), .A2(new_n4862_), .A3(new_n4687_), .ZN(new_n4864_));
  INV_X1     g4815(.I(new_n4862_), .ZN(new_n4865_));
  AOI21_X1   g4816(.A1(new_n4684_), .A2(new_n4661_), .B(new_n4651_), .ZN(new_n4866_));
  NOR2_X1    g4817(.A1(new_n4662_), .A2(new_n4680_), .ZN(new_n4867_));
  OAI21_X1   g4818(.A1(new_n4867_), .A2(new_n4866_), .B(new_n4598_), .ZN(new_n4868_));
  INV_X1     g4819(.I(new_n4687_), .ZN(new_n4869_));
  AOI21_X1   g4820(.A1(new_n4868_), .A2(new_n4865_), .B(new_n4869_), .ZN(new_n4870_));
  OAI21_X1   g4821(.A1(new_n4870_), .A2(new_n4864_), .B(new_n4745_), .ZN(new_n4871_));
  XOR2_X1    g4822(.A1(new_n4871_), .A2(new_n4861_), .Z(new_n4872_));
  NAND2_X1   g4823(.A1(new_n4686_), .A2(new_n4869_), .ZN(new_n4873_));
  XOR2_X1    g4824(.A1(new_n4872_), .A2(new_n4873_), .Z(new_n4874_));
  INV_X1     g4825(.I(new_n3780_), .ZN(new_n4875_));
  INV_X1     g4826(.I(new_n470_), .ZN(new_n4876_));
  NOR4_X1    g4827(.A1(new_n2316_), .A2(new_n194_), .A3(new_n331_), .A4(new_n1091_), .ZN(new_n4877_));
  INV_X1     g4828(.I(new_n1077_), .ZN(new_n4878_));
  NOR3_X1    g4829(.A1(new_n4878_), .A2(new_n257_), .A3(new_n1699_), .ZN(new_n4879_));
  NAND4_X1   g4830(.A1(new_n4879_), .A2(new_n4876_), .A3(new_n4877_), .A4(new_n2382_), .ZN(new_n4880_));
  NOR4_X1    g4831(.A1(new_n301_), .A2(new_n1021_), .A3(new_n369_), .A4(new_n525_), .ZN(new_n4881_));
  NAND3_X1   g4832(.A1(new_n1086_), .A2(new_n418_), .A3(new_n813_), .ZN(new_n4882_));
  NOR4_X1    g4833(.A1(new_n4882_), .A2(new_n2311_), .A3(new_n3405_), .A4(new_n4881_), .ZN(new_n4883_));
  INV_X1     g4834(.I(new_n4883_), .ZN(new_n4884_));
  NOR3_X1    g4835(.A1(new_n4875_), .A2(new_n4880_), .A3(new_n4884_), .ZN(new_n4885_));
  INV_X1     g4836(.I(new_n4885_), .ZN(new_n4886_));
  NAND2_X1   g4837(.A1(new_n4874_), .A2(new_n4886_), .ZN(new_n4887_));
  XNOR2_X1   g4838(.A1(new_n4872_), .A2(new_n4873_), .ZN(new_n4888_));
  NAND2_X1   g4839(.A1(new_n4888_), .A2(new_n4885_), .ZN(new_n4889_));
  NAND2_X1   g4840(.A1(new_n4889_), .A2(new_n4887_), .ZN(new_n4890_));
  NOR2_X1    g4841(.A1(new_n4784_), .A2(new_n4890_), .ZN(new_n4891_));
  INV_X1     g4842(.I(new_n4890_), .ZN(new_n4892_));
  NOR2_X1    g4843(.A1(new_n4892_), .A2(new_n4783_), .ZN(new_n4893_));
  NOR2_X1    g4844(.A1(new_n4893_), .A2(new_n4891_), .ZN(new_n4894_));
  AOI21_X1   g4845(.A1(new_n4771_), .A2(new_n4767_), .B(new_n4671_), .ZN(new_n4895_));
  NOR3_X1    g4846(.A1(new_n4672_), .A2(new_n4781_), .A3(new_n4782_), .ZN(new_n4896_));
  OAI22_X1   g4847(.A1(new_n4896_), .A2(new_n4895_), .B1(new_n4667_), .B2(new_n4668_), .ZN(new_n4897_));
  NAND2_X1   g4848(.A1(new_n4897_), .A2(new_n4102_), .ZN(new_n4898_));
  XOR2_X1    g4849(.A1(new_n4894_), .A2(new_n4898_), .Z(\sin[6] ));
  INV_X1     g4850(.I(new_n4895_), .ZN(new_n4900_));
  NAND3_X1   g4851(.A1(new_n4671_), .A2(new_n4767_), .A3(new_n4771_), .ZN(new_n4901_));
  AOI21_X1   g4852(.A1(new_n4900_), .A2(new_n4901_), .B(new_n4777_), .ZN(new_n4902_));
  AOI21_X1   g4853(.A1(new_n4894_), .A2(new_n4902_), .B(new_n4585_), .ZN(new_n4903_));
  NOR2_X1    g4854(.A1(new_n4890_), .A2(new_n4783_), .ZN(new_n4904_));
  XOR2_X1    g4855(.A1(new_n4792_), .A2(new_n943_), .Z(new_n4905_));
  INV_X1     g4856(.I(new_n4905_), .ZN(new_n4906_));
  NAND3_X1   g4857(.A1(new_n4839_), .A2(new_n4844_), .A3(new_n4906_), .ZN(new_n4907_));
  NAND2_X1   g4858(.A1(new_n4839_), .A2(new_n4844_), .ZN(new_n4908_));
  NAND2_X1   g4859(.A1(new_n4908_), .A2(new_n4905_), .ZN(new_n4909_));
  AOI22_X1   g4860(.A1(new_n4791_), .A2(new_n4906_), .B1(new_n4907_), .B2(new_n4909_), .ZN(new_n4910_));
  INV_X1     g4861(.I(new_n4843_), .ZN(new_n4911_));
  AOI21_X1   g4862(.A1(new_n4911_), .A2(new_n4801_), .B(new_n4842_), .ZN(new_n4912_));
  NOR2_X1    g4863(.A1(new_n4134_), .A2(new_n4136_), .ZN(new_n4913_));
  AOI22_X1   g4864(.A1(new_n4028_), .A2(new_n3009_), .B1(new_n2773_), .B2(new_n3895_), .ZN(new_n4914_));
  AOI21_X1   g4865(.A1(new_n2776_), .A2(new_n4131_), .B(new_n4914_), .ZN(new_n4915_));
  OR3_X2     g4866(.A1(new_n4913_), .A2(new_n2779_), .A3(new_n4915_), .Z(new_n4916_));
  XOR2_X1    g4867(.A1(new_n4916_), .A2(new_n1134_), .Z(new_n4917_));
  NOR2_X1    g4868(.A1(new_n4822_), .A2(new_n4806_), .ZN(new_n4918_));
  NOR2_X1    g4869(.A1(new_n4918_), .A2(new_n4824_), .ZN(new_n4919_));
  INV_X1     g4870(.I(new_n4709_), .ZN(new_n4920_));
  OAI21_X1   g4871(.A1(new_n4920_), .A2(new_n69_), .B(new_n4698_), .ZN(new_n4921_));
  OAI21_X1   g4872(.A1(new_n2739_), .A2(new_n4709_), .B(new_n4921_), .ZN(new_n4922_));
  OAI21_X1   g4873(.A1(new_n4922_), .A2(new_n69_), .B(new_n658_), .ZN(new_n4923_));
  AOI22_X1   g4874(.A1(new_n4923_), .A2(new_n2619_), .B1(new_n69_), .B2(new_n4922_), .ZN(new_n4924_));
  OAI22_X1   g4875(.A1(new_n2551_), .A2(new_n2791_), .B1(new_n2576_), .B2(new_n2830_), .ZN(new_n4925_));
  NAND2_X1   g4876(.A1(new_n2559_), .A2(new_n2795_), .ZN(new_n4926_));
  AOI21_X1   g4877(.A1(new_n4925_), .A2(new_n4926_), .B(new_n2796_), .ZN(new_n4927_));
  NAND2_X1   g4878(.A1(new_n3653_), .A2(new_n4927_), .ZN(new_n4928_));
  XOR2_X1    g4879(.A1(new_n4928_), .A2(new_n659_), .Z(new_n4929_));
  NOR2_X1    g4880(.A1(new_n2593_), .A2(new_n659_), .ZN(new_n4930_));
  NOR2_X1    g4881(.A1(new_n62_), .A2(new_n69_), .ZN(new_n4931_));
  NOR2_X1    g4882(.A1(new_n943_), .A2(new_n2739_), .ZN(new_n4932_));
  NOR2_X1    g4883(.A1(new_n4932_), .A2(new_n4931_), .ZN(new_n4933_));
  INV_X1     g4884(.I(new_n4933_), .ZN(new_n4934_));
  NOR2_X1    g4885(.A1(new_n4930_), .A2(new_n2740_), .ZN(new_n4935_));
  AOI21_X1   g4886(.A1(new_n4930_), .A2(new_n4934_), .B(new_n4935_), .ZN(new_n4936_));
  INV_X1     g4887(.I(new_n4936_), .ZN(new_n4937_));
  NAND2_X1   g4888(.A1(new_n4929_), .A2(new_n4937_), .ZN(new_n4938_));
  NOR2_X1    g4889(.A1(new_n4929_), .A2(new_n4937_), .ZN(new_n4939_));
  INV_X1     g4890(.I(new_n4939_), .ZN(new_n4940_));
  NAND2_X1   g4891(.A1(new_n4940_), .A2(new_n4938_), .ZN(new_n4941_));
  XOR2_X1    g4892(.A1(new_n4929_), .A2(new_n4936_), .Z(new_n4942_));
  NOR2_X1    g4893(.A1(new_n4924_), .A2(new_n4942_), .ZN(new_n4943_));
  AOI21_X1   g4894(.A1(new_n4924_), .A2(new_n4941_), .B(new_n4943_), .ZN(new_n4944_));
  OAI22_X1   g4895(.A1(new_n3449_), .A2(new_n2850_), .B1(new_n2882_), .B2(new_n3419_), .ZN(new_n4945_));
  NAND2_X1   g4896(.A1(new_n3414_), .A2(new_n2855_), .ZN(new_n4946_));
  AOI21_X1   g4897(.A1(new_n4945_), .A2(new_n4946_), .B(new_n2881_), .ZN(new_n4947_));
  NAND2_X1   g4898(.A1(new_n3464_), .A2(new_n4947_), .ZN(new_n4948_));
  XOR2_X1    g4899(.A1(new_n4948_), .A2(new_n576_), .Z(new_n4949_));
  INV_X1     g4900(.I(new_n4949_), .ZN(new_n4950_));
  NAND2_X1   g4901(.A1(new_n4944_), .A2(new_n4950_), .ZN(new_n4951_));
  NAND2_X1   g4902(.A1(new_n4924_), .A2(new_n4941_), .ZN(new_n4952_));
  OAI21_X1   g4903(.A1(new_n4924_), .A2(new_n4942_), .B(new_n4952_), .ZN(new_n4953_));
  NAND2_X1   g4904(.A1(new_n4953_), .A2(new_n4949_), .ZN(new_n4954_));
  AOI21_X1   g4905(.A1(new_n4951_), .A2(new_n4954_), .B(new_n4919_), .ZN(new_n4955_));
  INV_X1     g4906(.I(new_n4919_), .ZN(new_n4956_));
  NAND2_X1   g4907(.A1(new_n4953_), .A2(new_n4950_), .ZN(new_n4957_));
  NAND2_X1   g4908(.A1(new_n4944_), .A2(new_n4949_), .ZN(new_n4958_));
  AOI21_X1   g4909(.A1(new_n4958_), .A2(new_n4957_), .B(new_n4956_), .ZN(new_n4959_));
  NOR2_X1    g4910(.A1(new_n4955_), .A2(new_n4959_), .ZN(new_n4960_));
  INV_X1     g4911(.I(new_n4960_), .ZN(new_n4961_));
  NAND2_X1   g4912(.A1(new_n4961_), .A2(new_n4917_), .ZN(new_n4962_));
  INV_X1     g4913(.I(new_n4917_), .ZN(new_n4963_));
  NAND2_X1   g4914(.A1(new_n4960_), .A2(new_n4963_), .ZN(new_n4964_));
  AOI21_X1   g4915(.A1(new_n4962_), .A2(new_n4964_), .B(new_n4912_), .ZN(new_n4965_));
  INV_X1     g4916(.I(new_n4912_), .ZN(new_n4966_));
  NAND2_X1   g4917(.A1(new_n4961_), .A2(new_n4963_), .ZN(new_n4967_));
  NAND2_X1   g4918(.A1(new_n4960_), .A2(new_n4917_), .ZN(new_n4968_));
  AOI21_X1   g4919(.A1(new_n4967_), .A2(new_n4968_), .B(new_n4966_), .ZN(new_n4969_));
  NOR2_X1    g4920(.A1(new_n4965_), .A2(new_n4969_), .ZN(new_n4970_));
  XNOR2_X1   g4921(.A1(new_n4970_), .A2(new_n4910_), .ZN(new_n4971_));
  INV_X1     g4922(.I(new_n4971_), .ZN(new_n4972_));
  NOR3_X1    g4923(.A1(new_n443_), .A2(new_n524_), .A3(new_n643_), .ZN(new_n4973_));
  NOR2_X1    g4924(.A1(new_n764_), .A2(new_n815_), .ZN(new_n4974_));
  NAND4_X1   g4925(.A1(new_n312_), .A2(new_n727_), .A3(new_n930_), .A4(new_n950_), .ZN(new_n4975_));
  NAND4_X1   g4926(.A1(new_n4749_), .A2(new_n4973_), .A3(new_n4975_), .A4(new_n4974_), .ZN(new_n4976_));
  NOR3_X1    g4927(.A1(new_n2466_), .A2(new_n4880_), .A3(new_n4976_), .ZN(new_n4977_));
  NAND2_X1   g4928(.A1(new_n4857_), .A2(new_n4739_), .ZN(new_n4978_));
  NAND3_X1   g4929(.A1(new_n4857_), .A2(new_n4739_), .A3(new_n4859_), .ZN(new_n4979_));
  OAI21_X1   g4930(.A1(new_n4785_), .A2(new_n4786_), .B(new_n4855_), .ZN(new_n4980_));
  NAND2_X1   g4931(.A1(new_n4979_), .A2(new_n4980_), .ZN(new_n4981_));
  NOR2_X1    g4932(.A1(new_n4873_), .A2(new_n4981_), .ZN(new_n4982_));
  OAI22_X1   g4933(.A1(new_n4871_), .A2(new_n4982_), .B1(new_n4978_), .B2(new_n4859_), .ZN(new_n4983_));
  XNOR2_X1   g4934(.A1(new_n4983_), .A2(new_n4977_), .ZN(new_n4984_));
  NOR2_X1    g4935(.A1(new_n4984_), .A2(new_n4972_), .ZN(new_n4985_));
  INV_X1     g4936(.I(new_n4985_), .ZN(new_n4986_));
  NAND2_X1   g4937(.A1(new_n4984_), .A2(new_n4972_), .ZN(new_n4987_));
  NAND2_X1   g4938(.A1(new_n4986_), .A2(new_n4987_), .ZN(new_n4988_));
  NOR2_X1    g4939(.A1(new_n4888_), .A2(new_n4886_), .ZN(new_n4989_));
  INV_X1     g4940(.I(new_n4989_), .ZN(new_n4990_));
  NOR2_X1    g4941(.A1(new_n4990_), .A2(new_n4988_), .ZN(new_n4991_));
  AOI21_X1   g4942(.A1(new_n4986_), .A2(new_n4987_), .B(new_n4989_), .ZN(new_n4992_));
  OAI21_X1   g4943(.A1(new_n4991_), .A2(new_n4992_), .B(new_n4904_), .ZN(new_n4993_));
  INV_X1     g4944(.I(new_n4904_), .ZN(new_n4994_));
  NOR2_X1    g4945(.A1(new_n4991_), .A2(new_n4992_), .ZN(new_n4995_));
  NAND2_X1   g4946(.A1(new_n4995_), .A2(new_n4994_), .ZN(new_n4996_));
  NAND2_X1   g4947(.A1(new_n4996_), .A2(new_n4993_), .ZN(new_n4997_));
  NAND2_X1   g4948(.A1(new_n4903_), .A2(new_n4997_), .ZN(new_n4998_));
  XOR2_X1    g4949(.A1(new_n4995_), .A2(new_n4904_), .Z(new_n4999_));
  OAI21_X1   g4950(.A1(new_n4903_), .A2(new_n4999_), .B(new_n4998_), .ZN(\sin[7] ));
  INV_X1     g4951(.I(new_n4993_), .ZN(new_n5001_));
  NAND2_X1   g4952(.A1(new_n4970_), .A2(new_n4910_), .ZN(new_n5002_));
  INV_X1     g4953(.I(new_n5002_), .ZN(new_n5003_));
  INV_X1     g4954(.I(new_n4745_), .ZN(new_n5004_));
  NAND3_X1   g4955(.A1(new_n4868_), .A2(new_n4865_), .A3(new_n4869_), .ZN(new_n5005_));
  NAND2_X1   g4956(.A1(new_n4686_), .A2(new_n4687_), .ZN(new_n5006_));
  AOI21_X1   g4957(.A1(new_n5005_), .A2(new_n5006_), .B(new_n5004_), .ZN(new_n5007_));
  NAND3_X1   g4958(.A1(new_n4861_), .A2(new_n4686_), .A3(new_n4869_), .ZN(new_n5008_));
  XNOR2_X1   g4959(.A1(new_n4970_), .A2(new_n4910_), .ZN(new_n5009_));
  OAI21_X1   g4960(.A1(new_n4978_), .A2(new_n4859_), .B(new_n5009_), .ZN(new_n5010_));
  AOI21_X1   g4961(.A1(new_n5007_), .A2(new_n5008_), .B(new_n5010_), .ZN(new_n5011_));
  NOR2_X1    g4962(.A1(new_n5011_), .A2(new_n5003_), .ZN(new_n5012_));
  INV_X1     g4963(.I(new_n4964_), .ZN(new_n5013_));
  OAI21_X1   g4964(.A1(new_n4912_), .A2(new_n5013_), .B(new_n4962_), .ZN(new_n5014_));
  NAND2_X1   g4965(.A1(new_n4131_), .A2(new_n3009_), .ZN(new_n5015_));
  NAND2_X1   g4966(.A1(new_n4028_), .A2(new_n2773_), .ZN(new_n5016_));
  NAND4_X1   g4967(.A1(new_n4376_), .A2(new_n2778_), .A3(new_n5015_), .A4(new_n5016_), .ZN(new_n5017_));
  XOR2_X1    g4968(.A1(new_n5017_), .A2(new_n1134_), .Z(new_n5018_));
  AOI22_X1   g4969(.A1(new_n3668_), .A2(new_n2848_), .B1(new_n2851_), .B2(new_n3414_), .ZN(new_n5019_));
  AOI21_X1   g4970(.A1(new_n2855_), .A2(new_n3895_), .B(new_n5019_), .ZN(new_n5020_));
  OAI21_X1   g4971(.A1(new_n4718_), .A2(new_n2881_), .B(new_n5020_), .ZN(new_n5021_));
  AOI21_X1   g4972(.A1(new_n4924_), .A2(new_n4938_), .B(new_n4939_), .ZN(new_n5022_));
  OAI22_X1   g4973(.A1(new_n2551_), .A2(new_n2794_), .B1(new_n2558_), .B2(new_n2830_), .ZN(new_n5023_));
  NAND2_X1   g4974(.A1(new_n3418_), .A2(new_n2790_), .ZN(new_n5024_));
  AOI21_X1   g4975(.A1(new_n5024_), .A2(new_n5023_), .B(new_n2796_), .ZN(new_n5025_));
  NAND2_X1   g4976(.A1(new_n3472_), .A2(new_n5025_), .ZN(new_n5026_));
  XOR2_X1    g4977(.A1(new_n5026_), .A2(new_n658_), .Z(new_n5027_));
  NOR2_X1    g4978(.A1(new_n4930_), .A2(new_n4931_), .ZN(new_n5028_));
  NOR2_X1    g4979(.A1(new_n5028_), .A2(new_n4932_), .ZN(new_n5029_));
  NOR2_X1    g4980(.A1(new_n2576_), .A2(new_n659_), .ZN(new_n5030_));
  INV_X1     g4981(.I(new_n5030_), .ZN(new_n5031_));
  NOR2_X1    g4982(.A1(new_n5031_), .A2(new_n5029_), .ZN(new_n5032_));
  NOR3_X1    g4983(.A1(new_n5030_), .A2(new_n4932_), .A3(new_n5028_), .ZN(new_n5033_));
  OAI21_X1   g4984(.A1(new_n5032_), .A2(new_n5033_), .B(new_n5027_), .ZN(new_n5034_));
  XOR2_X1    g4985(.A1(new_n5030_), .A2(new_n5029_), .Z(new_n5035_));
  OAI21_X1   g4986(.A1(new_n5027_), .A2(new_n5035_), .B(new_n5034_), .ZN(new_n5036_));
  XOR2_X1    g4987(.A1(new_n5022_), .A2(new_n5036_), .Z(new_n5037_));
  XOR2_X1    g4988(.A1(new_n5037_), .A2(new_n790_), .Z(new_n5038_));
  XOR2_X1    g4989(.A1(new_n5038_), .A2(new_n5021_), .Z(new_n5039_));
  INV_X1     g4990(.I(new_n4951_), .ZN(new_n5040_));
  NOR2_X1    g4991(.A1(new_n4959_), .A2(new_n5040_), .ZN(new_n5041_));
  INV_X1     g4992(.I(new_n5041_), .ZN(new_n5042_));
  AND2_X2    g4993(.A1(new_n5039_), .A2(new_n5042_), .Z(new_n5043_));
  NOR2_X1    g4994(.A1(new_n5039_), .A2(new_n5042_), .ZN(new_n5044_));
  NOR2_X1    g4995(.A1(new_n5043_), .A2(new_n5044_), .ZN(new_n5045_));
  INV_X1     g4996(.I(new_n5045_), .ZN(new_n5046_));
  NAND2_X1   g4997(.A1(new_n5046_), .A2(new_n5018_), .ZN(new_n5047_));
  INV_X1     g4998(.I(new_n5018_), .ZN(new_n5048_));
  NAND2_X1   g4999(.A1(new_n5045_), .A2(new_n5048_), .ZN(new_n5049_));
  NAND2_X1   g5000(.A1(new_n5047_), .A2(new_n5049_), .ZN(new_n5050_));
  NOR2_X1    g5001(.A1(new_n5050_), .A2(new_n5014_), .ZN(new_n5051_));
  INV_X1     g5002(.I(new_n5051_), .ZN(new_n5052_));
  NAND2_X1   g5003(.A1(new_n5050_), .A2(new_n5014_), .ZN(new_n5053_));
  NAND2_X1   g5004(.A1(new_n5052_), .A2(new_n5053_), .ZN(new_n5054_));
  NOR4_X1    g5005(.A1(new_n608_), .A2(new_n533_), .A3(new_n974_), .A4(new_n595_), .ZN(new_n5055_));
  NOR4_X1    g5006(.A1(new_n1649_), .A2(new_n5055_), .A3(new_n534_), .A4(new_n889_), .ZN(new_n5056_));
  NAND3_X1   g5007(.A1(new_n2374_), .A2(new_n2294_), .A3(new_n5056_), .ZN(new_n5057_));
  INV_X1     g5008(.I(new_n5057_), .ZN(new_n5058_));
  INV_X1     g5009(.I(new_n1712_), .ZN(new_n5059_));
  NAND4_X1   g5010(.A1(new_n1088_), .A2(new_n223_), .A3(new_n412_), .A4(new_n504_), .ZN(new_n5060_));
  NOR4_X1    g5011(.A1(new_n3382_), .A2(new_n378_), .A3(new_n263_), .A4(new_n856_), .ZN(new_n5061_));
  NOR4_X1    g5012(.A1(new_n1078_), .A2(new_n5059_), .A3(new_n5060_), .A4(new_n5061_), .ZN(new_n5062_));
  NAND3_X1   g5013(.A1(new_n5058_), .A2(new_n3749_), .A3(new_n5062_), .ZN(new_n5063_));
  INV_X1     g5014(.I(new_n5063_), .ZN(new_n5064_));
  XOR2_X1    g5015(.A1(new_n5054_), .A2(new_n5064_), .Z(new_n5065_));
  NOR2_X1    g5016(.A1(new_n5065_), .A2(new_n5012_), .ZN(new_n5066_));
  XOR2_X1    g5017(.A1(new_n5054_), .A2(new_n5063_), .Z(new_n5067_));
  NOR3_X1    g5018(.A1(new_n5067_), .A2(new_n5003_), .A3(new_n5011_), .ZN(new_n5068_));
  AOI21_X1   g5019(.A1(new_n4983_), .A2(new_n4971_), .B(new_n4977_), .ZN(new_n5069_));
  OAI21_X1   g5020(.A1(new_n4971_), .A2(new_n4983_), .B(new_n5069_), .ZN(new_n5070_));
  NOR2_X1    g5021(.A1(new_n4989_), .A2(new_n5070_), .ZN(new_n5071_));
  NOR3_X1    g5022(.A1(new_n5071_), .A2(new_n5066_), .A3(new_n5068_), .ZN(new_n5072_));
  NOR2_X1    g5023(.A1(new_n5068_), .A2(new_n5066_), .ZN(new_n5073_));
  NOR3_X1    g5024(.A1(new_n5073_), .A2(new_n4989_), .A3(new_n5070_), .ZN(new_n5074_));
  NOR2_X1    g5025(.A1(new_n5072_), .A2(new_n5074_), .ZN(new_n5075_));
  INV_X1     g5026(.I(new_n5075_), .ZN(new_n5076_));
  OAI21_X1   g5027(.A1(new_n4893_), .A2(new_n4891_), .B(new_n4897_), .ZN(new_n5077_));
  OAI21_X1   g5028(.A1(new_n4991_), .A2(new_n4992_), .B(new_n4890_), .ZN(new_n5078_));
  INV_X1     g5029(.I(new_n5078_), .ZN(new_n5079_));
  NOR3_X1    g5030(.A1(new_n4991_), .A2(new_n4890_), .A3(new_n4992_), .ZN(new_n5080_));
  OAI21_X1   g5031(.A1(new_n5079_), .A2(new_n5080_), .B(new_n5077_), .ZN(new_n5081_));
  NAND2_X1   g5032(.A1(new_n5081_), .A2(new_n4102_), .ZN(new_n5082_));
  XOR2_X1    g5033(.A1(new_n5082_), .A2(new_n5076_), .Z(new_n5083_));
  XOR2_X1    g5034(.A1(new_n5083_), .A2(new_n5001_), .Z(\sin[8] ));
  AOI21_X1   g5035(.A1(new_n5048_), .A2(new_n5042_), .B(new_n5045_), .ZN(new_n5085_));
  XOR2_X1    g5036(.A1(new_n5021_), .A2(new_n576_), .Z(new_n5086_));
  XOR2_X1    g5037(.A1(new_n5086_), .A2(new_n5036_), .Z(new_n5087_));
  INV_X1     g5038(.I(new_n5087_), .ZN(new_n5088_));
  OAI21_X1   g5039(.A1(new_n5022_), .A2(new_n5086_), .B(new_n5088_), .ZN(new_n5089_));
  AOI22_X1   g5040(.A1(new_n3895_), .A2(new_n2851_), .B1(new_n2848_), .B2(new_n3414_), .ZN(new_n5090_));
  AOI21_X1   g5041(.A1(new_n2855_), .A2(new_n4028_), .B(new_n5090_), .ZN(new_n5091_));
  OR3_X2     g5042(.A1(new_n4794_), .A2(new_n2881_), .A3(new_n5091_), .Z(new_n5092_));
  XOR2_X1    g5043(.A1(new_n5092_), .A2(new_n576_), .Z(new_n5093_));
  INV_X1     g5044(.I(new_n5093_), .ZN(new_n5094_));
  NOR2_X1    g5045(.A1(new_n5027_), .A2(new_n5033_), .ZN(new_n5095_));
  NOR2_X1    g5046(.A1(new_n5095_), .A2(new_n5032_), .ZN(new_n5096_));
  OAI22_X1   g5047(.A1(new_n3419_), .A2(new_n2794_), .B1(new_n2551_), .B2(new_n2830_), .ZN(new_n5097_));
  NAND2_X1   g5048(.A1(new_n3668_), .A2(new_n2790_), .ZN(new_n5098_));
  AOI21_X1   g5049(.A1(new_n5098_), .A2(new_n5097_), .B(new_n2796_), .ZN(new_n5099_));
  NAND2_X1   g5050(.A1(new_n3994_), .A2(new_n5099_), .ZN(new_n5100_));
  XOR2_X1    g5051(.A1(new_n5100_), .A2(new_n658_), .Z(new_n5101_));
  NAND2_X1   g5052(.A1(new_n3142_), .A2(new_n658_), .ZN(new_n5102_));
  XNOR2_X1   g5053(.A1(new_n5101_), .A2(new_n5102_), .ZN(new_n5103_));
  XOR2_X1    g5054(.A1(new_n5103_), .A2(new_n5096_), .Z(new_n5104_));
  NAND2_X1   g5055(.A1(new_n5104_), .A2(new_n5094_), .ZN(new_n5105_));
  NOR2_X1    g5056(.A1(new_n5103_), .A2(new_n5096_), .ZN(new_n5106_));
  AND2_X2    g5057(.A1(new_n5103_), .A2(new_n5096_), .Z(new_n5107_));
  OAI21_X1   g5058(.A1(new_n5107_), .A2(new_n5106_), .B(new_n5093_), .ZN(new_n5108_));
  NAND2_X1   g5059(.A1(new_n5105_), .A2(new_n5108_), .ZN(new_n5109_));
  AOI22_X1   g5060(.A1(new_n4439_), .A2(new_n2778_), .B1(new_n2773_), .B2(new_n4131_), .ZN(new_n5110_));
  XOR2_X1    g5061(.A1(new_n5109_), .A2(new_n5110_), .Z(new_n5111_));
  XOR2_X1    g5062(.A1(new_n5111_), .A2(new_n1132_), .Z(new_n5112_));
  XOR2_X1    g5063(.A1(new_n5112_), .A2(new_n5089_), .Z(new_n5113_));
  INV_X1     g5064(.I(new_n5113_), .ZN(new_n5114_));
  NOR2_X1    g5065(.A1(new_n5114_), .A2(new_n5085_), .ZN(new_n5115_));
  INV_X1     g5066(.I(new_n5085_), .ZN(new_n5116_));
  NOR2_X1    g5067(.A1(new_n5116_), .A2(new_n5113_), .ZN(new_n5117_));
  NOR2_X1    g5068(.A1(new_n5115_), .A2(new_n5117_), .ZN(new_n5118_));
  INV_X1     g5069(.I(new_n5014_), .ZN(new_n5119_));
  AOI21_X1   g5070(.A1(new_n5012_), .A2(new_n5050_), .B(new_n5119_), .ZN(new_n5120_));
  AND2_X2    g5071(.A1(new_n5120_), .A2(new_n5118_), .Z(new_n5121_));
  NOR2_X1    g5072(.A1(new_n5120_), .A2(new_n5118_), .ZN(new_n5122_));
  NOR2_X1    g5073(.A1(new_n5121_), .A2(new_n5122_), .ZN(new_n5123_));
  NOR2_X1    g5074(.A1(new_n301_), .A2(new_n872_), .ZN(new_n5124_));
  NAND4_X1   g5075(.A1(new_n3393_), .A2(new_n469_), .A3(new_n3404_), .A4(new_n5124_), .ZN(new_n5125_));
  NOR4_X1    g5076(.A1(new_n741_), .A2(new_n172_), .A3(new_n239_), .A4(new_n1090_), .ZN(new_n5126_));
  NOR3_X1    g5077(.A1(new_n5125_), .A2(new_n3375_), .A3(new_n5126_), .ZN(new_n5127_));
  AND2_X2    g5078(.A1(new_n5127_), .A2(new_n725_), .Z(new_n5128_));
  NAND3_X1   g5079(.A1(new_n2385_), .A2(new_n5128_), .A3(new_n3783_), .ZN(new_n5129_));
  XOR2_X1    g5080(.A1(new_n5123_), .A2(new_n5129_), .Z(new_n5130_));
  OAI21_X1   g5081(.A1(new_n4993_), .A2(new_n5075_), .B(new_n5130_), .ZN(new_n5131_));
  NOR3_X1    g5082(.A1(new_n4993_), .A2(new_n5075_), .A3(new_n5130_), .ZN(new_n5132_));
  INV_X1     g5083(.I(new_n5132_), .ZN(new_n5133_));
  NAND2_X1   g5084(.A1(new_n5133_), .A2(new_n5131_), .ZN(new_n5134_));
  NOR2_X1    g5085(.A1(new_n4993_), .A2(new_n5075_), .ZN(new_n5135_));
  INV_X1     g5086(.I(new_n5135_), .ZN(new_n5136_));
  NAND2_X1   g5087(.A1(new_n4993_), .A2(new_n5075_), .ZN(new_n5137_));
  AOI21_X1   g5088(.A1(new_n5136_), .A2(new_n5137_), .B(new_n5081_), .ZN(new_n5138_));
  NOR2_X1    g5089(.A1(new_n5138_), .A2(new_n4585_), .ZN(new_n5139_));
  XOR2_X1    g5090(.A1(new_n5139_), .A2(new_n5134_), .Z(\sin[9] ));
  NAND2_X1   g5091(.A1(new_n4892_), .A2(new_n4783_), .ZN(new_n5141_));
  NAND2_X1   g5092(.A1(new_n4784_), .A2(new_n4890_), .ZN(new_n5142_));
  AOI21_X1   g5093(.A1(new_n5141_), .A2(new_n5142_), .B(new_n4902_), .ZN(new_n5143_));
  INV_X1     g5094(.I(new_n5080_), .ZN(new_n5144_));
  AOI21_X1   g5095(.A1(new_n5078_), .A2(new_n5144_), .B(new_n5143_), .ZN(new_n5145_));
  INV_X1     g5096(.I(new_n5137_), .ZN(new_n5146_));
  OAI21_X1   g5097(.A1(new_n5146_), .A2(new_n5135_), .B(new_n5145_), .ZN(new_n5147_));
  OAI21_X1   g5098(.A1(new_n5147_), .A2(new_n5134_), .B(new_n4102_), .ZN(new_n5148_));
  INV_X1     g5099(.I(new_n5130_), .ZN(new_n5149_));
  NOR3_X1    g5100(.A1(new_n4993_), .A2(new_n5149_), .A3(new_n5075_), .ZN(new_n5150_));
  INV_X1     g5101(.I(new_n5089_), .ZN(new_n5151_));
  XOR2_X1    g5102(.A1(new_n5110_), .A2(new_n1134_), .Z(new_n5152_));
  NOR3_X1    g5103(.A1(new_n5151_), .A2(new_n5109_), .A3(new_n5152_), .ZN(new_n5153_));
  AOI21_X1   g5104(.A1(new_n5151_), .A2(new_n5109_), .B(new_n5153_), .ZN(new_n5154_));
  XOR2_X1    g5105(.A1(new_n5101_), .A2(new_n2558_), .Z(new_n5155_));
  NAND2_X1   g5106(.A1(new_n5155_), .A2(new_n658_), .ZN(new_n5156_));
  AOI21_X1   g5107(.A1(new_n2576_), .A2(new_n5101_), .B(new_n5156_), .ZN(new_n5157_));
  NOR2_X1    g5108(.A1(new_n2551_), .A2(new_n659_), .ZN(new_n5158_));
  INV_X1     g5109(.I(new_n5158_), .ZN(new_n5159_));
  XOR2_X1    g5110(.A1(new_n5030_), .A2(new_n1132_), .Z(new_n5160_));
  NOR2_X1    g5111(.A1(new_n5159_), .A2(new_n5160_), .ZN(new_n5161_));
  NOR2_X1    g5112(.A1(new_n5031_), .A2(new_n1132_), .ZN(new_n5162_));
  NOR2_X1    g5113(.A1(new_n5030_), .A2(new_n1134_), .ZN(new_n5163_));
  NOR2_X1    g5114(.A1(new_n5162_), .A2(new_n5163_), .ZN(new_n5164_));
  NOR2_X1    g5115(.A1(new_n5158_), .A2(new_n5164_), .ZN(new_n5165_));
  NOR2_X1    g5116(.A1(new_n5161_), .A2(new_n5165_), .ZN(new_n5166_));
  INV_X1     g5117(.I(new_n5166_), .ZN(new_n5167_));
  XOR2_X1    g5118(.A1(new_n5157_), .A2(new_n5167_), .Z(new_n5168_));
  OAI22_X1   g5119(.A1(new_n3449_), .A2(new_n2794_), .B1(new_n2830_), .B2(new_n3419_), .ZN(new_n5169_));
  NAND2_X1   g5120(.A1(new_n3414_), .A2(new_n2790_), .ZN(new_n5170_));
  AOI21_X1   g5121(.A1(new_n5169_), .A2(new_n5170_), .B(new_n2796_), .ZN(new_n5171_));
  NAND2_X1   g5122(.A1(new_n3464_), .A2(new_n5171_), .ZN(new_n5172_));
  XOR2_X1    g5123(.A1(new_n5172_), .A2(new_n659_), .Z(new_n5173_));
  NAND2_X1   g5124(.A1(new_n5168_), .A2(new_n5173_), .ZN(new_n5174_));
  OR2_X2     g5125(.A1(new_n5168_), .A2(new_n5173_), .Z(new_n5175_));
  AND2_X2    g5126(.A1(new_n5175_), .A2(new_n5174_), .Z(new_n5176_));
  NOR2_X1    g5127(.A1(new_n5094_), .A2(new_n5107_), .ZN(new_n5177_));
  NOR2_X1    g5128(.A1(new_n5177_), .A2(new_n5106_), .ZN(new_n5178_));
  AOI22_X1   g5129(.A1(new_n4028_), .A2(new_n2851_), .B1(new_n2848_), .B2(new_n3895_), .ZN(new_n5179_));
  AOI21_X1   g5130(.A1(new_n2855_), .A2(new_n4131_), .B(new_n5179_), .ZN(new_n5180_));
  NOR3_X1    g5131(.A1(new_n4913_), .A2(new_n2881_), .A3(new_n5180_), .ZN(new_n5181_));
  XOR2_X1    g5132(.A1(new_n5181_), .A2(new_n790_), .Z(new_n5182_));
  XOR2_X1    g5133(.A1(new_n5178_), .A2(new_n5182_), .Z(new_n5183_));
  NOR2_X1    g5134(.A1(new_n5176_), .A2(new_n5183_), .ZN(new_n5184_));
  INV_X1     g5135(.I(new_n5176_), .ZN(new_n5185_));
  INV_X1     g5136(.I(new_n5178_), .ZN(new_n5186_));
  NOR2_X1    g5137(.A1(new_n5186_), .A2(new_n5182_), .ZN(new_n5187_));
  INV_X1     g5138(.I(new_n5187_), .ZN(new_n5188_));
  NAND2_X1   g5139(.A1(new_n5186_), .A2(new_n5182_), .ZN(new_n5189_));
  AOI21_X1   g5140(.A1(new_n5188_), .A2(new_n5189_), .B(new_n5185_), .ZN(new_n5190_));
  NOR2_X1    g5141(.A1(new_n5190_), .A2(new_n5184_), .ZN(new_n5191_));
  XOR2_X1    g5142(.A1(new_n5191_), .A2(new_n5154_), .Z(new_n5192_));
  INV_X1     g5143(.I(new_n5192_), .ZN(new_n5193_));
  NOR4_X1    g5144(.A1(new_n4878_), .A2(new_n3785_), .A3(new_n632_), .A4(new_n3405_), .ZN(new_n5194_));
  NAND2_X1   g5145(.A1(new_n330_), .A2(new_n619_), .ZN(new_n5195_));
  NAND2_X1   g5146(.A1(new_n153_), .A2(new_n613_), .ZN(new_n5196_));
  NOR4_X1    g5147(.A1(new_n3784_), .A2(new_n404_), .A3(new_n5195_), .A4(new_n5196_), .ZN(new_n5197_));
  NOR2_X1    g5148(.A1(new_n546_), .A2(new_n882_), .ZN(new_n5198_));
  NAND4_X1   g5149(.A1(new_n5198_), .A2(new_n3756_), .A3(new_n5194_), .A4(new_n5197_), .ZN(new_n5199_));
  NOR2_X1    g5150(.A1(new_n4978_), .A2(new_n4859_), .ZN(new_n5200_));
  XOR2_X1    g5151(.A1(new_n4970_), .A2(new_n4910_), .Z(new_n5201_));
  NOR2_X1    g5152(.A1(new_n5200_), .A2(new_n5201_), .ZN(new_n5202_));
  OAI21_X1   g5153(.A1(new_n4871_), .A2(new_n4982_), .B(new_n5202_), .ZN(new_n5203_));
  AOI21_X1   g5154(.A1(new_n5047_), .A2(new_n5049_), .B(new_n5014_), .ZN(new_n5204_));
  NAND3_X1   g5155(.A1(new_n5203_), .A2(new_n5002_), .A3(new_n5204_), .ZN(new_n5205_));
  NOR3_X1    g5156(.A1(new_n5115_), .A2(new_n5117_), .A3(new_n5204_), .ZN(new_n5206_));
  NAND2_X1   g5157(.A1(new_n5205_), .A2(new_n5206_), .ZN(new_n5207_));
  XOR2_X1    g5158(.A1(new_n5207_), .A2(new_n5199_), .Z(new_n5208_));
  NOR2_X1    g5159(.A1(new_n5208_), .A2(new_n5193_), .ZN(new_n5209_));
  INV_X1     g5160(.I(new_n5204_), .ZN(new_n5210_));
  NOR3_X1    g5161(.A1(new_n5011_), .A2(new_n5003_), .A3(new_n5210_), .ZN(new_n5211_));
  INV_X1     g5162(.I(new_n5206_), .ZN(new_n5212_));
  NOR2_X1    g5163(.A1(new_n5211_), .A2(new_n5212_), .ZN(new_n5213_));
  XOR2_X1    g5164(.A1(new_n5213_), .A2(new_n5199_), .Z(new_n5214_));
  NOR2_X1    g5165(.A1(new_n5214_), .A2(new_n5192_), .ZN(new_n5215_));
  NOR3_X1    g5166(.A1(new_n5121_), .A2(new_n5122_), .A3(new_n5129_), .ZN(new_n5216_));
  INV_X1     g5167(.I(new_n5216_), .ZN(new_n5217_));
  OR3_X2     g5168(.A1(new_n5217_), .A2(new_n5209_), .A3(new_n5215_), .Z(new_n5218_));
  OAI21_X1   g5169(.A1(new_n5209_), .A2(new_n5215_), .B(new_n5217_), .ZN(new_n5219_));
  NAND2_X1   g5170(.A1(new_n5218_), .A2(new_n5219_), .ZN(new_n5220_));
  NAND2_X1   g5171(.A1(new_n5150_), .A2(new_n5220_), .ZN(new_n5221_));
  INV_X1     g5172(.I(new_n5221_), .ZN(new_n5222_));
  NOR2_X1    g5173(.A1(new_n5150_), .A2(new_n5220_), .ZN(new_n5223_));
  NOR2_X1    g5174(.A1(new_n5222_), .A2(new_n5223_), .ZN(new_n5224_));
  XOR2_X1    g5175(.A1(new_n5150_), .A2(new_n5220_), .Z(new_n5225_));
  NAND2_X1   g5176(.A1(new_n5148_), .A2(new_n5225_), .ZN(new_n5226_));
  OAI21_X1   g5177(.A1(new_n5148_), .A2(new_n5224_), .B(new_n5226_), .ZN(\sin[10] ));
  INV_X1     g5178(.I(new_n5154_), .ZN(new_n5228_));
  OAI21_X1   g5179(.A1(new_n5211_), .A2(new_n5212_), .B(new_n5191_), .ZN(new_n5229_));
  INV_X1     g5180(.I(new_n5191_), .ZN(new_n5230_));
  NAND3_X1   g5181(.A1(new_n5205_), .A2(new_n5230_), .A3(new_n5206_), .ZN(new_n5231_));
  AOI22_X1   g5182(.A1(new_n5229_), .A2(new_n5231_), .B1(new_n5207_), .B2(new_n5228_), .ZN(new_n5232_));
  OAI21_X1   g5183(.A1(new_n5176_), .A2(new_n5187_), .B(new_n5189_), .ZN(new_n5233_));
  NAND2_X1   g5184(.A1(new_n4131_), .A2(new_n2851_), .ZN(new_n5234_));
  NAND2_X1   g5185(.A1(new_n4028_), .A2(new_n2848_), .ZN(new_n5235_));
  NAND4_X1   g5186(.A1(new_n4376_), .A2(new_n2858_), .A3(new_n5234_), .A4(new_n5235_), .ZN(new_n5236_));
  XOR2_X1    g5187(.A1(new_n5236_), .A2(new_n576_), .Z(new_n5237_));
  AOI22_X1   g5188(.A1(new_n3668_), .A2(new_n2829_), .B1(new_n2795_), .B2(new_n3414_), .ZN(new_n5238_));
  AOI21_X1   g5189(.A1(new_n2790_), .A2(new_n3895_), .B(new_n5238_), .ZN(new_n5239_));
  NOR3_X1    g5190(.A1(new_n4718_), .A2(new_n2796_), .A3(new_n5239_), .ZN(new_n5240_));
  XOR2_X1    g5191(.A1(new_n5240_), .A2(new_n658_), .Z(new_n5241_));
  INV_X1     g5192(.I(new_n5162_), .ZN(new_n5242_));
  AOI21_X1   g5193(.A1(new_n5159_), .A2(new_n5242_), .B(new_n5163_), .ZN(new_n5243_));
  INV_X1     g5194(.I(new_n5243_), .ZN(new_n5244_));
  NOR2_X1    g5195(.A1(new_n3419_), .A2(new_n659_), .ZN(new_n5245_));
  NAND2_X1   g5196(.A1(new_n5244_), .A2(new_n5245_), .ZN(new_n5246_));
  INV_X1     g5197(.I(new_n5245_), .ZN(new_n5247_));
  NAND2_X1   g5198(.A1(new_n5247_), .A2(new_n5243_), .ZN(new_n5248_));
  AOI21_X1   g5199(.A1(new_n5246_), .A2(new_n5248_), .B(new_n5241_), .ZN(new_n5249_));
  XNOR2_X1   g5200(.A1(new_n5243_), .A2(new_n5245_), .ZN(new_n5250_));
  AOI21_X1   g5201(.A1(new_n5241_), .A2(new_n5250_), .B(new_n5249_), .ZN(new_n5251_));
  OAI21_X1   g5202(.A1(new_n5157_), .A2(new_n5167_), .B(new_n5174_), .ZN(new_n5252_));
  XOR2_X1    g5203(.A1(new_n5252_), .A2(new_n5251_), .Z(new_n5253_));
  XNOR2_X1   g5204(.A1(new_n5253_), .A2(new_n5237_), .ZN(new_n5254_));
  XOR2_X1    g5205(.A1(new_n5254_), .A2(new_n5233_), .Z(new_n5255_));
  AND4_X2    g5206(.A1(new_n294_), .A2(new_n373_), .A3(new_n947_), .A4(new_n954_), .Z(new_n5256_));
  NAND4_X1   g5207(.A1(new_n538_), .A2(new_n644_), .A3(new_n4013_), .A4(new_n5256_), .ZN(new_n5257_));
  XOR2_X1    g5208(.A1(new_n5255_), .A2(new_n5257_), .Z(new_n5258_));
  XOR2_X1    g5209(.A1(new_n5255_), .A2(new_n5257_), .Z(new_n5259_));
  NOR2_X1    g5210(.A1(new_n5232_), .A2(new_n5259_), .ZN(new_n5260_));
  AOI21_X1   g5211(.A1(new_n5232_), .A2(new_n5258_), .B(new_n5260_), .ZN(new_n5261_));
  XOR2_X1    g5212(.A1(new_n5207_), .A2(new_n5193_), .Z(new_n5262_));
  NAND2_X1   g5213(.A1(new_n5262_), .A2(new_n5199_), .ZN(new_n5263_));
  NAND2_X1   g5214(.A1(new_n5217_), .A2(new_n5263_), .ZN(new_n5264_));
  XOR2_X1    g5215(.A1(new_n5264_), .A2(new_n5261_), .Z(new_n5265_));
  INV_X1     g5216(.I(new_n5265_), .ZN(new_n5266_));
  INV_X1     g5217(.I(new_n5131_), .ZN(new_n5267_));
  NOR2_X1    g5218(.A1(new_n5267_), .A2(new_n5132_), .ZN(new_n5268_));
  XOR2_X1    g5219(.A1(new_n5220_), .A2(new_n5130_), .Z(new_n5269_));
  OAI21_X1   g5220(.A1(new_n5138_), .A2(new_n5268_), .B(new_n5269_), .ZN(new_n5270_));
  NAND2_X1   g5221(.A1(new_n5270_), .A2(new_n4102_), .ZN(new_n5271_));
  XOR2_X1    g5222(.A1(new_n5271_), .A2(new_n5266_), .Z(new_n5272_));
  XOR2_X1    g5223(.A1(new_n5272_), .A2(new_n5222_), .Z(\sin[11] ));
  NAND3_X1   g5224(.A1(new_n5266_), .A2(new_n5150_), .A3(new_n5220_), .ZN(new_n5274_));
  NAND2_X1   g5225(.A1(new_n5251_), .A2(new_n5237_), .ZN(new_n5275_));
  NOR2_X1    g5226(.A1(new_n5251_), .A2(new_n5237_), .ZN(new_n5276_));
  OAI21_X1   g5227(.A1(new_n5252_), .A2(new_n5276_), .B(new_n5275_), .ZN(new_n5277_));
  AOI22_X1   g5228(.A1(new_n3895_), .A2(new_n2795_), .B1(new_n2829_), .B2(new_n3414_), .ZN(new_n5278_));
  AOI21_X1   g5229(.A1(new_n2790_), .A2(new_n4028_), .B(new_n5278_), .ZN(new_n5279_));
  OR3_X2     g5230(.A1(new_n4794_), .A2(new_n2796_), .A3(new_n5279_), .Z(new_n5280_));
  XOR2_X1    g5231(.A1(new_n5280_), .A2(new_n659_), .Z(new_n5281_));
  AOI22_X1   g5232(.A1(new_n4439_), .A2(new_n2858_), .B1(new_n2848_), .B2(new_n4131_), .ZN(new_n5282_));
  NAND2_X1   g5233(.A1(new_n5241_), .A2(new_n5248_), .ZN(new_n5283_));
  NOR3_X1    g5234(.A1(new_n3449_), .A2(new_n659_), .A3(new_n3418_), .ZN(new_n5284_));
  INV_X1     g5235(.I(new_n5284_), .ZN(new_n5285_));
  NOR2_X1    g5236(.A1(new_n3449_), .A2(new_n659_), .ZN(new_n5286_));
  NOR2_X1    g5237(.A1(new_n5247_), .A2(new_n5286_), .ZN(new_n5287_));
  INV_X1     g5238(.I(new_n5287_), .ZN(new_n5288_));
  AOI22_X1   g5239(.A1(new_n5283_), .A2(new_n5246_), .B1(new_n5285_), .B2(new_n5288_), .ZN(new_n5289_));
  NAND2_X1   g5240(.A1(new_n5283_), .A2(new_n5246_), .ZN(new_n5290_));
  XOR2_X1    g5241(.A1(new_n5286_), .A2(new_n5245_), .Z(new_n5291_));
  NOR2_X1    g5242(.A1(new_n5290_), .A2(new_n5291_), .ZN(new_n5292_));
  NOR2_X1    g5243(.A1(new_n5292_), .A2(new_n5289_), .ZN(new_n5293_));
  XOR2_X1    g5244(.A1(new_n5293_), .A2(new_n5282_), .Z(new_n5294_));
  XOR2_X1    g5245(.A1(new_n5294_), .A2(new_n576_), .Z(new_n5295_));
  XOR2_X1    g5246(.A1(new_n5295_), .A2(new_n5281_), .Z(new_n5296_));
  XOR2_X1    g5247(.A1(new_n5296_), .A2(new_n5277_), .Z(new_n5297_));
  INV_X1     g5248(.I(new_n5297_), .ZN(new_n5298_));
  INV_X1     g5249(.I(new_n5254_), .ZN(new_n5299_));
  NAND2_X1   g5250(.A1(new_n5213_), .A2(new_n5230_), .ZN(new_n5300_));
  AOI21_X1   g5251(.A1(new_n5205_), .A2(new_n5206_), .B(new_n5230_), .ZN(new_n5301_));
  NOR3_X1    g5252(.A1(new_n5211_), .A2(new_n5191_), .A3(new_n5212_), .ZN(new_n5302_));
  OAI21_X1   g5253(.A1(new_n5302_), .A2(new_n5301_), .B(new_n5154_), .ZN(new_n5303_));
  NAND3_X1   g5254(.A1(new_n5303_), .A2(new_n5300_), .A3(new_n5233_), .ZN(new_n5304_));
  INV_X1     g5255(.I(new_n5233_), .ZN(new_n5305_));
  NAND2_X1   g5256(.A1(new_n5232_), .A2(new_n5305_), .ZN(new_n5306_));
  AOI21_X1   g5257(.A1(new_n5306_), .A2(new_n5304_), .B(new_n5299_), .ZN(new_n5307_));
  NAND2_X1   g5258(.A1(new_n5307_), .A2(new_n5298_), .ZN(new_n5308_));
  NOR2_X1    g5259(.A1(new_n5207_), .A2(new_n5191_), .ZN(new_n5309_));
  AOI21_X1   g5260(.A1(new_n5229_), .A2(new_n5231_), .B(new_n5228_), .ZN(new_n5310_));
  NOR3_X1    g5261(.A1(new_n5310_), .A2(new_n5309_), .A3(new_n5305_), .ZN(new_n5311_));
  AOI21_X1   g5262(.A1(new_n5303_), .A2(new_n5300_), .B(new_n5233_), .ZN(new_n5312_));
  OAI21_X1   g5263(.A1(new_n5312_), .A2(new_n5311_), .B(new_n5254_), .ZN(new_n5313_));
  NAND2_X1   g5264(.A1(new_n5313_), .A2(new_n5297_), .ZN(new_n5314_));
  NAND2_X1   g5265(.A1(new_n5232_), .A2(new_n5233_), .ZN(new_n5315_));
  INV_X1     g5266(.I(new_n5315_), .ZN(new_n5316_));
  NAND3_X1   g5267(.A1(new_n5314_), .A2(new_n5308_), .A3(new_n5316_), .ZN(new_n5317_));
  AOI21_X1   g5268(.A1(new_n5314_), .A2(new_n5308_), .B(new_n5316_), .ZN(new_n5318_));
  INV_X1     g5269(.I(new_n5318_), .ZN(new_n5319_));
  NAND2_X1   g5270(.A1(new_n5319_), .A2(new_n5317_), .ZN(new_n5320_));
  NOR4_X1    g5271(.A1(new_n2425_), .A2(new_n267_), .A3(new_n533_), .A4(new_n715_), .ZN(new_n5321_));
  INV_X1     g5272(.I(new_n5321_), .ZN(new_n5322_));
  NAND2_X1   g5273(.A1(new_n319_), .A2(new_n342_), .ZN(new_n5323_));
  NOR4_X1    g5274(.A1(new_n5323_), .A2(new_n865_), .A3(new_n1090_), .A4(new_n597_), .ZN(new_n5324_));
  INV_X1     g5275(.I(new_n5324_), .ZN(new_n5325_));
  NOR4_X1    g5276(.A1(new_n5322_), .A2(new_n823_), .A3(new_n4403_), .A4(new_n5325_), .ZN(new_n5326_));
  NAND3_X1   g5277(.A1(new_n5326_), .A2(new_n248_), .A3(new_n1643_), .ZN(new_n5327_));
  INV_X1     g5278(.I(new_n5327_), .ZN(new_n5328_));
  NOR2_X1    g5279(.A1(new_n5320_), .A2(new_n5328_), .ZN(new_n5329_));
  INV_X1     g5280(.I(new_n5317_), .ZN(new_n5330_));
  NOR2_X1    g5281(.A1(new_n5330_), .A2(new_n5318_), .ZN(new_n5331_));
  NOR2_X1    g5282(.A1(new_n5331_), .A2(new_n5327_), .ZN(new_n5332_));
  NOR3_X1    g5283(.A1(new_n5329_), .A2(new_n5274_), .A3(new_n5332_), .ZN(new_n5333_));
  NOR2_X1    g5284(.A1(new_n5221_), .A2(new_n5265_), .ZN(new_n5334_));
  NAND2_X1   g5285(.A1(new_n5331_), .A2(new_n5327_), .ZN(new_n5335_));
  NAND2_X1   g5286(.A1(new_n5320_), .A2(new_n5328_), .ZN(new_n5336_));
  AOI21_X1   g5287(.A1(new_n5335_), .A2(new_n5336_), .B(new_n5334_), .ZN(new_n5337_));
  NOR2_X1    g5288(.A1(new_n5337_), .A2(new_n5333_), .ZN(new_n5338_));
  NAND2_X1   g5289(.A1(new_n5147_), .A2(new_n5134_), .ZN(new_n5339_));
  NAND2_X1   g5290(.A1(new_n5221_), .A2(new_n5265_), .ZN(new_n5340_));
  NAND2_X1   g5291(.A1(new_n5340_), .A2(new_n5274_), .ZN(new_n5341_));
  NAND3_X1   g5292(.A1(new_n5339_), .A2(new_n5341_), .A3(new_n5269_), .ZN(new_n5342_));
  NAND2_X1   g5293(.A1(new_n5342_), .A2(new_n4102_), .ZN(new_n5343_));
  XOR2_X1    g5294(.A1(new_n5343_), .A2(new_n5338_), .Z(\sin[12] ));
  NAND2_X1   g5295(.A1(new_n5290_), .A2(new_n5288_), .ZN(new_n5345_));
  NAND2_X1   g5296(.A1(new_n5345_), .A2(new_n5285_), .ZN(new_n5346_));
  AOI22_X1   g5297(.A1(new_n4028_), .A2(new_n2795_), .B1(new_n2829_), .B2(new_n3895_), .ZN(new_n5347_));
  AOI21_X1   g5298(.A1(new_n2790_), .A2(new_n4131_), .B(new_n5347_), .ZN(new_n5348_));
  OR3_X2     g5299(.A1(new_n4913_), .A2(new_n2796_), .A3(new_n5348_), .Z(new_n5349_));
  XOR2_X1    g5300(.A1(new_n5349_), .A2(new_n659_), .Z(new_n5350_));
  INV_X1     g5301(.I(new_n5350_), .ZN(new_n5351_));
  NOR3_X1    g5302(.A1(new_n3905_), .A2(new_n659_), .A3(new_n3897_), .ZN(new_n5352_));
  XOR2_X1    g5303(.A1(new_n5352_), .A2(new_n576_), .Z(new_n5353_));
  NOR2_X1    g5304(.A1(new_n5351_), .A2(new_n5353_), .ZN(new_n5354_));
  NAND2_X1   g5305(.A1(new_n5351_), .A2(new_n5353_), .ZN(new_n5355_));
  INV_X1     g5306(.I(new_n5355_), .ZN(new_n5356_));
  OAI21_X1   g5307(.A1(new_n5356_), .A2(new_n5354_), .B(new_n5346_), .ZN(new_n5357_));
  XOR2_X1    g5308(.A1(new_n5350_), .A2(new_n5353_), .Z(new_n5358_));
  OAI21_X1   g5309(.A1(new_n5346_), .A2(new_n5358_), .B(new_n5357_), .ZN(new_n5359_));
  NOR2_X1    g5310(.A1(new_n5293_), .A2(new_n5281_), .ZN(new_n5360_));
  INV_X1     g5311(.I(new_n5281_), .ZN(new_n5361_));
  XOR2_X1    g5312(.A1(new_n5282_), .A2(new_n576_), .Z(new_n5362_));
  NOR2_X1    g5313(.A1(new_n5361_), .A2(new_n5362_), .ZN(new_n5363_));
  AOI21_X1   g5314(.A1(new_n5293_), .A2(new_n5363_), .B(new_n5360_), .ZN(new_n5364_));
  XOR2_X1    g5315(.A1(new_n5359_), .A2(new_n5364_), .Z(new_n5365_));
  INV_X1     g5316(.I(new_n5365_), .ZN(new_n5366_));
  NAND3_X1   g5317(.A1(new_n5232_), .A2(new_n5233_), .A3(new_n5298_), .ZN(new_n5367_));
  NAND2_X1   g5318(.A1(new_n5307_), .A2(new_n5367_), .ZN(new_n5368_));
  NAND2_X1   g5319(.A1(new_n5296_), .A2(new_n5277_), .ZN(new_n5369_));
  AOI21_X1   g5320(.A1(new_n5368_), .A2(new_n5369_), .B(new_n5366_), .ZN(new_n5370_));
  NAND2_X1   g5321(.A1(new_n5369_), .A2(new_n5366_), .ZN(new_n5371_));
  AOI21_X1   g5322(.A1(new_n5307_), .A2(new_n5367_), .B(new_n5371_), .ZN(new_n5372_));
  NOR2_X1    g5323(.A1(new_n5370_), .A2(new_n5372_), .ZN(new_n5373_));
  NAND2_X1   g5324(.A1(new_n542_), .A2(new_n440_), .ZN(new_n5374_));
  NOR4_X1    g5325(.A1(new_n5374_), .A2(new_n483_), .A3(new_n488_), .A4(new_n832_), .ZN(new_n5375_));
  NAND2_X1   g5326(.A1(new_n131_), .A2(new_n288_), .ZN(new_n5376_));
  NOR4_X1    g5327(.A1(new_n5376_), .A2(new_n257_), .A3(new_n484_), .A4(new_n869_), .ZN(new_n5377_));
  NAND4_X1   g5328(.A1(new_n733_), .A2(new_n726_), .A3(new_n463_), .A4(new_n550_), .ZN(new_n5378_));
  NAND4_X1   g5329(.A1(new_n5377_), .A2(new_n5375_), .A3(new_n4226_), .A4(new_n5378_), .ZN(new_n5379_));
  NOR4_X1    g5330(.A1(new_n3734_), .A2(new_n5379_), .A3(new_n2520_), .A4(new_n353_), .ZN(new_n5380_));
  NAND3_X1   g5331(.A1(new_n5274_), .A2(new_n5331_), .A3(new_n5328_), .ZN(new_n5381_));
  NAND3_X1   g5332(.A1(new_n5334_), .A2(new_n5320_), .A3(new_n5327_), .ZN(new_n5382_));
  AOI21_X1   g5333(.A1(new_n5382_), .A2(new_n5381_), .B(new_n5380_), .ZN(new_n5383_));
  INV_X1     g5334(.I(new_n5380_), .ZN(new_n5384_));
  NOR3_X1    g5335(.A1(new_n5334_), .A2(new_n5320_), .A3(new_n5327_), .ZN(new_n5385_));
  NOR3_X1    g5336(.A1(new_n5274_), .A2(new_n5331_), .A3(new_n5328_), .ZN(new_n5386_));
  NOR3_X1    g5337(.A1(new_n5385_), .A2(new_n5386_), .A3(new_n5384_), .ZN(new_n5387_));
  OAI21_X1   g5338(.A1(new_n5387_), .A2(new_n5383_), .B(new_n5373_), .ZN(new_n5388_));
  INV_X1     g5339(.I(new_n5373_), .ZN(new_n5389_));
  OAI21_X1   g5340(.A1(new_n5385_), .A2(new_n5386_), .B(new_n5384_), .ZN(new_n5390_));
  NAND3_X1   g5341(.A1(new_n5382_), .A2(new_n5381_), .A3(new_n5380_), .ZN(new_n5391_));
  NAND3_X1   g5342(.A1(new_n5390_), .A2(new_n5391_), .A3(new_n5389_), .ZN(new_n5392_));
  NAND2_X1   g5343(.A1(new_n5388_), .A2(new_n5392_), .ZN(new_n5393_));
  NOR3_X1    g5344(.A1(new_n5342_), .A2(new_n5333_), .A3(new_n5337_), .ZN(new_n5394_));
  NOR2_X1    g5345(.A1(new_n5394_), .A2(new_n4585_), .ZN(new_n5395_));
  XOR2_X1    g5346(.A1(new_n5393_), .A2(new_n5395_), .Z(\sin[13] ));
  NAND3_X1   g5347(.A1(new_n5319_), .A2(new_n5317_), .A3(new_n5328_), .ZN(new_n5397_));
  OAI21_X1   g5348(.A1(new_n5373_), .A2(new_n5380_), .B(new_n5397_), .ZN(new_n5398_));
  NAND2_X1   g5349(.A1(new_n5397_), .A2(new_n5389_), .ZN(new_n5399_));
  NAND3_X1   g5350(.A1(new_n5331_), .A2(new_n5328_), .A3(new_n5373_), .ZN(new_n5400_));
  AOI21_X1   g5351(.A1(new_n5399_), .A2(new_n5400_), .B(new_n5380_), .ZN(new_n5401_));
  AOI21_X1   g5352(.A1(new_n5331_), .A2(new_n5328_), .B(new_n5373_), .ZN(new_n5402_));
  NOR2_X1    g5353(.A1(new_n5397_), .A2(new_n5389_), .ZN(new_n5403_));
  NOR3_X1    g5354(.A1(new_n5403_), .A2(new_n5402_), .A3(new_n5384_), .ZN(new_n5404_));
  OAI21_X1   g5355(.A1(new_n5404_), .A2(new_n5401_), .B(new_n5333_), .ZN(new_n5405_));
  INV_X1     g5356(.I(new_n5367_), .ZN(new_n5406_));
  INV_X1     g5357(.I(new_n5371_), .ZN(new_n5407_));
  OAI21_X1   g5358(.A1(new_n5313_), .A2(new_n5406_), .B(new_n5407_), .ZN(new_n5408_));
  NAND2_X1   g5359(.A1(new_n5359_), .A2(new_n5364_), .ZN(new_n5409_));
  NAND2_X1   g5360(.A1(new_n5408_), .A2(new_n5409_), .ZN(new_n5410_));
  AOI21_X1   g5361(.A1(new_n5285_), .A2(new_n5345_), .B(new_n5354_), .ZN(new_n5411_));
  NOR2_X1    g5362(.A1(new_n5411_), .A2(new_n5356_), .ZN(new_n5412_));
  NAND2_X1   g5363(.A1(new_n4131_), .A2(new_n2795_), .ZN(new_n5413_));
  NAND2_X1   g5364(.A1(new_n4028_), .A2(new_n2829_), .ZN(new_n5414_));
  NAND4_X1   g5365(.A1(new_n4376_), .A2(new_n2824_), .A3(new_n5413_), .A4(new_n5414_), .ZN(new_n5415_));
  XOR2_X1    g5366(.A1(new_n5415_), .A2(new_n659_), .Z(new_n5416_));
  NOR2_X1    g5367(.A1(new_n3894_), .A2(new_n659_), .ZN(new_n5417_));
  NOR3_X1    g5368(.A1(new_n3414_), .A2(new_n576_), .A3(new_n658_), .ZN(new_n5418_));
  XOR2_X1    g5369(.A1(new_n5417_), .A2(new_n5418_), .Z(new_n5419_));
  NOR2_X1    g5370(.A1(new_n5416_), .A2(new_n5419_), .ZN(new_n5420_));
  XNOR2_X1   g5371(.A1(new_n5417_), .A2(new_n5418_), .ZN(new_n5421_));
  INV_X1     g5372(.I(new_n5421_), .ZN(new_n5422_));
  AOI21_X1   g5373(.A1(new_n5416_), .A2(new_n5422_), .B(new_n5420_), .ZN(new_n5423_));
  XOR2_X1    g5374(.A1(new_n5412_), .A2(new_n5423_), .Z(new_n5424_));
  INV_X1     g5375(.I(new_n5424_), .ZN(new_n5425_));
  NAND2_X1   g5376(.A1(new_n5410_), .A2(new_n5425_), .ZN(new_n5426_));
  INV_X1     g5377(.I(new_n5409_), .ZN(new_n5427_));
  NOR2_X1    g5378(.A1(new_n5372_), .A2(new_n5427_), .ZN(new_n5428_));
  INV_X1     g5379(.I(new_n5423_), .ZN(new_n5429_));
  XOR2_X1    g5380(.A1(new_n5412_), .A2(new_n5429_), .Z(new_n5430_));
  INV_X1     g5381(.I(new_n5430_), .ZN(new_n5431_));
  NAND2_X1   g5382(.A1(new_n5428_), .A2(new_n5431_), .ZN(new_n5432_));
  NAND4_X1   g5383(.A1(new_n2424_), .A2(new_n392_), .A3(new_n2395_), .A4(new_n3404_), .ZN(new_n5433_));
  NOR4_X1    g5384(.A1(new_n293_), .A2(new_n189_), .A3(new_n424_), .A4(new_n603_), .ZN(new_n5434_));
  NAND3_X1   g5385(.A1(new_n359_), .A2(new_n288_), .A3(new_n634_), .ZN(new_n5435_));
  NOR4_X1    g5386(.A1(new_n5433_), .A2(new_n1067_), .A3(new_n5434_), .A4(new_n5435_), .ZN(new_n5436_));
  INV_X1     g5387(.I(new_n5436_), .ZN(new_n5437_));
  NOR4_X1    g5388(.A1(new_n5437_), .A2(new_n2296_), .A3(new_n1026_), .A4(new_n1094_), .ZN(new_n5438_));
  INV_X1     g5389(.I(new_n5438_), .ZN(new_n5439_));
  NAND3_X1   g5390(.A1(new_n5432_), .A2(new_n5426_), .A3(new_n5439_), .ZN(new_n5440_));
  NOR2_X1    g5391(.A1(new_n5428_), .A2(new_n5424_), .ZN(new_n5441_));
  NOR2_X1    g5392(.A1(new_n5410_), .A2(new_n5430_), .ZN(new_n5442_));
  OAI21_X1   g5393(.A1(new_n5441_), .A2(new_n5442_), .B(new_n5438_), .ZN(new_n5443_));
  NAND2_X1   g5394(.A1(new_n5443_), .A2(new_n5440_), .ZN(new_n5444_));
  NAND2_X1   g5395(.A1(new_n5405_), .A2(new_n5444_), .ZN(new_n5445_));
  NAND3_X1   g5396(.A1(new_n5334_), .A2(new_n5336_), .A3(new_n5335_), .ZN(new_n5446_));
  OAI21_X1   g5397(.A1(new_n5403_), .A2(new_n5402_), .B(new_n5384_), .ZN(new_n5447_));
  NAND3_X1   g5398(.A1(new_n5399_), .A2(new_n5400_), .A3(new_n5380_), .ZN(new_n5448_));
  AOI21_X1   g5399(.A1(new_n5447_), .A2(new_n5448_), .B(new_n5446_), .ZN(new_n5449_));
  NOR3_X1    g5400(.A1(new_n5441_), .A2(new_n5442_), .A3(new_n5438_), .ZN(new_n5450_));
  AOI21_X1   g5401(.A1(new_n5432_), .A2(new_n5426_), .B(new_n5439_), .ZN(new_n5451_));
  NOR2_X1    g5402(.A1(new_n5451_), .A2(new_n5450_), .ZN(new_n5452_));
  NAND2_X1   g5403(.A1(new_n5449_), .A2(new_n5452_), .ZN(new_n5453_));
  AOI21_X1   g5404(.A1(new_n5453_), .A2(new_n5445_), .B(new_n5398_), .ZN(new_n5454_));
  AOI22_X1   g5405(.A1(new_n5331_), .A2(new_n5328_), .B1(new_n5389_), .B2(new_n5384_), .ZN(new_n5455_));
  NAND2_X1   g5406(.A1(new_n5449_), .A2(new_n5444_), .ZN(new_n5456_));
  NAND2_X1   g5407(.A1(new_n5405_), .A2(new_n5452_), .ZN(new_n5457_));
  AOI21_X1   g5408(.A1(new_n5456_), .A2(new_n5457_), .B(new_n5455_), .ZN(new_n5458_));
  NOR2_X1    g5409(.A1(new_n5454_), .A2(new_n5458_), .ZN(new_n5459_));
  NAND3_X1   g5410(.A1(new_n5388_), .A2(new_n5394_), .A3(new_n5392_), .ZN(new_n5460_));
  NAND2_X1   g5411(.A1(new_n5460_), .A2(new_n4102_), .ZN(new_n5461_));
  XOR2_X1    g5412(.A1(new_n5459_), .A2(new_n5461_), .Z(\sin[14] ));
  AOI21_X1   g5413(.A1(new_n5390_), .A2(new_n5391_), .B(new_n5389_), .ZN(new_n5463_));
  NOR3_X1    g5414(.A1(new_n5387_), .A2(new_n5383_), .A3(new_n5373_), .ZN(new_n5464_));
  NAND4_X1   g5415(.A1(new_n5338_), .A2(new_n5339_), .A3(new_n5269_), .A4(new_n5341_), .ZN(new_n5465_));
  NOR3_X1    g5416(.A1(new_n5464_), .A2(new_n5465_), .A3(new_n5463_), .ZN(new_n5466_));
  AOI21_X1   g5417(.A1(new_n5459_), .A2(new_n5466_), .B(new_n4585_), .ZN(new_n5467_));
  XOR2_X1    g5418(.A1(new_n5455_), .A2(new_n5444_), .Z(new_n5468_));
  INV_X1     g5419(.I(new_n4439_), .ZN(new_n5469_));
  OAI22_X1   g5420(.A1(new_n5469_), .A2(new_n2796_), .B1(new_n2830_), .B2(new_n4129_), .ZN(new_n5470_));
  NAND2_X1   g5421(.A1(new_n4109_), .A2(new_n658_), .ZN(new_n5471_));
  XOR2_X1    g5422(.A1(new_n5470_), .A2(new_n5471_), .Z(new_n5472_));
  INV_X1     g5423(.I(new_n5417_), .ZN(new_n5473_));
  INV_X1     g5424(.I(new_n5418_), .ZN(new_n5474_));
  OAI21_X1   g5425(.A1(new_n5417_), .A2(new_n5418_), .B(new_n5416_), .ZN(new_n5475_));
  OAI21_X1   g5426(.A1(new_n5473_), .A2(new_n5474_), .B(new_n5475_), .ZN(new_n5476_));
  XOR2_X1    g5427(.A1(new_n5476_), .A2(new_n5472_), .Z(new_n5477_));
  INV_X1     g5428(.I(new_n5412_), .ZN(new_n5478_));
  NAND3_X1   g5429(.A1(new_n5408_), .A2(new_n5409_), .A3(new_n5478_), .ZN(new_n5479_));
  OAI21_X1   g5430(.A1(new_n5372_), .A2(new_n5427_), .B(new_n5412_), .ZN(new_n5480_));
  NAND2_X1   g5431(.A1(new_n5480_), .A2(new_n5479_), .ZN(new_n5481_));
  NAND3_X1   g5432(.A1(new_n5481_), .A2(new_n5423_), .A3(new_n5477_), .ZN(new_n5482_));
  INV_X1     g5433(.I(new_n5477_), .ZN(new_n5483_));
  NOR3_X1    g5434(.A1(new_n5372_), .A2(new_n5427_), .A3(new_n5412_), .ZN(new_n5484_));
  AOI21_X1   g5435(.A1(new_n5408_), .A2(new_n5409_), .B(new_n5478_), .ZN(new_n5485_));
  OAI21_X1   g5436(.A1(new_n5484_), .A2(new_n5485_), .B(new_n5423_), .ZN(new_n5486_));
  NAND2_X1   g5437(.A1(new_n5486_), .A2(new_n5483_), .ZN(new_n5487_));
  NOR2_X1    g5438(.A1(new_n5428_), .A2(new_n5412_), .ZN(new_n5488_));
  NAND3_X1   g5439(.A1(new_n5487_), .A2(new_n5482_), .A3(new_n5488_), .ZN(new_n5489_));
  NOR2_X1    g5440(.A1(new_n5486_), .A2(new_n5483_), .ZN(new_n5490_));
  AOI21_X1   g5441(.A1(new_n5481_), .A2(new_n5423_), .B(new_n5477_), .ZN(new_n5491_));
  INV_X1     g5442(.I(new_n5488_), .ZN(new_n5492_));
  OAI21_X1   g5443(.A1(new_n5490_), .A2(new_n5491_), .B(new_n5492_), .ZN(new_n5493_));
  NOR4_X1    g5444(.A1(new_n858_), .A2(new_n301_), .A3(new_n305_), .A4(new_n376_), .ZN(new_n5494_));
  NOR3_X1    g5445(.A1(new_n1702_), .A2(new_n620_), .A3(new_n393_), .ZN(new_n5495_));
  INV_X1     g5446(.I(new_n289_), .ZN(new_n5496_));
  NAND4_X1   g5447(.A1(new_n1086_), .A2(new_n5496_), .A3(new_n503_), .A4(new_n439_), .ZN(new_n5497_));
  NOR4_X1    g5448(.A1(new_n5497_), .A2(new_n5325_), .A3(new_n935_), .A4(new_n5495_), .ZN(new_n5498_));
  NAND3_X1   g5449(.A1(new_n2428_), .A2(new_n5494_), .A3(new_n5498_), .ZN(new_n5499_));
  AOI21_X1   g5450(.A1(new_n5493_), .A2(new_n5489_), .B(new_n5499_), .ZN(new_n5500_));
  NOR3_X1    g5451(.A1(new_n5490_), .A2(new_n5491_), .A3(new_n5492_), .ZN(new_n5501_));
  AOI21_X1   g5452(.A1(new_n5487_), .A2(new_n5482_), .B(new_n5488_), .ZN(new_n5502_));
  INV_X1     g5453(.I(new_n5499_), .ZN(new_n5503_));
  NOR3_X1    g5454(.A1(new_n5501_), .A2(new_n5502_), .A3(new_n5503_), .ZN(new_n5504_));
  OAI22_X1   g5455(.A1(new_n5468_), .A2(new_n5405_), .B1(new_n5500_), .B2(new_n5504_), .ZN(new_n5505_));
  NAND2_X1   g5456(.A1(new_n5398_), .A2(new_n5452_), .ZN(new_n5506_));
  NAND2_X1   g5457(.A1(new_n5455_), .A2(new_n5444_), .ZN(new_n5507_));
  NAND2_X1   g5458(.A1(new_n5506_), .A2(new_n5507_), .ZN(new_n5508_));
  OAI21_X1   g5459(.A1(new_n5501_), .A2(new_n5502_), .B(new_n5503_), .ZN(new_n5509_));
  NAND3_X1   g5460(.A1(new_n5493_), .A2(new_n5489_), .A3(new_n5499_), .ZN(new_n5510_));
  NAND4_X1   g5461(.A1(new_n5449_), .A2(new_n5508_), .A3(new_n5509_), .A4(new_n5510_), .ZN(new_n5511_));
  NAND2_X1   g5462(.A1(new_n5505_), .A2(new_n5511_), .ZN(new_n5512_));
  NAND2_X1   g5463(.A1(new_n5467_), .A2(new_n5512_), .ZN(new_n5513_));
  NAND2_X1   g5464(.A1(new_n5449_), .A2(new_n5508_), .ZN(new_n5514_));
  NOR2_X1    g5465(.A1(new_n5504_), .A2(new_n5500_), .ZN(new_n5515_));
  XOR2_X1    g5466(.A1(new_n5514_), .A2(new_n5515_), .Z(new_n5516_));
  OAI21_X1   g5467(.A1(new_n5467_), .A2(new_n5516_), .B(new_n5513_), .ZN(\sin[15] ));
  NOR3_X1    g5468(.A1(new_n5501_), .A2(new_n5502_), .A3(new_n5499_), .ZN(new_n5518_));
  NOR2_X1    g5469(.A1(new_n5470_), .A2(new_n4023_), .ZN(new_n5519_));
  NAND2_X1   g5470(.A1(new_n5470_), .A2(new_n4023_), .ZN(new_n5520_));
  NAND2_X1   g5471(.A1(new_n5520_), .A2(new_n4109_), .ZN(new_n5521_));
  OAI21_X1   g5472(.A1(new_n5521_), .A2(new_n5519_), .B(new_n658_), .ZN(new_n5522_));
  XNOR2_X1   g5473(.A1(new_n5522_), .A2(new_n5470_), .ZN(new_n5523_));
  NAND3_X1   g5474(.A1(new_n5410_), .A2(new_n5478_), .A3(new_n5477_), .ZN(new_n5524_));
  NAND3_X1   g5475(.A1(new_n5481_), .A2(new_n5524_), .A3(new_n5423_), .ZN(new_n5525_));
  INV_X1     g5476(.I(new_n5476_), .ZN(new_n5526_));
  NAND2_X1   g5477(.A1(new_n5526_), .A2(new_n5472_), .ZN(new_n5527_));
  NAND3_X1   g5478(.A1(new_n5525_), .A2(new_n5523_), .A3(new_n5527_), .ZN(new_n5528_));
  INV_X1     g5479(.I(new_n5523_), .ZN(new_n5529_));
  NOR3_X1    g5480(.A1(new_n5428_), .A2(new_n5412_), .A3(new_n5483_), .ZN(new_n5530_));
  OAI21_X1   g5481(.A1(new_n5486_), .A2(new_n5530_), .B(new_n5527_), .ZN(new_n5531_));
  NAND2_X1   g5482(.A1(new_n5531_), .A2(new_n5529_), .ZN(new_n5532_));
  NOR2_X1    g5483(.A1(new_n4131_), .A2(new_n3895_), .ZN(new_n5533_));
  NOR2_X1    g5484(.A1(new_n4129_), .A2(new_n3894_), .ZN(new_n5534_));
  OAI21_X1   g5485(.A1(new_n5533_), .A2(new_n5534_), .B(new_n658_), .ZN(new_n5535_));
  INV_X1     g5486(.I(new_n5535_), .ZN(new_n5536_));
  NAND3_X1   g5487(.A1(new_n5532_), .A2(new_n5528_), .A3(new_n5536_), .ZN(new_n5537_));
  NOR2_X1    g5488(.A1(new_n5531_), .A2(new_n5529_), .ZN(new_n5538_));
  AOI21_X1   g5489(.A1(new_n5525_), .A2(new_n5527_), .B(new_n5523_), .ZN(new_n5539_));
  OAI21_X1   g5490(.A1(new_n5538_), .A2(new_n5539_), .B(new_n5535_), .ZN(new_n5540_));
  INV_X1     g5491(.I(new_n1680_), .ZN(new_n5541_));
  NAND3_X1   g5492(.A1(new_n403_), .A2(new_n455_), .A3(new_n556_), .ZN(new_n5542_));
  NOR4_X1    g5493(.A1(new_n5542_), .A2(new_n369_), .A3(new_n603_), .A4(new_n878_), .ZN(new_n5543_));
  NAND4_X1   g5494(.A1(new_n5543_), .A2(new_n3770_), .A3(new_n1657_), .A4(new_n5375_), .ZN(new_n5544_));
  NOR3_X1    g5495(.A1(new_n5541_), .A2(new_n3736_), .A3(new_n5544_), .ZN(new_n5545_));
  INV_X1     g5496(.I(new_n5545_), .ZN(new_n5546_));
  AOI21_X1   g5497(.A1(new_n5540_), .A2(new_n5537_), .B(new_n5546_), .ZN(new_n5547_));
  NOR3_X1    g5498(.A1(new_n5538_), .A2(new_n5539_), .A3(new_n5535_), .ZN(new_n5548_));
  AOI21_X1   g5499(.A1(new_n5532_), .A2(new_n5528_), .B(new_n5536_), .ZN(new_n5549_));
  NOR3_X1    g5500(.A1(new_n5548_), .A2(new_n5549_), .A3(new_n5545_), .ZN(new_n5550_));
  OAI21_X1   g5501(.A1(new_n5550_), .A2(new_n5547_), .B(new_n5518_), .ZN(new_n5551_));
  NAND3_X1   g5502(.A1(new_n5493_), .A2(new_n5489_), .A3(new_n5503_), .ZN(new_n5552_));
  NOR3_X1    g5503(.A1(new_n5548_), .A2(new_n5549_), .A3(new_n5546_), .ZN(new_n5553_));
  AOI21_X1   g5504(.A1(new_n5540_), .A2(new_n5537_), .B(new_n5545_), .ZN(new_n5554_));
  OAI21_X1   g5505(.A1(new_n5553_), .A2(new_n5554_), .B(new_n5552_), .ZN(new_n5555_));
  NAND2_X1   g5506(.A1(new_n5551_), .A2(new_n5555_), .ZN(new_n5556_));
  XOR2_X1    g5507(.A1(new_n5556_), .A2(new_n5511_), .Z(new_n5557_));
  AOI22_X1   g5508(.A1(new_n5449_), .A2(new_n5508_), .B1(new_n5509_), .B2(new_n5510_), .ZN(new_n5558_));
  NOR4_X1    g5509(.A1(new_n5468_), .A2(new_n5405_), .A3(new_n5500_), .A4(new_n5504_), .ZN(new_n5559_));
  NOR2_X1    g5510(.A1(new_n5559_), .A2(new_n5558_), .ZN(new_n5560_));
  NOR4_X1    g5511(.A1(new_n5560_), .A2(new_n5454_), .A3(new_n5460_), .A4(new_n5458_), .ZN(new_n5561_));
  NOR2_X1    g5512(.A1(new_n5561_), .A2(new_n4585_), .ZN(new_n5562_));
  XOR2_X1    g5513(.A1(new_n5557_), .A2(new_n5562_), .Z(\sin[16] ));
  NOR2_X1    g5514(.A1(new_n5548_), .A2(new_n5549_), .ZN(new_n5564_));
  INV_X1     g5515(.I(new_n3380_), .ZN(new_n5565_));
  NOR2_X1    g5516(.A1(new_n869_), .A2(new_n534_), .ZN(new_n5566_));
  NAND4_X1   g5517(.A1(new_n5566_), .A2(new_n264_), .A3(new_n719_), .A4(new_n714_), .ZN(new_n5567_));
  INV_X1     g5518(.I(new_n5567_), .ZN(new_n5568_));
  NOR4_X1    g5519(.A1(new_n212_), .A2(new_n3382_), .A3(new_n192_), .A4(new_n747_), .ZN(new_n5569_));
  AND4_X2    g5520(.A1(new_n421_), .A2(new_n5568_), .A3(new_n739_), .A4(new_n5569_), .Z(new_n5570_));
  INV_X1     g5521(.I(new_n5570_), .ZN(new_n5571_));
  NOR3_X1    g5522(.A1(new_n5565_), .A2(new_n5571_), .A3(new_n466_), .ZN(new_n5572_));
  NOR3_X1    g5523(.A1(new_n5564_), .A2(new_n5552_), .A3(new_n5572_), .ZN(new_n5573_));
  NAND2_X1   g5524(.A1(new_n5540_), .A2(new_n5537_), .ZN(new_n5574_));
  INV_X1     g5525(.I(new_n5572_), .ZN(new_n5575_));
  AOI21_X1   g5526(.A1(new_n5574_), .A2(new_n5518_), .B(new_n5575_), .ZN(new_n5576_));
  AOI21_X1   g5527(.A1(new_n5537_), .A2(new_n5540_), .B(new_n5518_), .ZN(new_n5577_));
  NOR3_X1    g5528(.A1(new_n5552_), .A2(new_n5548_), .A3(new_n5549_), .ZN(new_n5578_));
  NOR2_X1    g5529(.A1(new_n5577_), .A2(new_n5578_), .ZN(new_n5579_));
  NOR4_X1    g5530(.A1(new_n5579_), .A2(new_n5546_), .A3(new_n5573_), .A4(new_n5576_), .ZN(new_n5580_));
  NAND3_X1   g5531(.A1(new_n5574_), .A2(new_n5518_), .A3(new_n5575_), .ZN(new_n5581_));
  OAI21_X1   g5532(.A1(new_n5564_), .A2(new_n5552_), .B(new_n5572_), .ZN(new_n5582_));
  OAI21_X1   g5533(.A1(new_n5548_), .A2(new_n5549_), .B(new_n5552_), .ZN(new_n5583_));
  NAND3_X1   g5534(.A1(new_n5518_), .A2(new_n5540_), .A3(new_n5537_), .ZN(new_n5584_));
  NAND2_X1   g5535(.A1(new_n5583_), .A2(new_n5584_), .ZN(new_n5585_));
  AOI22_X1   g5536(.A1(new_n5585_), .A2(new_n5545_), .B1(new_n5582_), .B2(new_n5581_), .ZN(new_n5586_));
  NOR2_X1    g5537(.A1(new_n5580_), .A2(new_n5586_), .ZN(new_n5587_));
  NAND3_X1   g5538(.A1(new_n5551_), .A2(new_n5555_), .A3(new_n5559_), .ZN(new_n5588_));
  NAND2_X1   g5539(.A1(new_n5587_), .A2(new_n5588_), .ZN(new_n5589_));
  OAI21_X1   g5540(.A1(new_n5548_), .A2(new_n5549_), .B(new_n5545_), .ZN(new_n5590_));
  NAND3_X1   g5541(.A1(new_n5540_), .A2(new_n5537_), .A3(new_n5546_), .ZN(new_n5591_));
  AOI21_X1   g5542(.A1(new_n5590_), .A2(new_n5591_), .B(new_n5552_), .ZN(new_n5592_));
  NAND3_X1   g5543(.A1(new_n5540_), .A2(new_n5537_), .A3(new_n5545_), .ZN(new_n5593_));
  OAI21_X1   g5544(.A1(new_n5548_), .A2(new_n5549_), .B(new_n5546_), .ZN(new_n5594_));
  AOI21_X1   g5545(.A1(new_n5594_), .A2(new_n5593_), .B(new_n5518_), .ZN(new_n5595_));
  NOR3_X1    g5546(.A1(new_n5592_), .A2(new_n5595_), .A3(new_n5511_), .ZN(new_n5596_));
  OAI21_X1   g5547(.A1(new_n5580_), .A2(new_n5586_), .B(new_n5596_), .ZN(new_n5597_));
  NAND2_X1   g5548(.A1(new_n5589_), .A2(new_n5597_), .ZN(new_n5598_));
  NOR2_X1    g5549(.A1(new_n5449_), .A2(new_n5452_), .ZN(new_n5599_));
  NOR2_X1    g5550(.A1(new_n5405_), .A2(new_n5444_), .ZN(new_n5600_));
  OAI21_X1   g5551(.A1(new_n5599_), .A2(new_n5600_), .B(new_n5455_), .ZN(new_n5601_));
  NOR2_X1    g5552(.A1(new_n5405_), .A2(new_n5452_), .ZN(new_n5602_));
  NOR2_X1    g5553(.A1(new_n5449_), .A2(new_n5444_), .ZN(new_n5603_));
  OAI21_X1   g5554(.A1(new_n5603_), .A2(new_n5602_), .B(new_n5398_), .ZN(new_n5604_));
  NAND4_X1   g5555(.A1(new_n5512_), .A2(new_n5466_), .A3(new_n5601_), .A4(new_n5604_), .ZN(new_n5605_));
  OAI21_X1   g5556(.A1(new_n5557_), .A2(new_n5605_), .B(new_n4102_), .ZN(new_n5606_));
  XOR2_X1    g5557(.A1(new_n5606_), .A2(new_n5598_), .Z(\sin[17] ));
  NAND4_X1   g5558(.A1(new_n5585_), .A2(new_n5582_), .A3(new_n5581_), .A4(new_n5545_), .ZN(new_n5608_));
  OAI22_X1   g5559(.A1(new_n5579_), .A2(new_n5546_), .B1(new_n5573_), .B2(new_n5576_), .ZN(new_n5609_));
  AOI21_X1   g5560(.A1(new_n5609_), .A2(new_n5608_), .B(new_n5588_), .ZN(new_n5610_));
  NOR2_X1    g5561(.A1(new_n2290_), .A2(new_n531_), .ZN(new_n5611_));
  NAND2_X1   g5562(.A1(new_n453_), .A2(new_n458_), .ZN(new_n5612_));
  NOR4_X1    g5563(.A1(new_n5612_), .A2(new_n3382_), .A3(new_n437_), .A4(new_n1091_), .ZN(new_n5613_));
  NAND4_X1   g5564(.A1(new_n5611_), .A2(new_n5613_), .A3(new_n2516_), .A4(new_n885_), .ZN(new_n5614_));
  NOR3_X1    g5565(.A1(new_n5614_), .A2(new_n952_), .A3(new_n3748_), .ZN(new_n5615_));
  AND2_X2    g5566(.A1(new_n5615_), .A2(new_n436_), .Z(new_n5616_));
  INV_X1     g5567(.I(new_n5616_), .ZN(new_n5617_));
  NAND2_X1   g5568(.A1(new_n5591_), .A2(new_n5518_), .ZN(new_n5618_));
  NOR2_X1    g5569(.A1(new_n5547_), .A2(new_n5572_), .ZN(new_n5619_));
  NAND2_X1   g5570(.A1(new_n5619_), .A2(new_n5618_), .ZN(new_n5620_));
  NOR2_X1    g5571(.A1(new_n5620_), .A2(new_n5617_), .ZN(new_n5621_));
  AOI21_X1   g5572(.A1(new_n5619_), .A2(new_n5618_), .B(new_n5616_), .ZN(new_n5622_));
  NOR3_X1    g5573(.A1(new_n5610_), .A2(new_n5621_), .A3(new_n5622_), .ZN(new_n5623_));
  AOI21_X1   g5574(.A1(new_n5610_), .A2(new_n5621_), .B(new_n5623_), .ZN(new_n5624_));
  OAI21_X1   g5575(.A1(new_n5580_), .A2(new_n5586_), .B(new_n5511_), .ZN(new_n5625_));
  NAND3_X1   g5576(.A1(new_n5609_), .A2(new_n5608_), .A3(new_n5559_), .ZN(new_n5626_));
  OAI21_X1   g5577(.A1(new_n5592_), .A2(new_n5595_), .B(new_n5511_), .ZN(new_n5627_));
  NAND2_X1   g5578(.A1(new_n5588_), .A2(new_n5627_), .ZN(new_n5628_));
  NAND4_X1   g5579(.A1(new_n5625_), .A2(new_n5626_), .A3(new_n5628_), .A4(new_n5561_), .ZN(new_n5629_));
  NAND2_X1   g5580(.A1(new_n5629_), .A2(new_n4102_), .ZN(new_n5630_));
  XOR2_X1    g5581(.A1(new_n5624_), .A2(new_n5630_), .Z(\sin[18] ));
  NOR2_X1    g5582(.A1(new_n5550_), .A2(new_n5552_), .ZN(new_n5632_));
  NAND2_X1   g5583(.A1(new_n5590_), .A2(new_n5575_), .ZN(new_n5633_));
  NOR2_X1    g5584(.A1(new_n5632_), .A2(new_n5633_), .ZN(new_n5634_));
  NAND2_X1   g5585(.A1(new_n5634_), .A2(new_n5616_), .ZN(new_n5635_));
  OAI21_X1   g5586(.A1(new_n5632_), .A2(new_n5633_), .B(new_n5617_), .ZN(new_n5636_));
  NAND4_X1   g5587(.A1(new_n213_), .A2(new_n455_), .A3(new_n468_), .A4(new_n363_), .ZN(new_n5637_));
  NAND4_X1   g5588(.A1(new_n4225_), .A2(new_n1083_), .A3(new_n419_), .A4(new_n646_), .ZN(new_n5638_));
  NAND2_X1   g5589(.A1(new_n4749_), .A2(new_n5638_), .ZN(new_n5639_));
  NOR4_X1    g5590(.A1(new_n819_), .A2(new_n2547_), .A3(new_n5637_), .A4(new_n5639_), .ZN(new_n5640_));
  NAND2_X1   g5591(.A1(new_n5640_), .A2(new_n5494_), .ZN(new_n5641_));
  NOR2_X1    g5592(.A1(new_n5616_), .A2(new_n5641_), .ZN(new_n5642_));
  AOI22_X1   g5593(.A1(new_n5636_), .A2(new_n5641_), .B1(new_n5620_), .B2(new_n5642_), .ZN(new_n5643_));
  AOI21_X1   g5594(.A1(new_n5610_), .A2(new_n5635_), .B(new_n5643_), .ZN(new_n5644_));
  INV_X1     g5595(.I(new_n5641_), .ZN(new_n5645_));
  INV_X1     g5596(.I(new_n5642_), .ZN(new_n5646_));
  OAI22_X1   g5597(.A1(new_n5622_), .A2(new_n5645_), .B1(new_n5634_), .B2(new_n5646_), .ZN(new_n5647_));
  NOR3_X1    g5598(.A1(new_n5597_), .A2(new_n5647_), .A3(new_n5621_), .ZN(new_n5648_));
  NOR2_X1    g5599(.A1(new_n5644_), .A2(new_n5648_), .ZN(new_n5649_));
  NAND2_X1   g5600(.A1(new_n5609_), .A2(new_n5608_), .ZN(new_n5650_));
  AOI22_X1   g5601(.A1(new_n5650_), .A2(new_n5596_), .B1(new_n5616_), .B2(new_n5634_), .ZN(new_n5651_));
  NOR2_X1    g5602(.A1(new_n5629_), .A2(new_n5651_), .ZN(new_n5652_));
  NOR2_X1    g5603(.A1(new_n5652_), .A2(new_n4585_), .ZN(new_n5653_));
  NAND2_X1   g5604(.A1(new_n5649_), .A2(new_n4102_), .ZN(new_n5654_));
  OAI22_X1   g5605(.A1(new_n5652_), .A2(new_n5654_), .B1(new_n5653_), .B2(new_n5649_), .ZN(\sin[19] ));
  NAND3_X1   g5606(.A1(new_n193_), .A2(new_n598_), .A3(new_n362_), .ZN(new_n5656_));
  NOR4_X1    g5607(.A1(new_n563_), .A2(new_n324_), .A3(new_n472_), .A4(new_n832_), .ZN(new_n5657_));
  NAND3_X1   g5608(.A1(new_n2545_), .A2(new_n619_), .A3(new_n452_), .ZN(new_n5658_));
  NOR4_X1    g5609(.A1(new_n649_), .A2(new_n5656_), .A3(new_n5657_), .A4(new_n5658_), .ZN(new_n5659_));
  NAND3_X1   g5610(.A1(new_n5058_), .A2(new_n1076_), .A3(new_n5659_), .ZN(new_n5660_));
  INV_X1     g5611(.I(new_n5660_), .ZN(new_n5661_));
  NOR2_X1    g5612(.A1(new_n5616_), .A2(new_n5645_), .ZN(new_n5662_));
  NOR3_X1    g5613(.A1(new_n5620_), .A2(new_n5661_), .A3(new_n5662_), .ZN(new_n5663_));
  NOR4_X1    g5614(.A1(new_n5597_), .A2(new_n5621_), .A3(new_n5643_), .A4(new_n5663_), .ZN(new_n5664_));
  NOR3_X1    g5615(.A1(new_n5597_), .A2(new_n5621_), .A3(new_n5643_), .ZN(new_n5665_));
  INV_X1     g5616(.I(new_n5662_), .ZN(new_n5666_));
  AOI21_X1   g5617(.A1(new_n5634_), .A2(new_n5666_), .B(new_n5660_), .ZN(new_n5667_));
  NOR2_X1    g5618(.A1(new_n5667_), .A2(new_n5663_), .ZN(new_n5668_));
  INV_X1     g5619(.I(new_n5668_), .ZN(new_n5669_));
  NOR3_X1    g5620(.A1(new_n5664_), .A2(new_n5665_), .A3(new_n5669_), .ZN(new_n5670_));
  AOI21_X1   g5621(.A1(new_n5649_), .A2(new_n5652_), .B(new_n4585_), .ZN(new_n5671_));
  XOR2_X1    g5622(.A1(new_n5671_), .A2(new_n5670_), .Z(\sin[20] ));
  NOR3_X1    g5623(.A1(new_n5661_), .A2(new_n5616_), .A3(new_n5645_), .ZN(new_n5673_));
  INV_X1     g5624(.I(new_n2474_), .ZN(new_n5674_));
  INV_X1     g5625(.I(new_n3888_), .ZN(new_n5675_));
  NOR4_X1    g5626(.A1(new_n627_), .A2(new_n414_), .A3(new_n5674_), .A4(new_n5675_), .ZN(new_n5676_));
  AOI21_X1   g5627(.A1(new_n5620_), .A2(new_n5673_), .B(new_n5676_), .ZN(new_n5677_));
  INV_X1     g5628(.I(new_n5673_), .ZN(new_n5678_));
  INV_X1     g5629(.I(new_n5676_), .ZN(new_n5679_));
  NOR3_X1    g5630(.A1(new_n5634_), .A2(new_n5678_), .A3(new_n5679_), .ZN(new_n5680_));
  NOR2_X1    g5631(.A1(new_n5680_), .A2(new_n5677_), .ZN(new_n5681_));
  NOR2_X1    g5632(.A1(new_n5664_), .A2(new_n5681_), .ZN(new_n5682_));
  NAND3_X1   g5633(.A1(new_n5634_), .A2(new_n5660_), .A3(new_n5666_), .ZN(new_n5683_));
  NAND4_X1   g5634(.A1(new_n5610_), .A2(new_n5647_), .A3(new_n5635_), .A4(new_n5683_), .ZN(new_n5684_));
  OAI21_X1   g5635(.A1(new_n5634_), .A2(new_n5678_), .B(new_n5679_), .ZN(new_n5685_));
  NAND3_X1   g5636(.A1(new_n5620_), .A2(new_n5673_), .A3(new_n5676_), .ZN(new_n5686_));
  NAND2_X1   g5637(.A1(new_n5685_), .A2(new_n5686_), .ZN(new_n5687_));
  NOR2_X1    g5638(.A1(new_n5684_), .A2(new_n5687_), .ZN(new_n5688_));
  NOR2_X1    g5639(.A1(new_n5682_), .A2(new_n5688_), .ZN(new_n5689_));
  OAI21_X1   g5640(.A1(new_n5597_), .A2(new_n5621_), .B(new_n5647_), .ZN(new_n5690_));
  NAND3_X1   g5641(.A1(new_n5610_), .A2(new_n5635_), .A3(new_n5643_), .ZN(new_n5691_));
  NAND2_X1   g5642(.A1(new_n5690_), .A2(new_n5691_), .ZN(new_n5692_));
  AOI21_X1   g5643(.A1(new_n5650_), .A2(new_n5511_), .B(new_n5605_), .ZN(new_n5693_));
  OAI22_X1   g5644(.A1(new_n5587_), .A2(new_n5588_), .B1(new_n5617_), .B2(new_n5620_), .ZN(new_n5694_));
  NAND4_X1   g5645(.A1(new_n5694_), .A2(new_n5693_), .A3(new_n5626_), .A4(new_n5628_), .ZN(new_n5695_));
  NOR3_X1    g5646(.A1(new_n5670_), .A2(new_n5695_), .A3(new_n5692_), .ZN(new_n5696_));
  NOR2_X1    g5647(.A1(new_n5696_), .A2(new_n4585_), .ZN(new_n5697_));
  NAND2_X1   g5648(.A1(new_n5689_), .A2(new_n4102_), .ZN(new_n5698_));
  OAI22_X1   g5649(.A1(new_n5697_), .A2(new_n5689_), .B1(new_n5698_), .B2(new_n5696_), .ZN(\sin[21] ));
  NOR2_X1    g5650(.A1(new_n383_), .A2(new_n637_), .ZN(new_n5700_));
  NAND2_X1   g5651(.A1(new_n628_), .A2(new_n5700_), .ZN(new_n5701_));
  NAND3_X1   g5652(.A1(new_n5664_), .A2(new_n5687_), .A3(new_n5701_), .ZN(new_n5702_));
  INV_X1     g5653(.I(new_n5701_), .ZN(new_n5703_));
  OAI21_X1   g5654(.A1(new_n5684_), .A2(new_n5681_), .B(new_n5703_), .ZN(new_n5704_));
  NOR3_X1    g5655(.A1(new_n5634_), .A2(new_n5678_), .A3(new_n5676_), .ZN(new_n5705_));
  NOR3_X1    g5656(.A1(new_n5684_), .A2(new_n5681_), .A3(new_n5705_), .ZN(new_n5706_));
  AOI21_X1   g5657(.A1(new_n5704_), .A2(new_n5702_), .B(new_n5706_), .ZN(new_n5707_));
  NAND2_X1   g5658(.A1(new_n5684_), .A2(new_n5687_), .ZN(new_n5708_));
  NAND2_X1   g5659(.A1(new_n5664_), .A2(new_n5681_), .ZN(new_n5709_));
  NAND2_X1   g5660(.A1(new_n5709_), .A2(new_n5708_), .ZN(new_n5710_));
  NAND3_X1   g5661(.A1(new_n5610_), .A2(new_n5647_), .A3(new_n5635_), .ZN(new_n5711_));
  NAND3_X1   g5662(.A1(new_n5684_), .A2(new_n5711_), .A3(new_n5668_), .ZN(new_n5712_));
  NAND3_X1   g5663(.A1(new_n5712_), .A2(new_n5649_), .A3(new_n5652_), .ZN(new_n5713_));
  OAI21_X1   g5664(.A1(new_n5713_), .A2(new_n5710_), .B(new_n4102_), .ZN(new_n5714_));
  XOR2_X1    g5665(.A1(new_n5714_), .A2(new_n5707_), .Z(\sin[22] ));
  NOR3_X1    g5666(.A1(new_n101_), .A2(\a[21] ), .A3(\a[22] ), .ZN(new_n5716_));
  INV_X1     g5667(.I(new_n5705_), .ZN(new_n5717_));
  NOR2_X1    g5668(.A1(new_n5705_), .A2(new_n5701_), .ZN(new_n5718_));
  NOR4_X1    g5669(.A1(new_n5634_), .A2(new_n5678_), .A3(new_n5676_), .A4(new_n5703_), .ZN(new_n5719_));
  OAI21_X1   g5670(.A1(new_n5718_), .A2(new_n5719_), .B(new_n5687_), .ZN(new_n5720_));
  OAI22_X1   g5671(.A1(new_n5720_), .A2(new_n5664_), .B1(new_n5703_), .B2(new_n5717_), .ZN(new_n5721_));
  NOR4_X1    g5672(.A1(new_n5684_), .A2(new_n5681_), .A3(new_n5703_), .A4(new_n5717_), .ZN(new_n5722_));
  NOR2_X1    g5673(.A1(new_n5721_), .A2(new_n5722_), .ZN(new_n5723_));
  INV_X1     g5674(.I(new_n5723_), .ZN(new_n5724_));
  NOR3_X1    g5675(.A1(new_n5707_), .A2(new_n5713_), .A3(new_n5710_), .ZN(new_n5725_));
  OAI21_X1   g5676(.A1(new_n5725_), .A2(new_n4585_), .B(new_n5724_), .ZN(new_n5726_));
  NAND2_X1   g5677(.A1(new_n5647_), .A2(new_n5635_), .ZN(new_n5727_));
  NAND2_X1   g5678(.A1(new_n5610_), .A2(new_n5683_), .ZN(new_n5728_));
  NOR4_X1    g5679(.A1(new_n5728_), .A2(new_n5727_), .A3(new_n5681_), .A4(new_n5703_), .ZN(new_n5729_));
  AOI21_X1   g5680(.A1(new_n5664_), .A2(new_n5687_), .B(new_n5701_), .ZN(new_n5730_));
  NOR2_X1    g5681(.A1(new_n5643_), .A2(new_n5621_), .ZN(new_n5731_));
  NOR2_X1    g5682(.A1(new_n5597_), .A2(new_n5663_), .ZN(new_n5732_));
  NAND4_X1   g5683(.A1(new_n5732_), .A2(new_n5731_), .A3(new_n5687_), .A4(new_n5717_), .ZN(new_n5733_));
  OAI21_X1   g5684(.A1(new_n5730_), .A2(new_n5729_), .B(new_n5733_), .ZN(new_n5734_));
  NAND3_X1   g5685(.A1(new_n5696_), .A2(new_n5734_), .A3(new_n5689_), .ZN(new_n5735_));
  NAND3_X1   g5686(.A1(new_n5735_), .A2(new_n4102_), .A3(new_n5723_), .ZN(new_n5736_));
  AOI21_X1   g5687(.A1(new_n5726_), .A2(new_n5736_), .B(new_n5716_), .ZN(\sin[23] ));
  OAI21_X1   g5688(.A1(new_n5707_), .A2(new_n5710_), .B(new_n5713_), .ZN(new_n5738_));
  NOR3_X1    g5689(.A1(new_n5713_), .A2(new_n5710_), .A3(new_n5721_), .ZN(new_n5739_));
  OR2_X2     g5690(.A1(new_n5722_), .A2(new_n5716_), .Z(new_n5740_));
  AOI21_X1   g5691(.A1(new_n5739_), .A2(new_n5734_), .B(new_n5740_), .ZN(new_n5741_));
  AOI21_X1   g5692(.A1(new_n5741_), .A2(new_n5738_), .B(new_n4585_), .ZN(\sin[24] ));
endmodule


