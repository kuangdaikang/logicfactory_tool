// Benchmark "adder" written by ABC on Fri Sep 15 11:19:37 2023

module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n403_, new_n404_, new_n405_, new_n406_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n432_, new_n433_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n470_, new_n471_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n489_, new_n490_, new_n491_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n512_, new_n513_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n553_, new_n554_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n575_, new_n576_,
    new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1024_, new_n1025_, new_n1026_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1048_, new_n1049_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1073_, new_n1074_, new_n1075_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1098_,
    new_n1099_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1122_, new_n1123_, new_n1124_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1146_,
    new_n1147_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1171_, new_n1172_, new_n1173_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1196_, new_n1197_, new_n1198_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1226_, new_n1227_,
    new_n1228_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1283_, new_n1284_, new_n1285_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1310_, new_n1311_, new_n1312_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1340_, new_n1341_,
    new_n1342_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1368_,
    new_n1369_, new_n1370_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1396_, new_n1397_, new_n1398_;
  XOR2_X1    g0000(.A1(\a[0] ), .A2(\b[0] ), .Z(\f[0] ));
  XNOR2_X1   g0001(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n387_));
  NAND2_X1   g0002(.A1(\a[0] ), .A2(\b[0] ), .ZN(new_n388_));
  XOR2_X1    g0003(.A1(new_n387_), .A2(new_n388_), .Z(\f[1] ));
  INV_X1     g0004(.I(\a[1] ), .ZN(new_n390_));
  AOI21_X1   g0005(.A1(\a[0] ), .A2(\b[0] ), .B(\b[1] ), .ZN(new_n391_));
  NAND3_X1   g0006(.A1(\a[0] ), .A2(\b[0] ), .A3(\b[1] ), .ZN(new_n392_));
  OAI21_X1   g0007(.A1(new_n390_), .A2(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1    g0008(.A1(\a[2] ), .A2(\b[2] ), .Z(new_n394_));
  XOR2_X1    g0009(.A1(new_n393_), .A2(new_n394_), .Z(\f[2] ));
  XNOR2_X1   g0010(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n396_));
  INV_X1     g0011(.I(\a[2] ), .ZN(new_n397_));
  INV_X1     g0012(.I(\b[2] ), .ZN(new_n398_));
  NOR2_X1    g0013(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1   g0014(.A1(new_n397_), .A2(new_n398_), .ZN(new_n400_));
  AOI21_X1   g0015(.A1(new_n393_), .A2(new_n400_), .B(new_n399_), .ZN(new_n401_));
  XOR2_X1    g0016(.A1(new_n401_), .A2(new_n396_), .Z(\f[3] ));
  NAND2_X1   g0017(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n403_));
  NOR2_X1    g0018(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n404_));
  OAI21_X1   g0019(.A1(new_n401_), .A2(new_n404_), .B(new_n403_), .ZN(new_n405_));
  XOR2_X1    g0020(.A1(new_n405_), .A2(\b[4] ), .Z(new_n406_));
  XOR2_X1    g0021(.A1(new_n406_), .A2(\a[4] ), .Z(\f[4] ));
  NOR2_X1    g0022(.A1(new_n405_), .A2(\b[4] ), .ZN(new_n408_));
  AOI21_X1   g0023(.A1(new_n405_), .A2(\b[4] ), .B(\a[4] ), .ZN(new_n409_));
  OR2_X2     g0024(.A1(new_n409_), .A2(new_n408_), .Z(new_n410_));
  XNOR2_X1   g0025(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n411_));
  XOR2_X1    g0026(.A1(new_n410_), .A2(new_n411_), .Z(\f[5] ));
  NOR2_X1    g0027(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n413_));
  INV_X1     g0028(.I(new_n413_), .ZN(new_n414_));
  NAND2_X1   g0029(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n415_));
  OAI21_X1   g0030(.A1(new_n409_), .A2(new_n408_), .B(new_n415_), .ZN(new_n416_));
  NAND2_X1   g0031(.A1(new_n416_), .A2(new_n414_), .ZN(new_n417_));
  XNOR2_X1   g0032(.A1(\a[6] ), .A2(\b[6] ), .ZN(new_n418_));
  XOR2_X1    g0033(.A1(new_n417_), .A2(new_n418_), .Z(\f[6] ));
  INV_X1     g0034(.I(\b[7] ), .ZN(new_n420_));
  INV_X1     g0035(.I(\a[6] ), .ZN(new_n421_));
  INV_X1     g0036(.I(\b[6] ), .ZN(new_n422_));
  NOR2_X1    g0037(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1     g0038(.I(new_n423_), .ZN(new_n424_));
  NAND2_X1   g0039(.A1(new_n421_), .A2(new_n422_), .ZN(new_n425_));
  NAND3_X1   g0040(.A1(new_n416_), .A2(new_n414_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1   g0041(.A1(new_n426_), .A2(new_n424_), .B(new_n420_), .ZN(new_n427_));
  NAND3_X1   g0042(.A1(new_n426_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n428_));
  INV_X1     g0043(.I(new_n428_), .ZN(new_n429_));
  NOR2_X1    g0044(.A1(new_n429_), .A2(new_n427_), .ZN(new_n430_));
  XOR2_X1    g0045(.A1(new_n430_), .A2(\a[7] ), .Z(\f[7] ));
  OAI21_X1   g0046(.A1(\a[7] ), .A2(new_n427_), .B(new_n428_), .ZN(new_n432_));
  XNOR2_X1   g0047(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n433_));
  XOR2_X1    g0048(.A1(new_n432_), .A2(new_n433_), .Z(\f[8] ));
  NOR2_X1    g0049(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n435_));
  NAND2_X1   g0050(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n436_));
  AOI21_X1   g0051(.A1(new_n432_), .A2(new_n436_), .B(new_n435_), .ZN(new_n437_));
  XOR2_X1    g0052(.A1(\a[9] ), .A2(\b[9] ), .Z(new_n438_));
  XOR2_X1    g0053(.A1(new_n437_), .A2(new_n438_), .Z(\f[9] ));
  INV_X1     g0054(.I(\b[10] ), .ZN(new_n440_));
  INV_X1     g0055(.I(\a[9] ), .ZN(new_n441_));
  INV_X1     g0056(.I(\b[9] ), .ZN(new_n442_));
  NOR2_X1    g0057(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1   g0058(.A1(new_n441_), .A2(new_n442_), .ZN(new_n444_));
  AOI21_X1   g0059(.A1(new_n437_), .A2(new_n444_), .B(new_n443_), .ZN(new_n445_));
  XOR2_X1    g0060(.A1(new_n445_), .A2(new_n440_), .Z(new_n446_));
  XOR2_X1    g0061(.A1(new_n446_), .A2(\a[10] ), .Z(\f[10] ));
  NAND2_X1   g0062(.A1(new_n445_), .A2(new_n440_), .ZN(new_n448_));
  INV_X1     g0063(.I(\a[10] ), .ZN(new_n449_));
  OAI21_X1   g0064(.A1(new_n445_), .A2(new_n440_), .B(new_n449_), .ZN(new_n450_));
  NAND2_X1   g0065(.A1(new_n450_), .A2(new_n448_), .ZN(new_n451_));
  XNOR2_X1   g0066(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n452_));
  XOR2_X1    g0067(.A1(new_n451_), .A2(new_n452_), .Z(\f[11] ));
  NOR2_X1    g0068(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n454_));
  NAND2_X1   g0069(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n455_));
  INV_X1     g0070(.I(new_n455_), .ZN(new_n456_));
  AOI21_X1   g0071(.A1(new_n450_), .A2(new_n448_), .B(new_n456_), .ZN(new_n457_));
  NOR2_X1    g0072(.A1(new_n457_), .A2(new_n454_), .ZN(new_n458_));
  XOR2_X1    g0073(.A1(\a[12] ), .A2(\b[12] ), .Z(new_n459_));
  XOR2_X1    g0074(.A1(new_n458_), .A2(new_n459_), .Z(\f[12] ));
  INV_X1     g0075(.I(\a[13] ), .ZN(new_n461_));
  AND2_X2    g0076(.A1(\a[12] ), .A2(\b[12] ), .Z(new_n462_));
  NOR2_X1    g0077(.A1(\a[12] ), .A2(\b[12] ), .ZN(new_n463_));
  NOR3_X1    g0078(.A1(new_n457_), .A2(new_n454_), .A3(new_n463_), .ZN(new_n464_));
  OAI21_X1   g0079(.A1(new_n464_), .A2(new_n462_), .B(\b[13] ), .ZN(new_n465_));
  NOR3_X1    g0080(.A1(new_n464_), .A2(\b[13] ), .A3(new_n462_), .ZN(new_n466_));
  INV_X1     g0081(.I(new_n466_), .ZN(new_n467_));
  NAND2_X1   g0082(.A1(new_n467_), .A2(new_n465_), .ZN(new_n468_));
  XOR2_X1    g0083(.A1(new_n468_), .A2(new_n461_), .Z(\f[13] ));
  AOI21_X1   g0084(.A1(new_n461_), .A2(new_n465_), .B(new_n466_), .ZN(new_n470_));
  XOR2_X1    g0085(.A1(\a[14] ), .A2(\b[14] ), .Z(new_n471_));
  XOR2_X1    g0086(.A1(new_n470_), .A2(new_n471_), .Z(\f[14] ));
  NOR2_X1    g0087(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n473_));
  INV_X1     g0088(.I(new_n473_), .ZN(new_n474_));
  NAND2_X1   g0089(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n475_));
  INV_X1     g0090(.I(new_n475_), .ZN(new_n476_));
  OAI21_X1   g0091(.A1(new_n470_), .A2(new_n476_), .B(new_n474_), .ZN(new_n477_));
  XNOR2_X1   g0092(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n478_));
  XOR2_X1    g0093(.A1(new_n477_), .A2(new_n478_), .Z(\f[15] ));
  AND2_X2    g0094(.A1(\a[15] ), .A2(\b[15] ), .Z(new_n480_));
  INV_X1     g0095(.I(new_n480_), .ZN(new_n481_));
  NOR2_X1    g0096(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n482_));
  OAI21_X1   g0097(.A1(new_n477_), .A2(new_n482_), .B(new_n481_), .ZN(new_n483_));
  NAND2_X1   g0098(.A1(new_n483_), .A2(\b[16] ), .ZN(new_n484_));
  NOR2_X1    g0099(.A1(new_n483_), .A2(\b[16] ), .ZN(new_n485_));
  INV_X1     g0100(.I(new_n485_), .ZN(new_n486_));
  NAND2_X1   g0101(.A1(new_n486_), .A2(new_n484_), .ZN(new_n487_));
  XNOR2_X1   g0102(.A1(new_n487_), .A2(\a[16] ), .ZN(\f[16] ));
  AOI21_X1   g0103(.A1(new_n483_), .A2(\b[16] ), .B(\a[16] ), .ZN(new_n489_));
  NOR2_X1    g0104(.A1(new_n489_), .A2(new_n485_), .ZN(new_n490_));
  XOR2_X1    g0105(.A1(\a[17] ), .A2(\b[17] ), .Z(new_n491_));
  XOR2_X1    g0106(.A1(new_n490_), .A2(new_n491_), .Z(\f[17] ));
  NOR2_X1    g0107(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n493_));
  INV_X1     g0108(.I(new_n493_), .ZN(new_n494_));
  NAND2_X1   g0109(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n495_));
  OAI21_X1   g0110(.A1(new_n489_), .A2(new_n485_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1   g0111(.A1(new_n496_), .A2(new_n494_), .ZN(new_n497_));
  XNOR2_X1   g0112(.A1(\a[18] ), .A2(\b[18] ), .ZN(new_n498_));
  XOR2_X1    g0113(.A1(new_n497_), .A2(new_n498_), .Z(\f[18] ));
  INV_X1     g0114(.I(\b[19] ), .ZN(new_n500_));
  INV_X1     g0115(.I(\a[18] ), .ZN(new_n501_));
  INV_X1     g0116(.I(\b[18] ), .ZN(new_n502_));
  NOR2_X1    g0117(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1     g0118(.I(new_n503_), .ZN(new_n504_));
  NAND2_X1   g0119(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  NAND3_X1   g0120(.A1(new_n496_), .A2(new_n494_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1   g0121(.A1(new_n506_), .A2(new_n504_), .B(new_n500_), .ZN(new_n507_));
  NAND3_X1   g0122(.A1(new_n506_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n508_));
  INV_X1     g0123(.I(new_n508_), .ZN(new_n509_));
  NOR2_X1    g0124(.A1(new_n509_), .A2(new_n507_), .ZN(new_n510_));
  XOR2_X1    g0125(.A1(new_n510_), .A2(\a[19] ), .Z(\f[19] ));
  OAI21_X1   g0126(.A1(\a[19] ), .A2(new_n507_), .B(new_n508_), .ZN(new_n512_));
  XNOR2_X1   g0127(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n513_));
  XOR2_X1    g0128(.A1(new_n512_), .A2(new_n513_), .Z(\f[20] ));
  NOR2_X1    g0129(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n515_));
  NAND2_X1   g0130(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n516_));
  AOI21_X1   g0131(.A1(new_n512_), .A2(new_n516_), .B(new_n515_), .ZN(new_n517_));
  XOR2_X1    g0132(.A1(\a[21] ), .A2(\b[21] ), .Z(new_n518_));
  XOR2_X1    g0133(.A1(new_n517_), .A2(new_n518_), .Z(\f[21] ));
  INV_X1     g0134(.I(\b[22] ), .ZN(new_n520_));
  INV_X1     g0135(.I(\a[21] ), .ZN(new_n521_));
  INV_X1     g0136(.I(\b[21] ), .ZN(new_n522_));
  NOR2_X1    g0137(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1    g0138(.A1(\a[21] ), .A2(\b[21] ), .ZN(new_n524_));
  INV_X1     g0139(.I(new_n524_), .ZN(new_n525_));
  AOI21_X1   g0140(.A1(new_n517_), .A2(new_n525_), .B(new_n523_), .ZN(new_n526_));
  NOR2_X1    g0141(.A1(new_n526_), .A2(new_n520_), .ZN(new_n527_));
  NAND2_X1   g0142(.A1(new_n526_), .A2(new_n520_), .ZN(new_n528_));
  INV_X1     g0143(.I(new_n528_), .ZN(new_n529_));
  NOR2_X1    g0144(.A1(new_n529_), .A2(new_n527_), .ZN(new_n530_));
  XOR2_X1    g0145(.A1(new_n530_), .A2(\a[22] ), .Z(\f[22] ));
  INV_X1     g0146(.I(\a[22] ), .ZN(new_n532_));
  OAI21_X1   g0147(.A1(new_n526_), .A2(new_n520_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1   g0148(.A1(new_n533_), .A2(new_n528_), .ZN(new_n534_));
  XNOR2_X1   g0149(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n535_));
  XOR2_X1    g0150(.A1(new_n534_), .A2(new_n535_), .Z(\f[23] ));
  NOR2_X1    g0151(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n537_));
  NAND2_X1   g0152(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n538_));
  INV_X1     g0153(.I(new_n538_), .ZN(new_n539_));
  AOI21_X1   g0154(.A1(new_n533_), .A2(new_n528_), .B(new_n539_), .ZN(new_n540_));
  NOR2_X1    g0155(.A1(new_n540_), .A2(new_n537_), .ZN(new_n541_));
  XOR2_X1    g0156(.A1(\a[24] ), .A2(\b[24] ), .Z(new_n542_));
  XOR2_X1    g0157(.A1(new_n541_), .A2(new_n542_), .Z(\f[24] ));
  INV_X1     g0158(.I(\a[25] ), .ZN(new_n544_));
  AND2_X2    g0159(.A1(\a[24] ), .A2(\b[24] ), .Z(new_n545_));
  NOR2_X1    g0160(.A1(\a[24] ), .A2(\b[24] ), .ZN(new_n546_));
  NOR3_X1    g0161(.A1(new_n540_), .A2(new_n537_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1   g0162(.A1(new_n547_), .A2(new_n545_), .B(\b[25] ), .ZN(new_n548_));
  NOR3_X1    g0163(.A1(new_n547_), .A2(\b[25] ), .A3(new_n545_), .ZN(new_n549_));
  INV_X1     g0164(.I(new_n549_), .ZN(new_n550_));
  NAND2_X1   g0165(.A1(new_n550_), .A2(new_n548_), .ZN(new_n551_));
  XOR2_X1    g0166(.A1(new_n551_), .A2(new_n544_), .Z(\f[25] ));
  AOI21_X1   g0167(.A1(new_n544_), .A2(new_n548_), .B(new_n549_), .ZN(new_n553_));
  XOR2_X1    g0168(.A1(\a[26] ), .A2(\b[26] ), .Z(new_n554_));
  XOR2_X1    g0169(.A1(new_n553_), .A2(new_n554_), .Z(\f[26] ));
  NOR2_X1    g0170(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n556_));
  INV_X1     g0171(.I(new_n556_), .ZN(new_n557_));
  NAND2_X1   g0172(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n558_));
  INV_X1     g0173(.I(new_n558_), .ZN(new_n559_));
  OAI21_X1   g0174(.A1(new_n553_), .A2(new_n559_), .B(new_n557_), .ZN(new_n560_));
  XNOR2_X1   g0175(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n561_));
  XOR2_X1    g0176(.A1(new_n560_), .A2(new_n561_), .Z(\f[27] ));
  INV_X1     g0177(.I(\a[28] ), .ZN(new_n563_));
  INV_X1     g0178(.I(\a[27] ), .ZN(new_n564_));
  INV_X1     g0179(.I(\b[27] ), .ZN(new_n565_));
  NOR2_X1    g0180(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1     g0181(.I(new_n566_), .ZN(new_n567_));
  NOR2_X1    g0182(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n568_));
  OAI21_X1   g0183(.A1(new_n560_), .A2(new_n568_), .B(new_n567_), .ZN(new_n569_));
  NAND2_X1   g0184(.A1(new_n569_), .A2(\b[28] ), .ZN(new_n570_));
  NOR2_X1    g0185(.A1(new_n569_), .A2(\b[28] ), .ZN(new_n571_));
  INV_X1     g0186(.I(new_n571_), .ZN(new_n572_));
  NAND2_X1   g0187(.A1(new_n572_), .A2(new_n570_), .ZN(new_n573_));
  XOR2_X1    g0188(.A1(new_n573_), .A2(new_n563_), .Z(\f[28] ));
  AOI21_X1   g0189(.A1(new_n569_), .A2(\b[28] ), .B(\a[28] ), .ZN(new_n575_));
  NOR2_X1    g0190(.A1(new_n575_), .A2(new_n571_), .ZN(new_n576_));
  XOR2_X1    g0191(.A1(\a[29] ), .A2(\b[29] ), .Z(new_n577_));
  XOR2_X1    g0192(.A1(new_n576_), .A2(new_n577_), .Z(\f[29] ));
  NOR2_X1    g0193(.A1(\a[29] ), .A2(\b[29] ), .ZN(new_n579_));
  INV_X1     g0194(.I(new_n579_), .ZN(new_n580_));
  INV_X1     g0195(.I(\a[29] ), .ZN(new_n581_));
  INV_X1     g0196(.I(\b[29] ), .ZN(new_n582_));
  NOR2_X1    g0197(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1     g0198(.I(new_n583_), .ZN(new_n584_));
  OAI21_X1   g0199(.A1(new_n575_), .A2(new_n571_), .B(new_n584_), .ZN(new_n585_));
  NAND2_X1   g0200(.A1(new_n585_), .A2(new_n580_), .ZN(new_n586_));
  XNOR2_X1   g0201(.A1(\a[30] ), .A2(\b[30] ), .ZN(new_n587_));
  XOR2_X1    g0202(.A1(new_n586_), .A2(new_n587_), .Z(\f[30] ));
  INV_X1     g0203(.I(\b[31] ), .ZN(new_n589_));
  AND2_X2    g0204(.A1(\a[30] ), .A2(\b[30] ), .Z(new_n590_));
  INV_X1     g0205(.I(new_n590_), .ZN(new_n591_));
  NOR2_X1    g0206(.A1(\a[30] ), .A2(\b[30] ), .ZN(new_n592_));
  INV_X1     g0207(.I(new_n592_), .ZN(new_n593_));
  NAND3_X1   g0208(.A1(new_n585_), .A2(new_n580_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1   g0209(.A1(new_n594_), .A2(new_n591_), .B(new_n589_), .ZN(new_n595_));
  NAND3_X1   g0210(.A1(new_n594_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n596_));
  INV_X1     g0211(.I(new_n596_), .ZN(new_n597_));
  NOR2_X1    g0212(.A1(new_n597_), .A2(new_n595_), .ZN(new_n598_));
  XOR2_X1    g0213(.A1(new_n598_), .A2(\a[31] ), .Z(\f[31] ));
  OAI21_X1   g0214(.A1(\a[31] ), .A2(new_n595_), .B(new_n596_), .ZN(new_n600_));
  XNOR2_X1   g0215(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n601_));
  XOR2_X1    g0216(.A1(new_n600_), .A2(new_n601_), .Z(\f[32] ));
  NOR2_X1    g0217(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n603_));
  NAND2_X1   g0218(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n604_));
  AOI21_X1   g0219(.A1(new_n600_), .A2(new_n604_), .B(new_n603_), .ZN(new_n605_));
  XOR2_X1    g0220(.A1(\a[33] ), .A2(\b[33] ), .Z(new_n606_));
  XOR2_X1    g0221(.A1(new_n605_), .A2(new_n606_), .Z(\f[33] ));
  INV_X1     g0222(.I(\b[34] ), .ZN(new_n608_));
  INV_X1     g0223(.I(\a[33] ), .ZN(new_n609_));
  INV_X1     g0224(.I(\b[33] ), .ZN(new_n610_));
  NOR2_X1    g0225(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1   g0226(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  AOI21_X1   g0227(.A1(new_n605_), .A2(new_n612_), .B(new_n611_), .ZN(new_n613_));
  NOR2_X1    g0228(.A1(new_n613_), .A2(new_n608_), .ZN(new_n614_));
  NAND2_X1   g0229(.A1(new_n613_), .A2(new_n608_), .ZN(new_n615_));
  INV_X1     g0230(.I(new_n615_), .ZN(new_n616_));
  NOR2_X1    g0231(.A1(new_n616_), .A2(new_n614_), .ZN(new_n617_));
  XOR2_X1    g0232(.A1(new_n617_), .A2(\a[34] ), .Z(\f[34] ));
  INV_X1     g0233(.I(\a[34] ), .ZN(new_n619_));
  OAI21_X1   g0234(.A1(new_n613_), .A2(new_n608_), .B(new_n619_), .ZN(new_n620_));
  NAND2_X1   g0235(.A1(new_n620_), .A2(new_n615_), .ZN(new_n621_));
  XNOR2_X1   g0236(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n622_));
  XOR2_X1    g0237(.A1(new_n621_), .A2(new_n622_), .Z(\f[35] ));
  NOR2_X1    g0238(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n624_));
  NAND2_X1   g0239(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n625_));
  INV_X1     g0240(.I(new_n625_), .ZN(new_n626_));
  AOI21_X1   g0241(.A1(new_n620_), .A2(new_n615_), .B(new_n626_), .ZN(new_n627_));
  NOR2_X1    g0242(.A1(new_n627_), .A2(new_n624_), .ZN(new_n628_));
  XOR2_X1    g0243(.A1(\a[36] ), .A2(\b[36] ), .Z(new_n629_));
  XOR2_X1    g0244(.A1(new_n628_), .A2(new_n629_), .Z(\f[36] ));
  INV_X1     g0245(.I(\a[37] ), .ZN(new_n631_));
  AND2_X2    g0246(.A1(\a[36] ), .A2(\b[36] ), .Z(new_n632_));
  NOR2_X1    g0247(.A1(\a[36] ), .A2(\b[36] ), .ZN(new_n633_));
  NOR3_X1    g0248(.A1(new_n627_), .A2(new_n624_), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1   g0249(.A1(new_n634_), .A2(new_n632_), .B(\b[37] ), .ZN(new_n635_));
  NOR3_X1    g0250(.A1(new_n634_), .A2(\b[37] ), .A3(new_n632_), .ZN(new_n636_));
  INV_X1     g0251(.I(new_n636_), .ZN(new_n637_));
  NAND2_X1   g0252(.A1(new_n637_), .A2(new_n635_), .ZN(new_n638_));
  XOR2_X1    g0253(.A1(new_n638_), .A2(new_n631_), .Z(\f[37] ));
  AOI21_X1   g0254(.A1(new_n631_), .A2(new_n635_), .B(new_n636_), .ZN(new_n640_));
  XOR2_X1    g0255(.A1(\a[38] ), .A2(\b[38] ), .Z(new_n641_));
  XOR2_X1    g0256(.A1(new_n640_), .A2(new_n641_), .Z(\f[38] ));
  NOR2_X1    g0257(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n643_));
  INV_X1     g0258(.I(new_n643_), .ZN(new_n644_));
  NAND2_X1   g0259(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n645_));
  INV_X1     g0260(.I(new_n645_), .ZN(new_n646_));
  OAI21_X1   g0261(.A1(new_n640_), .A2(new_n646_), .B(new_n644_), .ZN(new_n647_));
  XNOR2_X1   g0262(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n648_));
  XOR2_X1    g0263(.A1(new_n647_), .A2(new_n648_), .Z(\f[39] ));
  INV_X1     g0264(.I(\a[40] ), .ZN(new_n650_));
  INV_X1     g0265(.I(\a[39] ), .ZN(new_n651_));
  INV_X1     g0266(.I(\b[39] ), .ZN(new_n652_));
  NOR2_X1    g0267(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1     g0268(.I(new_n653_), .ZN(new_n654_));
  NOR2_X1    g0269(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n655_));
  OAI21_X1   g0270(.A1(new_n647_), .A2(new_n655_), .B(new_n654_), .ZN(new_n656_));
  NAND2_X1   g0271(.A1(new_n656_), .A2(\b[40] ), .ZN(new_n657_));
  NOR2_X1    g0272(.A1(new_n656_), .A2(\b[40] ), .ZN(new_n658_));
  INV_X1     g0273(.I(new_n658_), .ZN(new_n659_));
  NAND2_X1   g0274(.A1(new_n659_), .A2(new_n657_), .ZN(new_n660_));
  XOR2_X1    g0275(.A1(new_n660_), .A2(new_n650_), .Z(\f[40] ));
  AOI21_X1   g0276(.A1(new_n656_), .A2(\b[40] ), .B(\a[40] ), .ZN(new_n662_));
  NOR2_X1    g0277(.A1(new_n662_), .A2(new_n658_), .ZN(new_n663_));
  XOR2_X1    g0278(.A1(\a[41] ), .A2(\b[41] ), .Z(new_n664_));
  XOR2_X1    g0279(.A1(new_n663_), .A2(new_n664_), .Z(\f[41] ));
  NOR2_X1    g0280(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n666_));
  INV_X1     g0281(.I(new_n666_), .ZN(new_n667_));
  NAND2_X1   g0282(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n668_));
  OAI21_X1   g0283(.A1(new_n662_), .A2(new_n658_), .B(new_n668_), .ZN(new_n669_));
  NAND2_X1   g0284(.A1(new_n669_), .A2(new_n667_), .ZN(new_n670_));
  XNOR2_X1   g0285(.A1(\a[42] ), .A2(\b[42] ), .ZN(new_n671_));
  XOR2_X1    g0286(.A1(new_n670_), .A2(new_n671_), .Z(\f[42] ));
  INV_X1     g0287(.I(\b[43] ), .ZN(new_n673_));
  AND2_X2    g0288(.A1(\a[42] ), .A2(\b[42] ), .Z(new_n674_));
  INV_X1     g0289(.I(new_n674_), .ZN(new_n675_));
  NOR2_X1    g0290(.A1(\a[42] ), .A2(\b[42] ), .ZN(new_n676_));
  INV_X1     g0291(.I(new_n676_), .ZN(new_n677_));
  NAND3_X1   g0292(.A1(new_n669_), .A2(new_n667_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1   g0293(.A1(new_n678_), .A2(new_n675_), .B(new_n673_), .ZN(new_n679_));
  NAND3_X1   g0294(.A1(new_n678_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n680_));
  INV_X1     g0295(.I(new_n680_), .ZN(new_n681_));
  NOR2_X1    g0296(.A1(new_n681_), .A2(new_n679_), .ZN(new_n682_));
  XOR2_X1    g0297(.A1(new_n682_), .A2(\a[43] ), .Z(\f[43] ));
  OAI21_X1   g0298(.A1(\a[43] ), .A2(new_n679_), .B(new_n680_), .ZN(new_n684_));
  XNOR2_X1   g0299(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n685_));
  XOR2_X1    g0300(.A1(new_n684_), .A2(new_n685_), .Z(\f[44] ));
  NOR2_X1    g0301(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n687_));
  NAND2_X1   g0302(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n688_));
  AOI21_X1   g0303(.A1(new_n684_), .A2(new_n688_), .B(new_n687_), .ZN(new_n689_));
  XOR2_X1    g0304(.A1(\a[45] ), .A2(\b[45] ), .Z(new_n690_));
  XOR2_X1    g0305(.A1(new_n689_), .A2(new_n690_), .Z(\f[45] ));
  INV_X1     g0306(.I(\b[46] ), .ZN(new_n692_));
  INV_X1     g0307(.I(\a[45] ), .ZN(new_n693_));
  INV_X1     g0308(.I(\b[45] ), .ZN(new_n694_));
  NOR2_X1    g0309(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1     g0310(.I(new_n695_), .ZN(new_n696_));
  INV_X1     g0311(.I(new_n687_), .ZN(new_n697_));
  NAND2_X1   g0312(.A1(new_n678_), .A2(new_n675_), .ZN(new_n698_));
  AOI21_X1   g0313(.A1(new_n698_), .A2(\b[43] ), .B(\a[43] ), .ZN(new_n699_));
  OAI21_X1   g0314(.A1(new_n699_), .A2(new_n681_), .B(new_n688_), .ZN(new_n700_));
  NOR2_X1    g0315(.A1(\a[45] ), .A2(\b[45] ), .ZN(new_n701_));
  INV_X1     g0316(.I(new_n701_), .ZN(new_n702_));
  NAND3_X1   g0317(.A1(new_n700_), .A2(new_n697_), .A3(new_n702_), .ZN(new_n703_));
  AOI21_X1   g0318(.A1(new_n703_), .A2(new_n696_), .B(new_n692_), .ZN(new_n704_));
  NAND3_X1   g0319(.A1(new_n703_), .A2(new_n692_), .A3(new_n696_), .ZN(new_n705_));
  INV_X1     g0320(.I(new_n705_), .ZN(new_n706_));
  NOR2_X1    g0321(.A1(new_n706_), .A2(new_n704_), .ZN(new_n707_));
  XOR2_X1    g0322(.A1(new_n707_), .A2(\a[46] ), .Z(\f[46] ));
  OAI21_X1   g0323(.A1(\a[46] ), .A2(new_n704_), .B(new_n705_), .ZN(new_n709_));
  XNOR2_X1   g0324(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n710_));
  XOR2_X1    g0325(.A1(new_n709_), .A2(new_n710_), .Z(\f[47] ));
  NOR2_X1    g0326(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n712_));
  NAND2_X1   g0327(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n713_));
  AOI21_X1   g0328(.A1(new_n709_), .A2(new_n713_), .B(new_n712_), .ZN(new_n714_));
  XOR2_X1    g0329(.A1(\a[48] ), .A2(\b[48] ), .Z(new_n715_));
  XOR2_X1    g0330(.A1(new_n714_), .A2(new_n715_), .Z(\f[48] ));
  INV_X1     g0331(.I(\a[49] ), .ZN(new_n717_));
  AND2_X2    g0332(.A1(\a[48] ), .A2(\b[48] ), .Z(new_n718_));
  INV_X1     g0333(.I(\a[46] ), .ZN(new_n719_));
  AOI21_X1   g0334(.A1(new_n689_), .A2(new_n702_), .B(new_n695_), .ZN(new_n720_));
  OAI21_X1   g0335(.A1(new_n720_), .A2(new_n692_), .B(new_n719_), .ZN(new_n721_));
  AOI22_X1   g0336(.A1(new_n721_), .A2(new_n705_), .B1(\a[47] ), .B2(\b[47] ), .ZN(new_n722_));
  NOR2_X1    g0337(.A1(\a[48] ), .A2(\b[48] ), .ZN(new_n723_));
  NOR3_X1    g0338(.A1(new_n722_), .A2(new_n712_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1   g0339(.A1(new_n724_), .A2(new_n718_), .B(\b[49] ), .ZN(new_n725_));
  INV_X1     g0340(.I(\b[49] ), .ZN(new_n726_));
  INV_X1     g0341(.I(new_n723_), .ZN(new_n727_));
  AOI21_X1   g0342(.A1(new_n714_), .A2(new_n727_), .B(new_n718_), .ZN(new_n728_));
  NAND2_X1   g0343(.A1(new_n728_), .A2(new_n726_), .ZN(new_n729_));
  NAND2_X1   g0344(.A1(new_n729_), .A2(new_n725_), .ZN(new_n730_));
  XOR2_X1    g0345(.A1(new_n730_), .A2(new_n717_), .Z(\f[49] ));
  NOR3_X1    g0346(.A1(new_n724_), .A2(\b[49] ), .A3(new_n718_), .ZN(new_n732_));
  AOI21_X1   g0347(.A1(new_n717_), .A2(new_n725_), .B(new_n732_), .ZN(new_n733_));
  XOR2_X1    g0348(.A1(\a[50] ), .A2(\b[50] ), .Z(new_n734_));
  XOR2_X1    g0349(.A1(new_n733_), .A2(new_n734_), .Z(\f[50] ));
  NOR2_X1    g0350(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n736_));
  INV_X1     g0351(.I(new_n736_), .ZN(new_n737_));
  NAND2_X1   g0352(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n738_));
  INV_X1     g0353(.I(new_n738_), .ZN(new_n739_));
  OAI21_X1   g0354(.A1(new_n733_), .A2(new_n739_), .B(new_n737_), .ZN(new_n740_));
  XNOR2_X1   g0355(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n741_));
  XOR2_X1    g0356(.A1(new_n740_), .A2(new_n741_), .Z(\f[51] ));
  INV_X1     g0357(.I(\a[52] ), .ZN(new_n743_));
  INV_X1     g0358(.I(\a[51] ), .ZN(new_n744_));
  INV_X1     g0359(.I(\b[51] ), .ZN(new_n745_));
  NOR2_X1    g0360(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1   g0361(.A1(new_n728_), .A2(new_n726_), .B(new_n717_), .ZN(new_n747_));
  AOI21_X1   g0362(.A1(new_n747_), .A2(new_n729_), .B(new_n739_), .ZN(new_n748_));
  NOR2_X1    g0363(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n749_));
  NOR3_X1    g0364(.A1(new_n748_), .A2(new_n736_), .A3(new_n749_), .ZN(new_n750_));
  OAI21_X1   g0365(.A1(new_n750_), .A2(new_n746_), .B(\b[52] ), .ZN(new_n751_));
  NOR3_X1    g0366(.A1(new_n750_), .A2(\b[52] ), .A3(new_n746_), .ZN(new_n752_));
  INV_X1     g0367(.I(new_n752_), .ZN(new_n753_));
  NAND2_X1   g0368(.A1(new_n753_), .A2(new_n751_), .ZN(new_n754_));
  XOR2_X1    g0369(.A1(new_n754_), .A2(new_n743_), .Z(\f[52] ));
  AOI21_X1   g0370(.A1(new_n743_), .A2(new_n751_), .B(new_n752_), .ZN(new_n756_));
  XOR2_X1    g0371(.A1(\a[53] ), .A2(\b[53] ), .Z(new_n757_));
  XOR2_X1    g0372(.A1(new_n756_), .A2(new_n757_), .Z(\f[53] ));
  NOR2_X1    g0373(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n759_));
  INV_X1     g0374(.I(new_n759_), .ZN(new_n760_));
  NAND2_X1   g0375(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n761_));
  INV_X1     g0376(.I(new_n761_), .ZN(new_n762_));
  OAI21_X1   g0377(.A1(new_n756_), .A2(new_n762_), .B(new_n760_), .ZN(new_n763_));
  XNOR2_X1   g0378(.A1(\a[54] ), .A2(\b[54] ), .ZN(new_n764_));
  XOR2_X1    g0379(.A1(new_n763_), .A2(new_n764_), .Z(\f[54] ));
  INV_X1     g0380(.I(\b[55] ), .ZN(new_n766_));
  AND2_X2    g0381(.A1(\a[54] ), .A2(\b[54] ), .Z(new_n767_));
  INV_X1     g0382(.I(new_n767_), .ZN(new_n768_));
  INV_X1     g0383(.I(new_n746_), .ZN(new_n769_));
  OAI21_X1   g0384(.A1(new_n740_), .A2(new_n749_), .B(new_n769_), .ZN(new_n770_));
  AOI21_X1   g0385(.A1(new_n770_), .A2(\b[52] ), .B(\a[52] ), .ZN(new_n771_));
  OAI21_X1   g0386(.A1(new_n771_), .A2(new_n752_), .B(new_n761_), .ZN(new_n772_));
  NOR2_X1    g0387(.A1(\a[54] ), .A2(\b[54] ), .ZN(new_n773_));
  INV_X1     g0388(.I(new_n773_), .ZN(new_n774_));
  NAND3_X1   g0389(.A1(new_n772_), .A2(new_n760_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1   g0390(.A1(new_n775_), .A2(new_n768_), .B(new_n766_), .ZN(new_n776_));
  OAI21_X1   g0391(.A1(new_n763_), .A2(new_n773_), .B(new_n768_), .ZN(new_n777_));
  NOR2_X1    g0392(.A1(new_n777_), .A2(\b[55] ), .ZN(new_n778_));
  NOR2_X1    g0393(.A1(new_n778_), .A2(new_n776_), .ZN(new_n779_));
  XOR2_X1    g0394(.A1(new_n779_), .A2(\a[55] ), .Z(\f[55] ));
  NAND3_X1   g0395(.A1(new_n775_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n781_));
  OAI21_X1   g0396(.A1(\a[55] ), .A2(new_n776_), .B(new_n781_), .ZN(new_n782_));
  XNOR2_X1   g0397(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n783_));
  XOR2_X1    g0398(.A1(new_n782_), .A2(new_n783_), .Z(\f[56] ));
  NOR2_X1    g0399(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n785_));
  NAND2_X1   g0400(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n786_));
  AOI21_X1   g0401(.A1(new_n782_), .A2(new_n786_), .B(new_n785_), .ZN(new_n787_));
  XOR2_X1    g0402(.A1(\a[57] ), .A2(\b[57] ), .Z(new_n788_));
  XOR2_X1    g0403(.A1(new_n787_), .A2(new_n788_), .Z(\f[57] ));
  INV_X1     g0404(.I(\b[58] ), .ZN(new_n790_));
  INV_X1     g0405(.I(\a[57] ), .ZN(new_n791_));
  INV_X1     g0406(.I(\b[57] ), .ZN(new_n792_));
  NOR2_X1    g0407(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1     g0408(.I(new_n793_), .ZN(new_n794_));
  INV_X1     g0409(.I(new_n785_), .ZN(new_n795_));
  AOI21_X1   g0410(.A1(new_n777_), .A2(\b[55] ), .B(\a[55] ), .ZN(new_n796_));
  OAI21_X1   g0411(.A1(new_n796_), .A2(new_n778_), .B(new_n786_), .ZN(new_n797_));
  NOR2_X1    g0412(.A1(\a[57] ), .A2(\b[57] ), .ZN(new_n798_));
  INV_X1     g0413(.I(new_n798_), .ZN(new_n799_));
  NAND3_X1   g0414(.A1(new_n797_), .A2(new_n795_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1   g0415(.A1(new_n800_), .A2(new_n794_), .B(new_n790_), .ZN(new_n801_));
  NAND3_X1   g0416(.A1(new_n800_), .A2(new_n790_), .A3(new_n794_), .ZN(new_n802_));
  INV_X1     g0417(.I(new_n802_), .ZN(new_n803_));
  NOR2_X1    g0418(.A1(new_n803_), .A2(new_n801_), .ZN(new_n804_));
  XOR2_X1    g0419(.A1(new_n804_), .A2(\a[58] ), .Z(\f[58] ));
  OAI21_X1   g0420(.A1(\a[58] ), .A2(new_n801_), .B(new_n802_), .ZN(new_n806_));
  XNOR2_X1   g0421(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n807_));
  XOR2_X1    g0422(.A1(new_n806_), .A2(new_n807_), .Z(\f[59] ));
  NOR2_X1    g0423(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n809_));
  NAND2_X1   g0424(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n810_));
  AOI21_X1   g0425(.A1(new_n806_), .A2(new_n810_), .B(new_n809_), .ZN(new_n811_));
  XOR2_X1    g0426(.A1(\a[60] ), .A2(\b[60] ), .Z(new_n812_));
  XOR2_X1    g0427(.A1(new_n811_), .A2(new_n812_), .Z(\f[60] ));
  INV_X1     g0428(.I(\a[61] ), .ZN(new_n814_));
  AND2_X2    g0429(.A1(\a[60] ), .A2(\b[60] ), .Z(new_n815_));
  INV_X1     g0430(.I(\a[58] ), .ZN(new_n816_));
  AOI21_X1   g0431(.A1(new_n787_), .A2(new_n799_), .B(new_n793_), .ZN(new_n817_));
  OAI21_X1   g0432(.A1(new_n817_), .A2(new_n790_), .B(new_n816_), .ZN(new_n818_));
  AOI22_X1   g0433(.A1(new_n818_), .A2(new_n802_), .B1(\a[59] ), .B2(\b[59] ), .ZN(new_n819_));
  NOR2_X1    g0434(.A1(\a[60] ), .A2(\b[60] ), .ZN(new_n820_));
  NOR3_X1    g0435(.A1(new_n819_), .A2(new_n809_), .A3(new_n820_), .ZN(new_n821_));
  OAI21_X1   g0436(.A1(new_n821_), .A2(new_n815_), .B(\b[61] ), .ZN(new_n822_));
  INV_X1     g0437(.I(\b[61] ), .ZN(new_n823_));
  INV_X1     g0438(.I(new_n820_), .ZN(new_n824_));
  AOI21_X1   g0439(.A1(new_n811_), .A2(new_n824_), .B(new_n815_), .ZN(new_n825_));
  NAND2_X1   g0440(.A1(new_n825_), .A2(new_n823_), .ZN(new_n826_));
  NAND2_X1   g0441(.A1(new_n826_), .A2(new_n822_), .ZN(new_n827_));
  XOR2_X1    g0442(.A1(new_n827_), .A2(new_n814_), .Z(\f[61] ));
  NOR3_X1    g0443(.A1(new_n821_), .A2(\b[61] ), .A3(new_n815_), .ZN(new_n829_));
  AOI21_X1   g0444(.A1(new_n814_), .A2(new_n822_), .B(new_n829_), .ZN(new_n830_));
  XOR2_X1    g0445(.A1(\a[62] ), .A2(\b[62] ), .Z(new_n831_));
  XOR2_X1    g0446(.A1(new_n830_), .A2(new_n831_), .Z(\f[62] ));
  NOR2_X1    g0447(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n833_));
  INV_X1     g0448(.I(new_n833_), .ZN(new_n834_));
  NAND2_X1   g0449(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n835_));
  INV_X1     g0450(.I(new_n835_), .ZN(new_n836_));
  OAI21_X1   g0451(.A1(new_n830_), .A2(new_n836_), .B(new_n834_), .ZN(new_n837_));
  XNOR2_X1   g0452(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n838_));
  XOR2_X1    g0453(.A1(new_n837_), .A2(new_n838_), .Z(\f[63] ));
  INV_X1     g0454(.I(\a[64] ), .ZN(new_n840_));
  INV_X1     g0455(.I(\a[63] ), .ZN(new_n841_));
  INV_X1     g0456(.I(\b[63] ), .ZN(new_n842_));
  NOR2_X1    g0457(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1   g0458(.A1(new_n825_), .A2(new_n823_), .B(new_n814_), .ZN(new_n844_));
  AOI21_X1   g0459(.A1(new_n844_), .A2(new_n826_), .B(new_n836_), .ZN(new_n845_));
  NOR2_X1    g0460(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n846_));
  NOR3_X1    g0461(.A1(new_n845_), .A2(new_n833_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1   g0462(.A1(new_n847_), .A2(new_n843_), .B(\b[64] ), .ZN(new_n848_));
  NOR3_X1    g0463(.A1(new_n847_), .A2(\b[64] ), .A3(new_n843_), .ZN(new_n849_));
  INV_X1     g0464(.I(new_n849_), .ZN(new_n850_));
  NAND2_X1   g0465(.A1(new_n850_), .A2(new_n848_), .ZN(new_n851_));
  XOR2_X1    g0466(.A1(new_n851_), .A2(new_n840_), .Z(\f[64] ));
  AOI21_X1   g0467(.A1(new_n840_), .A2(new_n848_), .B(new_n849_), .ZN(new_n853_));
  XOR2_X1    g0468(.A1(\a[65] ), .A2(\b[65] ), .Z(new_n854_));
  XOR2_X1    g0469(.A1(new_n853_), .A2(new_n854_), .Z(\f[65] ));
  NOR2_X1    g0470(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n856_));
  INV_X1     g0471(.I(new_n856_), .ZN(new_n857_));
  NAND2_X1   g0472(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n858_));
  INV_X1     g0473(.I(new_n858_), .ZN(new_n859_));
  OAI21_X1   g0474(.A1(new_n853_), .A2(new_n859_), .B(new_n857_), .ZN(new_n860_));
  XNOR2_X1   g0475(.A1(\a[66] ), .A2(\b[66] ), .ZN(new_n861_));
  XOR2_X1    g0476(.A1(new_n860_), .A2(new_n861_), .Z(\f[66] ));
  INV_X1     g0477(.I(\b[67] ), .ZN(new_n863_));
  AND2_X2    g0478(.A1(\a[66] ), .A2(\b[66] ), .Z(new_n864_));
  INV_X1     g0479(.I(new_n864_), .ZN(new_n865_));
  INV_X1     g0480(.I(new_n843_), .ZN(new_n866_));
  OAI21_X1   g0481(.A1(new_n837_), .A2(new_n846_), .B(new_n866_), .ZN(new_n867_));
  AOI21_X1   g0482(.A1(new_n867_), .A2(\b[64] ), .B(\a[64] ), .ZN(new_n868_));
  OAI21_X1   g0483(.A1(new_n868_), .A2(new_n849_), .B(new_n858_), .ZN(new_n869_));
  NOR2_X1    g0484(.A1(\a[66] ), .A2(\b[66] ), .ZN(new_n870_));
  INV_X1     g0485(.I(new_n870_), .ZN(new_n871_));
  NAND3_X1   g0486(.A1(new_n869_), .A2(new_n857_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1   g0487(.A1(new_n872_), .A2(new_n865_), .B(new_n863_), .ZN(new_n873_));
  OAI21_X1   g0488(.A1(new_n860_), .A2(new_n870_), .B(new_n865_), .ZN(new_n874_));
  NOR2_X1    g0489(.A1(new_n874_), .A2(\b[67] ), .ZN(new_n875_));
  NOR2_X1    g0490(.A1(new_n875_), .A2(new_n873_), .ZN(new_n876_));
  XOR2_X1    g0491(.A1(new_n876_), .A2(\a[67] ), .Z(\f[67] ));
  NAND3_X1   g0492(.A1(new_n872_), .A2(new_n863_), .A3(new_n865_), .ZN(new_n878_));
  OAI21_X1   g0493(.A1(\a[67] ), .A2(new_n873_), .B(new_n878_), .ZN(new_n879_));
  XNOR2_X1   g0494(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n880_));
  XOR2_X1    g0495(.A1(new_n879_), .A2(new_n880_), .Z(\f[68] ));
  NOR2_X1    g0496(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n882_));
  NAND2_X1   g0497(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n883_));
  AOI21_X1   g0498(.A1(new_n879_), .A2(new_n883_), .B(new_n882_), .ZN(new_n884_));
  XOR2_X1    g0499(.A1(\a[69] ), .A2(\b[69] ), .Z(new_n885_));
  XOR2_X1    g0500(.A1(new_n884_), .A2(new_n885_), .Z(\f[69] ));
  INV_X1     g0501(.I(\b[70] ), .ZN(new_n887_));
  INV_X1     g0502(.I(\a[69] ), .ZN(new_n888_));
  INV_X1     g0503(.I(\b[69] ), .ZN(new_n889_));
  NOR2_X1    g0504(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1     g0505(.I(new_n890_), .ZN(new_n891_));
  INV_X1     g0506(.I(new_n882_), .ZN(new_n892_));
  AOI21_X1   g0507(.A1(new_n874_), .A2(\b[67] ), .B(\a[67] ), .ZN(new_n893_));
  OAI21_X1   g0508(.A1(new_n893_), .A2(new_n875_), .B(new_n883_), .ZN(new_n894_));
  NOR2_X1    g0509(.A1(\a[69] ), .A2(\b[69] ), .ZN(new_n895_));
  INV_X1     g0510(.I(new_n895_), .ZN(new_n896_));
  NAND3_X1   g0511(.A1(new_n894_), .A2(new_n892_), .A3(new_n896_), .ZN(new_n897_));
  AOI21_X1   g0512(.A1(new_n897_), .A2(new_n891_), .B(new_n887_), .ZN(new_n898_));
  NAND3_X1   g0513(.A1(new_n897_), .A2(new_n887_), .A3(new_n891_), .ZN(new_n899_));
  INV_X1     g0514(.I(new_n899_), .ZN(new_n900_));
  NOR2_X1    g0515(.A1(new_n900_), .A2(new_n898_), .ZN(new_n901_));
  XOR2_X1    g0516(.A1(new_n901_), .A2(\a[70] ), .Z(\f[70] ));
  OAI21_X1   g0517(.A1(\a[70] ), .A2(new_n898_), .B(new_n899_), .ZN(new_n903_));
  XNOR2_X1   g0518(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n904_));
  XOR2_X1    g0519(.A1(new_n903_), .A2(new_n904_), .Z(\f[71] ));
  NOR2_X1    g0520(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n906_));
  NAND2_X1   g0521(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n907_));
  AOI21_X1   g0522(.A1(new_n903_), .A2(new_n907_), .B(new_n906_), .ZN(new_n908_));
  XOR2_X1    g0523(.A1(\a[72] ), .A2(\b[72] ), .Z(new_n909_));
  XOR2_X1    g0524(.A1(new_n908_), .A2(new_n909_), .Z(\f[72] ));
  INV_X1     g0525(.I(\a[73] ), .ZN(new_n911_));
  AND2_X2    g0526(.A1(\a[72] ), .A2(\b[72] ), .Z(new_n912_));
  INV_X1     g0527(.I(\a[70] ), .ZN(new_n913_));
  AOI21_X1   g0528(.A1(new_n884_), .A2(new_n896_), .B(new_n890_), .ZN(new_n914_));
  OAI21_X1   g0529(.A1(new_n914_), .A2(new_n887_), .B(new_n913_), .ZN(new_n915_));
  AOI22_X1   g0530(.A1(new_n915_), .A2(new_n899_), .B1(\a[71] ), .B2(\b[71] ), .ZN(new_n916_));
  NOR2_X1    g0531(.A1(\a[72] ), .A2(\b[72] ), .ZN(new_n917_));
  NOR3_X1    g0532(.A1(new_n916_), .A2(new_n906_), .A3(new_n917_), .ZN(new_n918_));
  OAI21_X1   g0533(.A1(new_n918_), .A2(new_n912_), .B(\b[73] ), .ZN(new_n919_));
  INV_X1     g0534(.I(\b[73] ), .ZN(new_n920_));
  INV_X1     g0535(.I(new_n917_), .ZN(new_n921_));
  AOI21_X1   g0536(.A1(new_n908_), .A2(new_n921_), .B(new_n912_), .ZN(new_n922_));
  NAND2_X1   g0537(.A1(new_n922_), .A2(new_n920_), .ZN(new_n923_));
  NAND2_X1   g0538(.A1(new_n923_), .A2(new_n919_), .ZN(new_n924_));
  XOR2_X1    g0539(.A1(new_n924_), .A2(new_n911_), .Z(\f[73] ));
  NOR3_X1    g0540(.A1(new_n918_), .A2(\b[73] ), .A3(new_n912_), .ZN(new_n926_));
  AOI21_X1   g0541(.A1(new_n911_), .A2(new_n919_), .B(new_n926_), .ZN(new_n927_));
  XOR2_X1    g0542(.A1(\a[74] ), .A2(\b[74] ), .Z(new_n928_));
  XOR2_X1    g0543(.A1(new_n927_), .A2(new_n928_), .Z(\f[74] ));
  NOR2_X1    g0544(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n930_));
  INV_X1     g0545(.I(new_n930_), .ZN(new_n931_));
  NAND2_X1   g0546(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n932_));
  INV_X1     g0547(.I(new_n932_), .ZN(new_n933_));
  OAI21_X1   g0548(.A1(new_n927_), .A2(new_n933_), .B(new_n931_), .ZN(new_n934_));
  XNOR2_X1   g0549(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n935_));
  XOR2_X1    g0550(.A1(new_n934_), .A2(new_n935_), .Z(\f[75] ));
  INV_X1     g0551(.I(\a[76] ), .ZN(new_n937_));
  INV_X1     g0552(.I(\a[75] ), .ZN(new_n938_));
  INV_X1     g0553(.I(\b[75] ), .ZN(new_n939_));
  NOR2_X1    g0554(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  OAI21_X1   g0555(.A1(new_n922_), .A2(new_n920_), .B(new_n911_), .ZN(new_n941_));
  AOI21_X1   g0556(.A1(new_n941_), .A2(new_n923_), .B(new_n933_), .ZN(new_n942_));
  NOR2_X1    g0557(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n943_));
  NOR3_X1    g0558(.A1(new_n942_), .A2(new_n930_), .A3(new_n943_), .ZN(new_n944_));
  OAI21_X1   g0559(.A1(new_n944_), .A2(new_n940_), .B(\b[76] ), .ZN(new_n945_));
  NOR3_X1    g0560(.A1(new_n944_), .A2(\b[76] ), .A3(new_n940_), .ZN(new_n946_));
  INV_X1     g0561(.I(new_n946_), .ZN(new_n947_));
  NAND2_X1   g0562(.A1(new_n947_), .A2(new_n945_), .ZN(new_n948_));
  XOR2_X1    g0563(.A1(new_n948_), .A2(new_n937_), .Z(\f[76] ));
  AOI21_X1   g0564(.A1(new_n937_), .A2(new_n945_), .B(new_n946_), .ZN(new_n950_));
  XOR2_X1    g0565(.A1(\a[77] ), .A2(\b[77] ), .Z(new_n951_));
  XOR2_X1    g0566(.A1(new_n950_), .A2(new_n951_), .Z(\f[77] ));
  NOR2_X1    g0567(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n953_));
  INV_X1     g0568(.I(new_n953_), .ZN(new_n954_));
  NAND2_X1   g0569(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n955_));
  INV_X1     g0570(.I(new_n955_), .ZN(new_n956_));
  OAI21_X1   g0571(.A1(new_n950_), .A2(new_n956_), .B(new_n954_), .ZN(new_n957_));
  XNOR2_X1   g0572(.A1(\a[78] ), .A2(\b[78] ), .ZN(new_n958_));
  XOR2_X1    g0573(.A1(new_n957_), .A2(new_n958_), .Z(\f[78] ));
  INV_X1     g0574(.I(\b[79] ), .ZN(new_n960_));
  AND2_X2    g0575(.A1(\a[78] ), .A2(\b[78] ), .Z(new_n961_));
  INV_X1     g0576(.I(new_n961_), .ZN(new_n962_));
  INV_X1     g0577(.I(new_n940_), .ZN(new_n963_));
  OAI21_X1   g0578(.A1(new_n934_), .A2(new_n943_), .B(new_n963_), .ZN(new_n964_));
  AOI21_X1   g0579(.A1(new_n964_), .A2(\b[76] ), .B(\a[76] ), .ZN(new_n965_));
  OAI21_X1   g0580(.A1(new_n965_), .A2(new_n946_), .B(new_n955_), .ZN(new_n966_));
  NOR2_X1    g0581(.A1(\a[78] ), .A2(\b[78] ), .ZN(new_n967_));
  INV_X1     g0582(.I(new_n967_), .ZN(new_n968_));
  NAND3_X1   g0583(.A1(new_n966_), .A2(new_n954_), .A3(new_n968_), .ZN(new_n969_));
  AOI21_X1   g0584(.A1(new_n969_), .A2(new_n962_), .B(new_n960_), .ZN(new_n970_));
  OAI21_X1   g0585(.A1(new_n957_), .A2(new_n967_), .B(new_n962_), .ZN(new_n971_));
  NOR2_X1    g0586(.A1(new_n971_), .A2(\b[79] ), .ZN(new_n972_));
  NOR2_X1    g0587(.A1(new_n972_), .A2(new_n970_), .ZN(new_n973_));
  XOR2_X1    g0588(.A1(new_n973_), .A2(\a[79] ), .Z(\f[79] ));
  NAND3_X1   g0589(.A1(new_n969_), .A2(new_n960_), .A3(new_n962_), .ZN(new_n975_));
  OAI21_X1   g0590(.A1(\a[79] ), .A2(new_n970_), .B(new_n975_), .ZN(new_n976_));
  XNOR2_X1   g0591(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n977_));
  XOR2_X1    g0592(.A1(new_n976_), .A2(new_n977_), .Z(\f[80] ));
  NOR2_X1    g0593(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n979_));
  NAND2_X1   g0594(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n980_));
  AOI21_X1   g0595(.A1(new_n976_), .A2(new_n980_), .B(new_n979_), .ZN(new_n981_));
  XOR2_X1    g0596(.A1(\a[81] ), .A2(\b[81] ), .Z(new_n982_));
  XOR2_X1    g0597(.A1(new_n981_), .A2(new_n982_), .Z(\f[81] ));
  INV_X1     g0598(.I(\b[82] ), .ZN(new_n984_));
  INV_X1     g0599(.I(\a[81] ), .ZN(new_n985_));
  INV_X1     g0600(.I(\b[81] ), .ZN(new_n986_));
  NOR2_X1    g0601(.A1(new_n985_), .A2(new_n986_), .ZN(new_n987_));
  INV_X1     g0602(.I(new_n987_), .ZN(new_n988_));
  INV_X1     g0603(.I(new_n979_), .ZN(new_n989_));
  AOI21_X1   g0604(.A1(new_n971_), .A2(\b[79] ), .B(\a[79] ), .ZN(new_n990_));
  OAI21_X1   g0605(.A1(new_n990_), .A2(new_n972_), .B(new_n980_), .ZN(new_n991_));
  NOR2_X1    g0606(.A1(\a[81] ), .A2(\b[81] ), .ZN(new_n992_));
  INV_X1     g0607(.I(new_n992_), .ZN(new_n993_));
  NAND3_X1   g0608(.A1(new_n991_), .A2(new_n989_), .A3(new_n993_), .ZN(new_n994_));
  AOI21_X1   g0609(.A1(new_n994_), .A2(new_n988_), .B(new_n984_), .ZN(new_n995_));
  NAND3_X1   g0610(.A1(new_n994_), .A2(new_n984_), .A3(new_n988_), .ZN(new_n996_));
  INV_X1     g0611(.I(new_n996_), .ZN(new_n997_));
  NOR2_X1    g0612(.A1(new_n997_), .A2(new_n995_), .ZN(new_n998_));
  XOR2_X1    g0613(.A1(new_n998_), .A2(\a[82] ), .Z(\f[82] ));
  OAI21_X1   g0614(.A1(\a[82] ), .A2(new_n995_), .B(new_n996_), .ZN(new_n1000_));
  XNOR2_X1   g0615(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1001_));
  XOR2_X1    g0616(.A1(new_n1000_), .A2(new_n1001_), .Z(\f[83] ));
  NOR2_X1    g0617(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1003_));
  NAND2_X1   g0618(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1004_));
  AOI21_X1   g0619(.A1(new_n1000_), .A2(new_n1004_), .B(new_n1003_), .ZN(new_n1005_));
  XOR2_X1    g0620(.A1(\a[84] ), .A2(\b[84] ), .Z(new_n1006_));
  XOR2_X1    g0621(.A1(new_n1005_), .A2(new_n1006_), .Z(\f[84] ));
  INV_X1     g0622(.I(\a[85] ), .ZN(new_n1008_));
  AND2_X2    g0623(.A1(\a[84] ), .A2(\b[84] ), .Z(new_n1009_));
  INV_X1     g0624(.I(\a[82] ), .ZN(new_n1010_));
  AOI21_X1   g0625(.A1(new_n981_), .A2(new_n993_), .B(new_n987_), .ZN(new_n1011_));
  OAI21_X1   g0626(.A1(new_n1011_), .A2(new_n984_), .B(new_n1010_), .ZN(new_n1012_));
  INV_X1     g0627(.I(new_n1004_), .ZN(new_n1013_));
  AOI21_X1   g0628(.A1(new_n1012_), .A2(new_n996_), .B(new_n1013_), .ZN(new_n1014_));
  NOR2_X1    g0629(.A1(\a[84] ), .A2(\b[84] ), .ZN(new_n1015_));
  NOR3_X1    g0630(.A1(new_n1014_), .A2(new_n1003_), .A3(new_n1015_), .ZN(new_n1016_));
  OAI21_X1   g0631(.A1(new_n1016_), .A2(new_n1009_), .B(\b[85] ), .ZN(new_n1017_));
  INV_X1     g0632(.I(\b[85] ), .ZN(new_n1018_));
  INV_X1     g0633(.I(new_n1015_), .ZN(new_n1019_));
  AOI21_X1   g0634(.A1(new_n1005_), .A2(new_n1019_), .B(new_n1009_), .ZN(new_n1020_));
  NAND2_X1   g0635(.A1(new_n1020_), .A2(new_n1018_), .ZN(new_n1021_));
  NAND2_X1   g0636(.A1(new_n1021_), .A2(new_n1017_), .ZN(new_n1022_));
  XOR2_X1    g0637(.A1(new_n1022_), .A2(new_n1008_), .Z(\f[85] ));
  NOR3_X1    g0638(.A1(new_n1016_), .A2(\b[85] ), .A3(new_n1009_), .ZN(new_n1024_));
  AOI21_X1   g0639(.A1(new_n1008_), .A2(new_n1017_), .B(new_n1024_), .ZN(new_n1025_));
  XOR2_X1    g0640(.A1(\a[86] ), .A2(\b[86] ), .Z(new_n1026_));
  XOR2_X1    g0641(.A1(new_n1025_), .A2(new_n1026_), .Z(\f[86] ));
  NOR2_X1    g0642(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n1028_));
  INV_X1     g0643(.I(new_n1028_), .ZN(new_n1029_));
  NAND2_X1   g0644(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n1030_));
  INV_X1     g0645(.I(new_n1030_), .ZN(new_n1031_));
  OAI21_X1   g0646(.A1(new_n1025_), .A2(new_n1031_), .B(new_n1029_), .ZN(new_n1032_));
  XNOR2_X1   g0647(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n1033_));
  XOR2_X1    g0648(.A1(new_n1032_), .A2(new_n1033_), .Z(\f[87] ));
  INV_X1     g0649(.I(\a[88] ), .ZN(new_n1035_));
  INV_X1     g0650(.I(\a[87] ), .ZN(new_n1036_));
  INV_X1     g0651(.I(\b[87] ), .ZN(new_n1037_));
  NOR2_X1    g0652(.A1(new_n1036_), .A2(new_n1037_), .ZN(new_n1038_));
  OAI21_X1   g0653(.A1(new_n1020_), .A2(new_n1018_), .B(new_n1008_), .ZN(new_n1039_));
  AOI21_X1   g0654(.A1(new_n1039_), .A2(new_n1021_), .B(new_n1031_), .ZN(new_n1040_));
  NOR2_X1    g0655(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n1041_));
  NOR3_X1    g0656(.A1(new_n1040_), .A2(new_n1028_), .A3(new_n1041_), .ZN(new_n1042_));
  OAI21_X1   g0657(.A1(new_n1042_), .A2(new_n1038_), .B(\b[88] ), .ZN(new_n1043_));
  NOR3_X1    g0658(.A1(new_n1042_), .A2(\b[88] ), .A3(new_n1038_), .ZN(new_n1044_));
  INV_X1     g0659(.I(new_n1044_), .ZN(new_n1045_));
  NAND2_X1   g0660(.A1(new_n1045_), .A2(new_n1043_), .ZN(new_n1046_));
  XOR2_X1    g0661(.A1(new_n1046_), .A2(new_n1035_), .Z(\f[88] ));
  AOI21_X1   g0662(.A1(new_n1035_), .A2(new_n1043_), .B(new_n1044_), .ZN(new_n1048_));
  XOR2_X1    g0663(.A1(\a[89] ), .A2(\b[89] ), .Z(new_n1049_));
  XOR2_X1    g0664(.A1(new_n1048_), .A2(new_n1049_), .Z(\f[89] ));
  NOR2_X1    g0665(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n1051_));
  INV_X1     g0666(.I(new_n1051_), .ZN(new_n1052_));
  NAND2_X1   g0667(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n1053_));
  INV_X1     g0668(.I(new_n1053_), .ZN(new_n1054_));
  OAI21_X1   g0669(.A1(new_n1048_), .A2(new_n1054_), .B(new_n1052_), .ZN(new_n1055_));
  XNOR2_X1   g0670(.A1(\a[90] ), .A2(\b[90] ), .ZN(new_n1056_));
  XOR2_X1    g0671(.A1(new_n1055_), .A2(new_n1056_), .Z(\f[90] ));
  INV_X1     g0672(.I(\b[91] ), .ZN(new_n1058_));
  AND2_X2    g0673(.A1(\a[90] ), .A2(\b[90] ), .Z(new_n1059_));
  INV_X1     g0674(.I(new_n1059_), .ZN(new_n1060_));
  INV_X1     g0675(.I(new_n1038_), .ZN(new_n1061_));
  OAI21_X1   g0676(.A1(new_n1032_), .A2(new_n1041_), .B(new_n1061_), .ZN(new_n1062_));
  AOI21_X1   g0677(.A1(new_n1062_), .A2(\b[88] ), .B(\a[88] ), .ZN(new_n1063_));
  OAI21_X1   g0678(.A1(new_n1063_), .A2(new_n1044_), .B(new_n1053_), .ZN(new_n1064_));
  NOR2_X1    g0679(.A1(\a[90] ), .A2(\b[90] ), .ZN(new_n1065_));
  INV_X1     g0680(.I(new_n1065_), .ZN(new_n1066_));
  NAND3_X1   g0681(.A1(new_n1064_), .A2(new_n1052_), .A3(new_n1066_), .ZN(new_n1067_));
  AOI21_X1   g0682(.A1(new_n1067_), .A2(new_n1060_), .B(new_n1058_), .ZN(new_n1068_));
  OAI21_X1   g0683(.A1(new_n1055_), .A2(new_n1065_), .B(new_n1060_), .ZN(new_n1069_));
  NOR2_X1    g0684(.A1(new_n1069_), .A2(\b[91] ), .ZN(new_n1070_));
  NOR2_X1    g0685(.A1(new_n1070_), .A2(new_n1068_), .ZN(new_n1071_));
  XOR2_X1    g0686(.A1(new_n1071_), .A2(\a[91] ), .Z(\f[91] ));
  NAND3_X1   g0687(.A1(new_n1067_), .A2(new_n1058_), .A3(new_n1060_), .ZN(new_n1073_));
  OAI21_X1   g0688(.A1(\a[91] ), .A2(new_n1068_), .B(new_n1073_), .ZN(new_n1074_));
  XNOR2_X1   g0689(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n1075_));
  XOR2_X1    g0690(.A1(new_n1074_), .A2(new_n1075_), .Z(\f[92] ));
  NOR2_X1    g0691(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n1077_));
  NAND2_X1   g0692(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n1078_));
  AOI21_X1   g0693(.A1(new_n1074_), .A2(new_n1078_), .B(new_n1077_), .ZN(new_n1079_));
  XOR2_X1    g0694(.A1(\a[93] ), .A2(\b[93] ), .Z(new_n1080_));
  XOR2_X1    g0695(.A1(new_n1079_), .A2(new_n1080_), .Z(\f[93] ));
  INV_X1     g0696(.I(\b[94] ), .ZN(new_n1082_));
  INV_X1     g0697(.I(\a[93] ), .ZN(new_n1083_));
  INV_X1     g0698(.I(\b[93] ), .ZN(new_n1084_));
  NOR2_X1    g0699(.A1(new_n1083_), .A2(new_n1084_), .ZN(new_n1085_));
  INV_X1     g0700(.I(new_n1085_), .ZN(new_n1086_));
  INV_X1     g0701(.I(new_n1077_), .ZN(new_n1087_));
  AOI21_X1   g0702(.A1(new_n1069_), .A2(\b[91] ), .B(\a[91] ), .ZN(new_n1088_));
  OAI21_X1   g0703(.A1(new_n1088_), .A2(new_n1070_), .B(new_n1078_), .ZN(new_n1089_));
  NOR2_X1    g0704(.A1(\a[93] ), .A2(\b[93] ), .ZN(new_n1090_));
  INV_X1     g0705(.I(new_n1090_), .ZN(new_n1091_));
  NAND3_X1   g0706(.A1(new_n1089_), .A2(new_n1087_), .A3(new_n1091_), .ZN(new_n1092_));
  AOI21_X1   g0707(.A1(new_n1092_), .A2(new_n1086_), .B(new_n1082_), .ZN(new_n1093_));
  NAND3_X1   g0708(.A1(new_n1092_), .A2(new_n1082_), .A3(new_n1086_), .ZN(new_n1094_));
  INV_X1     g0709(.I(new_n1094_), .ZN(new_n1095_));
  NOR2_X1    g0710(.A1(new_n1095_), .A2(new_n1093_), .ZN(new_n1096_));
  XOR2_X1    g0711(.A1(new_n1096_), .A2(\a[94] ), .Z(\f[94] ));
  OAI21_X1   g0712(.A1(\a[94] ), .A2(new_n1093_), .B(new_n1094_), .ZN(new_n1098_));
  XNOR2_X1   g0713(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1099_));
  XOR2_X1    g0714(.A1(new_n1098_), .A2(new_n1099_), .Z(\f[95] ));
  NOR2_X1    g0715(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1101_));
  NAND2_X1   g0716(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1102_));
  AOI21_X1   g0717(.A1(new_n1098_), .A2(new_n1102_), .B(new_n1101_), .ZN(new_n1103_));
  XOR2_X1    g0718(.A1(\a[96] ), .A2(\b[96] ), .Z(new_n1104_));
  XOR2_X1    g0719(.A1(new_n1103_), .A2(new_n1104_), .Z(\f[96] ));
  INV_X1     g0720(.I(\a[97] ), .ZN(new_n1106_));
  AND2_X2    g0721(.A1(\a[96] ), .A2(\b[96] ), .Z(new_n1107_));
  INV_X1     g0722(.I(\a[94] ), .ZN(new_n1108_));
  AOI21_X1   g0723(.A1(new_n1079_), .A2(new_n1091_), .B(new_n1085_), .ZN(new_n1109_));
  OAI21_X1   g0724(.A1(new_n1109_), .A2(new_n1082_), .B(new_n1108_), .ZN(new_n1110_));
  INV_X1     g0725(.I(new_n1102_), .ZN(new_n1111_));
  AOI21_X1   g0726(.A1(new_n1110_), .A2(new_n1094_), .B(new_n1111_), .ZN(new_n1112_));
  NOR2_X1    g0727(.A1(\a[96] ), .A2(\b[96] ), .ZN(new_n1113_));
  NOR3_X1    g0728(.A1(new_n1112_), .A2(new_n1101_), .A3(new_n1113_), .ZN(new_n1114_));
  OAI21_X1   g0729(.A1(new_n1114_), .A2(new_n1107_), .B(\b[97] ), .ZN(new_n1115_));
  INV_X1     g0730(.I(\b[97] ), .ZN(new_n1116_));
  INV_X1     g0731(.I(new_n1113_), .ZN(new_n1117_));
  AOI21_X1   g0732(.A1(new_n1103_), .A2(new_n1117_), .B(new_n1107_), .ZN(new_n1118_));
  NAND2_X1   g0733(.A1(new_n1118_), .A2(new_n1116_), .ZN(new_n1119_));
  NAND2_X1   g0734(.A1(new_n1119_), .A2(new_n1115_), .ZN(new_n1120_));
  XOR2_X1    g0735(.A1(new_n1120_), .A2(new_n1106_), .Z(\f[97] ));
  NOR3_X1    g0736(.A1(new_n1114_), .A2(\b[97] ), .A3(new_n1107_), .ZN(new_n1122_));
  AOI21_X1   g0737(.A1(new_n1106_), .A2(new_n1115_), .B(new_n1122_), .ZN(new_n1123_));
  XOR2_X1    g0738(.A1(\a[98] ), .A2(\b[98] ), .Z(new_n1124_));
  XOR2_X1    g0739(.A1(new_n1123_), .A2(new_n1124_), .Z(\f[98] ));
  NOR2_X1    g0740(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n1126_));
  INV_X1     g0741(.I(new_n1126_), .ZN(new_n1127_));
  NAND2_X1   g0742(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n1128_));
  INV_X1     g0743(.I(new_n1128_), .ZN(new_n1129_));
  OAI21_X1   g0744(.A1(new_n1123_), .A2(new_n1129_), .B(new_n1127_), .ZN(new_n1130_));
  XNOR2_X1   g0745(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n1131_));
  XOR2_X1    g0746(.A1(new_n1130_), .A2(new_n1131_), .Z(\f[99] ));
  INV_X1     g0747(.I(\a[100] ), .ZN(new_n1133_));
  INV_X1     g0748(.I(\a[99] ), .ZN(new_n1134_));
  INV_X1     g0749(.I(\b[99] ), .ZN(new_n1135_));
  NOR2_X1    g0750(.A1(new_n1134_), .A2(new_n1135_), .ZN(new_n1136_));
  OAI21_X1   g0751(.A1(new_n1118_), .A2(new_n1116_), .B(new_n1106_), .ZN(new_n1137_));
  AOI21_X1   g0752(.A1(new_n1137_), .A2(new_n1119_), .B(new_n1129_), .ZN(new_n1138_));
  NOR2_X1    g0753(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n1139_));
  NOR3_X1    g0754(.A1(new_n1138_), .A2(new_n1126_), .A3(new_n1139_), .ZN(new_n1140_));
  OAI21_X1   g0755(.A1(new_n1140_), .A2(new_n1136_), .B(\b[100] ), .ZN(new_n1141_));
  NOR3_X1    g0756(.A1(new_n1140_), .A2(\b[100] ), .A3(new_n1136_), .ZN(new_n1142_));
  INV_X1     g0757(.I(new_n1142_), .ZN(new_n1143_));
  NAND2_X1   g0758(.A1(new_n1143_), .A2(new_n1141_), .ZN(new_n1144_));
  XOR2_X1    g0759(.A1(new_n1144_), .A2(new_n1133_), .Z(\f[100] ));
  AOI21_X1   g0760(.A1(new_n1133_), .A2(new_n1141_), .B(new_n1142_), .ZN(new_n1146_));
  XOR2_X1    g0761(.A1(\a[101] ), .A2(\b[101] ), .Z(new_n1147_));
  XOR2_X1    g0762(.A1(new_n1146_), .A2(new_n1147_), .Z(\f[101] ));
  NOR2_X1    g0763(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n1149_));
  INV_X1     g0764(.I(new_n1149_), .ZN(new_n1150_));
  NAND2_X1   g0765(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n1151_));
  INV_X1     g0766(.I(new_n1151_), .ZN(new_n1152_));
  OAI21_X1   g0767(.A1(new_n1146_), .A2(new_n1152_), .B(new_n1150_), .ZN(new_n1153_));
  XNOR2_X1   g0768(.A1(\a[102] ), .A2(\b[102] ), .ZN(new_n1154_));
  XOR2_X1    g0769(.A1(new_n1153_), .A2(new_n1154_), .Z(\f[102] ));
  INV_X1     g0770(.I(\b[103] ), .ZN(new_n1156_));
  AND2_X2    g0771(.A1(\a[102] ), .A2(\b[102] ), .Z(new_n1157_));
  INV_X1     g0772(.I(new_n1157_), .ZN(new_n1158_));
  INV_X1     g0773(.I(new_n1136_), .ZN(new_n1159_));
  OAI21_X1   g0774(.A1(new_n1130_), .A2(new_n1139_), .B(new_n1159_), .ZN(new_n1160_));
  AOI21_X1   g0775(.A1(new_n1160_), .A2(\b[100] ), .B(\a[100] ), .ZN(new_n1161_));
  OAI21_X1   g0776(.A1(new_n1161_), .A2(new_n1142_), .B(new_n1151_), .ZN(new_n1162_));
  NOR2_X1    g0777(.A1(\a[102] ), .A2(\b[102] ), .ZN(new_n1163_));
  INV_X1     g0778(.I(new_n1163_), .ZN(new_n1164_));
  NAND3_X1   g0779(.A1(new_n1162_), .A2(new_n1150_), .A3(new_n1164_), .ZN(new_n1165_));
  AOI21_X1   g0780(.A1(new_n1165_), .A2(new_n1158_), .B(new_n1156_), .ZN(new_n1166_));
  OAI21_X1   g0781(.A1(new_n1153_), .A2(new_n1163_), .B(new_n1158_), .ZN(new_n1167_));
  NOR2_X1    g0782(.A1(new_n1167_), .A2(\b[103] ), .ZN(new_n1168_));
  NOR2_X1    g0783(.A1(new_n1168_), .A2(new_n1166_), .ZN(new_n1169_));
  XOR2_X1    g0784(.A1(new_n1169_), .A2(\a[103] ), .Z(\f[103] ));
  NAND3_X1   g0785(.A1(new_n1165_), .A2(new_n1156_), .A3(new_n1158_), .ZN(new_n1171_));
  OAI21_X1   g0786(.A1(\a[103] ), .A2(new_n1166_), .B(new_n1171_), .ZN(new_n1172_));
  XNOR2_X1   g0787(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1173_));
  XOR2_X1    g0788(.A1(new_n1172_), .A2(new_n1173_), .Z(\f[104] ));
  NOR2_X1    g0789(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1175_));
  NAND2_X1   g0790(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1176_));
  AOI21_X1   g0791(.A1(new_n1172_), .A2(new_n1176_), .B(new_n1175_), .ZN(new_n1177_));
  XOR2_X1    g0792(.A1(\a[105] ), .A2(\b[105] ), .Z(new_n1178_));
  XOR2_X1    g0793(.A1(new_n1177_), .A2(new_n1178_), .Z(\f[105] ));
  INV_X1     g0794(.I(\b[106] ), .ZN(new_n1180_));
  INV_X1     g0795(.I(\a[105] ), .ZN(new_n1181_));
  INV_X1     g0796(.I(\b[105] ), .ZN(new_n1182_));
  NOR2_X1    g0797(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1183_));
  NAND2_X1   g0798(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1184_));
  AOI21_X1   g0799(.A1(new_n1177_), .A2(new_n1184_), .B(new_n1183_), .ZN(new_n1185_));
  NOR2_X1    g0800(.A1(new_n1185_), .A2(new_n1180_), .ZN(new_n1186_));
  INV_X1     g0801(.I(new_n1183_), .ZN(new_n1187_));
  INV_X1     g0802(.I(new_n1175_), .ZN(new_n1188_));
  AOI21_X1   g0803(.A1(new_n1167_), .A2(\b[103] ), .B(\a[103] ), .ZN(new_n1189_));
  OAI21_X1   g0804(.A1(new_n1189_), .A2(new_n1168_), .B(new_n1176_), .ZN(new_n1190_));
  NAND3_X1   g0805(.A1(new_n1190_), .A2(new_n1188_), .A3(new_n1184_), .ZN(new_n1191_));
  NAND2_X1   g0806(.A1(new_n1191_), .A2(new_n1187_), .ZN(new_n1192_));
  NOR2_X1    g0807(.A1(new_n1192_), .A2(\b[106] ), .ZN(new_n1193_));
  NOR2_X1    g0808(.A1(new_n1186_), .A2(new_n1193_), .ZN(new_n1194_));
  XOR2_X1    g0809(.A1(new_n1194_), .A2(\a[106] ), .Z(\f[106] ));
  AOI21_X1   g0810(.A1(new_n1192_), .A2(\b[106] ), .B(\a[106] ), .ZN(new_n1196_));
  NOR2_X1    g0811(.A1(new_n1196_), .A2(new_n1193_), .ZN(new_n1197_));
  XOR2_X1    g0812(.A1(\a[107] ), .A2(\b[107] ), .Z(new_n1198_));
  XOR2_X1    g0813(.A1(new_n1197_), .A2(new_n1198_), .Z(\f[107] ));
  NOR2_X1    g0814(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1200_));
  INV_X1     g0815(.I(new_n1200_), .ZN(new_n1201_));
  NAND2_X1   g0816(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1202_));
  OAI21_X1   g0817(.A1(new_n1196_), .A2(new_n1193_), .B(new_n1202_), .ZN(new_n1203_));
  NAND2_X1   g0818(.A1(new_n1203_), .A2(new_n1201_), .ZN(new_n1204_));
  XNOR2_X1   g0819(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1205_));
  XOR2_X1    g0820(.A1(new_n1204_), .A2(new_n1205_), .Z(\f[108] ));
  INV_X1     g0821(.I(\a[109] ), .ZN(new_n1207_));
  INV_X1     g0822(.I(\a[108] ), .ZN(new_n1208_));
  INV_X1     g0823(.I(\b[108] ), .ZN(new_n1209_));
  NOR2_X1    g0824(.A1(new_n1208_), .A2(new_n1209_), .ZN(new_n1210_));
  NAND2_X1   g0825(.A1(new_n1185_), .A2(new_n1180_), .ZN(new_n1211_));
  INV_X1     g0826(.I(\a[106] ), .ZN(new_n1212_));
  OAI21_X1   g0827(.A1(new_n1185_), .A2(new_n1180_), .B(new_n1212_), .ZN(new_n1213_));
  INV_X1     g0828(.I(new_n1202_), .ZN(new_n1214_));
  AOI21_X1   g0829(.A1(new_n1213_), .A2(new_n1211_), .B(new_n1214_), .ZN(new_n1215_));
  NOR2_X1    g0830(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1216_));
  NOR3_X1    g0831(.A1(new_n1215_), .A2(new_n1200_), .A3(new_n1216_), .ZN(new_n1217_));
  OAI21_X1   g0832(.A1(new_n1217_), .A2(new_n1210_), .B(\b[109] ), .ZN(new_n1218_));
  INV_X1     g0833(.I(\b[109] ), .ZN(new_n1219_));
  INV_X1     g0834(.I(new_n1210_), .ZN(new_n1220_));
  INV_X1     g0835(.I(new_n1216_), .ZN(new_n1221_));
  NAND3_X1   g0836(.A1(new_n1203_), .A2(new_n1201_), .A3(new_n1221_), .ZN(new_n1222_));
  NAND3_X1   g0837(.A1(new_n1222_), .A2(new_n1219_), .A3(new_n1220_), .ZN(new_n1223_));
  NAND2_X1   g0838(.A1(new_n1218_), .A2(new_n1223_), .ZN(new_n1224_));
  XOR2_X1    g0839(.A1(new_n1224_), .A2(new_n1207_), .Z(\f[109] ));
  AOI21_X1   g0840(.A1(new_n1222_), .A2(new_n1220_), .B(new_n1219_), .ZN(new_n1226_));
  OAI21_X1   g0841(.A1(\a[109] ), .A2(new_n1226_), .B(new_n1223_), .ZN(new_n1227_));
  XNOR2_X1   g0842(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1228_));
  XOR2_X1    g0843(.A1(new_n1227_), .A2(new_n1228_), .Z(\f[110] ));
  NOR2_X1    g0844(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1230_));
  NAND2_X1   g0845(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1231_));
  AOI21_X1   g0846(.A1(new_n1227_), .A2(new_n1231_), .B(new_n1230_), .ZN(new_n1232_));
  XOR2_X1    g0847(.A1(\a[111] ), .A2(\b[111] ), .Z(new_n1233_));
  XOR2_X1    g0848(.A1(new_n1232_), .A2(new_n1233_), .Z(\f[111] ));
  INV_X1     g0849(.I(\b[112] ), .ZN(new_n1235_));
  INV_X1     g0850(.I(\a[111] ), .ZN(new_n1236_));
  INV_X1     g0851(.I(\b[111] ), .ZN(new_n1237_));
  NOR2_X1    g0852(.A1(new_n1236_), .A2(new_n1237_), .ZN(new_n1238_));
  NOR2_X1    g0853(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1239_));
  INV_X1     g0854(.I(new_n1239_), .ZN(new_n1240_));
  AOI21_X1   g0855(.A1(new_n1232_), .A2(new_n1240_), .B(new_n1238_), .ZN(new_n1241_));
  NOR2_X1    g0856(.A1(new_n1241_), .A2(new_n1235_), .ZN(new_n1242_));
  NOR3_X1    g0857(.A1(new_n1217_), .A2(\b[109] ), .A3(new_n1210_), .ZN(new_n1243_));
  AOI21_X1   g0858(.A1(new_n1207_), .A2(new_n1218_), .B(new_n1243_), .ZN(new_n1244_));
  INV_X1     g0859(.I(new_n1230_), .ZN(new_n1245_));
  INV_X1     g0860(.I(new_n1231_), .ZN(new_n1246_));
  OAI21_X1   g0861(.A1(new_n1244_), .A2(new_n1246_), .B(new_n1245_), .ZN(new_n1247_));
  INV_X1     g0862(.I(new_n1238_), .ZN(new_n1248_));
  OAI21_X1   g0863(.A1(new_n1247_), .A2(new_n1239_), .B(new_n1248_), .ZN(new_n1249_));
  NOR2_X1    g0864(.A1(new_n1249_), .A2(\b[112] ), .ZN(new_n1250_));
  NOR2_X1    g0865(.A1(new_n1250_), .A2(new_n1242_), .ZN(new_n1251_));
  XOR2_X1    g0866(.A1(new_n1251_), .A2(\a[112] ), .Z(\f[112] ));
  NAND2_X1   g0867(.A1(new_n1241_), .A2(new_n1235_), .ZN(new_n1253_));
  INV_X1     g0868(.I(\a[112] ), .ZN(new_n1254_));
  OAI21_X1   g0869(.A1(new_n1241_), .A2(new_n1235_), .B(new_n1254_), .ZN(new_n1255_));
  NAND2_X1   g0870(.A1(new_n1255_), .A2(new_n1253_), .ZN(new_n1256_));
  XNOR2_X1   g0871(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1257_));
  XOR2_X1    g0872(.A1(new_n1256_), .A2(new_n1257_), .Z(\f[113] ));
  NOR2_X1    g0873(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1259_));
  NAND2_X1   g0874(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1260_));
  INV_X1     g0875(.I(new_n1260_), .ZN(new_n1261_));
  AOI21_X1   g0876(.A1(new_n1255_), .A2(new_n1253_), .B(new_n1261_), .ZN(new_n1262_));
  NOR2_X1    g0877(.A1(new_n1262_), .A2(new_n1259_), .ZN(new_n1263_));
  XOR2_X1    g0878(.A1(\a[114] ), .A2(\b[114] ), .Z(new_n1264_));
  XOR2_X1    g0879(.A1(new_n1263_), .A2(new_n1264_), .Z(\f[114] ));
  INV_X1     g0880(.I(\a[115] ), .ZN(new_n1266_));
  INV_X1     g0881(.I(\a[114] ), .ZN(new_n1267_));
  INV_X1     g0882(.I(\b[114] ), .ZN(new_n1268_));
  NOR2_X1    g0883(.A1(new_n1267_), .A2(new_n1268_), .ZN(new_n1269_));
  NOR2_X1    g0884(.A1(\a[114] ), .A2(\b[114] ), .ZN(new_n1270_));
  NOR3_X1    g0885(.A1(new_n1262_), .A2(new_n1259_), .A3(new_n1270_), .ZN(new_n1271_));
  OAI21_X1   g0886(.A1(new_n1271_), .A2(new_n1269_), .B(\b[115] ), .ZN(new_n1272_));
  INV_X1     g0887(.I(\b[115] ), .ZN(new_n1273_));
  INV_X1     g0888(.I(new_n1269_), .ZN(new_n1274_));
  INV_X1     g0889(.I(new_n1259_), .ZN(new_n1275_));
  AOI21_X1   g0890(.A1(new_n1249_), .A2(\b[112] ), .B(\a[112] ), .ZN(new_n1276_));
  OAI21_X1   g0891(.A1(new_n1276_), .A2(new_n1250_), .B(new_n1260_), .ZN(new_n1277_));
  INV_X1     g0892(.I(new_n1270_), .ZN(new_n1278_));
  NAND3_X1   g0893(.A1(new_n1277_), .A2(new_n1275_), .A3(new_n1278_), .ZN(new_n1279_));
  NAND3_X1   g0894(.A1(new_n1279_), .A2(new_n1273_), .A3(new_n1274_), .ZN(new_n1280_));
  NAND2_X1   g0895(.A1(new_n1280_), .A2(new_n1272_), .ZN(new_n1281_));
  XOR2_X1    g0896(.A1(new_n1281_), .A2(new_n1266_), .Z(\f[115] ));
  NOR3_X1    g0897(.A1(new_n1271_), .A2(\b[115] ), .A3(new_n1269_), .ZN(new_n1283_));
  AOI21_X1   g0898(.A1(new_n1266_), .A2(new_n1272_), .B(new_n1283_), .ZN(new_n1284_));
  XOR2_X1    g0899(.A1(\a[116] ), .A2(\b[116] ), .Z(new_n1285_));
  XOR2_X1    g0900(.A1(new_n1284_), .A2(new_n1285_), .Z(\f[116] ));
  NOR2_X1    g0901(.A1(\a[116] ), .A2(\b[116] ), .ZN(new_n1287_));
  INV_X1     g0902(.I(new_n1287_), .ZN(new_n1288_));
  NAND2_X1   g0903(.A1(\a[116] ), .A2(\b[116] ), .ZN(new_n1289_));
  INV_X1     g0904(.I(new_n1289_), .ZN(new_n1290_));
  OAI21_X1   g0905(.A1(new_n1284_), .A2(new_n1290_), .B(new_n1288_), .ZN(new_n1291_));
  XNOR2_X1   g0906(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1292_));
  XOR2_X1    g0907(.A1(new_n1291_), .A2(new_n1292_), .Z(\f[117] ));
  INV_X1     g0908(.I(\b[118] ), .ZN(new_n1294_));
  AOI21_X1   g0909(.A1(new_n1279_), .A2(new_n1274_), .B(new_n1273_), .ZN(new_n1295_));
  OAI21_X1   g0910(.A1(\a[115] ), .A2(new_n1295_), .B(new_n1280_), .ZN(new_n1296_));
  AOI21_X1   g0911(.A1(new_n1296_), .A2(new_n1289_), .B(new_n1287_), .ZN(new_n1297_));
  INV_X1     g0912(.I(\a[117] ), .ZN(new_n1298_));
  INV_X1     g0913(.I(\b[117] ), .ZN(new_n1299_));
  NOR2_X1    g0914(.A1(new_n1298_), .A2(new_n1299_), .ZN(new_n1300_));
  NOR2_X1    g0915(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1301_));
  INV_X1     g0916(.I(new_n1301_), .ZN(new_n1302_));
  AOI21_X1   g0917(.A1(new_n1297_), .A2(new_n1302_), .B(new_n1300_), .ZN(new_n1303_));
  NOR2_X1    g0918(.A1(new_n1303_), .A2(new_n1294_), .ZN(new_n1304_));
  INV_X1     g0919(.I(new_n1300_), .ZN(new_n1305_));
  OAI21_X1   g0920(.A1(new_n1291_), .A2(new_n1301_), .B(new_n1305_), .ZN(new_n1306_));
  NOR2_X1    g0921(.A1(new_n1306_), .A2(\b[118] ), .ZN(new_n1307_));
  NOR2_X1    g0922(.A1(new_n1304_), .A2(new_n1307_), .ZN(new_n1308_));
  XOR2_X1    g0923(.A1(new_n1308_), .A2(\a[118] ), .Z(\f[118] ));
  AOI21_X1   g0924(.A1(new_n1306_), .A2(\b[118] ), .B(\a[118] ), .ZN(new_n1310_));
  NOR2_X1    g0925(.A1(new_n1310_), .A2(new_n1307_), .ZN(new_n1311_));
  XOR2_X1    g0926(.A1(\a[119] ), .A2(\b[119] ), .Z(new_n1312_));
  XOR2_X1    g0927(.A1(new_n1311_), .A2(new_n1312_), .Z(\f[119] ));
  NOR2_X1    g0928(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1314_));
  INV_X1     g0929(.I(new_n1314_), .ZN(new_n1315_));
  NAND2_X1   g0930(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1316_));
  OAI21_X1   g0931(.A1(new_n1310_), .A2(new_n1307_), .B(new_n1316_), .ZN(new_n1317_));
  NAND2_X1   g0932(.A1(new_n1317_), .A2(new_n1315_), .ZN(new_n1318_));
  XNOR2_X1   g0933(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1319_));
  XOR2_X1    g0934(.A1(new_n1318_), .A2(new_n1319_), .Z(\f[120] ));
  INV_X1     g0935(.I(\a[121] ), .ZN(new_n1321_));
  INV_X1     g0936(.I(\a[120] ), .ZN(new_n1322_));
  INV_X1     g0937(.I(\b[120] ), .ZN(new_n1323_));
  NOR2_X1    g0938(.A1(new_n1322_), .A2(new_n1323_), .ZN(new_n1324_));
  NAND2_X1   g0939(.A1(new_n1303_), .A2(new_n1294_), .ZN(new_n1325_));
  INV_X1     g0940(.I(\a[118] ), .ZN(new_n1326_));
  OAI21_X1   g0941(.A1(new_n1303_), .A2(new_n1294_), .B(new_n1326_), .ZN(new_n1327_));
  INV_X1     g0942(.I(new_n1316_), .ZN(new_n1328_));
  AOI21_X1   g0943(.A1(new_n1327_), .A2(new_n1325_), .B(new_n1328_), .ZN(new_n1329_));
  NOR2_X1    g0944(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1330_));
  NOR3_X1    g0945(.A1(new_n1329_), .A2(new_n1314_), .A3(new_n1330_), .ZN(new_n1331_));
  OAI21_X1   g0946(.A1(new_n1331_), .A2(new_n1324_), .B(\b[121] ), .ZN(new_n1332_));
  INV_X1     g0947(.I(\b[121] ), .ZN(new_n1333_));
  INV_X1     g0948(.I(new_n1324_), .ZN(new_n1334_));
  INV_X1     g0949(.I(new_n1330_), .ZN(new_n1335_));
  NAND3_X1   g0950(.A1(new_n1317_), .A2(new_n1315_), .A3(new_n1335_), .ZN(new_n1336_));
  NAND3_X1   g0951(.A1(new_n1336_), .A2(new_n1333_), .A3(new_n1334_), .ZN(new_n1337_));
  NAND2_X1   g0952(.A1(new_n1332_), .A2(new_n1337_), .ZN(new_n1338_));
  XOR2_X1    g0953(.A1(new_n1338_), .A2(new_n1321_), .Z(\f[121] ));
  AOI21_X1   g0954(.A1(new_n1336_), .A2(new_n1334_), .B(new_n1333_), .ZN(new_n1340_));
  OAI21_X1   g0955(.A1(\a[121] ), .A2(new_n1340_), .B(new_n1337_), .ZN(new_n1341_));
  XNOR2_X1   g0956(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1342_));
  XOR2_X1    g0957(.A1(new_n1341_), .A2(new_n1342_), .Z(\f[122] ));
  NOR2_X1    g0958(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1344_));
  NAND2_X1   g0959(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1345_));
  AOI21_X1   g0960(.A1(new_n1341_), .A2(new_n1345_), .B(new_n1344_), .ZN(new_n1346_));
  XOR2_X1    g0961(.A1(\a[123] ), .A2(\b[123] ), .Z(new_n1347_));
  XOR2_X1    g0962(.A1(new_n1346_), .A2(new_n1347_), .Z(\f[123] ));
  INV_X1     g0963(.I(\a[124] ), .ZN(new_n1349_));
  NOR3_X1    g0964(.A1(new_n1331_), .A2(\b[121] ), .A3(new_n1324_), .ZN(new_n1350_));
  AOI21_X1   g0965(.A1(new_n1321_), .A2(new_n1332_), .B(new_n1350_), .ZN(new_n1351_));
  INV_X1     g0966(.I(new_n1344_), .ZN(new_n1352_));
  INV_X1     g0967(.I(new_n1345_), .ZN(new_n1353_));
  OAI21_X1   g0968(.A1(new_n1351_), .A2(new_n1353_), .B(new_n1352_), .ZN(new_n1354_));
  INV_X1     g0969(.I(\a[123] ), .ZN(new_n1355_));
  INV_X1     g0970(.I(\b[123] ), .ZN(new_n1356_));
  NOR2_X1    g0971(.A1(new_n1355_), .A2(new_n1356_), .ZN(new_n1357_));
  INV_X1     g0972(.I(new_n1357_), .ZN(new_n1358_));
  NOR2_X1    g0973(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1359_));
  OAI21_X1   g0974(.A1(new_n1354_), .A2(new_n1359_), .B(new_n1358_), .ZN(new_n1360_));
  NAND2_X1   g0975(.A1(new_n1360_), .A2(\b[124] ), .ZN(new_n1361_));
  INV_X1     g0976(.I(\b[124] ), .ZN(new_n1362_));
  INV_X1     g0977(.I(new_n1359_), .ZN(new_n1363_));
  AOI21_X1   g0978(.A1(new_n1346_), .A2(new_n1363_), .B(new_n1357_), .ZN(new_n1364_));
  NAND2_X1   g0979(.A1(new_n1364_), .A2(new_n1362_), .ZN(new_n1365_));
  NAND2_X1   g0980(.A1(new_n1361_), .A2(new_n1365_), .ZN(new_n1366_));
  XOR2_X1    g0981(.A1(new_n1366_), .A2(new_n1349_), .Z(\f[124] ));
  OAI21_X1   g0982(.A1(new_n1364_), .A2(new_n1362_), .B(new_n1349_), .ZN(new_n1368_));
  NAND2_X1   g0983(.A1(new_n1368_), .A2(new_n1365_), .ZN(new_n1369_));
  XNOR2_X1   g0984(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1370_));
  XOR2_X1    g0985(.A1(new_n1369_), .A2(new_n1370_), .Z(\f[125] ));
  NOR2_X1    g0986(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1372_));
  NAND2_X1   g0987(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1373_));
  INV_X1     g0988(.I(new_n1373_), .ZN(new_n1374_));
  AOI21_X1   g0989(.A1(new_n1368_), .A2(new_n1365_), .B(new_n1374_), .ZN(new_n1375_));
  NOR2_X1    g0990(.A1(new_n1375_), .A2(new_n1372_), .ZN(new_n1376_));
  XOR2_X1    g0991(.A1(\a[126] ), .A2(\b[126] ), .Z(new_n1377_));
  XOR2_X1    g0992(.A1(new_n1376_), .A2(new_n1377_), .Z(\f[126] ));
  INV_X1     g0993(.I(\a[126] ), .ZN(new_n1379_));
  INV_X1     g0994(.I(\b[126] ), .ZN(new_n1380_));
  NOR2_X1    g0995(.A1(new_n1379_), .A2(new_n1380_), .ZN(new_n1381_));
  NOR2_X1    g0996(.A1(\a[126] ), .A2(\b[126] ), .ZN(new_n1382_));
  NOR3_X1    g0997(.A1(new_n1375_), .A2(new_n1372_), .A3(new_n1382_), .ZN(new_n1383_));
  XNOR2_X1   g0998(.A1(\a[127] ), .A2(\b[127] ), .ZN(new_n1384_));
  INV_X1     g0999(.I(new_n1384_), .ZN(new_n1385_));
  NOR3_X1    g1000(.A1(new_n1383_), .A2(new_n1381_), .A3(new_n1385_), .ZN(new_n1386_));
  INV_X1     g1001(.I(new_n1381_), .ZN(new_n1387_));
  INV_X1     g1002(.I(new_n1372_), .ZN(new_n1388_));
  NOR2_X1    g1003(.A1(new_n1360_), .A2(\b[124] ), .ZN(new_n1389_));
  AOI21_X1   g1004(.A1(new_n1360_), .A2(\b[124] ), .B(\a[124] ), .ZN(new_n1390_));
  OAI21_X1   g1005(.A1(new_n1390_), .A2(new_n1389_), .B(new_n1373_), .ZN(new_n1391_));
  INV_X1     g1006(.I(new_n1382_), .ZN(new_n1392_));
  NAND3_X1   g1007(.A1(new_n1391_), .A2(new_n1388_), .A3(new_n1392_), .ZN(new_n1393_));
  AOI21_X1   g1008(.A1(new_n1393_), .A2(new_n1387_), .B(new_n1384_), .ZN(new_n1394_));
  NOR2_X1    g1009(.A1(new_n1394_), .A2(new_n1386_), .ZN(\f[127] ));
  INV_X1     g1010(.I(\a[127] ), .ZN(new_n1396_));
  OAI21_X1   g1011(.A1(new_n1383_), .A2(new_n1381_), .B(\b[127] ), .ZN(new_n1397_));
  NOR3_X1    g1012(.A1(new_n1383_), .A2(\b[127] ), .A3(new_n1381_), .ZN(new_n1398_));
  AOI21_X1   g1013(.A1(new_n1396_), .A2(new_n1397_), .B(new_n1398_), .ZN(cOut));
endmodule


