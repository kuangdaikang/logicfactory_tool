// Benchmark "bar" written by ABC on Fri Sep 15 11:20:26 2023

module bar ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] ,
    \shift[3] , \shift[4] , \shift[5] , \shift[6] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] ,
    \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ;
  wire new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_,
    new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_,
    new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_,
    new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_,
    new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_,
    new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_,
    new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_,
    new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_,
    new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_,
    new_n1580_, new_n1581_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_,
    new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_,
    new_n1778_, new_n1779_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2080_, new_n2081_, new_n2082_, new_n2083_,
    new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_,
    new_n2090_, new_n2091_, new_n2092_, new_n2093_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2146_, new_n2147_, new_n2148_,
    new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2183_, new_n2184_, new_n2186_, new_n2187_, new_n2189_,
    new_n2190_, new_n2192_, new_n2193_, new_n2195_, new_n2196_, new_n2198_,
    new_n2199_, new_n2201_, new_n2202_, new_n2204_, new_n2205_, new_n2207_,
    new_n2208_, new_n2210_, new_n2211_, new_n2213_, new_n2214_, new_n2216_,
    new_n2217_, new_n2219_, new_n2220_, new_n2222_, new_n2223_, new_n2225_,
    new_n2226_, new_n2228_, new_n2229_, new_n2231_, new_n2232_, new_n2234_,
    new_n2235_, new_n2237_, new_n2238_, new_n2240_, new_n2241_, new_n2243_,
    new_n2244_, new_n2246_, new_n2247_, new_n2249_, new_n2250_, new_n2252_,
    new_n2253_, new_n2255_, new_n2256_, new_n2258_, new_n2259_, new_n2261_,
    new_n2262_, new_n2264_, new_n2265_, new_n2267_, new_n2268_, new_n2270_,
    new_n2271_, new_n2273_, new_n2274_, new_n2276_, new_n2277_, new_n2279_,
    new_n2280_, new_n2282_, new_n2283_, new_n2285_, new_n2286_, new_n2288_,
    new_n2289_, new_n2291_, new_n2292_, new_n2294_, new_n2295_, new_n2297_,
    new_n2298_, new_n2300_, new_n2301_, new_n2303_, new_n2304_, new_n2306_,
    new_n2307_, new_n2309_, new_n2310_, new_n2312_, new_n2313_, new_n2315_,
    new_n2316_, new_n2318_, new_n2319_, new_n2321_, new_n2322_, new_n2324_,
    new_n2325_, new_n2327_, new_n2328_, new_n2330_, new_n2331_, new_n2333_,
    new_n2334_, new_n2336_, new_n2337_, new_n2339_, new_n2340_, new_n2342_,
    new_n2343_, new_n2345_, new_n2346_, new_n2348_, new_n2349_, new_n2351_,
    new_n2352_, new_n2354_, new_n2355_, new_n2357_, new_n2358_, new_n2360_,
    new_n2361_, new_n2363_, new_n2364_, new_n2366_, new_n2367_, new_n2369_,
    new_n2370_, new_n2372_, new_n2373_;
  INV_X1     g0000(.I(\shift[6] ), .ZN(new_n264_));
  INV_X1     g0001(.I(\shift[5] ), .ZN(new_n265_));
  INV_X1     g0002(.I(\shift[2] ), .ZN(new_n266_));
  NAND2_X1   g0003(.A1(\a[67] ), .A2(\shift[0] ), .ZN(new_n267_));
  INV_X1     g0004(.I(\shift[0] ), .ZN(new_n268_));
  NAND2_X1   g0005(.A1(new_n268_), .A2(\a[68] ), .ZN(new_n269_));
  AOI21_X1   g0006(.A1(new_n269_), .A2(new_n267_), .B(\shift[1] ), .ZN(new_n270_));
  INV_X1     g0007(.I(\shift[1] ), .ZN(new_n271_));
  NAND2_X1   g0008(.A1(\a[65] ), .A2(\shift[0] ), .ZN(new_n272_));
  NAND2_X1   g0009(.A1(new_n268_), .A2(\a[66] ), .ZN(new_n273_));
  AOI21_X1   g0010(.A1(new_n273_), .A2(new_n272_), .B(new_n271_), .ZN(new_n274_));
  OAI21_X1   g0011(.A1(new_n270_), .A2(new_n274_), .B(\shift[3] ), .ZN(new_n275_));
  INV_X1     g0012(.I(\shift[3] ), .ZN(new_n276_));
  NAND2_X1   g0013(.A1(\a[75] ), .A2(\shift[0] ), .ZN(new_n277_));
  NAND2_X1   g0014(.A1(new_n268_), .A2(\a[76] ), .ZN(new_n278_));
  AOI21_X1   g0015(.A1(new_n278_), .A2(new_n277_), .B(\shift[1] ), .ZN(new_n279_));
  NAND2_X1   g0016(.A1(\a[73] ), .A2(\shift[0] ), .ZN(new_n280_));
  NAND2_X1   g0017(.A1(new_n268_), .A2(\a[74] ), .ZN(new_n281_));
  AOI21_X1   g0018(.A1(new_n281_), .A2(new_n280_), .B(new_n271_), .ZN(new_n282_));
  OAI21_X1   g0019(.A1(new_n279_), .A2(new_n282_), .B(new_n276_), .ZN(new_n283_));
  AOI21_X1   g0020(.A1(new_n275_), .A2(new_n283_), .B(new_n266_), .ZN(new_n284_));
  NAND2_X1   g0021(.A1(\a[79] ), .A2(\shift[0] ), .ZN(new_n285_));
  NAND2_X1   g0022(.A1(new_n268_), .A2(\a[80] ), .ZN(new_n286_));
  AOI21_X1   g0023(.A1(new_n286_), .A2(new_n285_), .B(\shift[1] ), .ZN(new_n287_));
  NAND2_X1   g0024(.A1(\a[77] ), .A2(\shift[0] ), .ZN(new_n288_));
  NAND2_X1   g0025(.A1(new_n268_), .A2(\a[78] ), .ZN(new_n289_));
  AOI21_X1   g0026(.A1(new_n289_), .A2(new_n288_), .B(new_n271_), .ZN(new_n290_));
  OAI21_X1   g0027(.A1(new_n287_), .A2(new_n290_), .B(new_n276_), .ZN(new_n291_));
  NAND2_X1   g0028(.A1(\a[71] ), .A2(\shift[0] ), .ZN(new_n292_));
  NAND2_X1   g0029(.A1(new_n268_), .A2(\a[72] ), .ZN(new_n293_));
  AOI21_X1   g0030(.A1(new_n293_), .A2(new_n292_), .B(\shift[1] ), .ZN(new_n294_));
  NAND2_X1   g0031(.A1(\a[69] ), .A2(\shift[0] ), .ZN(new_n295_));
  NAND2_X1   g0032(.A1(new_n268_), .A2(\a[70] ), .ZN(new_n296_));
  AOI21_X1   g0033(.A1(new_n296_), .A2(new_n295_), .B(new_n271_), .ZN(new_n297_));
  OAI21_X1   g0034(.A1(new_n294_), .A2(new_n297_), .B(\shift[3] ), .ZN(new_n298_));
  AOI21_X1   g0035(.A1(new_n291_), .A2(new_n298_), .B(\shift[2] ), .ZN(new_n299_));
  OAI21_X1   g0036(.A1(new_n284_), .A2(new_n299_), .B(\shift[4] ), .ZN(new_n300_));
  INV_X1     g0037(.I(\shift[4] ), .ZN(new_n301_));
  NAND2_X1   g0038(.A1(\a[83] ), .A2(\shift[0] ), .ZN(new_n302_));
  NAND2_X1   g0039(.A1(new_n268_), .A2(\a[84] ), .ZN(new_n303_));
  AOI21_X1   g0040(.A1(new_n303_), .A2(new_n302_), .B(\shift[1] ), .ZN(new_n304_));
  NAND2_X1   g0041(.A1(\a[81] ), .A2(\shift[0] ), .ZN(new_n305_));
  NAND2_X1   g0042(.A1(new_n268_), .A2(\a[82] ), .ZN(new_n306_));
  AOI21_X1   g0043(.A1(new_n306_), .A2(new_n305_), .B(new_n271_), .ZN(new_n307_));
  OAI21_X1   g0044(.A1(new_n304_), .A2(new_n307_), .B(\shift[3] ), .ZN(new_n308_));
  NAND2_X1   g0045(.A1(\a[91] ), .A2(\shift[0] ), .ZN(new_n309_));
  NAND2_X1   g0046(.A1(new_n268_), .A2(\a[92] ), .ZN(new_n310_));
  AOI21_X1   g0047(.A1(new_n310_), .A2(new_n309_), .B(\shift[1] ), .ZN(new_n311_));
  NAND2_X1   g0048(.A1(\a[89] ), .A2(\shift[0] ), .ZN(new_n312_));
  NAND2_X1   g0049(.A1(new_n268_), .A2(\a[90] ), .ZN(new_n313_));
  AOI21_X1   g0050(.A1(new_n313_), .A2(new_n312_), .B(new_n271_), .ZN(new_n314_));
  OAI21_X1   g0051(.A1(new_n311_), .A2(new_n314_), .B(new_n276_), .ZN(new_n315_));
  AOI21_X1   g0052(.A1(new_n308_), .A2(new_n315_), .B(new_n266_), .ZN(new_n316_));
  NAND2_X1   g0053(.A1(\a[95] ), .A2(\shift[0] ), .ZN(new_n317_));
  NAND2_X1   g0054(.A1(new_n268_), .A2(\a[96] ), .ZN(new_n318_));
  AOI21_X1   g0055(.A1(new_n318_), .A2(new_n317_), .B(\shift[1] ), .ZN(new_n319_));
  NAND2_X1   g0056(.A1(\a[93] ), .A2(\shift[0] ), .ZN(new_n320_));
  NAND2_X1   g0057(.A1(new_n268_), .A2(\a[94] ), .ZN(new_n321_));
  AOI21_X1   g0058(.A1(new_n321_), .A2(new_n320_), .B(new_n271_), .ZN(new_n322_));
  OAI21_X1   g0059(.A1(new_n319_), .A2(new_n322_), .B(new_n276_), .ZN(new_n323_));
  NAND2_X1   g0060(.A1(\a[87] ), .A2(\shift[0] ), .ZN(new_n324_));
  NAND2_X1   g0061(.A1(new_n268_), .A2(\a[88] ), .ZN(new_n325_));
  AOI21_X1   g0062(.A1(new_n325_), .A2(new_n324_), .B(\shift[1] ), .ZN(new_n326_));
  NAND2_X1   g0063(.A1(\a[85] ), .A2(\shift[0] ), .ZN(new_n327_));
  NAND2_X1   g0064(.A1(new_n268_), .A2(\a[86] ), .ZN(new_n328_));
  AOI21_X1   g0065(.A1(new_n328_), .A2(new_n327_), .B(new_n271_), .ZN(new_n329_));
  OAI21_X1   g0066(.A1(new_n326_), .A2(new_n329_), .B(\shift[3] ), .ZN(new_n330_));
  AOI21_X1   g0067(.A1(new_n323_), .A2(new_n330_), .B(\shift[2] ), .ZN(new_n331_));
  OAI21_X1   g0068(.A1(new_n316_), .A2(new_n331_), .B(new_n301_), .ZN(new_n332_));
  AOI21_X1   g0069(.A1(new_n300_), .A2(new_n332_), .B(new_n265_), .ZN(new_n333_));
  NAND2_X1   g0070(.A1(\a[99] ), .A2(\shift[0] ), .ZN(new_n334_));
  NAND2_X1   g0071(.A1(new_n268_), .A2(\a[100] ), .ZN(new_n335_));
  AOI21_X1   g0072(.A1(new_n335_), .A2(new_n334_), .B(\shift[1] ), .ZN(new_n336_));
  NAND2_X1   g0073(.A1(\a[97] ), .A2(\shift[0] ), .ZN(new_n337_));
  NAND2_X1   g0074(.A1(new_n268_), .A2(\a[98] ), .ZN(new_n338_));
  AOI21_X1   g0075(.A1(new_n338_), .A2(new_n337_), .B(new_n271_), .ZN(new_n339_));
  OAI21_X1   g0076(.A1(new_n336_), .A2(new_n339_), .B(\shift[3] ), .ZN(new_n340_));
  NAND2_X1   g0077(.A1(\a[107] ), .A2(\shift[0] ), .ZN(new_n341_));
  NAND2_X1   g0078(.A1(new_n268_), .A2(\a[108] ), .ZN(new_n342_));
  AOI21_X1   g0079(.A1(new_n342_), .A2(new_n341_), .B(\shift[1] ), .ZN(new_n343_));
  NAND2_X1   g0080(.A1(\a[105] ), .A2(\shift[0] ), .ZN(new_n344_));
  NAND2_X1   g0081(.A1(new_n268_), .A2(\a[106] ), .ZN(new_n345_));
  AOI21_X1   g0082(.A1(new_n345_), .A2(new_n344_), .B(new_n271_), .ZN(new_n346_));
  OAI21_X1   g0083(.A1(new_n343_), .A2(new_n346_), .B(new_n276_), .ZN(new_n347_));
  AOI21_X1   g0084(.A1(new_n340_), .A2(new_n347_), .B(new_n266_), .ZN(new_n348_));
  NAND2_X1   g0085(.A1(\a[111] ), .A2(\shift[0] ), .ZN(new_n349_));
  NAND2_X1   g0086(.A1(new_n268_), .A2(\a[112] ), .ZN(new_n350_));
  AOI21_X1   g0087(.A1(new_n350_), .A2(new_n349_), .B(\shift[1] ), .ZN(new_n351_));
  NAND2_X1   g0088(.A1(\a[109] ), .A2(\shift[0] ), .ZN(new_n352_));
  NAND2_X1   g0089(.A1(new_n268_), .A2(\a[110] ), .ZN(new_n353_));
  AOI21_X1   g0090(.A1(new_n353_), .A2(new_n352_), .B(new_n271_), .ZN(new_n354_));
  OAI21_X1   g0091(.A1(new_n351_), .A2(new_n354_), .B(new_n276_), .ZN(new_n355_));
  NAND2_X1   g0092(.A1(\a[103] ), .A2(\shift[0] ), .ZN(new_n356_));
  NAND2_X1   g0093(.A1(new_n268_), .A2(\a[104] ), .ZN(new_n357_));
  AOI21_X1   g0094(.A1(new_n357_), .A2(new_n356_), .B(\shift[1] ), .ZN(new_n358_));
  NAND2_X1   g0095(.A1(\a[101] ), .A2(\shift[0] ), .ZN(new_n359_));
  NAND2_X1   g0096(.A1(new_n268_), .A2(\a[102] ), .ZN(new_n360_));
  AOI21_X1   g0097(.A1(new_n360_), .A2(new_n359_), .B(new_n271_), .ZN(new_n361_));
  OAI21_X1   g0098(.A1(new_n358_), .A2(new_n361_), .B(\shift[3] ), .ZN(new_n362_));
  AOI21_X1   g0099(.A1(new_n355_), .A2(new_n362_), .B(\shift[2] ), .ZN(new_n363_));
  OAI21_X1   g0100(.A1(new_n348_), .A2(new_n363_), .B(\shift[4] ), .ZN(new_n364_));
  NAND2_X1   g0101(.A1(\a[115] ), .A2(\shift[0] ), .ZN(new_n365_));
  NAND2_X1   g0102(.A1(new_n268_), .A2(\a[116] ), .ZN(new_n366_));
  AOI21_X1   g0103(.A1(new_n366_), .A2(new_n365_), .B(\shift[1] ), .ZN(new_n367_));
  NAND2_X1   g0104(.A1(\a[113] ), .A2(\shift[0] ), .ZN(new_n368_));
  NAND2_X1   g0105(.A1(new_n268_), .A2(\a[114] ), .ZN(new_n369_));
  AOI21_X1   g0106(.A1(new_n369_), .A2(new_n368_), .B(new_n271_), .ZN(new_n370_));
  OAI21_X1   g0107(.A1(new_n367_), .A2(new_n370_), .B(\shift[3] ), .ZN(new_n371_));
  NAND2_X1   g0108(.A1(\a[123] ), .A2(\shift[0] ), .ZN(new_n372_));
  NAND2_X1   g0109(.A1(new_n268_), .A2(\a[124] ), .ZN(new_n373_));
  AOI21_X1   g0110(.A1(new_n373_), .A2(new_n372_), .B(\shift[1] ), .ZN(new_n374_));
  NAND2_X1   g0111(.A1(\a[121] ), .A2(\shift[0] ), .ZN(new_n375_));
  NAND2_X1   g0112(.A1(new_n268_), .A2(\a[122] ), .ZN(new_n376_));
  AOI21_X1   g0113(.A1(new_n376_), .A2(new_n375_), .B(new_n271_), .ZN(new_n377_));
  OAI21_X1   g0114(.A1(new_n374_), .A2(new_n377_), .B(new_n276_), .ZN(new_n378_));
  AOI21_X1   g0115(.A1(new_n371_), .A2(new_n378_), .B(new_n266_), .ZN(new_n379_));
  NAND2_X1   g0116(.A1(\a[127] ), .A2(\shift[0] ), .ZN(new_n380_));
  NAND2_X1   g0117(.A1(new_n268_), .A2(\a[0] ), .ZN(new_n381_));
  AOI21_X1   g0118(.A1(new_n381_), .A2(new_n380_), .B(\shift[1] ), .ZN(new_n382_));
  NAND2_X1   g0119(.A1(\a[125] ), .A2(\shift[0] ), .ZN(new_n383_));
  NAND2_X1   g0120(.A1(new_n268_), .A2(\a[126] ), .ZN(new_n384_));
  AOI21_X1   g0121(.A1(new_n384_), .A2(new_n383_), .B(new_n271_), .ZN(new_n385_));
  OAI21_X1   g0122(.A1(new_n382_), .A2(new_n385_), .B(new_n276_), .ZN(new_n386_));
  NAND2_X1   g0123(.A1(\a[119] ), .A2(\shift[0] ), .ZN(new_n387_));
  NAND2_X1   g0124(.A1(new_n268_), .A2(\a[120] ), .ZN(new_n388_));
  AOI21_X1   g0125(.A1(new_n388_), .A2(new_n387_), .B(\shift[1] ), .ZN(new_n389_));
  NAND2_X1   g0126(.A1(\a[117] ), .A2(\shift[0] ), .ZN(new_n390_));
  NAND2_X1   g0127(.A1(new_n268_), .A2(\a[118] ), .ZN(new_n391_));
  AOI21_X1   g0128(.A1(new_n391_), .A2(new_n390_), .B(new_n271_), .ZN(new_n392_));
  OAI21_X1   g0129(.A1(new_n389_), .A2(new_n392_), .B(\shift[3] ), .ZN(new_n393_));
  AOI21_X1   g0130(.A1(new_n386_), .A2(new_n393_), .B(\shift[2] ), .ZN(new_n394_));
  OAI21_X1   g0131(.A1(new_n379_), .A2(new_n394_), .B(new_n301_), .ZN(new_n395_));
  AOI21_X1   g0132(.A1(new_n364_), .A2(new_n395_), .B(\shift[5] ), .ZN(new_n396_));
  OAI21_X1   g0133(.A1(new_n333_), .A2(new_n396_), .B(new_n264_), .ZN(new_n397_));
  NAND2_X1   g0134(.A1(\a[3] ), .A2(\shift[0] ), .ZN(new_n398_));
  NAND2_X1   g0135(.A1(new_n268_), .A2(\a[4] ), .ZN(new_n399_));
  AOI21_X1   g0136(.A1(new_n399_), .A2(new_n398_), .B(\shift[1] ), .ZN(new_n400_));
  NAND2_X1   g0137(.A1(\a[1] ), .A2(\shift[0] ), .ZN(new_n401_));
  NAND2_X1   g0138(.A1(new_n268_), .A2(\a[2] ), .ZN(new_n402_));
  AOI21_X1   g0139(.A1(new_n402_), .A2(new_n401_), .B(new_n271_), .ZN(new_n403_));
  OAI21_X1   g0140(.A1(new_n400_), .A2(new_n403_), .B(\shift[3] ), .ZN(new_n404_));
  NAND2_X1   g0141(.A1(\a[11] ), .A2(\shift[0] ), .ZN(new_n405_));
  NAND2_X1   g0142(.A1(new_n268_), .A2(\a[12] ), .ZN(new_n406_));
  AOI21_X1   g0143(.A1(new_n406_), .A2(new_n405_), .B(\shift[1] ), .ZN(new_n407_));
  NAND2_X1   g0144(.A1(\a[9] ), .A2(\shift[0] ), .ZN(new_n408_));
  NAND2_X1   g0145(.A1(new_n268_), .A2(\a[10] ), .ZN(new_n409_));
  AOI21_X1   g0146(.A1(new_n409_), .A2(new_n408_), .B(new_n271_), .ZN(new_n410_));
  OAI21_X1   g0147(.A1(new_n407_), .A2(new_n410_), .B(new_n276_), .ZN(new_n411_));
  AOI21_X1   g0148(.A1(new_n404_), .A2(new_n411_), .B(new_n266_), .ZN(new_n412_));
  NAND2_X1   g0149(.A1(\a[15] ), .A2(\shift[0] ), .ZN(new_n413_));
  NAND2_X1   g0150(.A1(new_n268_), .A2(\a[16] ), .ZN(new_n414_));
  AOI21_X1   g0151(.A1(new_n414_), .A2(new_n413_), .B(\shift[1] ), .ZN(new_n415_));
  NAND2_X1   g0152(.A1(\a[13] ), .A2(\shift[0] ), .ZN(new_n416_));
  NAND2_X1   g0153(.A1(new_n268_), .A2(\a[14] ), .ZN(new_n417_));
  AOI21_X1   g0154(.A1(new_n417_), .A2(new_n416_), .B(new_n271_), .ZN(new_n418_));
  OAI21_X1   g0155(.A1(new_n415_), .A2(new_n418_), .B(new_n276_), .ZN(new_n419_));
  NAND2_X1   g0156(.A1(\a[7] ), .A2(\shift[0] ), .ZN(new_n420_));
  NAND2_X1   g0157(.A1(new_n268_), .A2(\a[8] ), .ZN(new_n421_));
  AOI21_X1   g0158(.A1(new_n421_), .A2(new_n420_), .B(\shift[1] ), .ZN(new_n422_));
  NAND2_X1   g0159(.A1(\a[5] ), .A2(\shift[0] ), .ZN(new_n423_));
  NAND2_X1   g0160(.A1(new_n268_), .A2(\a[6] ), .ZN(new_n424_));
  AOI21_X1   g0161(.A1(new_n424_), .A2(new_n423_), .B(new_n271_), .ZN(new_n425_));
  OAI21_X1   g0162(.A1(new_n422_), .A2(new_n425_), .B(\shift[3] ), .ZN(new_n426_));
  AOI21_X1   g0163(.A1(new_n419_), .A2(new_n426_), .B(\shift[2] ), .ZN(new_n427_));
  OAI21_X1   g0164(.A1(new_n412_), .A2(new_n427_), .B(\shift[4] ), .ZN(new_n428_));
  NAND2_X1   g0165(.A1(\a[19] ), .A2(\shift[0] ), .ZN(new_n429_));
  NAND2_X1   g0166(.A1(new_n268_), .A2(\a[20] ), .ZN(new_n430_));
  AOI21_X1   g0167(.A1(new_n430_), .A2(new_n429_), .B(\shift[1] ), .ZN(new_n431_));
  NAND2_X1   g0168(.A1(\a[17] ), .A2(\shift[0] ), .ZN(new_n432_));
  NAND2_X1   g0169(.A1(new_n268_), .A2(\a[18] ), .ZN(new_n433_));
  AOI21_X1   g0170(.A1(new_n433_), .A2(new_n432_), .B(new_n271_), .ZN(new_n434_));
  OAI21_X1   g0171(.A1(new_n431_), .A2(new_n434_), .B(\shift[3] ), .ZN(new_n435_));
  NAND2_X1   g0172(.A1(\a[27] ), .A2(\shift[0] ), .ZN(new_n436_));
  NAND2_X1   g0173(.A1(new_n268_), .A2(\a[28] ), .ZN(new_n437_));
  AOI21_X1   g0174(.A1(new_n437_), .A2(new_n436_), .B(\shift[1] ), .ZN(new_n438_));
  NAND2_X1   g0175(.A1(\a[25] ), .A2(\shift[0] ), .ZN(new_n439_));
  NAND2_X1   g0176(.A1(new_n268_), .A2(\a[26] ), .ZN(new_n440_));
  AOI21_X1   g0177(.A1(new_n440_), .A2(new_n439_), .B(new_n271_), .ZN(new_n441_));
  OAI21_X1   g0178(.A1(new_n438_), .A2(new_n441_), .B(new_n276_), .ZN(new_n442_));
  AOI21_X1   g0179(.A1(new_n435_), .A2(new_n442_), .B(new_n266_), .ZN(new_n443_));
  NAND2_X1   g0180(.A1(\a[31] ), .A2(\shift[0] ), .ZN(new_n444_));
  NAND2_X1   g0181(.A1(new_n268_), .A2(\a[32] ), .ZN(new_n445_));
  AOI21_X1   g0182(.A1(new_n445_), .A2(new_n444_), .B(\shift[1] ), .ZN(new_n446_));
  NAND2_X1   g0183(.A1(\a[29] ), .A2(\shift[0] ), .ZN(new_n447_));
  NAND2_X1   g0184(.A1(new_n268_), .A2(\a[30] ), .ZN(new_n448_));
  AOI21_X1   g0185(.A1(new_n448_), .A2(new_n447_), .B(new_n271_), .ZN(new_n449_));
  OAI21_X1   g0186(.A1(new_n446_), .A2(new_n449_), .B(new_n276_), .ZN(new_n450_));
  NAND2_X1   g0187(.A1(\a[23] ), .A2(\shift[0] ), .ZN(new_n451_));
  NAND2_X1   g0188(.A1(new_n268_), .A2(\a[24] ), .ZN(new_n452_));
  AOI21_X1   g0189(.A1(new_n452_), .A2(new_n451_), .B(\shift[1] ), .ZN(new_n453_));
  NAND2_X1   g0190(.A1(\a[21] ), .A2(\shift[0] ), .ZN(new_n454_));
  NAND2_X1   g0191(.A1(new_n268_), .A2(\a[22] ), .ZN(new_n455_));
  AOI21_X1   g0192(.A1(new_n455_), .A2(new_n454_), .B(new_n271_), .ZN(new_n456_));
  OAI21_X1   g0193(.A1(new_n453_), .A2(new_n456_), .B(\shift[3] ), .ZN(new_n457_));
  AOI21_X1   g0194(.A1(new_n450_), .A2(new_n457_), .B(\shift[2] ), .ZN(new_n458_));
  OAI21_X1   g0195(.A1(new_n443_), .A2(new_n458_), .B(new_n301_), .ZN(new_n459_));
  AOI21_X1   g0196(.A1(new_n428_), .A2(new_n459_), .B(new_n265_), .ZN(new_n460_));
  NAND2_X1   g0197(.A1(\a[35] ), .A2(\shift[0] ), .ZN(new_n461_));
  NAND2_X1   g0198(.A1(new_n268_), .A2(\a[36] ), .ZN(new_n462_));
  AOI21_X1   g0199(.A1(new_n462_), .A2(new_n461_), .B(\shift[1] ), .ZN(new_n463_));
  NAND2_X1   g0200(.A1(\a[33] ), .A2(\shift[0] ), .ZN(new_n464_));
  NAND2_X1   g0201(.A1(new_n268_), .A2(\a[34] ), .ZN(new_n465_));
  AOI21_X1   g0202(.A1(new_n465_), .A2(new_n464_), .B(new_n271_), .ZN(new_n466_));
  OAI21_X1   g0203(.A1(new_n463_), .A2(new_n466_), .B(\shift[3] ), .ZN(new_n467_));
  NAND2_X1   g0204(.A1(\a[43] ), .A2(\shift[0] ), .ZN(new_n468_));
  NAND2_X1   g0205(.A1(new_n268_), .A2(\a[44] ), .ZN(new_n469_));
  AOI21_X1   g0206(.A1(new_n469_), .A2(new_n468_), .B(\shift[1] ), .ZN(new_n470_));
  NAND2_X1   g0207(.A1(\a[41] ), .A2(\shift[0] ), .ZN(new_n471_));
  NAND2_X1   g0208(.A1(new_n268_), .A2(\a[42] ), .ZN(new_n472_));
  AOI21_X1   g0209(.A1(new_n472_), .A2(new_n471_), .B(new_n271_), .ZN(new_n473_));
  OAI21_X1   g0210(.A1(new_n470_), .A2(new_n473_), .B(new_n276_), .ZN(new_n474_));
  AOI21_X1   g0211(.A1(new_n467_), .A2(new_n474_), .B(new_n266_), .ZN(new_n475_));
  NAND2_X1   g0212(.A1(\a[47] ), .A2(\shift[0] ), .ZN(new_n476_));
  NAND2_X1   g0213(.A1(new_n268_), .A2(\a[48] ), .ZN(new_n477_));
  AOI21_X1   g0214(.A1(new_n477_), .A2(new_n476_), .B(\shift[1] ), .ZN(new_n478_));
  NAND2_X1   g0215(.A1(\a[45] ), .A2(\shift[0] ), .ZN(new_n479_));
  NAND2_X1   g0216(.A1(new_n268_), .A2(\a[46] ), .ZN(new_n480_));
  AOI21_X1   g0217(.A1(new_n480_), .A2(new_n479_), .B(new_n271_), .ZN(new_n481_));
  OAI21_X1   g0218(.A1(new_n478_), .A2(new_n481_), .B(new_n276_), .ZN(new_n482_));
  INV_X1     g0219(.I(\a[38] ), .ZN(new_n483_));
  INV_X1     g0220(.I(\a[39] ), .ZN(new_n484_));
  NAND2_X1   g0221(.A1(new_n268_), .A2(\shift[1] ), .ZN(new_n485_));
  NAND2_X1   g0222(.A1(new_n271_), .A2(\shift[0] ), .ZN(new_n486_));
  OAI22_X1   g0223(.A1(new_n483_), .A2(new_n485_), .B1(new_n486_), .B2(new_n484_), .ZN(new_n487_));
  INV_X1     g0224(.I(\a[37] ), .ZN(new_n488_));
  INV_X1     g0225(.I(\a[40] ), .ZN(new_n489_));
  OR2_X2     g0226(.A1(\shift[0] ), .A2(\shift[1] ), .Z(new_n490_));
  NAND2_X1   g0227(.A1(\shift[0] ), .A2(\shift[1] ), .ZN(new_n491_));
  OAI22_X1   g0228(.A1(new_n490_), .A2(new_n489_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1   g0229(.A1(new_n487_), .A2(new_n492_), .B(\shift[3] ), .ZN(new_n493_));
  AOI21_X1   g0230(.A1(new_n493_), .A2(new_n482_), .B(\shift[2] ), .ZN(new_n494_));
  OAI21_X1   g0231(.A1(new_n494_), .A2(new_n475_), .B(\shift[4] ), .ZN(new_n495_));
  NAND2_X1   g0232(.A1(\a[51] ), .A2(\shift[0] ), .ZN(new_n496_));
  NAND2_X1   g0233(.A1(new_n268_), .A2(\a[52] ), .ZN(new_n497_));
  AOI21_X1   g0234(.A1(new_n497_), .A2(new_n496_), .B(\shift[1] ), .ZN(new_n498_));
  NAND2_X1   g0235(.A1(\a[49] ), .A2(\shift[0] ), .ZN(new_n499_));
  NAND2_X1   g0236(.A1(new_n268_), .A2(\a[50] ), .ZN(new_n500_));
  AOI21_X1   g0237(.A1(new_n500_), .A2(new_n499_), .B(new_n271_), .ZN(new_n501_));
  OAI21_X1   g0238(.A1(new_n498_), .A2(new_n501_), .B(\shift[3] ), .ZN(new_n502_));
  NAND2_X1   g0239(.A1(\a[59] ), .A2(\shift[0] ), .ZN(new_n503_));
  NAND2_X1   g0240(.A1(new_n268_), .A2(\a[60] ), .ZN(new_n504_));
  AOI21_X1   g0241(.A1(new_n504_), .A2(new_n503_), .B(\shift[1] ), .ZN(new_n505_));
  NAND2_X1   g0242(.A1(\a[57] ), .A2(\shift[0] ), .ZN(new_n506_));
  NAND2_X1   g0243(.A1(new_n268_), .A2(\a[58] ), .ZN(new_n507_));
  AOI21_X1   g0244(.A1(new_n507_), .A2(new_n506_), .B(new_n271_), .ZN(new_n508_));
  OAI21_X1   g0245(.A1(new_n505_), .A2(new_n508_), .B(new_n276_), .ZN(new_n509_));
  AOI21_X1   g0246(.A1(new_n502_), .A2(new_n509_), .B(new_n266_), .ZN(new_n510_));
  NAND2_X1   g0247(.A1(\a[63] ), .A2(\shift[0] ), .ZN(new_n511_));
  NAND2_X1   g0248(.A1(new_n268_), .A2(\a[64] ), .ZN(new_n512_));
  AOI21_X1   g0249(.A1(new_n512_), .A2(new_n511_), .B(\shift[1] ), .ZN(new_n513_));
  NAND2_X1   g0250(.A1(\a[61] ), .A2(\shift[0] ), .ZN(new_n514_));
  NAND2_X1   g0251(.A1(new_n268_), .A2(\a[62] ), .ZN(new_n515_));
  AOI21_X1   g0252(.A1(new_n515_), .A2(new_n514_), .B(new_n271_), .ZN(new_n516_));
  OAI21_X1   g0253(.A1(new_n513_), .A2(new_n516_), .B(new_n276_), .ZN(new_n517_));
  NAND2_X1   g0254(.A1(\a[55] ), .A2(\shift[0] ), .ZN(new_n518_));
  NAND2_X1   g0255(.A1(new_n268_), .A2(\a[56] ), .ZN(new_n519_));
  AOI21_X1   g0256(.A1(new_n519_), .A2(new_n518_), .B(\shift[1] ), .ZN(new_n520_));
  NAND2_X1   g0257(.A1(\a[53] ), .A2(\shift[0] ), .ZN(new_n521_));
  NAND2_X1   g0258(.A1(new_n268_), .A2(\a[54] ), .ZN(new_n522_));
  AOI21_X1   g0259(.A1(new_n522_), .A2(new_n521_), .B(new_n271_), .ZN(new_n523_));
  OAI21_X1   g0260(.A1(new_n520_), .A2(new_n523_), .B(\shift[3] ), .ZN(new_n524_));
  AOI21_X1   g0261(.A1(new_n517_), .A2(new_n524_), .B(\shift[2] ), .ZN(new_n525_));
  OAI21_X1   g0262(.A1(new_n510_), .A2(new_n525_), .B(new_n301_), .ZN(new_n526_));
  AOI21_X1   g0263(.A1(new_n495_), .A2(new_n526_), .B(\shift[5] ), .ZN(new_n527_));
  OAI21_X1   g0264(.A1(new_n460_), .A2(new_n527_), .B(\shift[6] ), .ZN(new_n528_));
  NAND2_X1   g0265(.A1(new_n397_), .A2(new_n528_), .ZN(\result[0] ));
  INV_X1     g0266(.I(\a[67] ), .ZN(new_n530_));
  INV_X1     g0267(.I(\a[68] ), .ZN(new_n531_));
  OAI22_X1   g0268(.A1(new_n530_), .A2(new_n485_), .B1(new_n486_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1     g0269(.I(\a[66] ), .ZN(new_n533_));
  INV_X1     g0270(.I(\a[69] ), .ZN(new_n534_));
  OAI22_X1   g0271(.A1(new_n490_), .A2(new_n534_), .B1(new_n533_), .B2(new_n491_), .ZN(new_n535_));
  OAI21_X1   g0272(.A1(new_n532_), .A2(new_n535_), .B(\shift[3] ), .ZN(new_n536_));
  NAND3_X1   g0273(.A1(new_n268_), .A2(\a[75] ), .A3(\shift[1] ), .ZN(new_n537_));
  NAND3_X1   g0274(.A1(new_n271_), .A2(\a[76] ), .A3(\shift[0] ), .ZN(new_n538_));
  NAND2_X1   g0275(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1     g0276(.I(\a[74] ), .ZN(new_n540_));
  INV_X1     g0277(.I(\a[77] ), .ZN(new_n541_));
  OAI22_X1   g0278(.A1(new_n490_), .A2(new_n541_), .B1(new_n540_), .B2(new_n491_), .ZN(new_n542_));
  OAI21_X1   g0279(.A1(new_n542_), .A2(new_n539_), .B(new_n276_), .ZN(new_n543_));
  AOI21_X1   g0280(.A1(new_n536_), .A2(new_n543_), .B(new_n266_), .ZN(new_n544_));
  INV_X1     g0281(.I(\a[79] ), .ZN(new_n545_));
  INV_X1     g0282(.I(\a[80] ), .ZN(new_n546_));
  OAI22_X1   g0283(.A1(new_n545_), .A2(new_n485_), .B1(new_n486_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1     g0284(.I(\a[78] ), .ZN(new_n548_));
  INV_X1     g0285(.I(\a[81] ), .ZN(new_n549_));
  OAI22_X1   g0286(.A1(new_n490_), .A2(new_n549_), .B1(new_n548_), .B2(new_n491_), .ZN(new_n550_));
  OAI21_X1   g0287(.A1(new_n547_), .A2(new_n550_), .B(new_n276_), .ZN(new_n551_));
  INV_X1     g0288(.I(\a[71] ), .ZN(new_n552_));
  INV_X1     g0289(.I(\a[72] ), .ZN(new_n553_));
  OAI22_X1   g0290(.A1(new_n552_), .A2(new_n485_), .B1(new_n486_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1     g0291(.I(\a[70] ), .ZN(new_n555_));
  INV_X1     g0292(.I(\a[73] ), .ZN(new_n556_));
  OAI22_X1   g0293(.A1(new_n490_), .A2(new_n556_), .B1(new_n555_), .B2(new_n491_), .ZN(new_n557_));
  OAI21_X1   g0294(.A1(new_n554_), .A2(new_n557_), .B(\shift[3] ), .ZN(new_n558_));
  AOI21_X1   g0295(.A1(new_n551_), .A2(new_n558_), .B(\shift[2] ), .ZN(new_n559_));
  OAI21_X1   g0296(.A1(new_n559_), .A2(new_n544_), .B(\shift[4] ), .ZN(new_n560_));
  INV_X1     g0297(.I(\a[83] ), .ZN(new_n561_));
  INV_X1     g0298(.I(\a[84] ), .ZN(new_n562_));
  OAI22_X1   g0299(.A1(new_n561_), .A2(new_n485_), .B1(new_n486_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1     g0300(.I(\a[82] ), .ZN(new_n564_));
  INV_X1     g0301(.I(\a[85] ), .ZN(new_n565_));
  OAI22_X1   g0302(.A1(new_n490_), .A2(new_n565_), .B1(new_n564_), .B2(new_n491_), .ZN(new_n566_));
  OAI21_X1   g0303(.A1(new_n563_), .A2(new_n566_), .B(\shift[3] ), .ZN(new_n567_));
  NAND3_X1   g0304(.A1(new_n268_), .A2(\a[91] ), .A3(\shift[1] ), .ZN(new_n568_));
  NAND3_X1   g0305(.A1(new_n271_), .A2(\a[92] ), .A3(\shift[0] ), .ZN(new_n569_));
  NAND2_X1   g0306(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1     g0307(.I(\a[90] ), .ZN(new_n571_));
  INV_X1     g0308(.I(\a[93] ), .ZN(new_n572_));
  OAI22_X1   g0309(.A1(new_n490_), .A2(new_n572_), .B1(new_n571_), .B2(new_n491_), .ZN(new_n573_));
  OAI21_X1   g0310(.A1(new_n573_), .A2(new_n570_), .B(new_n276_), .ZN(new_n574_));
  AOI21_X1   g0311(.A1(new_n567_), .A2(new_n574_), .B(new_n266_), .ZN(new_n575_));
  NAND3_X1   g0312(.A1(new_n268_), .A2(\a[95] ), .A3(\shift[1] ), .ZN(new_n576_));
  NAND3_X1   g0313(.A1(new_n271_), .A2(\a[96] ), .A3(\shift[0] ), .ZN(new_n577_));
  NAND2_X1   g0314(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1     g0315(.I(\a[94] ), .ZN(new_n579_));
  INV_X1     g0316(.I(\a[97] ), .ZN(new_n580_));
  OAI22_X1   g0317(.A1(new_n490_), .A2(new_n580_), .B1(new_n579_), .B2(new_n491_), .ZN(new_n581_));
  OAI21_X1   g0318(.A1(new_n581_), .A2(new_n578_), .B(new_n276_), .ZN(new_n582_));
  INV_X1     g0319(.I(\a[87] ), .ZN(new_n583_));
  INV_X1     g0320(.I(\a[88] ), .ZN(new_n584_));
  OAI22_X1   g0321(.A1(new_n583_), .A2(new_n485_), .B1(new_n486_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1     g0322(.I(\a[86] ), .ZN(new_n586_));
  INV_X1     g0323(.I(\a[89] ), .ZN(new_n587_));
  OAI22_X1   g0324(.A1(new_n490_), .A2(new_n587_), .B1(new_n586_), .B2(new_n491_), .ZN(new_n588_));
  OAI21_X1   g0325(.A1(new_n585_), .A2(new_n588_), .B(\shift[3] ), .ZN(new_n589_));
  AOI21_X1   g0326(.A1(new_n589_), .A2(new_n582_), .B(\shift[2] ), .ZN(new_n590_));
  OAI21_X1   g0327(.A1(new_n575_), .A2(new_n590_), .B(new_n301_), .ZN(new_n591_));
  AOI21_X1   g0328(.A1(new_n560_), .A2(new_n591_), .B(new_n265_), .ZN(new_n592_));
  INV_X1     g0329(.I(\a[99] ), .ZN(new_n593_));
  INV_X1     g0330(.I(\a[100] ), .ZN(new_n594_));
  OAI22_X1   g0331(.A1(new_n593_), .A2(new_n485_), .B1(new_n486_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1     g0332(.I(\a[98] ), .ZN(new_n596_));
  INV_X1     g0333(.I(\a[101] ), .ZN(new_n597_));
  OAI22_X1   g0334(.A1(new_n490_), .A2(new_n597_), .B1(new_n596_), .B2(new_n491_), .ZN(new_n598_));
  OAI21_X1   g0335(.A1(new_n595_), .A2(new_n598_), .B(\shift[3] ), .ZN(new_n599_));
  INV_X1     g0336(.I(\a[107] ), .ZN(new_n600_));
  INV_X1     g0337(.I(\a[108] ), .ZN(new_n601_));
  OAI22_X1   g0338(.A1(new_n600_), .A2(new_n485_), .B1(new_n486_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1     g0339(.I(\a[106] ), .ZN(new_n603_));
  INV_X1     g0340(.I(\a[109] ), .ZN(new_n604_));
  OAI22_X1   g0341(.A1(new_n490_), .A2(new_n604_), .B1(new_n603_), .B2(new_n491_), .ZN(new_n605_));
  OAI21_X1   g0342(.A1(new_n602_), .A2(new_n605_), .B(new_n276_), .ZN(new_n606_));
  AOI21_X1   g0343(.A1(new_n599_), .A2(new_n606_), .B(new_n266_), .ZN(new_n607_));
  NAND3_X1   g0344(.A1(new_n268_), .A2(\a[111] ), .A3(\shift[1] ), .ZN(new_n608_));
  NAND3_X1   g0345(.A1(new_n271_), .A2(\a[112] ), .A3(\shift[0] ), .ZN(new_n609_));
  NAND2_X1   g0346(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1     g0347(.I(\a[110] ), .ZN(new_n611_));
  INV_X1     g0348(.I(\a[113] ), .ZN(new_n612_));
  OAI22_X1   g0349(.A1(new_n490_), .A2(new_n612_), .B1(new_n611_), .B2(new_n491_), .ZN(new_n613_));
  OAI21_X1   g0350(.A1(new_n613_), .A2(new_n610_), .B(new_n276_), .ZN(new_n614_));
  NAND3_X1   g0351(.A1(new_n268_), .A2(\a[103] ), .A3(\shift[1] ), .ZN(new_n615_));
  NAND3_X1   g0352(.A1(new_n271_), .A2(\a[104] ), .A3(\shift[0] ), .ZN(new_n616_));
  NAND2_X1   g0353(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1     g0354(.I(\a[105] ), .ZN(new_n618_));
  NAND3_X1   g0355(.A1(\a[102] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n619_));
  OAI21_X1   g0356(.A1(new_n490_), .A2(new_n618_), .B(new_n619_), .ZN(new_n620_));
  OAI21_X1   g0357(.A1(new_n617_), .A2(new_n620_), .B(\shift[3] ), .ZN(new_n621_));
  AOI21_X1   g0358(.A1(new_n614_), .A2(new_n621_), .B(\shift[2] ), .ZN(new_n622_));
  OAI21_X1   g0359(.A1(new_n607_), .A2(new_n622_), .B(\shift[4] ), .ZN(new_n623_));
  INV_X1     g0360(.I(\a[115] ), .ZN(new_n624_));
  INV_X1     g0361(.I(\a[116] ), .ZN(new_n625_));
  OAI22_X1   g0362(.A1(new_n624_), .A2(new_n485_), .B1(new_n486_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1     g0363(.I(\a[114] ), .ZN(new_n627_));
  INV_X1     g0364(.I(\a[117] ), .ZN(new_n628_));
  OAI22_X1   g0365(.A1(new_n490_), .A2(new_n628_), .B1(new_n627_), .B2(new_n491_), .ZN(new_n629_));
  OAI21_X1   g0366(.A1(new_n626_), .A2(new_n629_), .B(\shift[3] ), .ZN(new_n630_));
  INV_X1     g0367(.I(\a[123] ), .ZN(new_n631_));
  INV_X1     g0368(.I(\a[124] ), .ZN(new_n632_));
  OAI22_X1   g0369(.A1(new_n631_), .A2(new_n485_), .B1(new_n486_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1     g0370(.I(\a[122] ), .ZN(new_n634_));
  INV_X1     g0371(.I(\a[125] ), .ZN(new_n635_));
  OAI22_X1   g0372(.A1(new_n490_), .A2(new_n635_), .B1(new_n634_), .B2(new_n491_), .ZN(new_n636_));
  OAI21_X1   g0373(.A1(new_n633_), .A2(new_n636_), .B(new_n276_), .ZN(new_n637_));
  AOI21_X1   g0374(.A1(new_n630_), .A2(new_n637_), .B(new_n266_), .ZN(new_n638_));
  NAND3_X1   g0375(.A1(new_n271_), .A2(\a[0] ), .A3(\shift[0] ), .ZN(new_n639_));
  NAND3_X1   g0376(.A1(new_n268_), .A2(\a[127] ), .A3(\shift[1] ), .ZN(new_n640_));
  NAND2_X1   g0377(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1     g0378(.I(\a[1] ), .ZN(new_n642_));
  INV_X1     g0379(.I(\a[126] ), .ZN(new_n643_));
  OAI22_X1   g0380(.A1(new_n490_), .A2(new_n642_), .B1(new_n643_), .B2(new_n491_), .ZN(new_n644_));
  OAI21_X1   g0381(.A1(new_n644_), .A2(new_n641_), .B(new_n276_), .ZN(new_n645_));
  NAND3_X1   g0382(.A1(new_n268_), .A2(\a[119] ), .A3(\shift[1] ), .ZN(new_n646_));
  NAND3_X1   g0383(.A1(new_n271_), .A2(\a[120] ), .A3(\shift[0] ), .ZN(new_n647_));
  NAND2_X1   g0384(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1     g0385(.I(\a[121] ), .ZN(new_n649_));
  NAND3_X1   g0386(.A1(\a[118] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n650_));
  OAI21_X1   g0387(.A1(new_n490_), .A2(new_n649_), .B(new_n650_), .ZN(new_n651_));
  OAI21_X1   g0388(.A1(new_n648_), .A2(new_n651_), .B(\shift[3] ), .ZN(new_n652_));
  AOI21_X1   g0389(.A1(new_n645_), .A2(new_n652_), .B(\shift[2] ), .ZN(new_n653_));
  OAI21_X1   g0390(.A1(new_n638_), .A2(new_n653_), .B(new_n301_), .ZN(new_n654_));
  AOI21_X1   g0391(.A1(new_n623_), .A2(new_n654_), .B(\shift[5] ), .ZN(new_n655_));
  OAI21_X1   g0392(.A1(new_n592_), .A2(new_n655_), .B(new_n264_), .ZN(new_n656_));
  NOR2_X1    g0393(.A1(\shift[4] ), .A2(\shift[5] ), .ZN(new_n657_));
  NAND3_X1   g0394(.A1(new_n268_), .A2(\a[51] ), .A3(\shift[1] ), .ZN(new_n658_));
  NAND3_X1   g0395(.A1(new_n271_), .A2(\a[52] ), .A3(\shift[0] ), .ZN(new_n659_));
  NAND2_X1   g0396(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1     g0397(.I(\a[50] ), .ZN(new_n661_));
  INV_X1     g0398(.I(\a[53] ), .ZN(new_n662_));
  OAI22_X1   g0399(.A1(new_n490_), .A2(new_n662_), .B1(new_n661_), .B2(new_n491_), .ZN(new_n663_));
  OAI21_X1   g0400(.A1(new_n663_), .A2(new_n660_), .B(\shift[3] ), .ZN(new_n664_));
  NAND3_X1   g0401(.A1(new_n268_), .A2(\a[59] ), .A3(\shift[1] ), .ZN(new_n665_));
  NAND3_X1   g0402(.A1(new_n271_), .A2(\a[60] ), .A3(\shift[0] ), .ZN(new_n666_));
  NAND2_X1   g0403(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1     g0404(.I(\a[58] ), .ZN(new_n668_));
  INV_X1     g0405(.I(\a[61] ), .ZN(new_n669_));
  OAI22_X1   g0406(.A1(new_n490_), .A2(new_n669_), .B1(new_n668_), .B2(new_n491_), .ZN(new_n670_));
  OAI21_X1   g0407(.A1(new_n670_), .A2(new_n667_), .B(new_n276_), .ZN(new_n671_));
  AOI21_X1   g0408(.A1(new_n664_), .A2(new_n671_), .B(new_n266_), .ZN(new_n672_));
  NAND3_X1   g0409(.A1(new_n268_), .A2(\a[63] ), .A3(\shift[1] ), .ZN(new_n673_));
  NAND3_X1   g0410(.A1(new_n271_), .A2(\a[64] ), .A3(\shift[0] ), .ZN(new_n674_));
  NAND2_X1   g0411(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1     g0412(.I(\a[62] ), .ZN(new_n676_));
  INV_X1     g0413(.I(\a[65] ), .ZN(new_n677_));
  OAI22_X1   g0414(.A1(new_n490_), .A2(new_n677_), .B1(new_n676_), .B2(new_n491_), .ZN(new_n678_));
  OAI21_X1   g0415(.A1(new_n678_), .A2(new_n675_), .B(new_n276_), .ZN(new_n679_));
  INV_X1     g0416(.I(\a[55] ), .ZN(new_n680_));
  INV_X1     g0417(.I(\a[56] ), .ZN(new_n681_));
  OAI22_X1   g0418(.A1(new_n680_), .A2(new_n485_), .B1(new_n486_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1     g0419(.I(\a[54] ), .ZN(new_n683_));
  INV_X1     g0420(.I(\a[57] ), .ZN(new_n684_));
  OAI22_X1   g0421(.A1(new_n490_), .A2(new_n684_), .B1(new_n683_), .B2(new_n491_), .ZN(new_n685_));
  OAI21_X1   g0422(.A1(new_n682_), .A2(new_n685_), .B(\shift[3] ), .ZN(new_n686_));
  AOI21_X1   g0423(.A1(new_n686_), .A2(new_n679_), .B(\shift[2] ), .ZN(new_n687_));
  OAI21_X1   g0424(.A1(new_n687_), .A2(new_n672_), .B(new_n657_), .ZN(new_n688_));
  NOR2_X1    g0425(.A1(new_n301_), .A2(new_n265_), .ZN(new_n689_));
  INV_X1     g0426(.I(\a[3] ), .ZN(new_n690_));
  INV_X1     g0427(.I(\a[4] ), .ZN(new_n691_));
  OAI22_X1   g0428(.A1(new_n690_), .A2(new_n485_), .B1(new_n486_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1     g0429(.I(\a[2] ), .ZN(new_n693_));
  INV_X1     g0430(.I(\a[5] ), .ZN(new_n694_));
  OAI22_X1   g0431(.A1(new_n490_), .A2(new_n694_), .B1(new_n693_), .B2(new_n491_), .ZN(new_n695_));
  OAI21_X1   g0432(.A1(new_n692_), .A2(new_n695_), .B(\shift[3] ), .ZN(new_n696_));
  INV_X1     g0433(.I(\a[11] ), .ZN(new_n697_));
  INV_X1     g0434(.I(\a[12] ), .ZN(new_n698_));
  OAI22_X1   g0435(.A1(new_n697_), .A2(new_n485_), .B1(new_n486_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1     g0436(.I(\a[10] ), .ZN(new_n700_));
  INV_X1     g0437(.I(\a[13] ), .ZN(new_n701_));
  OAI22_X1   g0438(.A1(new_n490_), .A2(new_n701_), .B1(new_n700_), .B2(new_n491_), .ZN(new_n702_));
  OAI21_X1   g0439(.A1(new_n699_), .A2(new_n702_), .B(new_n276_), .ZN(new_n703_));
  AOI21_X1   g0440(.A1(new_n696_), .A2(new_n703_), .B(new_n266_), .ZN(new_n704_));
  NAND3_X1   g0441(.A1(new_n268_), .A2(\a[15] ), .A3(\shift[1] ), .ZN(new_n705_));
  NAND3_X1   g0442(.A1(new_n271_), .A2(\a[16] ), .A3(\shift[0] ), .ZN(new_n706_));
  NAND2_X1   g0443(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1     g0444(.I(\a[14] ), .ZN(new_n708_));
  INV_X1     g0445(.I(\a[17] ), .ZN(new_n709_));
  OAI22_X1   g0446(.A1(new_n490_), .A2(new_n709_), .B1(new_n708_), .B2(new_n491_), .ZN(new_n710_));
  OAI21_X1   g0447(.A1(new_n710_), .A2(new_n707_), .B(new_n276_), .ZN(new_n711_));
  NAND3_X1   g0448(.A1(new_n268_), .A2(\a[7] ), .A3(\shift[1] ), .ZN(new_n712_));
  NAND3_X1   g0449(.A1(new_n271_), .A2(\a[8] ), .A3(\shift[0] ), .ZN(new_n713_));
  NAND2_X1   g0450(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1     g0451(.I(\a[6] ), .ZN(new_n715_));
  INV_X1     g0452(.I(\a[9] ), .ZN(new_n716_));
  OAI22_X1   g0453(.A1(new_n490_), .A2(new_n716_), .B1(new_n715_), .B2(new_n491_), .ZN(new_n717_));
  OAI21_X1   g0454(.A1(new_n717_), .A2(new_n714_), .B(\shift[3] ), .ZN(new_n718_));
  AOI21_X1   g0455(.A1(new_n711_), .A2(new_n718_), .B(\shift[2] ), .ZN(new_n719_));
  OAI21_X1   g0456(.A1(new_n704_), .A2(new_n719_), .B(new_n689_), .ZN(new_n720_));
  NAND2_X1   g0457(.A1(new_n688_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1    g0458(.A1(new_n301_), .A2(\shift[5] ), .ZN(new_n722_));
  NAND3_X1   g0459(.A1(new_n268_), .A2(\a[35] ), .A3(\shift[1] ), .ZN(new_n723_));
  NAND3_X1   g0460(.A1(new_n271_), .A2(\a[36] ), .A3(\shift[0] ), .ZN(new_n724_));
  NAND2_X1   g0461(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1   g0462(.A1(\a[34] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n726_));
  OAI21_X1   g0463(.A1(new_n490_), .A2(new_n488_), .B(new_n726_), .ZN(new_n727_));
  OAI21_X1   g0464(.A1(new_n725_), .A2(new_n727_), .B(\shift[3] ), .ZN(new_n728_));
  NAND2_X1   g0465(.A1(\a[44] ), .A2(\shift[0] ), .ZN(new_n729_));
  NAND2_X1   g0466(.A1(new_n268_), .A2(\a[45] ), .ZN(new_n730_));
  AOI21_X1   g0467(.A1(new_n730_), .A2(new_n729_), .B(\shift[1] ), .ZN(new_n731_));
  NAND2_X1   g0468(.A1(\a[42] ), .A2(\shift[0] ), .ZN(new_n732_));
  NAND2_X1   g0469(.A1(new_n268_), .A2(\a[43] ), .ZN(new_n733_));
  AOI21_X1   g0470(.A1(new_n733_), .A2(new_n732_), .B(new_n271_), .ZN(new_n734_));
  OAI21_X1   g0471(.A1(new_n731_), .A2(new_n734_), .B(new_n276_), .ZN(new_n735_));
  AOI21_X1   g0472(.A1(new_n728_), .A2(new_n735_), .B(new_n266_), .ZN(new_n736_));
  NAND3_X1   g0473(.A1(new_n268_), .A2(\a[47] ), .A3(\shift[1] ), .ZN(new_n737_));
  NAND3_X1   g0474(.A1(new_n271_), .A2(\a[48] ), .A3(\shift[0] ), .ZN(new_n738_));
  NAND2_X1   g0475(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1     g0476(.I(\a[46] ), .ZN(new_n740_));
  INV_X1     g0477(.I(\a[49] ), .ZN(new_n741_));
  OAI22_X1   g0478(.A1(new_n490_), .A2(new_n741_), .B1(new_n740_), .B2(new_n491_), .ZN(new_n742_));
  OAI21_X1   g0479(.A1(new_n742_), .A2(new_n739_), .B(new_n276_), .ZN(new_n743_));
  NAND2_X1   g0480(.A1(\a[38] ), .A2(\shift[0] ), .ZN(new_n744_));
  NAND2_X1   g0481(.A1(new_n268_), .A2(\a[39] ), .ZN(new_n745_));
  AOI21_X1   g0482(.A1(new_n745_), .A2(new_n744_), .B(new_n271_), .ZN(new_n746_));
  NAND2_X1   g0483(.A1(\a[40] ), .A2(\shift[0] ), .ZN(new_n747_));
  NAND2_X1   g0484(.A1(new_n268_), .A2(\a[41] ), .ZN(new_n748_));
  AOI21_X1   g0485(.A1(new_n748_), .A2(new_n747_), .B(\shift[1] ), .ZN(new_n749_));
  OAI21_X1   g0486(.A1(new_n746_), .A2(new_n749_), .B(\shift[3] ), .ZN(new_n750_));
  AOI21_X1   g0487(.A1(new_n743_), .A2(new_n750_), .B(\shift[2] ), .ZN(new_n751_));
  OAI21_X1   g0488(.A1(new_n736_), .A2(new_n751_), .B(new_n722_), .ZN(new_n752_));
  NOR2_X1    g0489(.A1(new_n265_), .A2(\shift[4] ), .ZN(new_n753_));
  INV_X1     g0490(.I(\a[19] ), .ZN(new_n754_));
  INV_X1     g0491(.I(\a[20] ), .ZN(new_n755_));
  OAI22_X1   g0492(.A1(new_n754_), .A2(new_n485_), .B1(new_n486_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1     g0493(.I(\a[18] ), .ZN(new_n757_));
  INV_X1     g0494(.I(\a[21] ), .ZN(new_n758_));
  OAI22_X1   g0495(.A1(new_n490_), .A2(new_n758_), .B1(new_n757_), .B2(new_n491_), .ZN(new_n759_));
  OAI21_X1   g0496(.A1(new_n756_), .A2(new_n759_), .B(\shift[3] ), .ZN(new_n760_));
  NAND3_X1   g0497(.A1(new_n268_), .A2(\a[27] ), .A3(\shift[1] ), .ZN(new_n761_));
  NAND3_X1   g0498(.A1(new_n271_), .A2(\a[28] ), .A3(\shift[0] ), .ZN(new_n762_));
  NAND2_X1   g0499(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1     g0500(.I(\a[26] ), .ZN(new_n764_));
  INV_X1     g0501(.I(\a[29] ), .ZN(new_n765_));
  OAI22_X1   g0502(.A1(new_n490_), .A2(new_n765_), .B1(new_n764_), .B2(new_n491_), .ZN(new_n766_));
  OAI21_X1   g0503(.A1(new_n766_), .A2(new_n763_), .B(new_n276_), .ZN(new_n767_));
  AOI21_X1   g0504(.A1(new_n760_), .A2(new_n767_), .B(new_n266_), .ZN(new_n768_));
  NAND3_X1   g0505(.A1(new_n268_), .A2(\a[31] ), .A3(\shift[1] ), .ZN(new_n769_));
  NAND3_X1   g0506(.A1(new_n271_), .A2(\a[32] ), .A3(\shift[0] ), .ZN(new_n770_));
  NAND2_X1   g0507(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1     g0508(.I(\a[30] ), .ZN(new_n772_));
  INV_X1     g0509(.I(\a[33] ), .ZN(new_n773_));
  OAI22_X1   g0510(.A1(new_n490_), .A2(new_n773_), .B1(new_n772_), .B2(new_n491_), .ZN(new_n774_));
  OAI21_X1   g0511(.A1(new_n774_), .A2(new_n771_), .B(new_n276_), .ZN(new_n775_));
  NAND3_X1   g0512(.A1(new_n268_), .A2(\a[23] ), .A3(\shift[1] ), .ZN(new_n776_));
  NAND3_X1   g0513(.A1(new_n271_), .A2(\a[24] ), .A3(\shift[0] ), .ZN(new_n777_));
  NAND2_X1   g0514(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1     g0515(.I(\a[22] ), .ZN(new_n779_));
  INV_X1     g0516(.I(\a[25] ), .ZN(new_n780_));
  OAI22_X1   g0517(.A1(new_n490_), .A2(new_n780_), .B1(new_n779_), .B2(new_n491_), .ZN(new_n781_));
  OAI21_X1   g0518(.A1(new_n781_), .A2(new_n778_), .B(\shift[3] ), .ZN(new_n782_));
  AOI21_X1   g0519(.A1(new_n775_), .A2(new_n782_), .B(\shift[2] ), .ZN(new_n783_));
  OAI21_X1   g0520(.A1(new_n768_), .A2(new_n783_), .B(new_n753_), .ZN(new_n784_));
  NAND2_X1   g0521(.A1(new_n784_), .A2(new_n752_), .ZN(new_n785_));
  OAI21_X1   g0522(.A1(new_n721_), .A2(new_n785_), .B(\shift[6] ), .ZN(new_n786_));
  NAND2_X1   g0523(.A1(new_n656_), .A2(new_n786_), .ZN(\result[1] ));
  AOI21_X1   g0524(.A1(new_n269_), .A2(new_n267_), .B(new_n271_), .ZN(new_n788_));
  AOI21_X1   g0525(.A1(new_n296_), .A2(new_n295_), .B(\shift[1] ), .ZN(new_n789_));
  OAI21_X1   g0526(.A1(new_n788_), .A2(new_n789_), .B(\shift[3] ), .ZN(new_n790_));
  AOI21_X1   g0527(.A1(new_n278_), .A2(new_n277_), .B(new_n271_), .ZN(new_n791_));
  AOI21_X1   g0528(.A1(new_n289_), .A2(new_n288_), .B(\shift[1] ), .ZN(new_n792_));
  OAI21_X1   g0529(.A1(new_n791_), .A2(new_n792_), .B(new_n276_), .ZN(new_n793_));
  AOI21_X1   g0530(.A1(new_n790_), .A2(new_n793_), .B(new_n266_), .ZN(new_n794_));
  AOI21_X1   g0531(.A1(new_n286_), .A2(new_n285_), .B(new_n271_), .ZN(new_n795_));
  AOI21_X1   g0532(.A1(new_n306_), .A2(new_n305_), .B(\shift[1] ), .ZN(new_n796_));
  OAI21_X1   g0533(.A1(new_n795_), .A2(new_n796_), .B(new_n276_), .ZN(new_n797_));
  AOI21_X1   g0534(.A1(new_n293_), .A2(new_n292_), .B(new_n271_), .ZN(new_n798_));
  AOI21_X1   g0535(.A1(new_n281_), .A2(new_n280_), .B(\shift[1] ), .ZN(new_n799_));
  OAI21_X1   g0536(.A1(new_n798_), .A2(new_n799_), .B(\shift[3] ), .ZN(new_n800_));
  AOI21_X1   g0537(.A1(new_n797_), .A2(new_n800_), .B(\shift[2] ), .ZN(new_n801_));
  OAI21_X1   g0538(.A1(new_n794_), .A2(new_n801_), .B(\shift[4] ), .ZN(new_n802_));
  AOI21_X1   g0539(.A1(new_n303_), .A2(new_n302_), .B(new_n271_), .ZN(new_n803_));
  AOI21_X1   g0540(.A1(new_n328_), .A2(new_n327_), .B(\shift[1] ), .ZN(new_n804_));
  OAI21_X1   g0541(.A1(new_n803_), .A2(new_n804_), .B(\shift[3] ), .ZN(new_n805_));
  AOI21_X1   g0542(.A1(new_n310_), .A2(new_n309_), .B(new_n271_), .ZN(new_n806_));
  AOI21_X1   g0543(.A1(new_n321_), .A2(new_n320_), .B(\shift[1] ), .ZN(new_n807_));
  OAI21_X1   g0544(.A1(new_n806_), .A2(new_n807_), .B(new_n276_), .ZN(new_n808_));
  AOI21_X1   g0545(.A1(new_n805_), .A2(new_n808_), .B(new_n266_), .ZN(new_n809_));
  AOI21_X1   g0546(.A1(new_n318_), .A2(new_n317_), .B(new_n271_), .ZN(new_n810_));
  AOI21_X1   g0547(.A1(new_n338_), .A2(new_n337_), .B(\shift[1] ), .ZN(new_n811_));
  OAI21_X1   g0548(.A1(new_n810_), .A2(new_n811_), .B(new_n276_), .ZN(new_n812_));
  AOI21_X1   g0549(.A1(new_n325_), .A2(new_n324_), .B(new_n271_), .ZN(new_n813_));
  AOI21_X1   g0550(.A1(new_n313_), .A2(new_n312_), .B(\shift[1] ), .ZN(new_n814_));
  OAI21_X1   g0551(.A1(new_n813_), .A2(new_n814_), .B(\shift[3] ), .ZN(new_n815_));
  AOI21_X1   g0552(.A1(new_n812_), .A2(new_n815_), .B(\shift[2] ), .ZN(new_n816_));
  OAI21_X1   g0553(.A1(new_n809_), .A2(new_n816_), .B(new_n301_), .ZN(new_n817_));
  AOI21_X1   g0554(.A1(new_n802_), .A2(new_n817_), .B(new_n265_), .ZN(new_n818_));
  AOI21_X1   g0555(.A1(new_n335_), .A2(new_n334_), .B(new_n271_), .ZN(new_n819_));
  AOI21_X1   g0556(.A1(new_n360_), .A2(new_n359_), .B(\shift[1] ), .ZN(new_n820_));
  OAI21_X1   g0557(.A1(new_n819_), .A2(new_n820_), .B(\shift[3] ), .ZN(new_n821_));
  AOI21_X1   g0558(.A1(new_n342_), .A2(new_n341_), .B(new_n271_), .ZN(new_n822_));
  AOI21_X1   g0559(.A1(new_n353_), .A2(new_n352_), .B(\shift[1] ), .ZN(new_n823_));
  OAI21_X1   g0560(.A1(new_n822_), .A2(new_n823_), .B(new_n276_), .ZN(new_n824_));
  AOI21_X1   g0561(.A1(new_n821_), .A2(new_n824_), .B(new_n266_), .ZN(new_n825_));
  AOI21_X1   g0562(.A1(new_n350_), .A2(new_n349_), .B(new_n271_), .ZN(new_n826_));
  AOI21_X1   g0563(.A1(new_n369_), .A2(new_n368_), .B(\shift[1] ), .ZN(new_n827_));
  OAI21_X1   g0564(.A1(new_n826_), .A2(new_n827_), .B(new_n276_), .ZN(new_n828_));
  AOI21_X1   g0565(.A1(new_n357_), .A2(new_n356_), .B(new_n271_), .ZN(new_n829_));
  AOI21_X1   g0566(.A1(new_n345_), .A2(new_n344_), .B(\shift[1] ), .ZN(new_n830_));
  OAI21_X1   g0567(.A1(new_n829_), .A2(new_n830_), .B(\shift[3] ), .ZN(new_n831_));
  AOI21_X1   g0568(.A1(new_n828_), .A2(new_n831_), .B(\shift[2] ), .ZN(new_n832_));
  OAI21_X1   g0569(.A1(new_n825_), .A2(new_n832_), .B(\shift[4] ), .ZN(new_n833_));
  AOI21_X1   g0570(.A1(new_n366_), .A2(new_n365_), .B(new_n271_), .ZN(new_n834_));
  AOI21_X1   g0571(.A1(new_n391_), .A2(new_n390_), .B(\shift[1] ), .ZN(new_n835_));
  OAI21_X1   g0572(.A1(new_n834_), .A2(new_n835_), .B(\shift[3] ), .ZN(new_n836_));
  AOI21_X1   g0573(.A1(new_n373_), .A2(new_n372_), .B(new_n271_), .ZN(new_n837_));
  AOI21_X1   g0574(.A1(new_n384_), .A2(new_n383_), .B(\shift[1] ), .ZN(new_n838_));
  OAI21_X1   g0575(.A1(new_n837_), .A2(new_n838_), .B(new_n276_), .ZN(new_n839_));
  AOI21_X1   g0576(.A1(new_n836_), .A2(new_n839_), .B(new_n266_), .ZN(new_n840_));
  AOI21_X1   g0577(.A1(new_n381_), .A2(new_n380_), .B(new_n271_), .ZN(new_n841_));
  AOI21_X1   g0578(.A1(new_n402_), .A2(new_n401_), .B(\shift[1] ), .ZN(new_n842_));
  OAI21_X1   g0579(.A1(new_n841_), .A2(new_n842_), .B(new_n276_), .ZN(new_n843_));
  AOI21_X1   g0580(.A1(new_n388_), .A2(new_n387_), .B(new_n271_), .ZN(new_n844_));
  AOI21_X1   g0581(.A1(new_n376_), .A2(new_n375_), .B(\shift[1] ), .ZN(new_n845_));
  OAI21_X1   g0582(.A1(new_n844_), .A2(new_n845_), .B(\shift[3] ), .ZN(new_n846_));
  AOI21_X1   g0583(.A1(new_n843_), .A2(new_n846_), .B(\shift[2] ), .ZN(new_n847_));
  OAI21_X1   g0584(.A1(new_n840_), .A2(new_n847_), .B(new_n301_), .ZN(new_n848_));
  AOI21_X1   g0585(.A1(new_n833_), .A2(new_n848_), .B(\shift[5] ), .ZN(new_n849_));
  OAI21_X1   g0586(.A1(new_n818_), .A2(new_n849_), .B(new_n264_), .ZN(new_n850_));
  INV_X1     g0587(.I(new_n657_), .ZN(new_n851_));
  INV_X1     g0588(.I(new_n689_), .ZN(new_n852_));
  AOI21_X1   g0589(.A1(new_n497_), .A2(new_n496_), .B(new_n271_), .ZN(new_n853_));
  AOI21_X1   g0590(.A1(new_n522_), .A2(new_n521_), .B(\shift[1] ), .ZN(new_n854_));
  OAI21_X1   g0591(.A1(new_n853_), .A2(new_n854_), .B(\shift[3] ), .ZN(new_n855_));
  AOI21_X1   g0592(.A1(new_n504_), .A2(new_n503_), .B(new_n271_), .ZN(new_n856_));
  AOI21_X1   g0593(.A1(new_n515_), .A2(new_n514_), .B(\shift[1] ), .ZN(new_n857_));
  OAI21_X1   g0594(.A1(new_n856_), .A2(new_n857_), .B(new_n276_), .ZN(new_n858_));
  AOI21_X1   g0595(.A1(new_n855_), .A2(new_n858_), .B(new_n266_), .ZN(new_n859_));
  AOI21_X1   g0596(.A1(new_n512_), .A2(new_n511_), .B(new_n271_), .ZN(new_n860_));
  AOI21_X1   g0597(.A1(new_n273_), .A2(new_n272_), .B(\shift[1] ), .ZN(new_n861_));
  OAI21_X1   g0598(.A1(new_n860_), .A2(new_n861_), .B(new_n276_), .ZN(new_n862_));
  AOI21_X1   g0599(.A1(new_n519_), .A2(new_n518_), .B(new_n271_), .ZN(new_n863_));
  AOI21_X1   g0600(.A1(new_n507_), .A2(new_n506_), .B(\shift[1] ), .ZN(new_n864_));
  OAI21_X1   g0601(.A1(new_n863_), .A2(new_n864_), .B(\shift[3] ), .ZN(new_n865_));
  AOI21_X1   g0602(.A1(new_n862_), .A2(new_n865_), .B(\shift[2] ), .ZN(new_n866_));
  NOR2_X1    g0603(.A1(new_n859_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1   g0604(.A1(new_n399_), .A2(new_n398_), .B(new_n271_), .ZN(new_n868_));
  AOI21_X1   g0605(.A1(new_n424_), .A2(new_n423_), .B(\shift[1] ), .ZN(new_n869_));
  OAI21_X1   g0606(.A1(new_n868_), .A2(new_n869_), .B(\shift[3] ), .ZN(new_n870_));
  AOI21_X1   g0607(.A1(new_n406_), .A2(new_n405_), .B(new_n271_), .ZN(new_n871_));
  AOI21_X1   g0608(.A1(new_n417_), .A2(new_n416_), .B(\shift[1] ), .ZN(new_n872_));
  OAI21_X1   g0609(.A1(new_n871_), .A2(new_n872_), .B(new_n276_), .ZN(new_n873_));
  AOI21_X1   g0610(.A1(new_n870_), .A2(new_n873_), .B(new_n266_), .ZN(new_n874_));
  AOI21_X1   g0611(.A1(new_n414_), .A2(new_n413_), .B(new_n271_), .ZN(new_n875_));
  AOI21_X1   g0612(.A1(new_n433_), .A2(new_n432_), .B(\shift[1] ), .ZN(new_n876_));
  OAI21_X1   g0613(.A1(new_n875_), .A2(new_n876_), .B(new_n276_), .ZN(new_n877_));
  AOI21_X1   g0614(.A1(new_n421_), .A2(new_n420_), .B(new_n271_), .ZN(new_n878_));
  AOI21_X1   g0615(.A1(new_n409_), .A2(new_n408_), .B(\shift[1] ), .ZN(new_n879_));
  OAI21_X1   g0616(.A1(new_n878_), .A2(new_n879_), .B(\shift[3] ), .ZN(new_n880_));
  AOI21_X1   g0617(.A1(new_n877_), .A2(new_n880_), .B(\shift[2] ), .ZN(new_n881_));
  NOR2_X1    g0618(.A1(new_n874_), .A2(new_n881_), .ZN(new_n882_));
  OAI22_X1   g0619(.A1(new_n851_), .A2(new_n867_), .B1(new_n882_), .B2(new_n852_), .ZN(new_n883_));
  AOI21_X1   g0620(.A1(new_n462_), .A2(new_n461_), .B(new_n271_), .ZN(new_n884_));
  NAND2_X1   g0621(.A1(\a[37] ), .A2(\shift[0] ), .ZN(new_n885_));
  NAND2_X1   g0622(.A1(new_n268_), .A2(\a[38] ), .ZN(new_n886_));
  AOI21_X1   g0623(.A1(new_n886_), .A2(new_n885_), .B(\shift[1] ), .ZN(new_n887_));
  OAI21_X1   g0624(.A1(new_n884_), .A2(new_n887_), .B(\shift[3] ), .ZN(new_n888_));
  AOI21_X1   g0625(.A1(new_n480_), .A2(new_n479_), .B(\shift[1] ), .ZN(new_n889_));
  AOI21_X1   g0626(.A1(new_n469_), .A2(new_n468_), .B(new_n271_), .ZN(new_n890_));
  OAI21_X1   g0627(.A1(new_n889_), .A2(new_n890_), .B(new_n276_), .ZN(new_n891_));
  AOI21_X1   g0628(.A1(new_n888_), .A2(new_n891_), .B(new_n266_), .ZN(new_n892_));
  AOI21_X1   g0629(.A1(new_n477_), .A2(new_n476_), .B(new_n271_), .ZN(new_n893_));
  AOI21_X1   g0630(.A1(new_n500_), .A2(new_n499_), .B(\shift[1] ), .ZN(new_n894_));
  OAI21_X1   g0631(.A1(new_n893_), .A2(new_n894_), .B(new_n276_), .ZN(new_n895_));
  NAND2_X1   g0632(.A1(\a[39] ), .A2(\shift[0] ), .ZN(new_n896_));
  NAND2_X1   g0633(.A1(new_n268_), .A2(\a[40] ), .ZN(new_n897_));
  AOI21_X1   g0634(.A1(new_n897_), .A2(new_n896_), .B(new_n271_), .ZN(new_n898_));
  AOI21_X1   g0635(.A1(new_n472_), .A2(new_n471_), .B(\shift[1] ), .ZN(new_n899_));
  OAI21_X1   g0636(.A1(new_n898_), .A2(new_n899_), .B(\shift[3] ), .ZN(new_n900_));
  AOI21_X1   g0637(.A1(new_n895_), .A2(new_n900_), .B(\shift[2] ), .ZN(new_n901_));
  OAI21_X1   g0638(.A1(new_n892_), .A2(new_n901_), .B(new_n722_), .ZN(new_n902_));
  AOI21_X1   g0639(.A1(new_n430_), .A2(new_n429_), .B(new_n271_), .ZN(new_n903_));
  AOI21_X1   g0640(.A1(new_n455_), .A2(new_n454_), .B(\shift[1] ), .ZN(new_n904_));
  OAI21_X1   g0641(.A1(new_n903_), .A2(new_n904_), .B(\shift[3] ), .ZN(new_n905_));
  AOI21_X1   g0642(.A1(new_n437_), .A2(new_n436_), .B(new_n271_), .ZN(new_n906_));
  AOI21_X1   g0643(.A1(new_n448_), .A2(new_n447_), .B(\shift[1] ), .ZN(new_n907_));
  OAI21_X1   g0644(.A1(new_n906_), .A2(new_n907_), .B(new_n276_), .ZN(new_n908_));
  AOI21_X1   g0645(.A1(new_n905_), .A2(new_n908_), .B(new_n266_), .ZN(new_n909_));
  AOI21_X1   g0646(.A1(new_n445_), .A2(new_n444_), .B(new_n271_), .ZN(new_n910_));
  AOI21_X1   g0647(.A1(new_n465_), .A2(new_n464_), .B(\shift[1] ), .ZN(new_n911_));
  OAI21_X1   g0648(.A1(new_n910_), .A2(new_n911_), .B(new_n276_), .ZN(new_n912_));
  AOI21_X1   g0649(.A1(new_n452_), .A2(new_n451_), .B(new_n271_), .ZN(new_n913_));
  AOI21_X1   g0650(.A1(new_n440_), .A2(new_n439_), .B(\shift[1] ), .ZN(new_n914_));
  OAI21_X1   g0651(.A1(new_n913_), .A2(new_n914_), .B(\shift[3] ), .ZN(new_n915_));
  AOI21_X1   g0652(.A1(new_n912_), .A2(new_n915_), .B(\shift[2] ), .ZN(new_n916_));
  OAI21_X1   g0653(.A1(new_n909_), .A2(new_n916_), .B(new_n753_), .ZN(new_n917_));
  NAND2_X1   g0654(.A1(new_n902_), .A2(new_n917_), .ZN(new_n918_));
  OAI21_X1   g0655(.A1(new_n883_), .A2(new_n918_), .B(\shift[6] ), .ZN(new_n919_));
  NAND2_X1   g0656(.A1(new_n850_), .A2(new_n919_), .ZN(\result[2] ));
  INV_X1     g0657(.I(\a[103] ), .ZN(new_n921_));
  OAI22_X1   g0658(.A1(new_n490_), .A2(new_n921_), .B1(new_n594_), .B2(new_n491_), .ZN(new_n922_));
  INV_X1     g0659(.I(\a[102] ), .ZN(new_n923_));
  OAI22_X1   g0660(.A1(new_n597_), .A2(new_n485_), .B1(new_n486_), .B2(new_n923_), .ZN(new_n924_));
  OAI21_X1   g0661(.A1(new_n924_), .A2(new_n922_), .B(\shift[3] ), .ZN(new_n925_));
  INV_X1     g0662(.I(\a[111] ), .ZN(new_n926_));
  OAI22_X1   g0663(.A1(new_n490_), .A2(new_n926_), .B1(new_n601_), .B2(new_n491_), .ZN(new_n927_));
  OAI22_X1   g0664(.A1(new_n604_), .A2(new_n485_), .B1(new_n486_), .B2(new_n611_), .ZN(new_n928_));
  OAI21_X1   g0665(.A1(new_n928_), .A2(new_n927_), .B(new_n276_), .ZN(new_n929_));
  AOI21_X1   g0666(.A1(new_n925_), .A2(new_n929_), .B(new_n266_), .ZN(new_n930_));
  INV_X1     g0667(.I(\a[112] ), .ZN(new_n931_));
  OAI22_X1   g0668(.A1(new_n490_), .A2(new_n624_), .B1(new_n931_), .B2(new_n491_), .ZN(new_n932_));
  OAI22_X1   g0669(.A1(new_n612_), .A2(new_n485_), .B1(new_n486_), .B2(new_n627_), .ZN(new_n933_));
  OAI21_X1   g0670(.A1(new_n933_), .A2(new_n932_), .B(new_n276_), .ZN(new_n934_));
  INV_X1     g0671(.I(\a[104] ), .ZN(new_n935_));
  OAI22_X1   g0672(.A1(new_n490_), .A2(new_n600_), .B1(new_n935_), .B2(new_n491_), .ZN(new_n936_));
  OAI22_X1   g0673(.A1(new_n618_), .A2(new_n485_), .B1(new_n486_), .B2(new_n603_), .ZN(new_n937_));
  OAI21_X1   g0674(.A1(new_n937_), .A2(new_n936_), .B(\shift[3] ), .ZN(new_n938_));
  AOI21_X1   g0675(.A1(new_n938_), .A2(new_n934_), .B(\shift[2] ), .ZN(new_n939_));
  OAI21_X1   g0676(.A1(new_n930_), .A2(new_n939_), .B(new_n722_), .ZN(new_n940_));
  OAI22_X1   g0677(.A1(new_n490_), .A2(new_n583_), .B1(new_n562_), .B2(new_n491_), .ZN(new_n941_));
  OAI22_X1   g0678(.A1(new_n565_), .A2(new_n485_), .B1(new_n486_), .B2(new_n586_), .ZN(new_n942_));
  OAI21_X1   g0679(.A1(new_n942_), .A2(new_n941_), .B(\shift[3] ), .ZN(new_n943_));
  INV_X1     g0680(.I(\a[92] ), .ZN(new_n944_));
  INV_X1     g0681(.I(\a[95] ), .ZN(new_n945_));
  OAI22_X1   g0682(.A1(new_n490_), .A2(new_n945_), .B1(new_n944_), .B2(new_n491_), .ZN(new_n946_));
  OAI22_X1   g0683(.A1(new_n572_), .A2(new_n485_), .B1(new_n486_), .B2(new_n579_), .ZN(new_n947_));
  OAI21_X1   g0684(.A1(new_n947_), .A2(new_n946_), .B(new_n276_), .ZN(new_n948_));
  AOI21_X1   g0685(.A1(new_n943_), .A2(new_n948_), .B(new_n266_), .ZN(new_n949_));
  NAND3_X1   g0686(.A1(\a[96] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n950_));
  OAI21_X1   g0687(.A1(new_n490_), .A2(new_n593_), .B(new_n950_), .ZN(new_n951_));
  NAND3_X1   g0688(.A1(new_n268_), .A2(\a[97] ), .A3(\shift[1] ), .ZN(new_n952_));
  NAND3_X1   g0689(.A1(new_n271_), .A2(\a[98] ), .A3(\shift[0] ), .ZN(new_n953_));
  NAND2_X1   g0690(.A1(new_n952_), .A2(new_n953_), .ZN(new_n954_));
  OAI21_X1   g0691(.A1(new_n954_), .A2(new_n951_), .B(new_n276_), .ZN(new_n955_));
  INV_X1     g0692(.I(\a[91] ), .ZN(new_n956_));
  OAI22_X1   g0693(.A1(new_n490_), .A2(new_n956_), .B1(new_n584_), .B2(new_n491_), .ZN(new_n957_));
  NAND3_X1   g0694(.A1(new_n268_), .A2(\a[89] ), .A3(\shift[1] ), .ZN(new_n958_));
  NAND3_X1   g0695(.A1(new_n271_), .A2(\a[90] ), .A3(\shift[0] ), .ZN(new_n959_));
  NAND2_X1   g0696(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  OAI21_X1   g0697(.A1(new_n957_), .A2(new_n960_), .B(\shift[3] ), .ZN(new_n961_));
  AOI21_X1   g0698(.A1(new_n961_), .A2(new_n955_), .B(\shift[2] ), .ZN(new_n962_));
  OAI21_X1   g0699(.A1(new_n949_), .A2(new_n962_), .B(new_n753_), .ZN(new_n963_));
  NAND2_X1   g0700(.A1(new_n940_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1     g0701(.I(\a[119] ), .ZN(new_n965_));
  OAI22_X1   g0702(.A1(new_n490_), .A2(new_n965_), .B1(new_n625_), .B2(new_n491_), .ZN(new_n966_));
  INV_X1     g0703(.I(\a[118] ), .ZN(new_n967_));
  OAI22_X1   g0704(.A1(new_n628_), .A2(new_n485_), .B1(new_n486_), .B2(new_n967_), .ZN(new_n968_));
  OAI21_X1   g0705(.A1(new_n968_), .A2(new_n966_), .B(\shift[3] ), .ZN(new_n969_));
  INV_X1     g0706(.I(\a[127] ), .ZN(new_n970_));
  OAI22_X1   g0707(.A1(new_n490_), .A2(new_n970_), .B1(new_n632_), .B2(new_n491_), .ZN(new_n971_));
  OAI22_X1   g0708(.A1(new_n635_), .A2(new_n485_), .B1(new_n486_), .B2(new_n643_), .ZN(new_n972_));
  OAI21_X1   g0709(.A1(new_n972_), .A2(new_n971_), .B(new_n276_), .ZN(new_n973_));
  AOI21_X1   g0710(.A1(new_n969_), .A2(new_n973_), .B(new_n266_), .ZN(new_n974_));
  NAND3_X1   g0711(.A1(\a[0] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n975_));
  OAI21_X1   g0712(.A1(new_n490_), .A2(new_n690_), .B(new_n975_), .ZN(new_n976_));
  NAND3_X1   g0713(.A1(new_n268_), .A2(\a[1] ), .A3(\shift[1] ), .ZN(new_n977_));
  NAND3_X1   g0714(.A1(new_n271_), .A2(\a[2] ), .A3(\shift[0] ), .ZN(new_n978_));
  NAND2_X1   g0715(.A1(new_n977_), .A2(new_n978_), .ZN(new_n979_));
  OAI21_X1   g0716(.A1(new_n979_), .A2(new_n976_), .B(new_n276_), .ZN(new_n980_));
  INV_X1     g0717(.I(\a[120] ), .ZN(new_n981_));
  OAI22_X1   g0718(.A1(new_n490_), .A2(new_n631_), .B1(new_n981_), .B2(new_n491_), .ZN(new_n982_));
  OAI22_X1   g0719(.A1(new_n649_), .A2(new_n485_), .B1(new_n486_), .B2(new_n634_), .ZN(new_n983_));
  OAI21_X1   g0720(.A1(new_n983_), .A2(new_n982_), .B(\shift[3] ), .ZN(new_n984_));
  AOI21_X1   g0721(.A1(new_n984_), .A2(new_n980_), .B(\shift[2] ), .ZN(new_n985_));
  OAI21_X1   g0722(.A1(new_n974_), .A2(new_n985_), .B(new_n657_), .ZN(new_n986_));
  OAI22_X1   g0723(.A1(new_n490_), .A2(new_n552_), .B1(new_n531_), .B2(new_n491_), .ZN(new_n987_));
  OAI22_X1   g0724(.A1(new_n534_), .A2(new_n485_), .B1(new_n486_), .B2(new_n555_), .ZN(new_n988_));
  OAI21_X1   g0725(.A1(new_n988_), .A2(new_n987_), .B(\shift[3] ), .ZN(new_n989_));
  INV_X1     g0726(.I(\a[76] ), .ZN(new_n990_));
  OAI22_X1   g0727(.A1(new_n490_), .A2(new_n545_), .B1(new_n990_), .B2(new_n491_), .ZN(new_n991_));
  OAI22_X1   g0728(.A1(new_n541_), .A2(new_n485_), .B1(new_n486_), .B2(new_n548_), .ZN(new_n992_));
  OAI21_X1   g0729(.A1(new_n992_), .A2(new_n991_), .B(new_n276_), .ZN(new_n993_));
  AOI21_X1   g0730(.A1(new_n989_), .A2(new_n993_), .B(new_n266_), .ZN(new_n994_));
  OAI22_X1   g0731(.A1(new_n490_), .A2(new_n561_), .B1(new_n546_), .B2(new_n491_), .ZN(new_n995_));
  OAI22_X1   g0732(.A1(new_n549_), .A2(new_n485_), .B1(new_n486_), .B2(new_n564_), .ZN(new_n996_));
  OAI21_X1   g0733(.A1(new_n996_), .A2(new_n995_), .B(new_n276_), .ZN(new_n997_));
  INV_X1     g0734(.I(\a[75] ), .ZN(new_n998_));
  OAI22_X1   g0735(.A1(new_n490_), .A2(new_n998_), .B1(new_n553_), .B2(new_n491_), .ZN(new_n999_));
  OAI22_X1   g0736(.A1(new_n556_), .A2(new_n485_), .B1(new_n486_), .B2(new_n540_), .ZN(new_n1000_));
  OAI21_X1   g0737(.A1(new_n1000_), .A2(new_n999_), .B(\shift[3] ), .ZN(new_n1001_));
  AOI21_X1   g0738(.A1(new_n997_), .A2(new_n1001_), .B(\shift[2] ), .ZN(new_n1002_));
  OAI21_X1   g0739(.A1(new_n994_), .A2(new_n1002_), .B(new_n689_), .ZN(new_n1003_));
  NAND2_X1   g0740(.A1(new_n1003_), .A2(new_n986_), .ZN(new_n1004_));
  OAI21_X1   g0741(.A1(new_n1004_), .A2(new_n964_), .B(new_n264_), .ZN(new_n1005_));
  NAND3_X1   g0742(.A1(\a[36] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1006_));
  OAI21_X1   g0743(.A1(new_n490_), .A2(new_n484_), .B(new_n1006_), .ZN(new_n1007_));
  NAND3_X1   g0744(.A1(new_n268_), .A2(\a[37] ), .A3(\shift[1] ), .ZN(new_n1008_));
  NAND3_X1   g0745(.A1(new_n271_), .A2(\a[38] ), .A3(\shift[0] ), .ZN(new_n1009_));
  NAND2_X1   g0746(.A1(new_n1008_), .A2(new_n1009_), .ZN(new_n1010_));
  OAI21_X1   g0747(.A1(new_n1010_), .A2(new_n1007_), .B(\shift[3] ), .ZN(new_n1011_));
  NAND2_X1   g0748(.A1(\a[46] ), .A2(\shift[0] ), .ZN(new_n1012_));
  NAND2_X1   g0749(.A1(new_n268_), .A2(\a[47] ), .ZN(new_n1013_));
  AOI21_X1   g0750(.A1(new_n1013_), .A2(new_n1012_), .B(\shift[1] ), .ZN(new_n1014_));
  AOI21_X1   g0751(.A1(new_n730_), .A2(new_n729_), .B(new_n271_), .ZN(new_n1015_));
  OAI21_X1   g0752(.A1(new_n1014_), .A2(new_n1015_), .B(new_n276_), .ZN(new_n1016_));
  AOI21_X1   g0753(.A1(new_n1011_), .A2(new_n1016_), .B(new_n266_), .ZN(new_n1017_));
  INV_X1     g0754(.I(\a[48] ), .ZN(new_n1018_));
  INV_X1     g0755(.I(\a[51] ), .ZN(new_n1019_));
  OAI22_X1   g0756(.A1(new_n490_), .A2(new_n1019_), .B1(new_n1018_), .B2(new_n491_), .ZN(new_n1020_));
  NAND3_X1   g0757(.A1(new_n268_), .A2(\a[49] ), .A3(\shift[1] ), .ZN(new_n1021_));
  NAND3_X1   g0758(.A1(new_n271_), .A2(\a[50] ), .A3(\shift[0] ), .ZN(new_n1022_));
  NAND2_X1   g0759(.A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1023_));
  OAI21_X1   g0760(.A1(new_n1020_), .A2(new_n1023_), .B(new_n276_), .ZN(new_n1024_));
  INV_X1     g0761(.I(\a[43] ), .ZN(new_n1025_));
  OAI22_X1   g0762(.A1(new_n490_), .A2(new_n1025_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n1026_));
  NAND3_X1   g0763(.A1(new_n268_), .A2(\a[41] ), .A3(\shift[1] ), .ZN(new_n1027_));
  NAND3_X1   g0764(.A1(new_n271_), .A2(\a[42] ), .A3(\shift[0] ), .ZN(new_n1028_));
  NAND2_X1   g0765(.A1(new_n1027_), .A2(new_n1028_), .ZN(new_n1029_));
  OAI21_X1   g0766(.A1(new_n1026_), .A2(new_n1029_), .B(\shift[3] ), .ZN(new_n1030_));
  AOI21_X1   g0767(.A1(new_n1024_), .A2(new_n1030_), .B(\shift[2] ), .ZN(new_n1031_));
  OAI21_X1   g0768(.A1(new_n1031_), .A2(new_n1017_), .B(\shift[4] ), .ZN(new_n1032_));
  NAND3_X1   g0769(.A1(\a[52] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1033_));
  OAI21_X1   g0770(.A1(new_n490_), .A2(new_n680_), .B(new_n1033_), .ZN(new_n1034_));
  NAND3_X1   g0771(.A1(new_n268_), .A2(\a[53] ), .A3(\shift[1] ), .ZN(new_n1035_));
  NAND3_X1   g0772(.A1(new_n271_), .A2(\a[54] ), .A3(\shift[0] ), .ZN(new_n1036_));
  NAND2_X1   g0773(.A1(new_n1035_), .A2(new_n1036_), .ZN(new_n1037_));
  OAI21_X1   g0774(.A1(new_n1037_), .A2(new_n1034_), .B(\shift[3] ), .ZN(new_n1038_));
  INV_X1     g0775(.I(\a[60] ), .ZN(new_n1039_));
  INV_X1     g0776(.I(\a[63] ), .ZN(new_n1040_));
  OAI22_X1   g0777(.A1(new_n490_), .A2(new_n1040_), .B1(new_n1039_), .B2(new_n491_), .ZN(new_n1041_));
  NAND3_X1   g0778(.A1(new_n268_), .A2(\a[61] ), .A3(\shift[1] ), .ZN(new_n1042_));
  NAND3_X1   g0779(.A1(new_n271_), .A2(\a[62] ), .A3(\shift[0] ), .ZN(new_n1043_));
  NAND2_X1   g0780(.A1(new_n1042_), .A2(new_n1043_), .ZN(new_n1044_));
  OAI21_X1   g0781(.A1(new_n1041_), .A2(new_n1044_), .B(new_n276_), .ZN(new_n1045_));
  AOI21_X1   g0782(.A1(new_n1045_), .A2(new_n1038_), .B(new_n266_), .ZN(new_n1046_));
  NAND3_X1   g0783(.A1(\a[64] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1047_));
  OAI21_X1   g0784(.A1(new_n490_), .A2(new_n530_), .B(new_n1047_), .ZN(new_n1048_));
  NAND3_X1   g0785(.A1(new_n268_), .A2(\a[65] ), .A3(\shift[1] ), .ZN(new_n1049_));
  NAND3_X1   g0786(.A1(new_n271_), .A2(\a[66] ), .A3(\shift[0] ), .ZN(new_n1050_));
  NAND2_X1   g0787(.A1(new_n1049_), .A2(new_n1050_), .ZN(new_n1051_));
  OAI21_X1   g0788(.A1(new_n1051_), .A2(new_n1048_), .B(new_n276_), .ZN(new_n1052_));
  INV_X1     g0789(.I(\a[59] ), .ZN(new_n1053_));
  OAI22_X1   g0790(.A1(new_n490_), .A2(new_n1053_), .B1(new_n681_), .B2(new_n491_), .ZN(new_n1054_));
  OAI22_X1   g0791(.A1(new_n684_), .A2(new_n485_), .B1(new_n486_), .B2(new_n668_), .ZN(new_n1055_));
  OAI21_X1   g0792(.A1(new_n1055_), .A2(new_n1054_), .B(\shift[3] ), .ZN(new_n1056_));
  AOI21_X1   g0793(.A1(new_n1056_), .A2(new_n1052_), .B(\shift[2] ), .ZN(new_n1057_));
  OAI21_X1   g0794(.A1(new_n1057_), .A2(new_n1046_), .B(new_n301_), .ZN(new_n1058_));
  AOI21_X1   g0795(.A1(new_n1058_), .A2(new_n1032_), .B(\shift[5] ), .ZN(new_n1059_));
  INV_X1     g0796(.I(\a[7] ), .ZN(new_n1060_));
  OAI22_X1   g0797(.A1(new_n490_), .A2(new_n1060_), .B1(new_n691_), .B2(new_n491_), .ZN(new_n1061_));
  OAI22_X1   g0798(.A1(new_n694_), .A2(new_n485_), .B1(new_n486_), .B2(new_n715_), .ZN(new_n1062_));
  OAI21_X1   g0799(.A1(new_n1062_), .A2(new_n1061_), .B(\shift[3] ), .ZN(new_n1063_));
  INV_X1     g0800(.I(\a[15] ), .ZN(new_n1064_));
  OAI22_X1   g0801(.A1(new_n490_), .A2(new_n1064_), .B1(new_n698_), .B2(new_n491_), .ZN(new_n1065_));
  OAI22_X1   g0802(.A1(new_n701_), .A2(new_n485_), .B1(new_n486_), .B2(new_n708_), .ZN(new_n1066_));
  OAI21_X1   g0803(.A1(new_n1066_), .A2(new_n1065_), .B(new_n276_), .ZN(new_n1067_));
  AOI21_X1   g0804(.A1(new_n1063_), .A2(new_n1067_), .B(new_n266_), .ZN(new_n1068_));
  NAND3_X1   g0805(.A1(\a[16] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1069_));
  OAI21_X1   g0806(.A1(new_n490_), .A2(new_n754_), .B(new_n1069_), .ZN(new_n1070_));
  NAND3_X1   g0807(.A1(new_n268_), .A2(\a[17] ), .A3(\shift[1] ), .ZN(new_n1071_));
  NAND3_X1   g0808(.A1(new_n271_), .A2(\a[18] ), .A3(\shift[0] ), .ZN(new_n1072_));
  NAND2_X1   g0809(.A1(new_n1071_), .A2(new_n1072_), .ZN(new_n1073_));
  OAI21_X1   g0810(.A1(new_n1073_), .A2(new_n1070_), .B(new_n276_), .ZN(new_n1074_));
  NAND3_X1   g0811(.A1(\a[8] ), .A2(\shift[0] ), .A3(\shift[1] ), .ZN(new_n1075_));
  OAI21_X1   g0812(.A1(new_n490_), .A2(new_n697_), .B(new_n1075_), .ZN(new_n1076_));
  NAND3_X1   g0813(.A1(new_n268_), .A2(\a[9] ), .A3(\shift[1] ), .ZN(new_n1077_));
  NAND3_X1   g0814(.A1(new_n271_), .A2(\a[10] ), .A3(\shift[0] ), .ZN(new_n1078_));
  NAND2_X1   g0815(.A1(new_n1077_), .A2(new_n1078_), .ZN(new_n1079_));
  OAI21_X1   g0816(.A1(new_n1079_), .A2(new_n1076_), .B(\shift[3] ), .ZN(new_n1080_));
  AOI21_X1   g0817(.A1(new_n1074_), .A2(new_n1080_), .B(\shift[2] ), .ZN(new_n1081_));
  OAI21_X1   g0818(.A1(new_n1068_), .A2(new_n1081_), .B(\shift[4] ), .ZN(new_n1082_));
  INV_X1     g0819(.I(\a[23] ), .ZN(new_n1083_));
  OAI22_X1   g0820(.A1(new_n490_), .A2(new_n1083_), .B1(new_n755_), .B2(new_n491_), .ZN(new_n1084_));
  OAI22_X1   g0821(.A1(new_n758_), .A2(new_n485_), .B1(new_n486_), .B2(new_n779_), .ZN(new_n1085_));
  OAI21_X1   g0822(.A1(new_n1085_), .A2(new_n1084_), .B(\shift[3] ), .ZN(new_n1086_));
  INV_X1     g0823(.I(\a[28] ), .ZN(new_n1087_));
  INV_X1     g0824(.I(\a[31] ), .ZN(new_n1088_));
  OAI22_X1   g0825(.A1(new_n490_), .A2(new_n1088_), .B1(new_n1087_), .B2(new_n491_), .ZN(new_n1089_));
  NAND3_X1   g0826(.A1(new_n268_), .A2(\a[29] ), .A3(\shift[1] ), .ZN(new_n1090_));
  NAND3_X1   g0827(.A1(new_n271_), .A2(\a[30] ), .A3(\shift[0] ), .ZN(new_n1091_));
  NAND2_X1   g0828(.A1(new_n1090_), .A2(new_n1091_), .ZN(new_n1092_));
  OAI21_X1   g0829(.A1(new_n1089_), .A2(new_n1092_), .B(new_n276_), .ZN(new_n1093_));
  AOI21_X1   g0830(.A1(new_n1086_), .A2(new_n1093_), .B(new_n266_), .ZN(new_n1094_));
  INV_X1     g0831(.I(\a[32] ), .ZN(new_n1095_));
  INV_X1     g0832(.I(\a[35] ), .ZN(new_n1096_));
  OAI22_X1   g0833(.A1(new_n490_), .A2(new_n1096_), .B1(new_n1095_), .B2(new_n491_), .ZN(new_n1097_));
  NAND3_X1   g0834(.A1(new_n268_), .A2(\a[33] ), .A3(\shift[1] ), .ZN(new_n1098_));
  NAND3_X1   g0835(.A1(new_n271_), .A2(\a[34] ), .A3(\shift[0] ), .ZN(new_n1099_));
  NAND2_X1   g0836(.A1(new_n1098_), .A2(new_n1099_), .ZN(new_n1100_));
  OAI21_X1   g0837(.A1(new_n1097_), .A2(new_n1100_), .B(new_n276_), .ZN(new_n1101_));
  INV_X1     g0838(.I(\a[24] ), .ZN(new_n1102_));
  INV_X1     g0839(.I(\a[27] ), .ZN(new_n1103_));
  OAI22_X1   g0840(.A1(new_n490_), .A2(new_n1103_), .B1(new_n1102_), .B2(new_n491_), .ZN(new_n1104_));
  NAND3_X1   g0841(.A1(new_n268_), .A2(\a[25] ), .A3(\shift[1] ), .ZN(new_n1105_));
  NAND3_X1   g0842(.A1(new_n271_), .A2(\a[26] ), .A3(\shift[0] ), .ZN(new_n1106_));
  NAND2_X1   g0843(.A1(new_n1105_), .A2(new_n1106_), .ZN(new_n1107_));
  OAI21_X1   g0844(.A1(new_n1104_), .A2(new_n1107_), .B(\shift[3] ), .ZN(new_n1108_));
  AOI21_X1   g0845(.A1(new_n1101_), .A2(new_n1108_), .B(\shift[2] ), .ZN(new_n1109_));
  OAI21_X1   g0846(.A1(new_n1094_), .A2(new_n1109_), .B(new_n301_), .ZN(new_n1110_));
  AOI21_X1   g0847(.A1(new_n1110_), .A2(new_n1082_), .B(new_n265_), .ZN(new_n1111_));
  OAI21_X1   g0848(.A1(new_n1111_), .A2(new_n1059_), .B(\shift[6] ), .ZN(new_n1112_));
  NAND2_X1   g0849(.A1(new_n1112_), .A2(new_n1005_), .ZN(\result[3] ));
  AOI21_X1   g0850(.A1(new_n291_), .A2(new_n298_), .B(new_n266_), .ZN(new_n1114_));
  OAI21_X1   g0851(.A1(new_n304_), .A2(new_n307_), .B(new_n276_), .ZN(new_n1115_));
  OAI21_X1   g0852(.A1(new_n279_), .A2(new_n282_), .B(\shift[3] ), .ZN(new_n1116_));
  AOI21_X1   g0853(.A1(new_n1115_), .A2(new_n1116_), .B(\shift[2] ), .ZN(new_n1117_));
  OAI21_X1   g0854(.A1(new_n1114_), .A2(new_n1117_), .B(\shift[4] ), .ZN(new_n1118_));
  AOI21_X1   g0855(.A1(new_n323_), .A2(new_n330_), .B(new_n266_), .ZN(new_n1119_));
  OAI21_X1   g0856(.A1(new_n336_), .A2(new_n339_), .B(new_n276_), .ZN(new_n1120_));
  OAI21_X1   g0857(.A1(new_n311_), .A2(new_n314_), .B(\shift[3] ), .ZN(new_n1121_));
  AOI21_X1   g0858(.A1(new_n1120_), .A2(new_n1121_), .B(\shift[2] ), .ZN(new_n1122_));
  OAI21_X1   g0859(.A1(new_n1119_), .A2(new_n1122_), .B(new_n301_), .ZN(new_n1123_));
  AOI21_X1   g0860(.A1(new_n1118_), .A2(new_n1123_), .B(new_n265_), .ZN(new_n1124_));
  AOI21_X1   g0861(.A1(new_n355_), .A2(new_n362_), .B(new_n266_), .ZN(new_n1125_));
  OAI21_X1   g0862(.A1(new_n367_), .A2(new_n370_), .B(new_n276_), .ZN(new_n1126_));
  OAI21_X1   g0863(.A1(new_n343_), .A2(new_n346_), .B(\shift[3] ), .ZN(new_n1127_));
  AOI21_X1   g0864(.A1(new_n1126_), .A2(new_n1127_), .B(\shift[2] ), .ZN(new_n1128_));
  OAI21_X1   g0865(.A1(new_n1125_), .A2(new_n1128_), .B(\shift[4] ), .ZN(new_n1129_));
  AOI21_X1   g0866(.A1(new_n386_), .A2(new_n393_), .B(new_n266_), .ZN(new_n1130_));
  OAI21_X1   g0867(.A1(new_n400_), .A2(new_n403_), .B(new_n276_), .ZN(new_n1131_));
  OAI21_X1   g0868(.A1(new_n374_), .A2(new_n377_), .B(\shift[3] ), .ZN(new_n1132_));
  AOI21_X1   g0869(.A1(new_n1131_), .A2(new_n1132_), .B(\shift[2] ), .ZN(new_n1133_));
  OAI21_X1   g0870(.A1(new_n1130_), .A2(new_n1133_), .B(new_n301_), .ZN(new_n1134_));
  AOI21_X1   g0871(.A1(new_n1129_), .A2(new_n1134_), .B(\shift[5] ), .ZN(new_n1135_));
  OAI21_X1   g0872(.A1(new_n1124_), .A2(new_n1135_), .B(new_n264_), .ZN(new_n1136_));
  AOI21_X1   g0873(.A1(new_n493_), .A2(new_n482_), .B(new_n266_), .ZN(new_n1137_));
  OAI21_X1   g0874(.A1(new_n498_), .A2(new_n501_), .B(new_n276_), .ZN(new_n1138_));
  OAI21_X1   g0875(.A1(new_n470_), .A2(new_n473_), .B(\shift[3] ), .ZN(new_n1139_));
  AOI21_X1   g0876(.A1(new_n1138_), .A2(new_n1139_), .B(\shift[2] ), .ZN(new_n1140_));
  OAI21_X1   g0877(.A1(new_n1137_), .A2(new_n1140_), .B(\shift[4] ), .ZN(new_n1141_));
  AOI21_X1   g0878(.A1(new_n517_), .A2(new_n524_), .B(new_n266_), .ZN(new_n1142_));
  OAI21_X1   g0879(.A1(new_n270_), .A2(new_n274_), .B(new_n276_), .ZN(new_n1143_));
  OAI21_X1   g0880(.A1(new_n505_), .A2(new_n508_), .B(\shift[3] ), .ZN(new_n1144_));
  AOI21_X1   g0881(.A1(new_n1143_), .A2(new_n1144_), .B(\shift[2] ), .ZN(new_n1145_));
  OAI21_X1   g0882(.A1(new_n1142_), .A2(new_n1145_), .B(new_n301_), .ZN(new_n1146_));
  AOI21_X1   g0883(.A1(new_n1141_), .A2(new_n1146_), .B(\shift[5] ), .ZN(new_n1147_));
  AOI21_X1   g0884(.A1(new_n450_), .A2(new_n457_), .B(new_n266_), .ZN(new_n1148_));
  OAI21_X1   g0885(.A1(new_n463_), .A2(new_n466_), .B(new_n276_), .ZN(new_n1149_));
  OAI21_X1   g0886(.A1(new_n438_), .A2(new_n441_), .B(\shift[3] ), .ZN(new_n1150_));
  AOI21_X1   g0887(.A1(new_n1149_), .A2(new_n1150_), .B(\shift[2] ), .ZN(new_n1151_));
  OAI21_X1   g0888(.A1(new_n1148_), .A2(new_n1151_), .B(new_n301_), .ZN(new_n1152_));
  AOI21_X1   g0889(.A1(new_n419_), .A2(new_n426_), .B(new_n266_), .ZN(new_n1153_));
  OAI21_X1   g0890(.A1(new_n431_), .A2(new_n434_), .B(new_n276_), .ZN(new_n1154_));
  OAI21_X1   g0891(.A1(new_n407_), .A2(new_n410_), .B(\shift[3] ), .ZN(new_n1155_));
  AOI21_X1   g0892(.A1(new_n1154_), .A2(new_n1155_), .B(\shift[2] ), .ZN(new_n1156_));
  OAI21_X1   g0893(.A1(new_n1153_), .A2(new_n1156_), .B(\shift[4] ), .ZN(new_n1157_));
  AOI21_X1   g0894(.A1(new_n1152_), .A2(new_n1157_), .B(new_n265_), .ZN(new_n1158_));
  OAI21_X1   g0895(.A1(new_n1147_), .A2(new_n1158_), .B(\shift[6] ), .ZN(new_n1159_));
  NAND2_X1   g0896(.A1(new_n1136_), .A2(new_n1159_), .ZN(\result[4] ));
  AOI21_X1   g0897(.A1(new_n551_), .A2(new_n558_), .B(new_n266_), .ZN(new_n1161_));
  OAI21_X1   g0898(.A1(new_n563_), .A2(new_n566_), .B(new_n276_), .ZN(new_n1162_));
  OAI21_X1   g0899(.A1(new_n542_), .A2(new_n539_), .B(\shift[3] ), .ZN(new_n1163_));
  AOI21_X1   g0900(.A1(new_n1162_), .A2(new_n1163_), .B(\shift[2] ), .ZN(new_n1164_));
  OAI21_X1   g0901(.A1(new_n1161_), .A2(new_n1164_), .B(\shift[4] ), .ZN(new_n1165_));
  AOI21_X1   g0902(.A1(new_n589_), .A2(new_n582_), .B(new_n266_), .ZN(new_n1166_));
  OAI21_X1   g0903(.A1(new_n595_), .A2(new_n598_), .B(new_n276_), .ZN(new_n1167_));
  OAI21_X1   g0904(.A1(new_n573_), .A2(new_n570_), .B(\shift[3] ), .ZN(new_n1168_));
  AOI21_X1   g0905(.A1(new_n1167_), .A2(new_n1168_), .B(\shift[2] ), .ZN(new_n1169_));
  OAI21_X1   g0906(.A1(new_n1166_), .A2(new_n1169_), .B(new_n301_), .ZN(new_n1170_));
  AOI21_X1   g0907(.A1(new_n1165_), .A2(new_n1170_), .B(new_n265_), .ZN(new_n1171_));
  AOI21_X1   g0908(.A1(new_n614_), .A2(new_n621_), .B(new_n266_), .ZN(new_n1172_));
  OAI21_X1   g0909(.A1(new_n626_), .A2(new_n629_), .B(new_n276_), .ZN(new_n1173_));
  OAI21_X1   g0910(.A1(new_n602_), .A2(new_n605_), .B(\shift[3] ), .ZN(new_n1174_));
  AOI21_X1   g0911(.A1(new_n1173_), .A2(new_n1174_), .B(\shift[2] ), .ZN(new_n1175_));
  OAI21_X1   g0912(.A1(new_n1175_), .A2(new_n1172_), .B(\shift[4] ), .ZN(new_n1176_));
  AOI21_X1   g0913(.A1(new_n645_), .A2(new_n652_), .B(new_n266_), .ZN(new_n1177_));
  OAI21_X1   g0914(.A1(new_n692_), .A2(new_n695_), .B(new_n276_), .ZN(new_n1178_));
  OAI21_X1   g0915(.A1(new_n633_), .A2(new_n636_), .B(\shift[3] ), .ZN(new_n1179_));
  AOI21_X1   g0916(.A1(new_n1178_), .A2(new_n1179_), .B(\shift[2] ), .ZN(new_n1180_));
  OAI21_X1   g0917(.A1(new_n1180_), .A2(new_n1177_), .B(new_n301_), .ZN(new_n1181_));
  AOI21_X1   g0918(.A1(new_n1176_), .A2(new_n1181_), .B(\shift[5] ), .ZN(new_n1182_));
  OAI21_X1   g0919(.A1(new_n1171_), .A2(new_n1182_), .B(new_n264_), .ZN(new_n1183_));
  AOI21_X1   g0920(.A1(new_n743_), .A2(new_n750_), .B(new_n266_), .ZN(new_n1184_));
  OAI21_X1   g0921(.A1(new_n663_), .A2(new_n660_), .B(new_n276_), .ZN(new_n1185_));
  OAI21_X1   g0922(.A1(new_n731_), .A2(new_n734_), .B(\shift[3] ), .ZN(new_n1186_));
  AOI21_X1   g0923(.A1(new_n1185_), .A2(new_n1186_), .B(\shift[2] ), .ZN(new_n1187_));
  OAI21_X1   g0924(.A1(new_n1184_), .A2(new_n1187_), .B(\shift[4] ), .ZN(new_n1188_));
  AOI21_X1   g0925(.A1(new_n686_), .A2(new_n679_), .B(new_n266_), .ZN(new_n1189_));
  OAI21_X1   g0926(.A1(new_n532_), .A2(new_n535_), .B(new_n276_), .ZN(new_n1190_));
  OAI21_X1   g0927(.A1(new_n670_), .A2(new_n667_), .B(\shift[3] ), .ZN(new_n1191_));
  AOI21_X1   g0928(.A1(new_n1190_), .A2(new_n1191_), .B(\shift[2] ), .ZN(new_n1192_));
  OAI21_X1   g0929(.A1(new_n1189_), .A2(new_n1192_), .B(new_n301_), .ZN(new_n1193_));
  AOI21_X1   g0930(.A1(new_n1193_), .A2(new_n1188_), .B(\shift[5] ), .ZN(new_n1194_));
  AOI21_X1   g0931(.A1(new_n775_), .A2(new_n782_), .B(new_n266_), .ZN(new_n1195_));
  OAI21_X1   g0932(.A1(new_n725_), .A2(new_n727_), .B(new_n276_), .ZN(new_n1196_));
  OAI21_X1   g0933(.A1(new_n766_), .A2(new_n763_), .B(\shift[3] ), .ZN(new_n1197_));
  AOI21_X1   g0934(.A1(new_n1197_), .A2(new_n1196_), .B(\shift[2] ), .ZN(new_n1198_));
  OAI21_X1   g0935(.A1(new_n1195_), .A2(new_n1198_), .B(new_n301_), .ZN(new_n1199_));
  AOI21_X1   g0936(.A1(new_n711_), .A2(new_n718_), .B(new_n266_), .ZN(new_n1200_));
  OAI21_X1   g0937(.A1(new_n756_), .A2(new_n759_), .B(new_n276_), .ZN(new_n1201_));
  OAI21_X1   g0938(.A1(new_n699_), .A2(new_n702_), .B(\shift[3] ), .ZN(new_n1202_));
  AOI21_X1   g0939(.A1(new_n1201_), .A2(new_n1202_), .B(\shift[2] ), .ZN(new_n1203_));
  OAI21_X1   g0940(.A1(new_n1203_), .A2(new_n1200_), .B(\shift[4] ), .ZN(new_n1204_));
  AOI21_X1   g0941(.A1(new_n1204_), .A2(new_n1199_), .B(new_n265_), .ZN(new_n1205_));
  OAI21_X1   g0942(.A1(new_n1205_), .A2(new_n1194_), .B(\shift[6] ), .ZN(new_n1206_));
  NAND2_X1   g0943(.A1(new_n1183_), .A2(new_n1206_), .ZN(\result[5] ));
  AOI21_X1   g0944(.A1(new_n797_), .A2(new_n800_), .B(new_n266_), .ZN(new_n1208_));
  OAI21_X1   g0945(.A1(new_n803_), .A2(new_n804_), .B(new_n276_), .ZN(new_n1209_));
  OAI21_X1   g0946(.A1(new_n791_), .A2(new_n792_), .B(\shift[3] ), .ZN(new_n1210_));
  AOI21_X1   g0947(.A1(new_n1209_), .A2(new_n1210_), .B(\shift[2] ), .ZN(new_n1211_));
  OAI21_X1   g0948(.A1(new_n1208_), .A2(new_n1211_), .B(\shift[4] ), .ZN(new_n1212_));
  AOI21_X1   g0949(.A1(new_n812_), .A2(new_n815_), .B(new_n266_), .ZN(new_n1213_));
  OAI21_X1   g0950(.A1(new_n819_), .A2(new_n820_), .B(new_n276_), .ZN(new_n1214_));
  OAI21_X1   g0951(.A1(new_n806_), .A2(new_n807_), .B(\shift[3] ), .ZN(new_n1215_));
  AOI21_X1   g0952(.A1(new_n1214_), .A2(new_n1215_), .B(\shift[2] ), .ZN(new_n1216_));
  OAI21_X1   g0953(.A1(new_n1213_), .A2(new_n1216_), .B(new_n301_), .ZN(new_n1217_));
  AOI21_X1   g0954(.A1(new_n1212_), .A2(new_n1217_), .B(new_n265_), .ZN(new_n1218_));
  AOI21_X1   g0955(.A1(new_n828_), .A2(new_n831_), .B(new_n266_), .ZN(new_n1219_));
  OAI21_X1   g0956(.A1(new_n834_), .A2(new_n835_), .B(new_n276_), .ZN(new_n1220_));
  OAI21_X1   g0957(.A1(new_n822_), .A2(new_n823_), .B(\shift[3] ), .ZN(new_n1221_));
  AOI21_X1   g0958(.A1(new_n1220_), .A2(new_n1221_), .B(\shift[2] ), .ZN(new_n1222_));
  OAI21_X1   g0959(.A1(new_n1219_), .A2(new_n1222_), .B(\shift[4] ), .ZN(new_n1223_));
  AOI21_X1   g0960(.A1(new_n843_), .A2(new_n846_), .B(new_n266_), .ZN(new_n1224_));
  OAI21_X1   g0961(.A1(new_n868_), .A2(new_n869_), .B(new_n276_), .ZN(new_n1225_));
  OAI21_X1   g0962(.A1(new_n837_), .A2(new_n838_), .B(\shift[3] ), .ZN(new_n1226_));
  AOI21_X1   g0963(.A1(new_n1225_), .A2(new_n1226_), .B(\shift[2] ), .ZN(new_n1227_));
  OAI21_X1   g0964(.A1(new_n1224_), .A2(new_n1227_), .B(new_n301_), .ZN(new_n1228_));
  AOI21_X1   g0965(.A1(new_n1223_), .A2(new_n1228_), .B(\shift[5] ), .ZN(new_n1229_));
  OAI21_X1   g0966(.A1(new_n1218_), .A2(new_n1229_), .B(new_n264_), .ZN(new_n1230_));
  AOI21_X1   g0967(.A1(new_n895_), .A2(new_n900_), .B(new_n266_), .ZN(new_n1231_));
  OAI21_X1   g0968(.A1(new_n853_), .A2(new_n854_), .B(new_n276_), .ZN(new_n1232_));
  OAI21_X1   g0969(.A1(new_n889_), .A2(new_n890_), .B(\shift[3] ), .ZN(new_n1233_));
  AOI21_X1   g0970(.A1(new_n1232_), .A2(new_n1233_), .B(\shift[2] ), .ZN(new_n1234_));
  OAI21_X1   g0971(.A1(new_n1231_), .A2(new_n1234_), .B(\shift[4] ), .ZN(new_n1235_));
  AOI21_X1   g0972(.A1(new_n862_), .A2(new_n865_), .B(new_n266_), .ZN(new_n1236_));
  OAI21_X1   g0973(.A1(new_n788_), .A2(new_n789_), .B(new_n276_), .ZN(new_n1237_));
  OAI21_X1   g0974(.A1(new_n856_), .A2(new_n857_), .B(\shift[3] ), .ZN(new_n1238_));
  AOI21_X1   g0975(.A1(new_n1237_), .A2(new_n1238_), .B(\shift[2] ), .ZN(new_n1239_));
  OAI21_X1   g0976(.A1(new_n1236_), .A2(new_n1239_), .B(new_n301_), .ZN(new_n1240_));
  AOI21_X1   g0977(.A1(new_n1235_), .A2(new_n1240_), .B(\shift[5] ), .ZN(new_n1241_));
  AOI21_X1   g0978(.A1(new_n912_), .A2(new_n915_), .B(new_n266_), .ZN(new_n1242_));
  OAI21_X1   g0979(.A1(new_n884_), .A2(new_n887_), .B(new_n276_), .ZN(new_n1243_));
  OAI21_X1   g0980(.A1(new_n906_), .A2(new_n907_), .B(\shift[3] ), .ZN(new_n1244_));
  AOI21_X1   g0981(.A1(new_n1243_), .A2(new_n1244_), .B(\shift[2] ), .ZN(new_n1245_));
  OAI21_X1   g0982(.A1(new_n1242_), .A2(new_n1245_), .B(new_n301_), .ZN(new_n1246_));
  AOI21_X1   g0983(.A1(new_n877_), .A2(new_n880_), .B(new_n266_), .ZN(new_n1247_));
  OAI21_X1   g0984(.A1(new_n903_), .A2(new_n904_), .B(new_n276_), .ZN(new_n1248_));
  OAI21_X1   g0985(.A1(new_n871_), .A2(new_n872_), .B(\shift[3] ), .ZN(new_n1249_));
  AOI21_X1   g0986(.A1(new_n1248_), .A2(new_n1249_), .B(\shift[2] ), .ZN(new_n1250_));
  OAI21_X1   g0987(.A1(new_n1247_), .A2(new_n1250_), .B(\shift[4] ), .ZN(new_n1251_));
  AOI21_X1   g0988(.A1(new_n1246_), .A2(new_n1251_), .B(new_n265_), .ZN(new_n1252_));
  OAI21_X1   g0989(.A1(new_n1241_), .A2(new_n1252_), .B(\shift[6] ), .ZN(new_n1253_));
  NAND2_X1   g0990(.A1(new_n1230_), .A2(new_n1253_), .ZN(\result[6] ));
  AOI21_X1   g0991(.A1(new_n997_), .A2(new_n1001_), .B(new_n266_), .ZN(new_n1255_));
  OAI21_X1   g0992(.A1(new_n942_), .A2(new_n941_), .B(new_n276_), .ZN(new_n1256_));
  OAI21_X1   g0993(.A1(new_n992_), .A2(new_n991_), .B(\shift[3] ), .ZN(new_n1257_));
  AOI21_X1   g0994(.A1(new_n1256_), .A2(new_n1257_), .B(\shift[2] ), .ZN(new_n1258_));
  OAI21_X1   g0995(.A1(new_n1255_), .A2(new_n1258_), .B(\shift[4] ), .ZN(new_n1259_));
  AOI21_X1   g0996(.A1(new_n961_), .A2(new_n955_), .B(new_n266_), .ZN(new_n1260_));
  OAI21_X1   g0997(.A1(new_n924_), .A2(new_n922_), .B(new_n276_), .ZN(new_n1261_));
  OAI21_X1   g0998(.A1(new_n947_), .A2(new_n946_), .B(\shift[3] ), .ZN(new_n1262_));
  AOI21_X1   g0999(.A1(new_n1261_), .A2(new_n1262_), .B(\shift[2] ), .ZN(new_n1263_));
  OAI21_X1   g1000(.A1(new_n1263_), .A2(new_n1260_), .B(new_n301_), .ZN(new_n1264_));
  AOI21_X1   g1001(.A1(new_n1259_), .A2(new_n1264_), .B(new_n265_), .ZN(new_n1265_));
  AOI21_X1   g1002(.A1(new_n938_), .A2(new_n934_), .B(new_n266_), .ZN(new_n1266_));
  OAI21_X1   g1003(.A1(new_n968_), .A2(new_n966_), .B(new_n276_), .ZN(new_n1267_));
  OAI21_X1   g1004(.A1(new_n928_), .A2(new_n927_), .B(\shift[3] ), .ZN(new_n1268_));
  AOI21_X1   g1005(.A1(new_n1267_), .A2(new_n1268_), .B(\shift[2] ), .ZN(new_n1269_));
  OAI21_X1   g1006(.A1(new_n1266_), .A2(new_n1269_), .B(\shift[4] ), .ZN(new_n1270_));
  AOI21_X1   g1007(.A1(new_n984_), .A2(new_n980_), .B(new_n266_), .ZN(new_n1271_));
  OAI21_X1   g1008(.A1(new_n1062_), .A2(new_n1061_), .B(new_n276_), .ZN(new_n1272_));
  OAI21_X1   g1009(.A1(new_n972_), .A2(new_n971_), .B(\shift[3] ), .ZN(new_n1273_));
  AOI21_X1   g1010(.A1(new_n1272_), .A2(new_n1273_), .B(\shift[2] ), .ZN(new_n1274_));
  OAI21_X1   g1011(.A1(new_n1274_), .A2(new_n1271_), .B(new_n301_), .ZN(new_n1275_));
  AOI21_X1   g1012(.A1(new_n1270_), .A2(new_n1275_), .B(\shift[5] ), .ZN(new_n1276_));
  OAI21_X1   g1013(.A1(new_n1276_), .A2(new_n1265_), .B(new_n264_), .ZN(new_n1277_));
  AOI21_X1   g1014(.A1(new_n1024_), .A2(new_n1030_), .B(new_n266_), .ZN(new_n1278_));
  OAI21_X1   g1015(.A1(new_n1014_), .A2(new_n1015_), .B(\shift[3] ), .ZN(new_n1279_));
  OAI21_X1   g1016(.A1(new_n1037_), .A2(new_n1034_), .B(new_n276_), .ZN(new_n1280_));
  AOI21_X1   g1017(.A1(new_n1280_), .A2(new_n1279_), .B(\shift[2] ), .ZN(new_n1281_));
  OAI21_X1   g1018(.A1(new_n1278_), .A2(new_n1281_), .B(\shift[4] ), .ZN(new_n1282_));
  AOI21_X1   g1019(.A1(new_n1056_), .A2(new_n1052_), .B(new_n266_), .ZN(new_n1283_));
  OAI21_X1   g1020(.A1(new_n988_), .A2(new_n987_), .B(new_n276_), .ZN(new_n1284_));
  OAI21_X1   g1021(.A1(new_n1041_), .A2(new_n1044_), .B(\shift[3] ), .ZN(new_n1285_));
  AOI21_X1   g1022(.A1(new_n1284_), .A2(new_n1285_), .B(\shift[2] ), .ZN(new_n1286_));
  OAI21_X1   g1023(.A1(new_n1286_), .A2(new_n1283_), .B(new_n301_), .ZN(new_n1287_));
  AOI21_X1   g1024(.A1(new_n1287_), .A2(new_n1282_), .B(\shift[5] ), .ZN(new_n1288_));
  AOI21_X1   g1025(.A1(new_n1101_), .A2(new_n1108_), .B(new_n266_), .ZN(new_n1289_));
  OAI21_X1   g1026(.A1(new_n1010_), .A2(new_n1007_), .B(new_n276_), .ZN(new_n1290_));
  OAI21_X1   g1027(.A1(new_n1089_), .A2(new_n1092_), .B(\shift[3] ), .ZN(new_n1291_));
  AOI21_X1   g1028(.A1(new_n1291_), .A2(new_n1290_), .B(\shift[2] ), .ZN(new_n1292_));
  OAI21_X1   g1029(.A1(new_n1289_), .A2(new_n1292_), .B(new_n301_), .ZN(new_n1293_));
  AOI21_X1   g1030(.A1(new_n1074_), .A2(new_n1080_), .B(new_n266_), .ZN(new_n1294_));
  OAI21_X1   g1031(.A1(new_n1085_), .A2(new_n1084_), .B(new_n276_), .ZN(new_n1295_));
  OAI21_X1   g1032(.A1(new_n1066_), .A2(new_n1065_), .B(\shift[3] ), .ZN(new_n1296_));
  AOI21_X1   g1033(.A1(new_n1295_), .A2(new_n1296_), .B(\shift[2] ), .ZN(new_n1297_));
  OAI21_X1   g1034(.A1(new_n1297_), .A2(new_n1294_), .B(\shift[4] ), .ZN(new_n1298_));
  AOI21_X1   g1035(.A1(new_n1298_), .A2(new_n1293_), .B(new_n265_), .ZN(new_n1299_));
  OAI21_X1   g1036(.A1(new_n1299_), .A2(new_n1288_), .B(\shift[6] ), .ZN(new_n1300_));
  NAND2_X1   g1037(.A1(new_n1277_), .A2(new_n1300_), .ZN(\result[7] ));
  AOI21_X1   g1038(.A1(new_n1115_), .A2(new_n1116_), .B(new_n266_), .ZN(new_n1302_));
  OAI21_X1   g1039(.A1(new_n326_), .A2(new_n329_), .B(new_n276_), .ZN(new_n1303_));
  OAI21_X1   g1040(.A1(new_n287_), .A2(new_n290_), .B(\shift[3] ), .ZN(new_n1304_));
  AOI21_X1   g1041(.A1(new_n1303_), .A2(new_n1304_), .B(\shift[2] ), .ZN(new_n1305_));
  OAI21_X1   g1042(.A1(new_n1302_), .A2(new_n1305_), .B(\shift[4] ), .ZN(new_n1306_));
  AOI21_X1   g1043(.A1(new_n1120_), .A2(new_n1121_), .B(new_n266_), .ZN(new_n1307_));
  OAI21_X1   g1044(.A1(new_n358_), .A2(new_n361_), .B(new_n276_), .ZN(new_n1308_));
  OAI21_X1   g1045(.A1(new_n319_), .A2(new_n322_), .B(\shift[3] ), .ZN(new_n1309_));
  AOI21_X1   g1046(.A1(new_n1308_), .A2(new_n1309_), .B(\shift[2] ), .ZN(new_n1310_));
  OAI21_X1   g1047(.A1(new_n1307_), .A2(new_n1310_), .B(new_n301_), .ZN(new_n1311_));
  AOI21_X1   g1048(.A1(new_n1306_), .A2(new_n1311_), .B(new_n265_), .ZN(new_n1312_));
  AOI21_X1   g1049(.A1(new_n1126_), .A2(new_n1127_), .B(new_n266_), .ZN(new_n1313_));
  OAI21_X1   g1050(.A1(new_n389_), .A2(new_n392_), .B(new_n276_), .ZN(new_n1314_));
  OAI21_X1   g1051(.A1(new_n351_), .A2(new_n354_), .B(\shift[3] ), .ZN(new_n1315_));
  AOI21_X1   g1052(.A1(new_n1314_), .A2(new_n1315_), .B(\shift[2] ), .ZN(new_n1316_));
  OAI21_X1   g1053(.A1(new_n1313_), .A2(new_n1316_), .B(\shift[4] ), .ZN(new_n1317_));
  AOI21_X1   g1054(.A1(new_n1131_), .A2(new_n1132_), .B(new_n266_), .ZN(new_n1318_));
  OAI21_X1   g1055(.A1(new_n422_), .A2(new_n425_), .B(new_n276_), .ZN(new_n1319_));
  OAI21_X1   g1056(.A1(new_n382_), .A2(new_n385_), .B(\shift[3] ), .ZN(new_n1320_));
  AOI21_X1   g1057(.A1(new_n1319_), .A2(new_n1320_), .B(\shift[2] ), .ZN(new_n1321_));
  OAI21_X1   g1058(.A1(new_n1318_), .A2(new_n1321_), .B(new_n301_), .ZN(new_n1322_));
  AOI21_X1   g1059(.A1(new_n1317_), .A2(new_n1322_), .B(\shift[5] ), .ZN(new_n1323_));
  OAI21_X1   g1060(.A1(new_n1312_), .A2(new_n1323_), .B(new_n264_), .ZN(new_n1324_));
  AOI21_X1   g1061(.A1(new_n1138_), .A2(new_n1139_), .B(new_n266_), .ZN(new_n1325_));
  OAI21_X1   g1062(.A1(new_n520_), .A2(new_n523_), .B(new_n276_), .ZN(new_n1326_));
  OAI21_X1   g1063(.A1(new_n478_), .A2(new_n481_), .B(\shift[3] ), .ZN(new_n1327_));
  AOI21_X1   g1064(.A1(new_n1326_), .A2(new_n1327_), .B(\shift[2] ), .ZN(new_n1328_));
  OAI21_X1   g1065(.A1(new_n1325_), .A2(new_n1328_), .B(\shift[4] ), .ZN(new_n1329_));
  AOI21_X1   g1066(.A1(new_n1143_), .A2(new_n1144_), .B(new_n266_), .ZN(new_n1330_));
  OAI21_X1   g1067(.A1(new_n294_), .A2(new_n297_), .B(new_n276_), .ZN(new_n1331_));
  OAI21_X1   g1068(.A1(new_n513_), .A2(new_n516_), .B(\shift[3] ), .ZN(new_n1332_));
  AOI21_X1   g1069(.A1(new_n1331_), .A2(new_n1332_), .B(\shift[2] ), .ZN(new_n1333_));
  OAI21_X1   g1070(.A1(new_n1330_), .A2(new_n1333_), .B(new_n301_), .ZN(new_n1334_));
  AOI21_X1   g1071(.A1(new_n1329_), .A2(new_n1334_), .B(\shift[5] ), .ZN(new_n1335_));
  AOI21_X1   g1072(.A1(new_n1149_), .A2(new_n1150_), .B(new_n266_), .ZN(new_n1336_));
  OAI21_X1   g1073(.A1(new_n487_), .A2(new_n492_), .B(new_n276_), .ZN(new_n1337_));
  OAI21_X1   g1074(.A1(new_n446_), .A2(new_n449_), .B(\shift[3] ), .ZN(new_n1338_));
  AOI21_X1   g1075(.A1(new_n1337_), .A2(new_n1338_), .B(\shift[2] ), .ZN(new_n1339_));
  OAI21_X1   g1076(.A1(new_n1339_), .A2(new_n1336_), .B(new_n301_), .ZN(new_n1340_));
  AOI21_X1   g1077(.A1(new_n1154_), .A2(new_n1155_), .B(new_n266_), .ZN(new_n1341_));
  OAI21_X1   g1078(.A1(new_n453_), .A2(new_n456_), .B(new_n276_), .ZN(new_n1342_));
  OAI21_X1   g1079(.A1(new_n415_), .A2(new_n418_), .B(\shift[3] ), .ZN(new_n1343_));
  AOI21_X1   g1080(.A1(new_n1342_), .A2(new_n1343_), .B(\shift[2] ), .ZN(new_n1344_));
  OAI21_X1   g1081(.A1(new_n1341_), .A2(new_n1344_), .B(\shift[4] ), .ZN(new_n1345_));
  AOI21_X1   g1082(.A1(new_n1340_), .A2(new_n1345_), .B(new_n265_), .ZN(new_n1346_));
  OAI21_X1   g1083(.A1(new_n1335_), .A2(new_n1346_), .B(\shift[6] ), .ZN(new_n1347_));
  NAND2_X1   g1084(.A1(new_n1324_), .A2(new_n1347_), .ZN(\result[8] ));
  AOI21_X1   g1085(.A1(new_n1162_), .A2(new_n1163_), .B(new_n266_), .ZN(new_n1349_));
  OAI21_X1   g1086(.A1(new_n585_), .A2(new_n588_), .B(new_n276_), .ZN(new_n1350_));
  OAI21_X1   g1087(.A1(new_n547_), .A2(new_n550_), .B(\shift[3] ), .ZN(new_n1351_));
  AOI21_X1   g1088(.A1(new_n1350_), .A2(new_n1351_), .B(\shift[2] ), .ZN(new_n1352_));
  OAI21_X1   g1089(.A1(new_n1352_), .A2(new_n1349_), .B(\shift[4] ), .ZN(new_n1353_));
  AOI21_X1   g1090(.A1(new_n1167_), .A2(new_n1168_), .B(new_n266_), .ZN(new_n1354_));
  OAI21_X1   g1091(.A1(new_n617_), .A2(new_n620_), .B(new_n276_), .ZN(new_n1355_));
  OAI21_X1   g1092(.A1(new_n581_), .A2(new_n578_), .B(\shift[3] ), .ZN(new_n1356_));
  AOI21_X1   g1093(.A1(new_n1356_), .A2(new_n1355_), .B(\shift[2] ), .ZN(new_n1357_));
  OAI21_X1   g1094(.A1(new_n1354_), .A2(new_n1357_), .B(new_n301_), .ZN(new_n1358_));
  AOI21_X1   g1095(.A1(new_n1353_), .A2(new_n1358_), .B(new_n265_), .ZN(new_n1359_));
  AOI21_X1   g1096(.A1(new_n1173_), .A2(new_n1174_), .B(new_n266_), .ZN(new_n1360_));
  OAI21_X1   g1097(.A1(new_n648_), .A2(new_n651_), .B(new_n276_), .ZN(new_n1361_));
  OAI21_X1   g1098(.A1(new_n613_), .A2(new_n610_), .B(\shift[3] ), .ZN(new_n1362_));
  AOI21_X1   g1099(.A1(new_n1362_), .A2(new_n1361_), .B(\shift[2] ), .ZN(new_n1363_));
  OAI21_X1   g1100(.A1(new_n1360_), .A2(new_n1363_), .B(\shift[4] ), .ZN(new_n1364_));
  AOI21_X1   g1101(.A1(new_n1178_), .A2(new_n1179_), .B(new_n266_), .ZN(new_n1365_));
  OAI21_X1   g1102(.A1(new_n717_), .A2(new_n714_), .B(new_n276_), .ZN(new_n1366_));
  OAI21_X1   g1103(.A1(new_n644_), .A2(new_n641_), .B(\shift[3] ), .ZN(new_n1367_));
  AOI21_X1   g1104(.A1(new_n1366_), .A2(new_n1367_), .B(\shift[2] ), .ZN(new_n1368_));
  OAI21_X1   g1105(.A1(new_n1365_), .A2(new_n1368_), .B(new_n301_), .ZN(new_n1369_));
  AOI21_X1   g1106(.A1(new_n1369_), .A2(new_n1364_), .B(\shift[5] ), .ZN(new_n1370_));
  OAI21_X1   g1107(.A1(new_n1370_), .A2(new_n1359_), .B(new_n264_), .ZN(new_n1371_));
  AOI21_X1   g1108(.A1(new_n1185_), .A2(new_n1186_), .B(new_n266_), .ZN(new_n1372_));
  OAI21_X1   g1109(.A1(new_n682_), .A2(new_n685_), .B(new_n276_), .ZN(new_n1373_));
  OAI21_X1   g1110(.A1(new_n742_), .A2(new_n739_), .B(\shift[3] ), .ZN(new_n1374_));
  AOI21_X1   g1111(.A1(new_n1373_), .A2(new_n1374_), .B(\shift[2] ), .ZN(new_n1375_));
  OAI21_X1   g1112(.A1(new_n1375_), .A2(new_n1372_), .B(\shift[4] ), .ZN(new_n1376_));
  AOI21_X1   g1113(.A1(new_n1190_), .A2(new_n1191_), .B(new_n266_), .ZN(new_n1377_));
  OAI21_X1   g1114(.A1(new_n554_), .A2(new_n557_), .B(new_n276_), .ZN(new_n1378_));
  OAI21_X1   g1115(.A1(new_n678_), .A2(new_n675_), .B(\shift[3] ), .ZN(new_n1379_));
  AOI21_X1   g1116(.A1(new_n1378_), .A2(new_n1379_), .B(\shift[2] ), .ZN(new_n1380_));
  OAI21_X1   g1117(.A1(new_n1377_), .A2(new_n1380_), .B(new_n301_), .ZN(new_n1381_));
  AOI21_X1   g1118(.A1(new_n1381_), .A2(new_n1376_), .B(\shift[5] ), .ZN(new_n1382_));
  AOI21_X1   g1119(.A1(new_n1197_), .A2(new_n1196_), .B(new_n266_), .ZN(new_n1383_));
  OAI21_X1   g1120(.A1(new_n746_), .A2(new_n749_), .B(new_n276_), .ZN(new_n1384_));
  OAI21_X1   g1121(.A1(new_n774_), .A2(new_n771_), .B(\shift[3] ), .ZN(new_n1385_));
  AOI21_X1   g1122(.A1(new_n1385_), .A2(new_n1384_), .B(\shift[2] ), .ZN(new_n1386_));
  OAI21_X1   g1123(.A1(new_n1383_), .A2(new_n1386_), .B(new_n301_), .ZN(new_n1387_));
  AOI21_X1   g1124(.A1(new_n1201_), .A2(new_n1202_), .B(new_n266_), .ZN(new_n1388_));
  OAI21_X1   g1125(.A1(new_n781_), .A2(new_n778_), .B(new_n276_), .ZN(new_n1389_));
  OAI21_X1   g1126(.A1(new_n710_), .A2(new_n707_), .B(\shift[3] ), .ZN(new_n1390_));
  AOI21_X1   g1127(.A1(new_n1389_), .A2(new_n1390_), .B(\shift[2] ), .ZN(new_n1391_));
  OAI21_X1   g1128(.A1(new_n1388_), .A2(new_n1391_), .B(\shift[4] ), .ZN(new_n1392_));
  AOI21_X1   g1129(.A1(new_n1392_), .A2(new_n1387_), .B(new_n265_), .ZN(new_n1393_));
  OAI21_X1   g1130(.A1(new_n1382_), .A2(new_n1393_), .B(\shift[6] ), .ZN(new_n1394_));
  NAND2_X1   g1131(.A1(new_n1371_), .A2(new_n1394_), .ZN(\result[9] ));
  AOI21_X1   g1132(.A1(new_n1209_), .A2(new_n1210_), .B(new_n266_), .ZN(new_n1396_));
  OAI21_X1   g1133(.A1(new_n813_), .A2(new_n814_), .B(new_n276_), .ZN(new_n1397_));
  OAI21_X1   g1134(.A1(new_n795_), .A2(new_n796_), .B(\shift[3] ), .ZN(new_n1398_));
  AOI21_X1   g1135(.A1(new_n1397_), .A2(new_n1398_), .B(\shift[2] ), .ZN(new_n1399_));
  OAI21_X1   g1136(.A1(new_n1396_), .A2(new_n1399_), .B(\shift[4] ), .ZN(new_n1400_));
  AOI21_X1   g1137(.A1(new_n1214_), .A2(new_n1215_), .B(new_n266_), .ZN(new_n1401_));
  OAI21_X1   g1138(.A1(new_n829_), .A2(new_n830_), .B(new_n276_), .ZN(new_n1402_));
  OAI21_X1   g1139(.A1(new_n810_), .A2(new_n811_), .B(\shift[3] ), .ZN(new_n1403_));
  AOI21_X1   g1140(.A1(new_n1402_), .A2(new_n1403_), .B(\shift[2] ), .ZN(new_n1404_));
  OAI21_X1   g1141(.A1(new_n1401_), .A2(new_n1404_), .B(new_n301_), .ZN(new_n1405_));
  AOI21_X1   g1142(.A1(new_n1400_), .A2(new_n1405_), .B(new_n265_), .ZN(new_n1406_));
  AOI21_X1   g1143(.A1(new_n1220_), .A2(new_n1221_), .B(new_n266_), .ZN(new_n1407_));
  OAI21_X1   g1144(.A1(new_n844_), .A2(new_n845_), .B(new_n276_), .ZN(new_n1408_));
  OAI21_X1   g1145(.A1(new_n826_), .A2(new_n827_), .B(\shift[3] ), .ZN(new_n1409_));
  AOI21_X1   g1146(.A1(new_n1408_), .A2(new_n1409_), .B(\shift[2] ), .ZN(new_n1410_));
  OAI21_X1   g1147(.A1(new_n1407_), .A2(new_n1410_), .B(\shift[4] ), .ZN(new_n1411_));
  AOI21_X1   g1148(.A1(new_n1225_), .A2(new_n1226_), .B(new_n266_), .ZN(new_n1412_));
  OAI21_X1   g1149(.A1(new_n878_), .A2(new_n879_), .B(new_n276_), .ZN(new_n1413_));
  OAI21_X1   g1150(.A1(new_n841_), .A2(new_n842_), .B(\shift[3] ), .ZN(new_n1414_));
  AOI21_X1   g1151(.A1(new_n1413_), .A2(new_n1414_), .B(\shift[2] ), .ZN(new_n1415_));
  OAI21_X1   g1152(.A1(new_n1412_), .A2(new_n1415_), .B(new_n301_), .ZN(new_n1416_));
  AOI21_X1   g1153(.A1(new_n1411_), .A2(new_n1416_), .B(\shift[5] ), .ZN(new_n1417_));
  OAI21_X1   g1154(.A1(new_n1406_), .A2(new_n1417_), .B(new_n264_), .ZN(new_n1418_));
  AOI21_X1   g1155(.A1(new_n1232_), .A2(new_n1233_), .B(new_n266_), .ZN(new_n1419_));
  OAI21_X1   g1156(.A1(new_n863_), .A2(new_n864_), .B(new_n276_), .ZN(new_n1420_));
  OAI21_X1   g1157(.A1(new_n893_), .A2(new_n894_), .B(\shift[3] ), .ZN(new_n1421_));
  AOI21_X1   g1158(.A1(new_n1420_), .A2(new_n1421_), .B(\shift[2] ), .ZN(new_n1422_));
  OAI21_X1   g1159(.A1(new_n1419_), .A2(new_n1422_), .B(\shift[4] ), .ZN(new_n1423_));
  AOI21_X1   g1160(.A1(new_n1237_), .A2(new_n1238_), .B(new_n266_), .ZN(new_n1424_));
  OAI21_X1   g1161(.A1(new_n798_), .A2(new_n799_), .B(new_n276_), .ZN(new_n1425_));
  OAI21_X1   g1162(.A1(new_n860_), .A2(new_n861_), .B(\shift[3] ), .ZN(new_n1426_));
  AOI21_X1   g1163(.A1(new_n1425_), .A2(new_n1426_), .B(\shift[2] ), .ZN(new_n1427_));
  OAI21_X1   g1164(.A1(new_n1424_), .A2(new_n1427_), .B(new_n301_), .ZN(new_n1428_));
  AOI21_X1   g1165(.A1(new_n1423_), .A2(new_n1428_), .B(\shift[5] ), .ZN(new_n1429_));
  AOI21_X1   g1166(.A1(new_n1243_), .A2(new_n1244_), .B(new_n266_), .ZN(new_n1430_));
  OAI21_X1   g1167(.A1(new_n898_), .A2(new_n899_), .B(new_n276_), .ZN(new_n1431_));
  OAI21_X1   g1168(.A1(new_n910_), .A2(new_n911_), .B(\shift[3] ), .ZN(new_n1432_));
  AOI21_X1   g1169(.A1(new_n1431_), .A2(new_n1432_), .B(\shift[2] ), .ZN(new_n1433_));
  OAI21_X1   g1170(.A1(new_n1430_), .A2(new_n1433_), .B(new_n301_), .ZN(new_n1434_));
  AOI21_X1   g1171(.A1(new_n1248_), .A2(new_n1249_), .B(new_n266_), .ZN(new_n1435_));
  OAI21_X1   g1172(.A1(new_n913_), .A2(new_n914_), .B(new_n276_), .ZN(new_n1436_));
  OAI21_X1   g1173(.A1(new_n875_), .A2(new_n876_), .B(\shift[3] ), .ZN(new_n1437_));
  AOI21_X1   g1174(.A1(new_n1436_), .A2(new_n1437_), .B(\shift[2] ), .ZN(new_n1438_));
  OAI21_X1   g1175(.A1(new_n1435_), .A2(new_n1438_), .B(\shift[4] ), .ZN(new_n1439_));
  AOI21_X1   g1176(.A1(new_n1434_), .A2(new_n1439_), .B(new_n265_), .ZN(new_n1440_));
  OAI21_X1   g1177(.A1(new_n1429_), .A2(new_n1440_), .B(\shift[6] ), .ZN(new_n1441_));
  NAND2_X1   g1178(.A1(new_n1418_), .A2(new_n1441_), .ZN(\result[10] ));
  AOI21_X1   g1179(.A1(new_n1256_), .A2(new_n1257_), .B(new_n266_), .ZN(new_n1443_));
  OAI21_X1   g1180(.A1(new_n957_), .A2(new_n960_), .B(new_n276_), .ZN(new_n1444_));
  OAI21_X1   g1181(.A1(new_n996_), .A2(new_n995_), .B(\shift[3] ), .ZN(new_n1445_));
  AOI21_X1   g1182(.A1(new_n1445_), .A2(new_n1444_), .B(\shift[2] ), .ZN(new_n1446_));
  OAI21_X1   g1183(.A1(new_n1443_), .A2(new_n1446_), .B(\shift[4] ), .ZN(new_n1447_));
  AOI21_X1   g1184(.A1(new_n1261_), .A2(new_n1262_), .B(new_n266_), .ZN(new_n1448_));
  OAI21_X1   g1185(.A1(new_n937_), .A2(new_n936_), .B(new_n276_), .ZN(new_n1449_));
  OAI21_X1   g1186(.A1(new_n954_), .A2(new_n951_), .B(\shift[3] ), .ZN(new_n1450_));
  AOI21_X1   g1187(.A1(new_n1449_), .A2(new_n1450_), .B(\shift[2] ), .ZN(new_n1451_));
  OAI21_X1   g1188(.A1(new_n1448_), .A2(new_n1451_), .B(new_n301_), .ZN(new_n1452_));
  AOI21_X1   g1189(.A1(new_n1447_), .A2(new_n1452_), .B(new_n265_), .ZN(new_n1453_));
  AOI21_X1   g1190(.A1(new_n1267_), .A2(new_n1268_), .B(new_n266_), .ZN(new_n1454_));
  OAI21_X1   g1191(.A1(new_n983_), .A2(new_n982_), .B(new_n276_), .ZN(new_n1455_));
  OAI21_X1   g1192(.A1(new_n933_), .A2(new_n932_), .B(\shift[3] ), .ZN(new_n1456_));
  AOI21_X1   g1193(.A1(new_n1455_), .A2(new_n1456_), .B(\shift[2] ), .ZN(new_n1457_));
  OAI21_X1   g1194(.A1(new_n1454_), .A2(new_n1457_), .B(\shift[4] ), .ZN(new_n1458_));
  AOI21_X1   g1195(.A1(new_n1272_), .A2(new_n1273_), .B(new_n266_), .ZN(new_n1459_));
  OAI21_X1   g1196(.A1(new_n1079_), .A2(new_n1076_), .B(new_n276_), .ZN(new_n1460_));
  OAI21_X1   g1197(.A1(new_n979_), .A2(new_n976_), .B(\shift[3] ), .ZN(new_n1461_));
  AOI21_X1   g1198(.A1(new_n1460_), .A2(new_n1461_), .B(\shift[2] ), .ZN(new_n1462_));
  OAI21_X1   g1199(.A1(new_n1459_), .A2(new_n1462_), .B(new_n301_), .ZN(new_n1463_));
  AOI21_X1   g1200(.A1(new_n1458_), .A2(new_n1463_), .B(\shift[5] ), .ZN(new_n1464_));
  OAI21_X1   g1201(.A1(new_n1453_), .A2(new_n1464_), .B(new_n264_), .ZN(new_n1465_));
  OAI21_X1   g1202(.A1(new_n1055_), .A2(new_n1054_), .B(new_n276_), .ZN(new_n1466_));
  OAI21_X1   g1203(.A1(new_n1020_), .A2(new_n1023_), .B(\shift[3] ), .ZN(new_n1467_));
  AOI21_X1   g1204(.A1(new_n1466_), .A2(new_n1467_), .B(\shift[2] ), .ZN(new_n1468_));
  AOI21_X1   g1205(.A1(new_n1280_), .A2(new_n1279_), .B(new_n266_), .ZN(new_n1469_));
  OAI21_X1   g1206(.A1(new_n1468_), .A2(new_n1469_), .B(\shift[4] ), .ZN(new_n1470_));
  AOI21_X1   g1207(.A1(new_n1284_), .A2(new_n1285_), .B(new_n266_), .ZN(new_n1471_));
  OAI21_X1   g1208(.A1(new_n1000_), .A2(new_n999_), .B(new_n276_), .ZN(new_n1472_));
  OAI21_X1   g1209(.A1(new_n1051_), .A2(new_n1048_), .B(\shift[3] ), .ZN(new_n1473_));
  AOI21_X1   g1210(.A1(new_n1472_), .A2(new_n1473_), .B(\shift[2] ), .ZN(new_n1474_));
  OAI21_X1   g1211(.A1(new_n1471_), .A2(new_n1474_), .B(new_n301_), .ZN(new_n1475_));
  AOI21_X1   g1212(.A1(new_n1475_), .A2(new_n1470_), .B(\shift[5] ), .ZN(new_n1476_));
  AOI21_X1   g1213(.A1(new_n1291_), .A2(new_n1290_), .B(new_n266_), .ZN(new_n1477_));
  OAI21_X1   g1214(.A1(new_n1026_), .A2(new_n1029_), .B(new_n276_), .ZN(new_n1478_));
  OAI21_X1   g1215(.A1(new_n1097_), .A2(new_n1100_), .B(\shift[3] ), .ZN(new_n1479_));
  AOI21_X1   g1216(.A1(new_n1478_), .A2(new_n1479_), .B(\shift[2] ), .ZN(new_n1480_));
  OAI21_X1   g1217(.A1(new_n1480_), .A2(new_n1477_), .B(new_n301_), .ZN(new_n1481_));
  AOI21_X1   g1218(.A1(new_n1295_), .A2(new_n1296_), .B(new_n266_), .ZN(new_n1482_));
  OAI21_X1   g1219(.A1(new_n1104_), .A2(new_n1107_), .B(new_n276_), .ZN(new_n1483_));
  OAI21_X1   g1220(.A1(new_n1073_), .A2(new_n1070_), .B(\shift[3] ), .ZN(new_n1484_));
  AOI21_X1   g1221(.A1(new_n1483_), .A2(new_n1484_), .B(\shift[2] ), .ZN(new_n1485_));
  OAI21_X1   g1222(.A1(new_n1482_), .A2(new_n1485_), .B(\shift[4] ), .ZN(new_n1486_));
  AOI21_X1   g1223(.A1(new_n1486_), .A2(new_n1481_), .B(new_n265_), .ZN(new_n1487_));
  OAI21_X1   g1224(.A1(new_n1487_), .A2(new_n1476_), .B(\shift[6] ), .ZN(new_n1488_));
  NAND2_X1   g1225(.A1(new_n1465_), .A2(new_n1488_), .ZN(\result[11] ));
  AOI21_X1   g1226(.A1(new_n1303_), .A2(new_n1304_), .B(new_n266_), .ZN(new_n1490_));
  AOI21_X1   g1227(.A1(new_n308_), .A2(new_n315_), .B(\shift[2] ), .ZN(new_n1491_));
  OAI21_X1   g1228(.A1(new_n1490_), .A2(new_n1491_), .B(\shift[4] ), .ZN(new_n1492_));
  AOI21_X1   g1229(.A1(new_n1308_), .A2(new_n1309_), .B(new_n266_), .ZN(new_n1493_));
  AOI21_X1   g1230(.A1(new_n340_), .A2(new_n347_), .B(\shift[2] ), .ZN(new_n1494_));
  OAI21_X1   g1231(.A1(new_n1493_), .A2(new_n1494_), .B(new_n301_), .ZN(new_n1495_));
  AOI21_X1   g1232(.A1(new_n1492_), .A2(new_n1495_), .B(new_n265_), .ZN(new_n1496_));
  AOI21_X1   g1233(.A1(new_n1314_), .A2(new_n1315_), .B(new_n266_), .ZN(new_n1497_));
  AOI21_X1   g1234(.A1(new_n371_), .A2(new_n378_), .B(\shift[2] ), .ZN(new_n1498_));
  OAI21_X1   g1235(.A1(new_n1497_), .A2(new_n1498_), .B(\shift[4] ), .ZN(new_n1499_));
  AOI21_X1   g1236(.A1(new_n1319_), .A2(new_n1320_), .B(new_n266_), .ZN(new_n1500_));
  AOI21_X1   g1237(.A1(new_n404_), .A2(new_n411_), .B(\shift[2] ), .ZN(new_n1501_));
  OAI21_X1   g1238(.A1(new_n1500_), .A2(new_n1501_), .B(new_n301_), .ZN(new_n1502_));
  AOI21_X1   g1239(.A1(new_n1499_), .A2(new_n1502_), .B(\shift[5] ), .ZN(new_n1503_));
  OAI21_X1   g1240(.A1(new_n1496_), .A2(new_n1503_), .B(new_n264_), .ZN(new_n1504_));
  AOI21_X1   g1241(.A1(new_n1326_), .A2(new_n1327_), .B(new_n266_), .ZN(new_n1505_));
  AOI21_X1   g1242(.A1(new_n502_), .A2(new_n509_), .B(\shift[2] ), .ZN(new_n1506_));
  OAI21_X1   g1243(.A1(new_n1505_), .A2(new_n1506_), .B(\shift[4] ), .ZN(new_n1507_));
  AOI21_X1   g1244(.A1(new_n1331_), .A2(new_n1332_), .B(new_n266_), .ZN(new_n1508_));
  AOI21_X1   g1245(.A1(new_n275_), .A2(new_n283_), .B(\shift[2] ), .ZN(new_n1509_));
  OAI21_X1   g1246(.A1(new_n1508_), .A2(new_n1509_), .B(new_n301_), .ZN(new_n1510_));
  AOI21_X1   g1247(.A1(new_n1507_), .A2(new_n1510_), .B(\shift[5] ), .ZN(new_n1511_));
  AOI21_X1   g1248(.A1(new_n1337_), .A2(new_n1338_), .B(new_n266_), .ZN(new_n1512_));
  AOI21_X1   g1249(.A1(new_n467_), .A2(new_n474_), .B(\shift[2] ), .ZN(new_n1513_));
  OAI21_X1   g1250(.A1(new_n1512_), .A2(new_n1513_), .B(new_n301_), .ZN(new_n1514_));
  AOI21_X1   g1251(.A1(new_n1342_), .A2(new_n1343_), .B(new_n266_), .ZN(new_n1515_));
  AOI21_X1   g1252(.A1(new_n435_), .A2(new_n442_), .B(\shift[2] ), .ZN(new_n1516_));
  OAI21_X1   g1253(.A1(new_n1515_), .A2(new_n1516_), .B(\shift[4] ), .ZN(new_n1517_));
  AOI21_X1   g1254(.A1(new_n1514_), .A2(new_n1517_), .B(new_n265_), .ZN(new_n1518_));
  OAI21_X1   g1255(.A1(new_n1511_), .A2(new_n1518_), .B(\shift[6] ), .ZN(new_n1519_));
  NAND2_X1   g1256(.A1(new_n1504_), .A2(new_n1519_), .ZN(\result[12] ));
  AOI21_X1   g1257(.A1(new_n1350_), .A2(new_n1351_), .B(new_n266_), .ZN(new_n1521_));
  AOI21_X1   g1258(.A1(new_n567_), .A2(new_n574_), .B(\shift[2] ), .ZN(new_n1522_));
  OAI21_X1   g1259(.A1(new_n1521_), .A2(new_n1522_), .B(\shift[4] ), .ZN(new_n1523_));
  AOI21_X1   g1260(.A1(new_n1356_), .A2(new_n1355_), .B(new_n266_), .ZN(new_n1524_));
  AOI21_X1   g1261(.A1(new_n599_), .A2(new_n606_), .B(\shift[2] ), .ZN(new_n1525_));
  OAI21_X1   g1262(.A1(new_n1525_), .A2(new_n1524_), .B(new_n301_), .ZN(new_n1526_));
  AOI21_X1   g1263(.A1(new_n1523_), .A2(new_n1526_), .B(new_n265_), .ZN(new_n1527_));
  AOI21_X1   g1264(.A1(new_n1362_), .A2(new_n1361_), .B(new_n266_), .ZN(new_n1528_));
  AOI21_X1   g1265(.A1(new_n630_), .A2(new_n637_), .B(\shift[2] ), .ZN(new_n1529_));
  OAI21_X1   g1266(.A1(new_n1529_), .A2(new_n1528_), .B(\shift[4] ), .ZN(new_n1530_));
  AOI21_X1   g1267(.A1(new_n1366_), .A2(new_n1367_), .B(new_n266_), .ZN(new_n1531_));
  AOI21_X1   g1268(.A1(new_n696_), .A2(new_n703_), .B(\shift[2] ), .ZN(new_n1532_));
  OAI21_X1   g1269(.A1(new_n1532_), .A2(new_n1531_), .B(new_n301_), .ZN(new_n1533_));
  AOI21_X1   g1270(.A1(new_n1533_), .A2(new_n1530_), .B(\shift[5] ), .ZN(new_n1534_));
  OAI21_X1   g1271(.A1(new_n1527_), .A2(new_n1534_), .B(new_n264_), .ZN(new_n1535_));
  AOI21_X1   g1272(.A1(new_n1373_), .A2(new_n1374_), .B(new_n266_), .ZN(new_n1536_));
  AOI21_X1   g1273(.A1(new_n664_), .A2(new_n671_), .B(\shift[2] ), .ZN(new_n1537_));
  OAI21_X1   g1274(.A1(new_n1536_), .A2(new_n1537_), .B(\shift[4] ), .ZN(new_n1538_));
  AOI21_X1   g1275(.A1(new_n1378_), .A2(new_n1379_), .B(new_n266_), .ZN(new_n1539_));
  AOI21_X1   g1276(.A1(new_n536_), .A2(new_n543_), .B(\shift[2] ), .ZN(new_n1540_));
  OAI21_X1   g1277(.A1(new_n1540_), .A2(new_n1539_), .B(new_n301_), .ZN(new_n1541_));
  AOI21_X1   g1278(.A1(new_n1538_), .A2(new_n1541_), .B(\shift[5] ), .ZN(new_n1542_));
  AOI21_X1   g1279(.A1(new_n1385_), .A2(new_n1384_), .B(new_n266_), .ZN(new_n1543_));
  AOI21_X1   g1280(.A1(new_n728_), .A2(new_n735_), .B(\shift[2] ), .ZN(new_n1544_));
  OAI21_X1   g1281(.A1(new_n1543_), .A2(new_n1544_), .B(new_n301_), .ZN(new_n1545_));
  AOI21_X1   g1282(.A1(new_n1389_), .A2(new_n1390_), .B(new_n266_), .ZN(new_n1546_));
  AOI21_X1   g1283(.A1(new_n760_), .A2(new_n767_), .B(\shift[2] ), .ZN(new_n1547_));
  OAI21_X1   g1284(.A1(new_n1547_), .A2(new_n1546_), .B(\shift[4] ), .ZN(new_n1548_));
  AOI21_X1   g1285(.A1(new_n1548_), .A2(new_n1545_), .B(new_n265_), .ZN(new_n1549_));
  OAI21_X1   g1286(.A1(new_n1542_), .A2(new_n1549_), .B(\shift[6] ), .ZN(new_n1550_));
  NAND2_X1   g1287(.A1(new_n1535_), .A2(new_n1550_), .ZN(\result[13] ));
  AOI21_X1   g1288(.A1(new_n1397_), .A2(new_n1398_), .B(new_n266_), .ZN(new_n1552_));
  AOI21_X1   g1289(.A1(new_n805_), .A2(new_n808_), .B(\shift[2] ), .ZN(new_n1553_));
  OAI21_X1   g1290(.A1(new_n1552_), .A2(new_n1553_), .B(\shift[4] ), .ZN(new_n1554_));
  AOI21_X1   g1291(.A1(new_n1402_), .A2(new_n1403_), .B(new_n266_), .ZN(new_n1555_));
  AOI21_X1   g1292(.A1(new_n821_), .A2(new_n824_), .B(\shift[2] ), .ZN(new_n1556_));
  OAI21_X1   g1293(.A1(new_n1555_), .A2(new_n1556_), .B(new_n301_), .ZN(new_n1557_));
  AOI21_X1   g1294(.A1(new_n1554_), .A2(new_n1557_), .B(new_n265_), .ZN(new_n1558_));
  AOI21_X1   g1295(.A1(new_n1408_), .A2(new_n1409_), .B(new_n266_), .ZN(new_n1559_));
  AOI21_X1   g1296(.A1(new_n836_), .A2(new_n839_), .B(\shift[2] ), .ZN(new_n1560_));
  OAI21_X1   g1297(.A1(new_n1559_), .A2(new_n1560_), .B(\shift[4] ), .ZN(new_n1561_));
  AOI21_X1   g1298(.A1(new_n1413_), .A2(new_n1414_), .B(new_n266_), .ZN(new_n1562_));
  AOI21_X1   g1299(.A1(new_n870_), .A2(new_n873_), .B(\shift[2] ), .ZN(new_n1563_));
  OAI21_X1   g1300(.A1(new_n1562_), .A2(new_n1563_), .B(new_n301_), .ZN(new_n1564_));
  AOI21_X1   g1301(.A1(new_n1561_), .A2(new_n1564_), .B(\shift[5] ), .ZN(new_n1565_));
  OAI21_X1   g1302(.A1(new_n1558_), .A2(new_n1565_), .B(new_n264_), .ZN(new_n1566_));
  AOI21_X1   g1303(.A1(new_n1420_), .A2(new_n1421_), .B(new_n266_), .ZN(new_n1567_));
  AOI21_X1   g1304(.A1(new_n855_), .A2(new_n858_), .B(\shift[2] ), .ZN(new_n1568_));
  OAI21_X1   g1305(.A1(new_n1567_), .A2(new_n1568_), .B(\shift[4] ), .ZN(new_n1569_));
  AOI21_X1   g1306(.A1(new_n1425_), .A2(new_n1426_), .B(new_n266_), .ZN(new_n1570_));
  AOI21_X1   g1307(.A1(new_n790_), .A2(new_n793_), .B(\shift[2] ), .ZN(new_n1571_));
  OAI21_X1   g1308(.A1(new_n1570_), .A2(new_n1571_), .B(new_n301_), .ZN(new_n1572_));
  AOI21_X1   g1309(.A1(new_n1569_), .A2(new_n1572_), .B(\shift[5] ), .ZN(new_n1573_));
  AOI21_X1   g1310(.A1(new_n1431_), .A2(new_n1432_), .B(new_n266_), .ZN(new_n1574_));
  AOI21_X1   g1311(.A1(new_n888_), .A2(new_n891_), .B(\shift[2] ), .ZN(new_n1575_));
  OAI21_X1   g1312(.A1(new_n1574_), .A2(new_n1575_), .B(new_n301_), .ZN(new_n1576_));
  AOI21_X1   g1313(.A1(new_n1436_), .A2(new_n1437_), .B(new_n266_), .ZN(new_n1577_));
  AOI21_X1   g1314(.A1(new_n905_), .A2(new_n908_), .B(\shift[2] ), .ZN(new_n1578_));
  OAI21_X1   g1315(.A1(new_n1577_), .A2(new_n1578_), .B(\shift[4] ), .ZN(new_n1579_));
  AOI21_X1   g1316(.A1(new_n1576_), .A2(new_n1579_), .B(new_n265_), .ZN(new_n1580_));
  OAI21_X1   g1317(.A1(new_n1573_), .A2(new_n1580_), .B(\shift[6] ), .ZN(new_n1581_));
  NAND2_X1   g1318(.A1(new_n1566_), .A2(new_n1581_), .ZN(\result[14] ));
  AOI21_X1   g1319(.A1(new_n1445_), .A2(new_n1444_), .B(new_n266_), .ZN(new_n1583_));
  AOI21_X1   g1320(.A1(new_n943_), .A2(new_n948_), .B(\shift[2] ), .ZN(new_n1584_));
  OAI21_X1   g1321(.A1(new_n1584_), .A2(new_n1583_), .B(\shift[4] ), .ZN(new_n1585_));
  AOI21_X1   g1322(.A1(new_n1449_), .A2(new_n1450_), .B(new_n266_), .ZN(new_n1586_));
  AOI21_X1   g1323(.A1(new_n925_), .A2(new_n929_), .B(\shift[2] ), .ZN(new_n1587_));
  OAI21_X1   g1324(.A1(new_n1587_), .A2(new_n1586_), .B(new_n301_), .ZN(new_n1588_));
  AOI21_X1   g1325(.A1(new_n1585_), .A2(new_n1588_), .B(new_n265_), .ZN(new_n1589_));
  AOI21_X1   g1326(.A1(new_n1455_), .A2(new_n1456_), .B(new_n266_), .ZN(new_n1590_));
  AOI21_X1   g1327(.A1(new_n969_), .A2(new_n973_), .B(\shift[2] ), .ZN(new_n1591_));
  OAI21_X1   g1328(.A1(new_n1590_), .A2(new_n1591_), .B(\shift[4] ), .ZN(new_n1592_));
  AOI21_X1   g1329(.A1(new_n1460_), .A2(new_n1461_), .B(new_n266_), .ZN(new_n1593_));
  AOI21_X1   g1330(.A1(new_n1063_), .A2(new_n1067_), .B(\shift[2] ), .ZN(new_n1594_));
  OAI21_X1   g1331(.A1(new_n1594_), .A2(new_n1593_), .B(new_n301_), .ZN(new_n1595_));
  AOI21_X1   g1332(.A1(new_n1592_), .A2(new_n1595_), .B(\shift[5] ), .ZN(new_n1596_));
  OAI21_X1   g1333(.A1(new_n1589_), .A2(new_n1596_), .B(new_n264_), .ZN(new_n1597_));
  AOI21_X1   g1334(.A1(new_n1466_), .A2(new_n1467_), .B(new_n266_), .ZN(new_n1598_));
  AOI21_X1   g1335(.A1(new_n1045_), .A2(new_n1038_), .B(\shift[2] ), .ZN(new_n1599_));
  OAI21_X1   g1336(.A1(new_n1598_), .A2(new_n1599_), .B(\shift[4] ), .ZN(new_n1600_));
  AOI21_X1   g1337(.A1(new_n1472_), .A2(new_n1473_), .B(new_n266_), .ZN(new_n1601_));
  AOI21_X1   g1338(.A1(new_n989_), .A2(new_n993_), .B(\shift[2] ), .ZN(new_n1602_));
  OAI21_X1   g1339(.A1(new_n1602_), .A2(new_n1601_), .B(new_n301_), .ZN(new_n1603_));
  AOI21_X1   g1340(.A1(new_n1603_), .A2(new_n1600_), .B(\shift[5] ), .ZN(new_n1604_));
  AOI21_X1   g1341(.A1(new_n1478_), .A2(new_n1479_), .B(new_n266_), .ZN(new_n1605_));
  AOI21_X1   g1342(.A1(new_n1011_), .A2(new_n1016_), .B(\shift[2] ), .ZN(new_n1606_));
  OAI21_X1   g1343(.A1(new_n1605_), .A2(new_n1606_), .B(new_n301_), .ZN(new_n1607_));
  AOI21_X1   g1344(.A1(new_n1483_), .A2(new_n1484_), .B(new_n266_), .ZN(new_n1608_));
  AOI21_X1   g1345(.A1(new_n1086_), .A2(new_n1093_), .B(\shift[2] ), .ZN(new_n1609_));
  OAI21_X1   g1346(.A1(new_n1609_), .A2(new_n1608_), .B(\shift[4] ), .ZN(new_n1610_));
  AOI21_X1   g1347(.A1(new_n1610_), .A2(new_n1607_), .B(new_n265_), .ZN(new_n1611_));
  OAI21_X1   g1348(.A1(new_n1604_), .A2(new_n1611_), .B(\shift[6] ), .ZN(new_n1612_));
  NAND2_X1   g1349(.A1(new_n1597_), .A2(new_n1612_), .ZN(\result[15] ));
  OAI21_X1   g1350(.A1(new_n316_), .A2(new_n331_), .B(\shift[4] ), .ZN(new_n1614_));
  OAI21_X1   g1351(.A1(new_n348_), .A2(new_n363_), .B(new_n301_), .ZN(new_n1615_));
  AOI21_X1   g1352(.A1(new_n1614_), .A2(new_n1615_), .B(new_n265_), .ZN(new_n1616_));
  OAI21_X1   g1353(.A1(new_n379_), .A2(new_n394_), .B(\shift[4] ), .ZN(new_n1617_));
  OAI21_X1   g1354(.A1(new_n412_), .A2(new_n427_), .B(new_n301_), .ZN(new_n1618_));
  AOI21_X1   g1355(.A1(new_n1617_), .A2(new_n1618_), .B(\shift[5] ), .ZN(new_n1619_));
  OAI21_X1   g1356(.A1(new_n1616_), .A2(new_n1619_), .B(new_n264_), .ZN(new_n1620_));
  NOR2_X1    g1357(.A1(new_n284_), .A2(new_n299_), .ZN(new_n1621_));
  NOR2_X1    g1358(.A1(new_n443_), .A2(new_n458_), .ZN(new_n1622_));
  OAI22_X1   g1359(.A1(new_n1621_), .A2(new_n851_), .B1(new_n1622_), .B2(new_n852_), .ZN(new_n1623_));
  OAI21_X1   g1360(.A1(new_n510_), .A2(new_n525_), .B(new_n722_), .ZN(new_n1624_));
  OAI21_X1   g1361(.A1(new_n494_), .A2(new_n475_), .B(new_n753_), .ZN(new_n1625_));
  NAND2_X1   g1362(.A1(new_n1624_), .A2(new_n1625_), .ZN(new_n1626_));
  OAI21_X1   g1363(.A1(new_n1623_), .A2(new_n1626_), .B(\shift[6] ), .ZN(new_n1627_));
  NAND2_X1   g1364(.A1(new_n1620_), .A2(new_n1627_), .ZN(\result[16] ));
  OAI21_X1   g1365(.A1(new_n575_), .A2(new_n590_), .B(\shift[4] ), .ZN(new_n1629_));
  OAI21_X1   g1366(.A1(new_n607_), .A2(new_n622_), .B(new_n301_), .ZN(new_n1630_));
  AOI21_X1   g1367(.A1(new_n1629_), .A2(new_n1630_), .B(new_n265_), .ZN(new_n1631_));
  OAI21_X1   g1368(.A1(new_n638_), .A2(new_n653_), .B(\shift[4] ), .ZN(new_n1632_));
  OAI21_X1   g1369(.A1(new_n704_), .A2(new_n719_), .B(new_n301_), .ZN(new_n1633_));
  AOI21_X1   g1370(.A1(new_n1633_), .A2(new_n1632_), .B(\shift[5] ), .ZN(new_n1634_));
  OAI21_X1   g1371(.A1(new_n1631_), .A2(new_n1634_), .B(new_n264_), .ZN(new_n1635_));
  OAI21_X1   g1372(.A1(new_n687_), .A2(new_n672_), .B(\shift[4] ), .ZN(new_n1636_));
  OAI21_X1   g1373(.A1(new_n559_), .A2(new_n544_), .B(new_n301_), .ZN(new_n1637_));
  AOI21_X1   g1374(.A1(new_n1637_), .A2(new_n1636_), .B(\shift[5] ), .ZN(new_n1638_));
  OAI21_X1   g1375(.A1(new_n736_), .A2(new_n751_), .B(new_n301_), .ZN(new_n1639_));
  OAI21_X1   g1376(.A1(new_n768_), .A2(new_n783_), .B(\shift[4] ), .ZN(new_n1640_));
  AOI21_X1   g1377(.A1(new_n1640_), .A2(new_n1639_), .B(new_n265_), .ZN(new_n1641_));
  OAI21_X1   g1378(.A1(new_n1638_), .A2(new_n1641_), .B(\shift[6] ), .ZN(new_n1642_));
  NAND2_X1   g1379(.A1(new_n1635_), .A2(new_n1642_), .ZN(\result[17] ));
  OAI21_X1   g1380(.A1(new_n809_), .A2(new_n816_), .B(\shift[4] ), .ZN(new_n1644_));
  OAI21_X1   g1381(.A1(new_n825_), .A2(new_n832_), .B(new_n301_), .ZN(new_n1645_));
  AOI21_X1   g1382(.A1(new_n1644_), .A2(new_n1645_), .B(new_n265_), .ZN(new_n1646_));
  OAI21_X1   g1383(.A1(new_n840_), .A2(new_n847_), .B(\shift[4] ), .ZN(new_n1647_));
  OAI21_X1   g1384(.A1(new_n874_), .A2(new_n881_), .B(new_n301_), .ZN(new_n1648_));
  AOI21_X1   g1385(.A1(new_n1647_), .A2(new_n1648_), .B(\shift[5] ), .ZN(new_n1649_));
  OAI21_X1   g1386(.A1(new_n1646_), .A2(new_n1649_), .B(new_n264_), .ZN(new_n1650_));
  OAI21_X1   g1387(.A1(new_n859_), .A2(new_n866_), .B(\shift[4] ), .ZN(new_n1651_));
  OAI21_X1   g1388(.A1(new_n794_), .A2(new_n801_), .B(new_n301_), .ZN(new_n1652_));
  AOI21_X1   g1389(.A1(new_n1651_), .A2(new_n1652_), .B(\shift[5] ), .ZN(new_n1653_));
  OAI21_X1   g1390(.A1(new_n892_), .A2(new_n901_), .B(new_n301_), .ZN(new_n1654_));
  OAI21_X1   g1391(.A1(new_n909_), .A2(new_n916_), .B(\shift[4] ), .ZN(new_n1655_));
  AOI21_X1   g1392(.A1(new_n1654_), .A2(new_n1655_), .B(new_n265_), .ZN(new_n1656_));
  OAI21_X1   g1393(.A1(new_n1653_), .A2(new_n1656_), .B(\shift[6] ), .ZN(new_n1657_));
  NAND2_X1   g1394(.A1(new_n1650_), .A2(new_n1657_), .ZN(\result[18] ));
  OAI21_X1   g1395(.A1(new_n930_), .A2(new_n939_), .B(new_n301_), .ZN(new_n1659_));
  OAI21_X1   g1396(.A1(new_n949_), .A2(new_n962_), .B(\shift[4] ), .ZN(new_n1660_));
  AOI21_X1   g1397(.A1(new_n1659_), .A2(new_n1660_), .B(new_n265_), .ZN(new_n1661_));
  OAI21_X1   g1398(.A1(new_n974_), .A2(new_n985_), .B(\shift[4] ), .ZN(new_n1662_));
  OAI21_X1   g1399(.A1(new_n1068_), .A2(new_n1081_), .B(new_n301_), .ZN(new_n1663_));
  AOI21_X1   g1400(.A1(new_n1662_), .A2(new_n1663_), .B(\shift[5] ), .ZN(new_n1664_));
  OAI21_X1   g1401(.A1(new_n1661_), .A2(new_n1664_), .B(new_n264_), .ZN(new_n1665_));
  OAI21_X1   g1402(.A1(new_n1057_), .A2(new_n1046_), .B(\shift[4] ), .ZN(new_n1666_));
  OAI21_X1   g1403(.A1(new_n994_), .A2(new_n1002_), .B(new_n301_), .ZN(new_n1667_));
  AOI21_X1   g1404(.A1(new_n1667_), .A2(new_n1666_), .B(\shift[5] ), .ZN(new_n1668_));
  OAI21_X1   g1405(.A1(new_n1031_), .A2(new_n1017_), .B(new_n301_), .ZN(new_n1669_));
  OAI21_X1   g1406(.A1(new_n1094_), .A2(new_n1109_), .B(\shift[4] ), .ZN(new_n1670_));
  AOI21_X1   g1407(.A1(new_n1670_), .A2(new_n1669_), .B(new_n265_), .ZN(new_n1671_));
  OAI21_X1   g1408(.A1(new_n1668_), .A2(new_n1671_), .B(\shift[6] ), .ZN(new_n1672_));
  NAND2_X1   g1409(.A1(new_n1665_), .A2(new_n1672_), .ZN(\result[19] ));
  OAI21_X1   g1410(.A1(new_n1119_), .A2(new_n1122_), .B(\shift[4] ), .ZN(new_n1674_));
  OAI21_X1   g1411(.A1(new_n1125_), .A2(new_n1128_), .B(new_n301_), .ZN(new_n1675_));
  AOI21_X1   g1412(.A1(new_n1674_), .A2(new_n1675_), .B(new_n265_), .ZN(new_n1676_));
  OAI21_X1   g1413(.A1(new_n1130_), .A2(new_n1133_), .B(\shift[4] ), .ZN(new_n1677_));
  OAI21_X1   g1414(.A1(new_n1153_), .A2(new_n1156_), .B(new_n301_), .ZN(new_n1678_));
  AOI21_X1   g1415(.A1(new_n1677_), .A2(new_n1678_), .B(\shift[5] ), .ZN(new_n1679_));
  OAI21_X1   g1416(.A1(new_n1676_), .A2(new_n1679_), .B(new_n264_), .ZN(new_n1680_));
  OAI21_X1   g1417(.A1(new_n1137_), .A2(new_n1140_), .B(\shift[5] ), .ZN(new_n1681_));
  OAI21_X1   g1418(.A1(new_n1114_), .A2(new_n1117_), .B(new_n265_), .ZN(new_n1682_));
  AOI21_X1   g1419(.A1(new_n1681_), .A2(new_n1682_), .B(\shift[4] ), .ZN(new_n1683_));
  OAI21_X1   g1420(.A1(new_n1142_), .A2(new_n1145_), .B(new_n265_), .ZN(new_n1684_));
  OAI21_X1   g1421(.A1(new_n1148_), .A2(new_n1151_), .B(\shift[5] ), .ZN(new_n1685_));
  AOI21_X1   g1422(.A1(new_n1684_), .A2(new_n1685_), .B(new_n301_), .ZN(new_n1686_));
  OAI21_X1   g1423(.A1(new_n1683_), .A2(new_n1686_), .B(\shift[6] ), .ZN(new_n1687_));
  NAND2_X1   g1424(.A1(new_n1680_), .A2(new_n1687_), .ZN(\result[20] ));
  OAI21_X1   g1425(.A1(new_n1166_), .A2(new_n1169_), .B(\shift[4] ), .ZN(new_n1689_));
  OAI21_X1   g1426(.A1(new_n1175_), .A2(new_n1172_), .B(new_n301_), .ZN(new_n1690_));
  AOI21_X1   g1427(.A1(new_n1689_), .A2(new_n1690_), .B(new_n265_), .ZN(new_n1691_));
  OAI21_X1   g1428(.A1(new_n1180_), .A2(new_n1177_), .B(\shift[4] ), .ZN(new_n1692_));
  OAI21_X1   g1429(.A1(new_n1203_), .A2(new_n1200_), .B(new_n301_), .ZN(new_n1693_));
  AOI21_X1   g1430(.A1(new_n1693_), .A2(new_n1692_), .B(\shift[5] ), .ZN(new_n1694_));
  OAI21_X1   g1431(.A1(new_n1691_), .A2(new_n1694_), .B(new_n264_), .ZN(new_n1695_));
  OAI21_X1   g1432(.A1(new_n1184_), .A2(new_n1187_), .B(\shift[5] ), .ZN(new_n1696_));
  OAI21_X1   g1433(.A1(new_n1161_), .A2(new_n1164_), .B(new_n265_), .ZN(new_n1697_));
  AOI21_X1   g1434(.A1(new_n1697_), .A2(new_n1696_), .B(\shift[4] ), .ZN(new_n1698_));
  OAI21_X1   g1435(.A1(new_n1189_), .A2(new_n1192_), .B(new_n265_), .ZN(new_n1699_));
  OAI21_X1   g1436(.A1(new_n1195_), .A2(new_n1198_), .B(\shift[5] ), .ZN(new_n1700_));
  AOI21_X1   g1437(.A1(new_n1699_), .A2(new_n1700_), .B(new_n301_), .ZN(new_n1701_));
  OAI21_X1   g1438(.A1(new_n1701_), .A2(new_n1698_), .B(\shift[6] ), .ZN(new_n1702_));
  NAND2_X1   g1439(.A1(new_n1695_), .A2(new_n1702_), .ZN(\result[21] ));
  OAI21_X1   g1440(.A1(new_n1213_), .A2(new_n1216_), .B(\shift[4] ), .ZN(new_n1704_));
  OAI21_X1   g1441(.A1(new_n1219_), .A2(new_n1222_), .B(new_n301_), .ZN(new_n1705_));
  AOI21_X1   g1442(.A1(new_n1704_), .A2(new_n1705_), .B(new_n265_), .ZN(new_n1706_));
  OAI21_X1   g1443(.A1(new_n1224_), .A2(new_n1227_), .B(\shift[4] ), .ZN(new_n1707_));
  OAI21_X1   g1444(.A1(new_n1247_), .A2(new_n1250_), .B(new_n301_), .ZN(new_n1708_));
  AOI21_X1   g1445(.A1(new_n1707_), .A2(new_n1708_), .B(\shift[5] ), .ZN(new_n1709_));
  OAI21_X1   g1446(.A1(new_n1706_), .A2(new_n1709_), .B(new_n264_), .ZN(new_n1710_));
  OAI21_X1   g1447(.A1(new_n1231_), .A2(new_n1234_), .B(\shift[5] ), .ZN(new_n1711_));
  OAI21_X1   g1448(.A1(new_n1208_), .A2(new_n1211_), .B(new_n265_), .ZN(new_n1712_));
  AOI21_X1   g1449(.A1(new_n1711_), .A2(new_n1712_), .B(\shift[4] ), .ZN(new_n1713_));
  OAI21_X1   g1450(.A1(new_n1236_), .A2(new_n1239_), .B(new_n265_), .ZN(new_n1714_));
  OAI21_X1   g1451(.A1(new_n1242_), .A2(new_n1245_), .B(\shift[5] ), .ZN(new_n1715_));
  AOI21_X1   g1452(.A1(new_n1714_), .A2(new_n1715_), .B(new_n301_), .ZN(new_n1716_));
  OAI21_X1   g1453(.A1(new_n1713_), .A2(new_n1716_), .B(\shift[6] ), .ZN(new_n1717_));
  NAND2_X1   g1454(.A1(new_n1710_), .A2(new_n1717_), .ZN(\result[22] ));
  OAI21_X1   g1455(.A1(new_n1297_), .A2(new_n1294_), .B(new_n657_), .ZN(new_n1719_));
  OAI21_X1   g1456(.A1(new_n1263_), .A2(new_n1260_), .B(new_n689_), .ZN(new_n1720_));
  NAND2_X1   g1457(.A1(new_n1719_), .A2(new_n1720_), .ZN(new_n1721_));
  INV_X1     g1458(.I(new_n722_), .ZN(new_n1722_));
  INV_X1     g1459(.I(new_n753_), .ZN(new_n1723_));
  NOR2_X1    g1460(.A1(new_n1266_), .A2(new_n1269_), .ZN(new_n1724_));
  NOR2_X1    g1461(.A1(new_n1274_), .A2(new_n1271_), .ZN(new_n1725_));
  OAI22_X1   g1462(.A1(new_n1724_), .A2(new_n1723_), .B1(new_n1725_), .B2(new_n1722_), .ZN(new_n1726_));
  OAI21_X1   g1463(.A1(new_n1726_), .A2(new_n1721_), .B(new_n264_), .ZN(new_n1727_));
  OAI21_X1   g1464(.A1(new_n1278_), .A2(new_n1281_), .B(new_n753_), .ZN(new_n1728_));
  OAI21_X1   g1465(.A1(new_n1286_), .A2(new_n1283_), .B(new_n722_), .ZN(new_n1729_));
  NAND2_X1   g1466(.A1(new_n1729_), .A2(new_n1728_), .ZN(new_n1730_));
  NOR2_X1    g1467(.A1(new_n1255_), .A2(new_n1258_), .ZN(new_n1731_));
  NOR2_X1    g1468(.A1(new_n1289_), .A2(new_n1292_), .ZN(new_n1732_));
  OAI22_X1   g1469(.A1(new_n1731_), .A2(new_n851_), .B1(new_n1732_), .B2(new_n852_), .ZN(new_n1733_));
  OAI21_X1   g1470(.A1(new_n1733_), .A2(new_n1730_), .B(\shift[6] ), .ZN(new_n1734_));
  NAND2_X1   g1471(.A1(new_n1727_), .A2(new_n1734_), .ZN(\result[23] ));
  NOR2_X1    g1472(.A1(new_n1307_), .A2(new_n1310_), .ZN(new_n1736_));
  NOR2_X1    g1473(.A1(new_n1341_), .A2(new_n1344_), .ZN(new_n1737_));
  OAI22_X1   g1474(.A1(new_n851_), .A2(new_n1737_), .B1(new_n1736_), .B2(new_n852_), .ZN(new_n1738_));
  NOR2_X1    g1475(.A1(new_n1313_), .A2(new_n1316_), .ZN(new_n1739_));
  NOR2_X1    g1476(.A1(new_n1318_), .A2(new_n1321_), .ZN(new_n1740_));
  OAI22_X1   g1477(.A1(new_n1722_), .A2(new_n1740_), .B1(new_n1739_), .B2(new_n1723_), .ZN(new_n1741_));
  OAI21_X1   g1478(.A1(new_n1738_), .A2(new_n1741_), .B(new_n264_), .ZN(new_n1742_));
  NOR2_X1    g1479(.A1(new_n1325_), .A2(new_n1328_), .ZN(new_n1743_));
  NOR2_X1    g1480(.A1(new_n1330_), .A2(new_n1333_), .ZN(new_n1744_));
  OAI22_X1   g1481(.A1(new_n1722_), .A2(new_n1744_), .B1(new_n1743_), .B2(new_n1723_), .ZN(new_n1745_));
  OAI21_X1   g1482(.A1(new_n1302_), .A2(new_n1305_), .B(new_n657_), .ZN(new_n1746_));
  OAI21_X1   g1483(.A1(new_n1339_), .A2(new_n1336_), .B(new_n689_), .ZN(new_n1747_));
  NAND2_X1   g1484(.A1(new_n1746_), .A2(new_n1747_), .ZN(new_n1748_));
  OAI21_X1   g1485(.A1(new_n1745_), .A2(new_n1748_), .B(\shift[6] ), .ZN(new_n1749_));
  NAND2_X1   g1486(.A1(new_n1742_), .A2(new_n1749_), .ZN(\result[24] ));
  NOR2_X1    g1487(.A1(new_n1354_), .A2(new_n1357_), .ZN(new_n1751_));
  NOR2_X1    g1488(.A1(new_n1388_), .A2(new_n1391_), .ZN(new_n1752_));
  OAI22_X1   g1489(.A1(new_n851_), .A2(new_n1752_), .B1(new_n1751_), .B2(new_n852_), .ZN(new_n1753_));
  OAI21_X1   g1490(.A1(new_n1365_), .A2(new_n1368_), .B(new_n722_), .ZN(new_n1754_));
  OAI21_X1   g1491(.A1(new_n1360_), .A2(new_n1363_), .B(new_n753_), .ZN(new_n1755_));
  NAND2_X1   g1492(.A1(new_n1754_), .A2(new_n1755_), .ZN(new_n1756_));
  OAI21_X1   g1493(.A1(new_n1753_), .A2(new_n1756_), .B(new_n264_), .ZN(new_n1757_));
  NOR2_X1    g1494(.A1(new_n1375_), .A2(new_n1372_), .ZN(new_n1758_));
  NOR2_X1    g1495(.A1(new_n1377_), .A2(new_n1380_), .ZN(new_n1759_));
  OAI22_X1   g1496(.A1(new_n1759_), .A2(new_n1722_), .B1(new_n1758_), .B2(new_n1723_), .ZN(new_n1760_));
  NOR2_X1    g1497(.A1(new_n1352_), .A2(new_n1349_), .ZN(new_n1761_));
  NOR2_X1    g1498(.A1(new_n1383_), .A2(new_n1386_), .ZN(new_n1762_));
  OAI22_X1   g1499(.A1(new_n1761_), .A2(new_n851_), .B1(new_n1762_), .B2(new_n852_), .ZN(new_n1763_));
  OAI21_X1   g1500(.A1(new_n1760_), .A2(new_n1763_), .B(\shift[6] ), .ZN(new_n1764_));
  NAND2_X1   g1501(.A1(new_n1764_), .A2(new_n1757_), .ZN(\result[25] ));
  OAI21_X1   g1502(.A1(new_n1401_), .A2(new_n1404_), .B(\shift[4] ), .ZN(new_n1766_));
  OAI21_X1   g1503(.A1(new_n1407_), .A2(new_n1410_), .B(new_n301_), .ZN(new_n1767_));
  AOI21_X1   g1504(.A1(new_n1766_), .A2(new_n1767_), .B(new_n265_), .ZN(new_n1768_));
  OAI21_X1   g1505(.A1(new_n1412_), .A2(new_n1415_), .B(\shift[4] ), .ZN(new_n1769_));
  OAI21_X1   g1506(.A1(new_n1435_), .A2(new_n1438_), .B(new_n301_), .ZN(new_n1770_));
  AOI21_X1   g1507(.A1(new_n1769_), .A2(new_n1770_), .B(\shift[5] ), .ZN(new_n1771_));
  OAI21_X1   g1508(.A1(new_n1768_), .A2(new_n1771_), .B(new_n264_), .ZN(new_n1772_));
  NOR2_X1    g1509(.A1(new_n1419_), .A2(new_n1422_), .ZN(new_n1773_));
  NOR2_X1    g1510(.A1(new_n1424_), .A2(new_n1427_), .ZN(new_n1774_));
  OAI22_X1   g1511(.A1(new_n1722_), .A2(new_n1774_), .B1(new_n1773_), .B2(new_n1723_), .ZN(new_n1775_));
  OAI21_X1   g1512(.A1(new_n1396_), .A2(new_n1399_), .B(new_n657_), .ZN(new_n1776_));
  OAI21_X1   g1513(.A1(new_n1430_), .A2(new_n1433_), .B(new_n689_), .ZN(new_n1777_));
  NAND2_X1   g1514(.A1(new_n1776_), .A2(new_n1777_), .ZN(new_n1778_));
  OAI21_X1   g1515(.A1(new_n1775_), .A2(new_n1778_), .B(\shift[6] ), .ZN(new_n1779_));
  NAND2_X1   g1516(.A1(new_n1772_), .A2(new_n1779_), .ZN(\result[26] ));
  OAI21_X1   g1517(.A1(new_n1448_), .A2(new_n1451_), .B(\shift[4] ), .ZN(new_n1781_));
  OAI21_X1   g1518(.A1(new_n1454_), .A2(new_n1457_), .B(new_n301_), .ZN(new_n1782_));
  AOI21_X1   g1519(.A1(new_n1782_), .A2(new_n1781_), .B(new_n265_), .ZN(new_n1783_));
  OAI21_X1   g1520(.A1(new_n1459_), .A2(new_n1462_), .B(\shift[4] ), .ZN(new_n1784_));
  OAI21_X1   g1521(.A1(new_n1482_), .A2(new_n1485_), .B(new_n301_), .ZN(new_n1785_));
  AOI21_X1   g1522(.A1(new_n1784_), .A2(new_n1785_), .B(\shift[5] ), .ZN(new_n1786_));
  OAI21_X1   g1523(.A1(new_n1783_), .A2(new_n1786_), .B(new_n264_), .ZN(new_n1787_));
  OAI21_X1   g1524(.A1(new_n1468_), .A2(new_n1469_), .B(new_n753_), .ZN(new_n1788_));
  OAI21_X1   g1525(.A1(new_n1471_), .A2(new_n1474_), .B(new_n722_), .ZN(new_n1789_));
  NAND2_X1   g1526(.A1(new_n1789_), .A2(new_n1788_), .ZN(new_n1790_));
  NOR2_X1    g1527(.A1(new_n1443_), .A2(new_n1446_), .ZN(new_n1791_));
  NOR2_X1    g1528(.A1(new_n1480_), .A2(new_n1477_), .ZN(new_n1792_));
  OAI22_X1   g1529(.A1(new_n851_), .A2(new_n1791_), .B1(new_n1792_), .B2(new_n852_), .ZN(new_n1793_));
  OAI21_X1   g1530(.A1(new_n1793_), .A2(new_n1790_), .B(\shift[6] ), .ZN(new_n1794_));
  NAND2_X1   g1531(.A1(new_n1787_), .A2(new_n1794_), .ZN(\result[27] ));
  OAI21_X1   g1532(.A1(new_n1493_), .A2(new_n1494_), .B(\shift[4] ), .ZN(new_n1796_));
  OAI21_X1   g1533(.A1(new_n1497_), .A2(new_n1498_), .B(new_n301_), .ZN(new_n1797_));
  AOI21_X1   g1534(.A1(new_n1796_), .A2(new_n1797_), .B(new_n265_), .ZN(new_n1798_));
  OAI21_X1   g1535(.A1(new_n1500_), .A2(new_n1501_), .B(\shift[4] ), .ZN(new_n1799_));
  OAI21_X1   g1536(.A1(new_n1515_), .A2(new_n1516_), .B(new_n301_), .ZN(new_n1800_));
  AOI21_X1   g1537(.A1(new_n1799_), .A2(new_n1800_), .B(\shift[5] ), .ZN(new_n1801_));
  OAI21_X1   g1538(.A1(new_n1798_), .A2(new_n1801_), .B(new_n264_), .ZN(new_n1802_));
  NOR2_X1    g1539(.A1(new_n1505_), .A2(new_n1506_), .ZN(new_n1803_));
  NOR2_X1    g1540(.A1(new_n1508_), .A2(new_n1509_), .ZN(new_n1804_));
  OAI22_X1   g1541(.A1(new_n1722_), .A2(new_n1804_), .B1(new_n1803_), .B2(new_n1723_), .ZN(new_n1805_));
  OAI21_X1   g1542(.A1(new_n1490_), .A2(new_n1491_), .B(new_n657_), .ZN(new_n1806_));
  OAI21_X1   g1543(.A1(new_n1512_), .A2(new_n1513_), .B(new_n689_), .ZN(new_n1807_));
  NAND2_X1   g1544(.A1(new_n1806_), .A2(new_n1807_), .ZN(new_n1808_));
  OAI21_X1   g1545(.A1(new_n1805_), .A2(new_n1808_), .B(\shift[6] ), .ZN(new_n1809_));
  NAND2_X1   g1546(.A1(new_n1802_), .A2(new_n1809_), .ZN(\result[28] ));
  OAI21_X1   g1547(.A1(new_n1525_), .A2(new_n1524_), .B(\shift[4] ), .ZN(new_n1811_));
  OAI21_X1   g1548(.A1(new_n1529_), .A2(new_n1528_), .B(new_n301_), .ZN(new_n1812_));
  AOI21_X1   g1549(.A1(new_n1811_), .A2(new_n1812_), .B(new_n265_), .ZN(new_n1813_));
  OAI21_X1   g1550(.A1(new_n1532_), .A2(new_n1531_), .B(\shift[4] ), .ZN(new_n1814_));
  OAI21_X1   g1551(.A1(new_n1547_), .A2(new_n1546_), .B(new_n301_), .ZN(new_n1815_));
  AOI21_X1   g1552(.A1(new_n1814_), .A2(new_n1815_), .B(\shift[5] ), .ZN(new_n1816_));
  OAI21_X1   g1553(.A1(new_n1816_), .A2(new_n1813_), .B(new_n264_), .ZN(new_n1817_));
  OAI21_X1   g1554(.A1(new_n1536_), .A2(new_n1537_), .B(new_n753_), .ZN(new_n1818_));
  OAI21_X1   g1555(.A1(new_n1540_), .A2(new_n1539_), .B(new_n722_), .ZN(new_n1819_));
  NAND2_X1   g1556(.A1(new_n1818_), .A2(new_n1819_), .ZN(new_n1820_));
  OAI21_X1   g1557(.A1(new_n1521_), .A2(new_n1522_), .B(new_n657_), .ZN(new_n1821_));
  OAI21_X1   g1558(.A1(new_n1543_), .A2(new_n1544_), .B(new_n689_), .ZN(new_n1822_));
  NAND2_X1   g1559(.A1(new_n1821_), .A2(new_n1822_), .ZN(new_n1823_));
  OAI21_X1   g1560(.A1(new_n1820_), .A2(new_n1823_), .B(\shift[6] ), .ZN(new_n1824_));
  NAND2_X1   g1561(.A1(new_n1817_), .A2(new_n1824_), .ZN(\result[29] ));
  OAI21_X1   g1562(.A1(new_n1555_), .A2(new_n1556_), .B(\shift[4] ), .ZN(new_n1826_));
  OAI21_X1   g1563(.A1(new_n1559_), .A2(new_n1560_), .B(new_n301_), .ZN(new_n1827_));
  AOI21_X1   g1564(.A1(new_n1826_), .A2(new_n1827_), .B(new_n265_), .ZN(new_n1828_));
  OAI21_X1   g1565(.A1(new_n1562_), .A2(new_n1563_), .B(\shift[4] ), .ZN(new_n1829_));
  OAI21_X1   g1566(.A1(new_n1577_), .A2(new_n1578_), .B(new_n301_), .ZN(new_n1830_));
  AOI21_X1   g1567(.A1(new_n1829_), .A2(new_n1830_), .B(\shift[5] ), .ZN(new_n1831_));
  OAI21_X1   g1568(.A1(new_n1828_), .A2(new_n1831_), .B(new_n264_), .ZN(new_n1832_));
  NOR2_X1    g1569(.A1(new_n1567_), .A2(new_n1568_), .ZN(new_n1833_));
  NOR2_X1    g1570(.A1(new_n1570_), .A2(new_n1571_), .ZN(new_n1834_));
  OAI22_X1   g1571(.A1(new_n1722_), .A2(new_n1834_), .B1(new_n1833_), .B2(new_n1723_), .ZN(new_n1835_));
  OAI21_X1   g1572(.A1(new_n1552_), .A2(new_n1553_), .B(new_n657_), .ZN(new_n1836_));
  OAI21_X1   g1573(.A1(new_n1574_), .A2(new_n1575_), .B(new_n689_), .ZN(new_n1837_));
  NAND2_X1   g1574(.A1(new_n1836_), .A2(new_n1837_), .ZN(new_n1838_));
  OAI21_X1   g1575(.A1(new_n1835_), .A2(new_n1838_), .B(\shift[6] ), .ZN(new_n1839_));
  NAND2_X1   g1576(.A1(new_n1832_), .A2(new_n1839_), .ZN(\result[30] ));
  OAI21_X1   g1577(.A1(new_n1587_), .A2(new_n1586_), .B(\shift[4] ), .ZN(new_n1841_));
  OAI21_X1   g1578(.A1(new_n1590_), .A2(new_n1591_), .B(new_n301_), .ZN(new_n1842_));
  AOI21_X1   g1579(.A1(new_n1842_), .A2(new_n1841_), .B(new_n265_), .ZN(new_n1843_));
  OAI21_X1   g1580(.A1(new_n1594_), .A2(new_n1593_), .B(\shift[4] ), .ZN(new_n1844_));
  OAI21_X1   g1581(.A1(new_n1609_), .A2(new_n1608_), .B(new_n301_), .ZN(new_n1845_));
  AOI21_X1   g1582(.A1(new_n1844_), .A2(new_n1845_), .B(\shift[5] ), .ZN(new_n1846_));
  OAI21_X1   g1583(.A1(new_n1843_), .A2(new_n1846_), .B(new_n264_), .ZN(new_n1847_));
  NOR2_X1    g1584(.A1(new_n1598_), .A2(new_n1599_), .ZN(new_n1848_));
  NOR2_X1    g1585(.A1(new_n1602_), .A2(new_n1601_), .ZN(new_n1849_));
  OAI22_X1   g1586(.A1(new_n1722_), .A2(new_n1849_), .B1(new_n1848_), .B2(new_n1723_), .ZN(new_n1850_));
  OAI21_X1   g1587(.A1(new_n1584_), .A2(new_n1583_), .B(new_n657_), .ZN(new_n1851_));
  OAI21_X1   g1588(.A1(new_n1605_), .A2(new_n1606_), .B(new_n689_), .ZN(new_n1852_));
  NAND2_X1   g1589(.A1(new_n1851_), .A2(new_n1852_), .ZN(new_n1853_));
  OAI21_X1   g1590(.A1(new_n1850_), .A2(new_n1853_), .B(\shift[6] ), .ZN(new_n1854_));
  NAND2_X1   g1591(.A1(new_n1847_), .A2(new_n1854_), .ZN(\result[31] ));
  AOI21_X1   g1592(.A1(new_n364_), .A2(new_n395_), .B(new_n265_), .ZN(new_n1856_));
  AOI21_X1   g1593(.A1(new_n428_), .A2(new_n459_), .B(\shift[5] ), .ZN(new_n1857_));
  OAI21_X1   g1594(.A1(new_n1856_), .A2(new_n1857_), .B(new_n264_), .ZN(new_n1858_));
  AOI21_X1   g1595(.A1(new_n300_), .A2(new_n332_), .B(\shift[5] ), .ZN(new_n1859_));
  AOI21_X1   g1596(.A1(new_n495_), .A2(new_n526_), .B(new_n265_), .ZN(new_n1860_));
  OAI21_X1   g1597(.A1(new_n1859_), .A2(new_n1860_), .B(\shift[6] ), .ZN(new_n1861_));
  NAND2_X1   g1598(.A1(new_n1858_), .A2(new_n1861_), .ZN(\result[32] ));
  AOI21_X1   g1599(.A1(new_n623_), .A2(new_n654_), .B(new_n265_), .ZN(new_n1863_));
  OAI21_X1   g1600(.A1(new_n704_), .A2(new_n719_), .B(\shift[4] ), .ZN(new_n1864_));
  OAI21_X1   g1601(.A1(new_n768_), .A2(new_n783_), .B(new_n301_), .ZN(new_n1865_));
  AOI21_X1   g1602(.A1(new_n1864_), .A2(new_n1865_), .B(\shift[5] ), .ZN(new_n1866_));
  OAI21_X1   g1603(.A1(new_n1866_), .A2(new_n1863_), .B(new_n264_), .ZN(new_n1867_));
  OAI21_X1   g1604(.A1(new_n559_), .A2(new_n544_), .B(new_n722_), .ZN(new_n1868_));
  OAI21_X1   g1605(.A1(new_n687_), .A2(new_n672_), .B(new_n753_), .ZN(new_n1869_));
  NAND2_X1   g1606(.A1(new_n1868_), .A2(new_n1869_), .ZN(new_n1870_));
  OAI21_X1   g1607(.A1(new_n575_), .A2(new_n590_), .B(new_n657_), .ZN(new_n1871_));
  OAI21_X1   g1608(.A1(new_n736_), .A2(new_n751_), .B(new_n689_), .ZN(new_n1872_));
  NAND2_X1   g1609(.A1(new_n1871_), .A2(new_n1872_), .ZN(new_n1873_));
  OAI21_X1   g1610(.A1(new_n1870_), .A2(new_n1873_), .B(\shift[6] ), .ZN(new_n1874_));
  NAND2_X1   g1611(.A1(new_n1867_), .A2(new_n1874_), .ZN(\result[33] ));
  AOI21_X1   g1612(.A1(new_n833_), .A2(new_n848_), .B(new_n265_), .ZN(new_n1876_));
  OAI21_X1   g1613(.A1(new_n874_), .A2(new_n881_), .B(\shift[4] ), .ZN(new_n1877_));
  OAI21_X1   g1614(.A1(new_n909_), .A2(new_n916_), .B(new_n301_), .ZN(new_n1878_));
  AOI21_X1   g1615(.A1(new_n1877_), .A2(new_n1878_), .B(\shift[5] ), .ZN(new_n1879_));
  OAI21_X1   g1616(.A1(new_n1876_), .A2(new_n1879_), .B(new_n264_), .ZN(new_n1880_));
  NOR2_X1    g1617(.A1(new_n794_), .A2(new_n801_), .ZN(new_n1881_));
  OAI22_X1   g1618(.A1(new_n1722_), .A2(new_n1881_), .B1(new_n867_), .B2(new_n1723_), .ZN(new_n1882_));
  OAI21_X1   g1619(.A1(new_n809_), .A2(new_n816_), .B(new_n657_), .ZN(new_n1883_));
  OAI21_X1   g1620(.A1(new_n892_), .A2(new_n901_), .B(new_n689_), .ZN(new_n1884_));
  NAND2_X1   g1621(.A1(new_n1883_), .A2(new_n1884_), .ZN(new_n1885_));
  OAI21_X1   g1622(.A1(new_n1882_), .A2(new_n1885_), .B(\shift[6] ), .ZN(new_n1886_));
  NAND2_X1   g1623(.A1(new_n1880_), .A2(new_n1886_), .ZN(\result[34] ));
  OAI21_X1   g1624(.A1(new_n1094_), .A2(new_n1109_), .B(new_n657_), .ZN(new_n1888_));
  OAI21_X1   g1625(.A1(new_n930_), .A2(new_n939_), .B(new_n689_), .ZN(new_n1889_));
  NAND2_X1   g1626(.A1(new_n1889_), .A2(new_n1888_), .ZN(new_n1890_));
  OAI21_X1   g1627(.A1(new_n974_), .A2(new_n985_), .B(new_n753_), .ZN(new_n1891_));
  OAI21_X1   g1628(.A1(new_n1068_), .A2(new_n1081_), .B(new_n722_), .ZN(new_n1892_));
  NAND2_X1   g1629(.A1(new_n1891_), .A2(new_n1892_), .ZN(new_n1893_));
  OAI21_X1   g1630(.A1(new_n1890_), .A2(new_n1893_), .B(new_n264_), .ZN(new_n1894_));
  OAI21_X1   g1631(.A1(new_n1057_), .A2(new_n1046_), .B(\shift[5] ), .ZN(new_n1895_));
  OAI21_X1   g1632(.A1(new_n949_), .A2(new_n962_), .B(new_n265_), .ZN(new_n1896_));
  AOI21_X1   g1633(.A1(new_n1896_), .A2(new_n1895_), .B(\shift[4] ), .ZN(new_n1897_));
  OAI21_X1   g1634(.A1(new_n994_), .A2(new_n1002_), .B(new_n265_), .ZN(new_n1898_));
  OAI21_X1   g1635(.A1(new_n1031_), .A2(new_n1017_), .B(\shift[5] ), .ZN(new_n1899_));
  AOI21_X1   g1636(.A1(new_n1898_), .A2(new_n1899_), .B(new_n301_), .ZN(new_n1900_));
  OAI21_X1   g1637(.A1(new_n1900_), .A2(new_n1897_), .B(\shift[6] ), .ZN(new_n1901_));
  NAND2_X1   g1638(.A1(new_n1901_), .A2(new_n1894_), .ZN(\result[35] ));
  AOI21_X1   g1639(.A1(new_n1129_), .A2(new_n1134_), .B(new_n265_), .ZN(new_n1903_));
  AOI21_X1   g1640(.A1(new_n1152_), .A2(new_n1157_), .B(\shift[5] ), .ZN(new_n1904_));
  OAI21_X1   g1641(.A1(new_n1903_), .A2(new_n1904_), .B(new_n264_), .ZN(new_n1905_));
  AOI21_X1   g1642(.A1(new_n1118_), .A2(new_n1123_), .B(\shift[5] ), .ZN(new_n1906_));
  AOI21_X1   g1643(.A1(new_n1141_), .A2(new_n1146_), .B(new_n265_), .ZN(new_n1907_));
  OAI21_X1   g1644(.A1(new_n1906_), .A2(new_n1907_), .B(\shift[6] ), .ZN(new_n1908_));
  NAND2_X1   g1645(.A1(new_n1905_), .A2(new_n1908_), .ZN(\result[36] ));
  AOI21_X1   g1646(.A1(new_n1176_), .A2(new_n1181_), .B(new_n265_), .ZN(new_n1910_));
  AOI21_X1   g1647(.A1(new_n1204_), .A2(new_n1199_), .B(\shift[5] ), .ZN(new_n1911_));
  OAI21_X1   g1648(.A1(new_n1910_), .A2(new_n1911_), .B(new_n264_), .ZN(new_n1912_));
  AOI21_X1   g1649(.A1(new_n1165_), .A2(new_n1170_), .B(\shift[5] ), .ZN(new_n1913_));
  AOI21_X1   g1650(.A1(new_n1193_), .A2(new_n1188_), .B(new_n265_), .ZN(new_n1914_));
  OAI21_X1   g1651(.A1(new_n1913_), .A2(new_n1914_), .B(\shift[6] ), .ZN(new_n1915_));
  NAND2_X1   g1652(.A1(new_n1912_), .A2(new_n1915_), .ZN(\result[37] ));
  AOI21_X1   g1653(.A1(new_n1223_), .A2(new_n1228_), .B(new_n265_), .ZN(new_n1917_));
  AOI21_X1   g1654(.A1(new_n1246_), .A2(new_n1251_), .B(\shift[5] ), .ZN(new_n1918_));
  OAI21_X1   g1655(.A1(new_n1917_), .A2(new_n1918_), .B(new_n264_), .ZN(new_n1919_));
  AOI21_X1   g1656(.A1(new_n1212_), .A2(new_n1217_), .B(\shift[5] ), .ZN(new_n1920_));
  AOI21_X1   g1657(.A1(new_n1235_), .A2(new_n1240_), .B(new_n265_), .ZN(new_n1921_));
  OAI21_X1   g1658(.A1(new_n1920_), .A2(new_n1921_), .B(\shift[6] ), .ZN(new_n1922_));
  NAND2_X1   g1659(.A1(new_n1919_), .A2(new_n1922_), .ZN(\result[38] ));
  AOI21_X1   g1660(.A1(new_n1298_), .A2(new_n1293_), .B(\shift[5] ), .ZN(new_n1924_));
  AOI21_X1   g1661(.A1(new_n1270_), .A2(new_n1275_), .B(new_n265_), .ZN(new_n1925_));
  OAI21_X1   g1662(.A1(new_n1925_), .A2(new_n1924_), .B(new_n264_), .ZN(new_n1926_));
  AOI21_X1   g1663(.A1(new_n1287_), .A2(new_n1282_), .B(new_n265_), .ZN(new_n1927_));
  AOI21_X1   g1664(.A1(new_n1259_), .A2(new_n1264_), .B(\shift[5] ), .ZN(new_n1928_));
  OAI21_X1   g1665(.A1(new_n1928_), .A2(new_n1927_), .B(\shift[6] ), .ZN(new_n1929_));
  NAND2_X1   g1666(.A1(new_n1926_), .A2(new_n1929_), .ZN(\result[39] ));
  AOI21_X1   g1667(.A1(new_n1340_), .A2(new_n1345_), .B(\shift[5] ), .ZN(new_n1931_));
  AOI21_X1   g1668(.A1(new_n1317_), .A2(new_n1322_), .B(new_n265_), .ZN(new_n1932_));
  OAI21_X1   g1669(.A1(new_n1931_), .A2(new_n1932_), .B(new_n264_), .ZN(new_n1933_));
  AOI21_X1   g1670(.A1(new_n1329_), .A2(new_n1334_), .B(new_n265_), .ZN(new_n1934_));
  AOI21_X1   g1671(.A1(new_n1306_), .A2(new_n1311_), .B(\shift[5] ), .ZN(new_n1935_));
  OAI21_X1   g1672(.A1(new_n1934_), .A2(new_n1935_), .B(\shift[6] ), .ZN(new_n1936_));
  NAND2_X1   g1673(.A1(new_n1933_), .A2(new_n1936_), .ZN(\result[40] ));
  AOI21_X1   g1674(.A1(new_n1392_), .A2(new_n1387_), .B(\shift[5] ), .ZN(new_n1938_));
  AOI21_X1   g1675(.A1(new_n1369_), .A2(new_n1364_), .B(new_n265_), .ZN(new_n1939_));
  OAI21_X1   g1676(.A1(new_n1939_), .A2(new_n1938_), .B(new_n264_), .ZN(new_n1940_));
  AOI21_X1   g1677(.A1(new_n1381_), .A2(new_n1376_), .B(new_n265_), .ZN(new_n1941_));
  AOI21_X1   g1678(.A1(new_n1353_), .A2(new_n1358_), .B(\shift[5] ), .ZN(new_n1942_));
  OAI21_X1   g1679(.A1(new_n1942_), .A2(new_n1941_), .B(\shift[6] ), .ZN(new_n1943_));
  NAND2_X1   g1680(.A1(new_n1940_), .A2(new_n1943_), .ZN(\result[41] ));
  AOI21_X1   g1681(.A1(new_n1411_), .A2(new_n1416_), .B(new_n265_), .ZN(new_n1945_));
  AOI21_X1   g1682(.A1(new_n1434_), .A2(new_n1439_), .B(\shift[5] ), .ZN(new_n1946_));
  OAI21_X1   g1683(.A1(new_n1945_), .A2(new_n1946_), .B(new_n264_), .ZN(new_n1947_));
  AOI21_X1   g1684(.A1(new_n1423_), .A2(new_n1428_), .B(new_n265_), .ZN(new_n1948_));
  AOI21_X1   g1685(.A1(new_n1400_), .A2(new_n1405_), .B(\shift[5] ), .ZN(new_n1949_));
  OAI21_X1   g1686(.A1(new_n1948_), .A2(new_n1949_), .B(\shift[6] ), .ZN(new_n1950_));
  NAND2_X1   g1687(.A1(new_n1947_), .A2(new_n1950_), .ZN(\result[42] ));
  AOI21_X1   g1688(.A1(new_n1458_), .A2(new_n1463_), .B(new_n265_), .ZN(new_n1952_));
  AOI21_X1   g1689(.A1(new_n1486_), .A2(new_n1481_), .B(\shift[5] ), .ZN(new_n1953_));
  OAI21_X1   g1690(.A1(new_n1952_), .A2(new_n1953_), .B(new_n264_), .ZN(new_n1954_));
  AOI21_X1   g1691(.A1(new_n1475_), .A2(new_n1470_), .B(new_n265_), .ZN(new_n1955_));
  AOI21_X1   g1692(.A1(new_n1447_), .A2(new_n1452_), .B(\shift[5] ), .ZN(new_n1956_));
  OAI21_X1   g1693(.A1(new_n1956_), .A2(new_n1955_), .B(\shift[6] ), .ZN(new_n1957_));
  NAND2_X1   g1694(.A1(new_n1954_), .A2(new_n1957_), .ZN(\result[43] ));
  AOI21_X1   g1695(.A1(new_n1499_), .A2(new_n1502_), .B(new_n265_), .ZN(new_n1959_));
  AOI21_X1   g1696(.A1(new_n1514_), .A2(new_n1517_), .B(\shift[5] ), .ZN(new_n1960_));
  OAI21_X1   g1697(.A1(new_n1959_), .A2(new_n1960_), .B(new_n264_), .ZN(new_n1961_));
  AOI21_X1   g1698(.A1(new_n1507_), .A2(new_n1510_), .B(new_n265_), .ZN(new_n1962_));
  AOI21_X1   g1699(.A1(new_n1492_), .A2(new_n1495_), .B(\shift[5] ), .ZN(new_n1963_));
  OAI21_X1   g1700(.A1(new_n1962_), .A2(new_n1963_), .B(\shift[6] ), .ZN(new_n1964_));
  NAND2_X1   g1701(.A1(new_n1961_), .A2(new_n1964_), .ZN(\result[44] ));
  AOI21_X1   g1702(.A1(new_n1533_), .A2(new_n1530_), .B(new_n265_), .ZN(new_n1966_));
  AOI21_X1   g1703(.A1(new_n1548_), .A2(new_n1545_), .B(\shift[5] ), .ZN(new_n1967_));
  OAI21_X1   g1704(.A1(new_n1966_), .A2(new_n1967_), .B(new_n264_), .ZN(new_n1968_));
  AOI21_X1   g1705(.A1(new_n1538_), .A2(new_n1541_), .B(new_n265_), .ZN(new_n1969_));
  AOI21_X1   g1706(.A1(new_n1523_), .A2(new_n1526_), .B(\shift[5] ), .ZN(new_n1970_));
  OAI21_X1   g1707(.A1(new_n1969_), .A2(new_n1970_), .B(\shift[6] ), .ZN(new_n1971_));
  NAND2_X1   g1708(.A1(new_n1971_), .A2(new_n1968_), .ZN(\result[45] ));
  AOI21_X1   g1709(.A1(new_n1561_), .A2(new_n1564_), .B(new_n265_), .ZN(new_n1973_));
  AOI21_X1   g1710(.A1(new_n1576_), .A2(new_n1579_), .B(\shift[5] ), .ZN(new_n1974_));
  OAI21_X1   g1711(.A1(new_n1973_), .A2(new_n1974_), .B(new_n264_), .ZN(new_n1975_));
  AOI21_X1   g1712(.A1(new_n1569_), .A2(new_n1572_), .B(new_n265_), .ZN(new_n1976_));
  AOI21_X1   g1713(.A1(new_n1554_), .A2(new_n1557_), .B(\shift[5] ), .ZN(new_n1977_));
  OAI21_X1   g1714(.A1(new_n1976_), .A2(new_n1977_), .B(\shift[6] ), .ZN(new_n1978_));
  NAND2_X1   g1715(.A1(new_n1975_), .A2(new_n1978_), .ZN(\result[46] ));
  AOI21_X1   g1716(.A1(new_n1592_), .A2(new_n1595_), .B(new_n265_), .ZN(new_n1980_));
  AOI21_X1   g1717(.A1(new_n1610_), .A2(new_n1607_), .B(\shift[5] ), .ZN(new_n1981_));
  OAI21_X1   g1718(.A1(new_n1980_), .A2(new_n1981_), .B(new_n264_), .ZN(new_n1982_));
  AOI21_X1   g1719(.A1(new_n1603_), .A2(new_n1600_), .B(new_n265_), .ZN(new_n1983_));
  AOI21_X1   g1720(.A1(new_n1585_), .A2(new_n1588_), .B(\shift[5] ), .ZN(new_n1984_));
  OAI21_X1   g1721(.A1(new_n1984_), .A2(new_n1983_), .B(\shift[6] ), .ZN(new_n1985_));
  NAND2_X1   g1722(.A1(new_n1985_), .A2(new_n1982_), .ZN(\result[47] ));
  AOI21_X1   g1723(.A1(new_n1617_), .A2(new_n1618_), .B(new_n265_), .ZN(new_n1987_));
  OAI21_X1   g1724(.A1(new_n443_), .A2(new_n458_), .B(\shift[4] ), .ZN(new_n1988_));
  OAI21_X1   g1725(.A1(new_n494_), .A2(new_n475_), .B(new_n301_), .ZN(new_n1989_));
  AOI21_X1   g1726(.A1(new_n1988_), .A2(new_n1989_), .B(\shift[5] ), .ZN(new_n1990_));
  OAI21_X1   g1727(.A1(new_n1987_), .A2(new_n1990_), .B(new_n264_), .ZN(new_n1991_));
  NOR2_X1    g1728(.A1(new_n316_), .A2(new_n331_), .ZN(new_n1992_));
  OAI22_X1   g1729(.A1(new_n1621_), .A2(new_n1723_), .B1(new_n1992_), .B2(new_n1722_), .ZN(new_n1993_));
  OAI21_X1   g1730(.A1(new_n348_), .A2(new_n363_), .B(new_n657_), .ZN(new_n1994_));
  OAI21_X1   g1731(.A1(new_n510_), .A2(new_n525_), .B(new_n689_), .ZN(new_n1995_));
  NAND2_X1   g1732(.A1(new_n1994_), .A2(new_n1995_), .ZN(new_n1996_));
  OAI21_X1   g1733(.A1(new_n1993_), .A2(new_n1996_), .B(\shift[6] ), .ZN(new_n1997_));
  NAND2_X1   g1734(.A1(new_n1991_), .A2(new_n1997_), .ZN(\result[48] ));
  AOI21_X1   g1735(.A1(new_n1633_), .A2(new_n1632_), .B(new_n265_), .ZN(new_n1999_));
  AOI21_X1   g1736(.A1(new_n1640_), .A2(new_n1639_), .B(\shift[5] ), .ZN(new_n2000_));
  OAI21_X1   g1737(.A1(new_n1999_), .A2(new_n2000_), .B(new_n264_), .ZN(new_n2001_));
  AOI21_X1   g1738(.A1(new_n1637_), .A2(new_n1636_), .B(new_n265_), .ZN(new_n2002_));
  AOI21_X1   g1739(.A1(new_n1629_), .A2(new_n1630_), .B(\shift[5] ), .ZN(new_n2003_));
  OAI21_X1   g1740(.A1(new_n2002_), .A2(new_n2003_), .B(\shift[6] ), .ZN(new_n2004_));
  NAND2_X1   g1741(.A1(new_n2004_), .A2(new_n2001_), .ZN(\result[49] ));
  AOI21_X1   g1742(.A1(new_n1647_), .A2(new_n1648_), .B(new_n265_), .ZN(new_n2006_));
  AOI21_X1   g1743(.A1(new_n1654_), .A2(new_n1655_), .B(\shift[5] ), .ZN(new_n2007_));
  OAI21_X1   g1744(.A1(new_n2006_), .A2(new_n2007_), .B(new_n264_), .ZN(new_n2008_));
  AOI21_X1   g1745(.A1(new_n1651_), .A2(new_n1652_), .B(new_n265_), .ZN(new_n2009_));
  AOI21_X1   g1746(.A1(new_n1644_), .A2(new_n1645_), .B(\shift[5] ), .ZN(new_n2010_));
  OAI21_X1   g1747(.A1(new_n2009_), .A2(new_n2010_), .B(\shift[6] ), .ZN(new_n2011_));
  NAND2_X1   g1748(.A1(new_n2008_), .A2(new_n2011_), .ZN(\result[50] ));
  AOI21_X1   g1749(.A1(new_n1670_), .A2(new_n1669_), .B(\shift[5] ), .ZN(new_n2013_));
  AOI21_X1   g1750(.A1(new_n1662_), .A2(new_n1663_), .B(new_n265_), .ZN(new_n2014_));
  OAI21_X1   g1751(.A1(new_n2014_), .A2(new_n2013_), .B(new_n264_), .ZN(new_n2015_));
  AOI21_X1   g1752(.A1(new_n1659_), .A2(new_n1895_), .B(new_n753_), .ZN(new_n2016_));
  AOI21_X1   g1753(.A1(new_n1667_), .A2(new_n1896_), .B(new_n657_), .ZN(new_n2017_));
  OAI21_X1   g1754(.A1(new_n2017_), .A2(new_n2016_), .B(\shift[6] ), .ZN(new_n2018_));
  NAND2_X1   g1755(.A1(new_n2018_), .A2(new_n2015_), .ZN(\result[51] ));
  NOR2_X1    g1756(.A1(new_n1130_), .A2(new_n1133_), .ZN(new_n2020_));
  NOR2_X1    g1757(.A1(new_n1137_), .A2(new_n1140_), .ZN(new_n2021_));
  OAI22_X1   g1758(.A1(new_n851_), .A2(new_n2021_), .B1(new_n2020_), .B2(new_n852_), .ZN(new_n2022_));
  NOR2_X1    g1759(.A1(new_n1148_), .A2(new_n1151_), .ZN(new_n2023_));
  NOR2_X1    g1760(.A1(new_n1153_), .A2(new_n1156_), .ZN(new_n2024_));
  OAI22_X1   g1761(.A1(new_n1722_), .A2(new_n2023_), .B1(new_n2024_), .B2(new_n1723_), .ZN(new_n2025_));
  OAI21_X1   g1762(.A1(new_n2022_), .A2(new_n2025_), .B(new_n264_), .ZN(new_n2026_));
  NOR2_X1    g1763(.A1(new_n1114_), .A2(new_n1117_), .ZN(new_n2027_));
  NOR2_X1    g1764(.A1(new_n1119_), .A2(new_n1122_), .ZN(new_n2028_));
  OAI22_X1   g1765(.A1(new_n1722_), .A2(new_n2028_), .B1(new_n2027_), .B2(new_n1723_), .ZN(new_n2029_));
  OAI21_X1   g1766(.A1(new_n1125_), .A2(new_n1128_), .B(new_n657_), .ZN(new_n2030_));
  OAI21_X1   g1767(.A1(new_n1142_), .A2(new_n1145_), .B(new_n689_), .ZN(new_n2031_));
  NAND2_X1   g1768(.A1(new_n2030_), .A2(new_n2031_), .ZN(new_n2032_));
  OAI21_X1   g1769(.A1(new_n2029_), .A2(new_n2032_), .B(\shift[6] ), .ZN(new_n2033_));
  NAND2_X1   g1770(.A1(new_n2026_), .A2(new_n2033_), .ZN(\result[52] ));
  OAI21_X1   g1771(.A1(new_n1184_), .A2(new_n1187_), .B(new_n657_), .ZN(new_n2035_));
  OAI21_X1   g1772(.A1(new_n1180_), .A2(new_n1177_), .B(new_n689_), .ZN(new_n2036_));
  NAND2_X1   g1773(.A1(new_n2036_), .A2(new_n2035_), .ZN(new_n2037_));
  NOR2_X1    g1774(.A1(new_n1195_), .A2(new_n1198_), .ZN(new_n2038_));
  NOR2_X1    g1775(.A1(new_n1203_), .A2(new_n1200_), .ZN(new_n2039_));
  OAI22_X1   g1776(.A1(new_n1723_), .A2(new_n2039_), .B1(new_n2038_), .B2(new_n1722_), .ZN(new_n2040_));
  OAI21_X1   g1777(.A1(new_n2040_), .A2(new_n2037_), .B(new_n264_), .ZN(new_n2041_));
  NOR2_X1    g1778(.A1(new_n1161_), .A2(new_n1164_), .ZN(new_n2042_));
  NOR2_X1    g1779(.A1(new_n1166_), .A2(new_n1169_), .ZN(new_n2043_));
  OAI22_X1   g1780(.A1(new_n1722_), .A2(new_n2043_), .B1(new_n2042_), .B2(new_n1723_), .ZN(new_n2044_));
  OAI21_X1   g1781(.A1(new_n1175_), .A2(new_n1172_), .B(new_n657_), .ZN(new_n2045_));
  OAI21_X1   g1782(.A1(new_n1189_), .A2(new_n1192_), .B(new_n689_), .ZN(new_n2046_));
  NAND2_X1   g1783(.A1(new_n2046_), .A2(new_n2045_), .ZN(new_n2047_));
  OAI21_X1   g1784(.A1(new_n2044_), .A2(new_n2047_), .B(\shift[6] ), .ZN(new_n2048_));
  NAND2_X1   g1785(.A1(new_n2048_), .A2(new_n2041_), .ZN(\result[53] ));
  NOR2_X1    g1786(.A1(new_n1224_), .A2(new_n1227_), .ZN(new_n2050_));
  NOR2_X1    g1787(.A1(new_n1231_), .A2(new_n1234_), .ZN(new_n2051_));
  OAI22_X1   g1788(.A1(new_n851_), .A2(new_n2051_), .B1(new_n2050_), .B2(new_n852_), .ZN(new_n2052_));
  NOR2_X1    g1789(.A1(new_n1242_), .A2(new_n1245_), .ZN(new_n2053_));
  NOR2_X1    g1790(.A1(new_n1247_), .A2(new_n1250_), .ZN(new_n2054_));
  OAI22_X1   g1791(.A1(new_n1722_), .A2(new_n2053_), .B1(new_n2054_), .B2(new_n1723_), .ZN(new_n2055_));
  OAI21_X1   g1792(.A1(new_n2052_), .A2(new_n2055_), .B(new_n264_), .ZN(new_n2056_));
  NOR2_X1    g1793(.A1(new_n1208_), .A2(new_n1211_), .ZN(new_n2057_));
  NOR2_X1    g1794(.A1(new_n1213_), .A2(new_n1216_), .ZN(new_n2058_));
  OAI22_X1   g1795(.A1(new_n1722_), .A2(new_n2058_), .B1(new_n2057_), .B2(new_n1723_), .ZN(new_n2059_));
  OAI21_X1   g1796(.A1(new_n1219_), .A2(new_n1222_), .B(new_n657_), .ZN(new_n2060_));
  OAI21_X1   g1797(.A1(new_n1236_), .A2(new_n1239_), .B(new_n689_), .ZN(new_n2061_));
  NAND2_X1   g1798(.A1(new_n2060_), .A2(new_n2061_), .ZN(new_n2062_));
  OAI21_X1   g1799(.A1(new_n2059_), .A2(new_n2062_), .B(\shift[6] ), .ZN(new_n2063_));
  NAND2_X1   g1800(.A1(new_n2056_), .A2(new_n2063_), .ZN(\result[54] ));
  OAI21_X1   g1801(.A1(new_n1297_), .A2(new_n1294_), .B(\shift[5] ), .ZN(new_n2065_));
  OAI21_X1   g1802(.A1(new_n1278_), .A2(new_n1281_), .B(new_n265_), .ZN(new_n2066_));
  AOI21_X1   g1803(.A1(new_n2065_), .A2(new_n2066_), .B(\shift[4] ), .ZN(new_n2067_));
  OAI21_X1   g1804(.A1(new_n1274_), .A2(new_n1271_), .B(\shift[5] ), .ZN(new_n2068_));
  OAI21_X1   g1805(.A1(new_n1289_), .A2(new_n1292_), .B(new_n265_), .ZN(new_n2069_));
  AOI21_X1   g1806(.A1(new_n2068_), .A2(new_n2069_), .B(new_n301_), .ZN(new_n2070_));
  OAI21_X1   g1807(.A1(new_n2070_), .A2(new_n2067_), .B(new_n264_), .ZN(new_n2071_));
  OAI21_X1   g1808(.A1(new_n1255_), .A2(new_n1258_), .B(new_n301_), .ZN(new_n2072_));
  OAI21_X1   g1809(.A1(new_n1286_), .A2(new_n1283_), .B(\shift[4] ), .ZN(new_n2073_));
  AOI21_X1   g1810(.A1(new_n2072_), .A2(new_n2073_), .B(new_n265_), .ZN(new_n2074_));
  OAI21_X1   g1811(.A1(new_n1263_), .A2(new_n1260_), .B(\shift[4] ), .ZN(new_n2075_));
  OAI21_X1   g1812(.A1(new_n1266_), .A2(new_n1269_), .B(new_n301_), .ZN(new_n2076_));
  AOI21_X1   g1813(.A1(new_n2076_), .A2(new_n2075_), .B(\shift[5] ), .ZN(new_n2077_));
  OAI21_X1   g1814(.A1(new_n2077_), .A2(new_n2074_), .B(\shift[6] ), .ZN(new_n2078_));
  NAND2_X1   g1815(.A1(new_n2078_), .A2(new_n2071_), .ZN(\result[55] ));
  OAI21_X1   g1816(.A1(new_n1341_), .A2(new_n1344_), .B(\shift[5] ), .ZN(new_n2080_));
  OAI21_X1   g1817(.A1(new_n1325_), .A2(new_n1328_), .B(new_n265_), .ZN(new_n2081_));
  AOI21_X1   g1818(.A1(new_n2080_), .A2(new_n2081_), .B(\shift[4] ), .ZN(new_n2082_));
  OAI21_X1   g1819(.A1(new_n1318_), .A2(new_n1321_), .B(\shift[5] ), .ZN(new_n2083_));
  OAI21_X1   g1820(.A1(new_n1339_), .A2(new_n1336_), .B(new_n265_), .ZN(new_n2084_));
  AOI21_X1   g1821(.A1(new_n2083_), .A2(new_n2084_), .B(new_n301_), .ZN(new_n2085_));
  OAI21_X1   g1822(.A1(new_n2082_), .A2(new_n2085_), .B(new_n264_), .ZN(new_n2086_));
  OAI21_X1   g1823(.A1(new_n1302_), .A2(new_n1305_), .B(new_n301_), .ZN(new_n2087_));
  OAI21_X1   g1824(.A1(new_n1330_), .A2(new_n1333_), .B(\shift[4] ), .ZN(new_n2088_));
  AOI21_X1   g1825(.A1(new_n2087_), .A2(new_n2088_), .B(new_n265_), .ZN(new_n2089_));
  OAI21_X1   g1826(.A1(new_n1307_), .A2(new_n1310_), .B(\shift[4] ), .ZN(new_n2090_));
  OAI21_X1   g1827(.A1(new_n1313_), .A2(new_n1316_), .B(new_n301_), .ZN(new_n2091_));
  AOI21_X1   g1828(.A1(new_n2090_), .A2(new_n2091_), .B(\shift[5] ), .ZN(new_n2092_));
  OAI21_X1   g1829(.A1(new_n2089_), .A2(new_n2092_), .B(\shift[6] ), .ZN(new_n2093_));
  NAND2_X1   g1830(.A1(new_n2086_), .A2(new_n2093_), .ZN(\result[56] ));
  OAI21_X1   g1831(.A1(new_n1388_), .A2(new_n1391_), .B(\shift[5] ), .ZN(new_n2095_));
  OAI21_X1   g1832(.A1(new_n1375_), .A2(new_n1372_), .B(new_n265_), .ZN(new_n2096_));
  AOI21_X1   g1833(.A1(new_n2095_), .A2(new_n2096_), .B(\shift[4] ), .ZN(new_n2097_));
  OAI21_X1   g1834(.A1(new_n1365_), .A2(new_n1368_), .B(\shift[5] ), .ZN(new_n2098_));
  OAI21_X1   g1835(.A1(new_n1383_), .A2(new_n1386_), .B(new_n265_), .ZN(new_n2099_));
  AOI21_X1   g1836(.A1(new_n2098_), .A2(new_n2099_), .B(new_n301_), .ZN(new_n2100_));
  OAI21_X1   g1837(.A1(new_n2097_), .A2(new_n2100_), .B(new_n264_), .ZN(new_n2101_));
  OAI21_X1   g1838(.A1(new_n1352_), .A2(new_n1349_), .B(new_n301_), .ZN(new_n2102_));
  OAI21_X1   g1839(.A1(new_n1377_), .A2(new_n1380_), .B(\shift[4] ), .ZN(new_n2103_));
  AOI21_X1   g1840(.A1(new_n2102_), .A2(new_n2103_), .B(new_n265_), .ZN(new_n2104_));
  OAI21_X1   g1841(.A1(new_n1354_), .A2(new_n1357_), .B(\shift[4] ), .ZN(new_n2105_));
  OAI21_X1   g1842(.A1(new_n1360_), .A2(new_n1363_), .B(new_n301_), .ZN(new_n2106_));
  AOI21_X1   g1843(.A1(new_n2106_), .A2(new_n2105_), .B(\shift[5] ), .ZN(new_n2107_));
  OAI21_X1   g1844(.A1(new_n2104_), .A2(new_n2107_), .B(\shift[6] ), .ZN(new_n2108_));
  NAND2_X1   g1845(.A1(new_n2108_), .A2(new_n2101_), .ZN(\result[57] ));
  NOR2_X1    g1846(.A1(new_n1412_), .A2(new_n1415_), .ZN(new_n2110_));
  OAI22_X1   g1847(.A1(new_n851_), .A2(new_n1773_), .B1(new_n2110_), .B2(new_n852_), .ZN(new_n2111_));
  OAI21_X1   g1848(.A1(new_n1430_), .A2(new_n1433_), .B(new_n722_), .ZN(new_n2112_));
  OAI21_X1   g1849(.A1(new_n1435_), .A2(new_n1438_), .B(new_n753_), .ZN(new_n2113_));
  NAND2_X1   g1850(.A1(new_n2112_), .A2(new_n2113_), .ZN(new_n2114_));
  OAI21_X1   g1851(.A1(new_n2111_), .A2(new_n2114_), .B(new_n264_), .ZN(new_n2115_));
  OAI21_X1   g1852(.A1(new_n1396_), .A2(new_n1399_), .B(new_n301_), .ZN(new_n2116_));
  OAI21_X1   g1853(.A1(new_n1424_), .A2(new_n1427_), .B(\shift[4] ), .ZN(new_n2117_));
  AOI21_X1   g1854(.A1(new_n2116_), .A2(new_n2117_), .B(new_n265_), .ZN(new_n2118_));
  AOI21_X1   g1855(.A1(new_n1766_), .A2(new_n1767_), .B(\shift[5] ), .ZN(new_n2119_));
  OAI21_X1   g1856(.A1(new_n2118_), .A2(new_n2119_), .B(\shift[6] ), .ZN(new_n2120_));
  NAND2_X1   g1857(.A1(new_n2120_), .A2(new_n2115_), .ZN(\result[58] ));
  OAI21_X1   g1858(.A1(new_n1468_), .A2(new_n1469_), .B(new_n657_), .ZN(new_n2122_));
  OAI21_X1   g1859(.A1(new_n1459_), .A2(new_n1462_), .B(new_n689_), .ZN(new_n2123_));
  NAND2_X1   g1860(.A1(new_n2123_), .A2(new_n2122_), .ZN(new_n2124_));
  NOR2_X1    g1861(.A1(new_n1482_), .A2(new_n1485_), .ZN(new_n2125_));
  OAI22_X1   g1862(.A1(new_n1723_), .A2(new_n2125_), .B1(new_n1792_), .B2(new_n1722_), .ZN(new_n2126_));
  OAI21_X1   g1863(.A1(new_n2126_), .A2(new_n2124_), .B(new_n264_), .ZN(new_n2127_));
  OAI21_X1   g1864(.A1(new_n1443_), .A2(new_n1446_), .B(new_n301_), .ZN(new_n2128_));
  OAI21_X1   g1865(.A1(new_n1471_), .A2(new_n1474_), .B(\shift[4] ), .ZN(new_n2129_));
  AOI21_X1   g1866(.A1(new_n2128_), .A2(new_n2129_), .B(new_n265_), .ZN(new_n2130_));
  AOI21_X1   g1867(.A1(new_n1782_), .A2(new_n1781_), .B(\shift[5] ), .ZN(new_n2131_));
  OAI21_X1   g1868(.A1(new_n2131_), .A2(new_n2130_), .B(\shift[6] ), .ZN(new_n2132_));
  NAND2_X1   g1869(.A1(new_n2132_), .A2(new_n2127_), .ZN(\result[59] ));
  NOR2_X1    g1870(.A1(new_n1500_), .A2(new_n1501_), .ZN(new_n2134_));
  OAI22_X1   g1871(.A1(new_n851_), .A2(new_n1803_), .B1(new_n2134_), .B2(new_n852_), .ZN(new_n2135_));
  OAI21_X1   g1872(.A1(new_n1512_), .A2(new_n1513_), .B(new_n722_), .ZN(new_n2136_));
  OAI21_X1   g1873(.A1(new_n1515_), .A2(new_n1516_), .B(new_n753_), .ZN(new_n2137_));
  NAND2_X1   g1874(.A1(new_n2136_), .A2(new_n2137_), .ZN(new_n2138_));
  OAI21_X1   g1875(.A1(new_n2135_), .A2(new_n2138_), .B(new_n264_), .ZN(new_n2139_));
  OAI21_X1   g1876(.A1(new_n1490_), .A2(new_n1491_), .B(new_n301_), .ZN(new_n2140_));
  OAI21_X1   g1877(.A1(new_n1508_), .A2(new_n1509_), .B(\shift[4] ), .ZN(new_n2141_));
  AOI21_X1   g1878(.A1(new_n2140_), .A2(new_n2141_), .B(new_n265_), .ZN(new_n2142_));
  AOI21_X1   g1879(.A1(new_n1796_), .A2(new_n1797_), .B(\shift[5] ), .ZN(new_n2143_));
  OAI21_X1   g1880(.A1(new_n2142_), .A2(new_n2143_), .B(\shift[6] ), .ZN(new_n2144_));
  NAND2_X1   g1881(.A1(new_n2144_), .A2(new_n2139_), .ZN(\result[60] ));
  OAI21_X1   g1882(.A1(new_n1536_), .A2(new_n1537_), .B(new_n657_), .ZN(new_n2146_));
  OAI21_X1   g1883(.A1(new_n1532_), .A2(new_n1531_), .B(new_n689_), .ZN(new_n2147_));
  NAND2_X1   g1884(.A1(new_n2146_), .A2(new_n2147_), .ZN(new_n2148_));
  OAI21_X1   g1885(.A1(new_n1543_), .A2(new_n1544_), .B(new_n722_), .ZN(new_n2149_));
  OAI21_X1   g1886(.A1(new_n1547_), .A2(new_n1546_), .B(new_n753_), .ZN(new_n2150_));
  NAND2_X1   g1887(.A1(new_n2150_), .A2(new_n2149_), .ZN(new_n2151_));
  OAI21_X1   g1888(.A1(new_n2148_), .A2(new_n2151_), .B(new_n264_), .ZN(new_n2152_));
  OAI21_X1   g1889(.A1(new_n1521_), .A2(new_n1522_), .B(new_n301_), .ZN(new_n2153_));
  OAI21_X1   g1890(.A1(new_n1540_), .A2(new_n1539_), .B(\shift[4] ), .ZN(new_n2154_));
  AOI21_X1   g1891(.A1(new_n2153_), .A2(new_n2154_), .B(new_n265_), .ZN(new_n2155_));
  AOI21_X1   g1892(.A1(new_n1811_), .A2(new_n1812_), .B(\shift[5] ), .ZN(new_n2156_));
  OAI21_X1   g1893(.A1(new_n2155_), .A2(new_n2156_), .B(\shift[6] ), .ZN(new_n2157_));
  NAND2_X1   g1894(.A1(new_n2157_), .A2(new_n2152_), .ZN(\result[61] ));
  NOR2_X1    g1895(.A1(new_n1562_), .A2(new_n1563_), .ZN(new_n2159_));
  OAI22_X1   g1896(.A1(new_n851_), .A2(new_n1833_), .B1(new_n2159_), .B2(new_n852_), .ZN(new_n2160_));
  OAI21_X1   g1897(.A1(new_n1574_), .A2(new_n1575_), .B(new_n722_), .ZN(new_n2161_));
  OAI21_X1   g1898(.A1(new_n1577_), .A2(new_n1578_), .B(new_n753_), .ZN(new_n2162_));
  NAND2_X1   g1899(.A1(new_n2161_), .A2(new_n2162_), .ZN(new_n2163_));
  OAI21_X1   g1900(.A1(new_n2160_), .A2(new_n2163_), .B(new_n264_), .ZN(new_n2164_));
  OAI21_X1   g1901(.A1(new_n1552_), .A2(new_n1553_), .B(new_n301_), .ZN(new_n2165_));
  OAI21_X1   g1902(.A1(new_n1570_), .A2(new_n1571_), .B(\shift[4] ), .ZN(new_n2166_));
  AOI21_X1   g1903(.A1(new_n2165_), .A2(new_n2166_), .B(new_n265_), .ZN(new_n2167_));
  AOI21_X1   g1904(.A1(new_n1826_), .A2(new_n1827_), .B(\shift[5] ), .ZN(new_n2168_));
  OAI21_X1   g1905(.A1(new_n2167_), .A2(new_n2168_), .B(\shift[6] ), .ZN(new_n2169_));
  NAND2_X1   g1906(.A1(new_n2169_), .A2(new_n2164_), .ZN(\result[62] ));
  NOR2_X1    g1907(.A1(new_n1594_), .A2(new_n1593_), .ZN(new_n2171_));
  OAI22_X1   g1908(.A1(new_n852_), .A2(new_n2171_), .B1(new_n1848_), .B2(new_n851_), .ZN(new_n2172_));
  OAI21_X1   g1909(.A1(new_n1605_), .A2(new_n1606_), .B(new_n722_), .ZN(new_n2173_));
  OAI21_X1   g1910(.A1(new_n1609_), .A2(new_n1608_), .B(new_n753_), .ZN(new_n2174_));
  NAND2_X1   g1911(.A1(new_n2174_), .A2(new_n2173_), .ZN(new_n2175_));
  OAI21_X1   g1912(.A1(new_n2172_), .A2(new_n2175_), .B(new_n264_), .ZN(new_n2176_));
  OAI21_X1   g1913(.A1(new_n1584_), .A2(new_n1583_), .B(new_n301_), .ZN(new_n2177_));
  OAI21_X1   g1914(.A1(new_n1602_), .A2(new_n1601_), .B(\shift[4] ), .ZN(new_n2178_));
  AOI21_X1   g1915(.A1(new_n2177_), .A2(new_n2178_), .B(new_n265_), .ZN(new_n2179_));
  AOI21_X1   g1916(.A1(new_n1842_), .A2(new_n1841_), .B(\shift[5] ), .ZN(new_n2180_));
  OAI21_X1   g1917(.A1(new_n2180_), .A2(new_n2179_), .B(\shift[6] ), .ZN(new_n2181_));
  NAND2_X1   g1918(.A1(new_n2181_), .A2(new_n2176_), .ZN(\result[63] ));
  OAI21_X1   g1919(.A1(new_n333_), .A2(new_n396_), .B(\shift[6] ), .ZN(new_n2183_));
  OAI21_X1   g1920(.A1(new_n460_), .A2(new_n527_), .B(new_n264_), .ZN(new_n2184_));
  NAND2_X1   g1921(.A1(new_n2183_), .A2(new_n2184_), .ZN(\result[64] ));
  OAI21_X1   g1922(.A1(new_n592_), .A2(new_n655_), .B(\shift[6] ), .ZN(new_n2186_));
  OAI21_X1   g1923(.A1(new_n721_), .A2(new_n785_), .B(new_n264_), .ZN(new_n2187_));
  NAND2_X1   g1924(.A1(new_n2186_), .A2(new_n2187_), .ZN(\result[65] ));
  OAI21_X1   g1925(.A1(new_n818_), .A2(new_n849_), .B(\shift[6] ), .ZN(new_n2189_));
  OAI21_X1   g1926(.A1(new_n883_), .A2(new_n918_), .B(new_n264_), .ZN(new_n2190_));
  NAND2_X1   g1927(.A1(new_n2189_), .A2(new_n2190_), .ZN(\result[66] ));
  OAI21_X1   g1928(.A1(new_n1004_), .A2(new_n964_), .B(\shift[6] ), .ZN(new_n2192_));
  OAI21_X1   g1929(.A1(new_n1111_), .A2(new_n1059_), .B(new_n264_), .ZN(new_n2193_));
  NAND2_X1   g1930(.A1(new_n2193_), .A2(new_n2192_), .ZN(\result[67] ));
  OAI21_X1   g1931(.A1(new_n1124_), .A2(new_n1135_), .B(\shift[6] ), .ZN(new_n2195_));
  OAI21_X1   g1932(.A1(new_n1147_), .A2(new_n1158_), .B(new_n264_), .ZN(new_n2196_));
  NAND2_X1   g1933(.A1(new_n2195_), .A2(new_n2196_), .ZN(\result[68] ));
  OAI21_X1   g1934(.A1(new_n1171_), .A2(new_n1182_), .B(\shift[6] ), .ZN(new_n2198_));
  OAI21_X1   g1935(.A1(new_n1205_), .A2(new_n1194_), .B(new_n264_), .ZN(new_n2199_));
  NAND2_X1   g1936(.A1(new_n2198_), .A2(new_n2199_), .ZN(\result[69] ));
  OAI21_X1   g1937(.A1(new_n1218_), .A2(new_n1229_), .B(\shift[6] ), .ZN(new_n2201_));
  OAI21_X1   g1938(.A1(new_n1241_), .A2(new_n1252_), .B(new_n264_), .ZN(new_n2202_));
  NAND2_X1   g1939(.A1(new_n2201_), .A2(new_n2202_), .ZN(\result[70] ));
  OAI21_X1   g1940(.A1(new_n1276_), .A2(new_n1265_), .B(\shift[6] ), .ZN(new_n2204_));
  OAI21_X1   g1941(.A1(new_n1299_), .A2(new_n1288_), .B(new_n264_), .ZN(new_n2205_));
  NAND2_X1   g1942(.A1(new_n2204_), .A2(new_n2205_), .ZN(\result[71] ));
  OAI21_X1   g1943(.A1(new_n1312_), .A2(new_n1323_), .B(\shift[6] ), .ZN(new_n2207_));
  OAI21_X1   g1944(.A1(new_n1335_), .A2(new_n1346_), .B(new_n264_), .ZN(new_n2208_));
  NAND2_X1   g1945(.A1(new_n2207_), .A2(new_n2208_), .ZN(\result[72] ));
  OAI21_X1   g1946(.A1(new_n1370_), .A2(new_n1359_), .B(\shift[6] ), .ZN(new_n2210_));
  OAI21_X1   g1947(.A1(new_n1382_), .A2(new_n1393_), .B(new_n264_), .ZN(new_n2211_));
  NAND2_X1   g1948(.A1(new_n2210_), .A2(new_n2211_), .ZN(\result[73] ));
  OAI21_X1   g1949(.A1(new_n1406_), .A2(new_n1417_), .B(\shift[6] ), .ZN(new_n2213_));
  OAI21_X1   g1950(.A1(new_n1429_), .A2(new_n1440_), .B(new_n264_), .ZN(new_n2214_));
  NAND2_X1   g1951(.A1(new_n2213_), .A2(new_n2214_), .ZN(\result[74] ));
  OAI21_X1   g1952(.A1(new_n1453_), .A2(new_n1464_), .B(\shift[6] ), .ZN(new_n2216_));
  OAI21_X1   g1953(.A1(new_n1487_), .A2(new_n1476_), .B(new_n264_), .ZN(new_n2217_));
  NAND2_X1   g1954(.A1(new_n2216_), .A2(new_n2217_), .ZN(\result[75] ));
  OAI21_X1   g1955(.A1(new_n1496_), .A2(new_n1503_), .B(\shift[6] ), .ZN(new_n2219_));
  OAI21_X1   g1956(.A1(new_n1511_), .A2(new_n1518_), .B(new_n264_), .ZN(new_n2220_));
  NAND2_X1   g1957(.A1(new_n2219_), .A2(new_n2220_), .ZN(\result[76] ));
  OAI21_X1   g1958(.A1(new_n1527_), .A2(new_n1534_), .B(\shift[6] ), .ZN(new_n2222_));
  OAI21_X1   g1959(.A1(new_n1542_), .A2(new_n1549_), .B(new_n264_), .ZN(new_n2223_));
  NAND2_X1   g1960(.A1(new_n2222_), .A2(new_n2223_), .ZN(\result[77] ));
  OAI21_X1   g1961(.A1(new_n1558_), .A2(new_n1565_), .B(\shift[6] ), .ZN(new_n2225_));
  OAI21_X1   g1962(.A1(new_n1573_), .A2(new_n1580_), .B(new_n264_), .ZN(new_n2226_));
  NAND2_X1   g1963(.A1(new_n2225_), .A2(new_n2226_), .ZN(\result[78] ));
  OAI21_X1   g1964(.A1(new_n1589_), .A2(new_n1596_), .B(\shift[6] ), .ZN(new_n2228_));
  OAI21_X1   g1965(.A1(new_n1604_), .A2(new_n1611_), .B(new_n264_), .ZN(new_n2229_));
  NAND2_X1   g1966(.A1(new_n2228_), .A2(new_n2229_), .ZN(\result[79] ));
  OAI21_X1   g1967(.A1(new_n1616_), .A2(new_n1619_), .B(\shift[6] ), .ZN(new_n2231_));
  OAI21_X1   g1968(.A1(new_n1623_), .A2(new_n1626_), .B(new_n264_), .ZN(new_n2232_));
  NAND2_X1   g1969(.A1(new_n2231_), .A2(new_n2232_), .ZN(\result[80] ));
  OAI21_X1   g1970(.A1(new_n1631_), .A2(new_n1634_), .B(\shift[6] ), .ZN(new_n2234_));
  OAI21_X1   g1971(.A1(new_n1638_), .A2(new_n1641_), .B(new_n264_), .ZN(new_n2235_));
  NAND2_X1   g1972(.A1(new_n2234_), .A2(new_n2235_), .ZN(\result[81] ));
  OAI21_X1   g1973(.A1(new_n1646_), .A2(new_n1649_), .B(\shift[6] ), .ZN(new_n2237_));
  OAI21_X1   g1974(.A1(new_n1653_), .A2(new_n1656_), .B(new_n264_), .ZN(new_n2238_));
  NAND2_X1   g1975(.A1(new_n2237_), .A2(new_n2238_), .ZN(\result[82] ));
  OAI21_X1   g1976(.A1(new_n1661_), .A2(new_n1664_), .B(\shift[6] ), .ZN(new_n2240_));
  OAI21_X1   g1977(.A1(new_n1668_), .A2(new_n1671_), .B(new_n264_), .ZN(new_n2241_));
  NAND2_X1   g1978(.A1(new_n2240_), .A2(new_n2241_), .ZN(\result[83] ));
  OAI21_X1   g1979(.A1(new_n1676_), .A2(new_n1679_), .B(\shift[6] ), .ZN(new_n2243_));
  OAI21_X1   g1980(.A1(new_n1683_), .A2(new_n1686_), .B(new_n264_), .ZN(new_n2244_));
  NAND2_X1   g1981(.A1(new_n2243_), .A2(new_n2244_), .ZN(\result[84] ));
  OAI21_X1   g1982(.A1(new_n1691_), .A2(new_n1694_), .B(\shift[6] ), .ZN(new_n2246_));
  OAI21_X1   g1983(.A1(new_n1701_), .A2(new_n1698_), .B(new_n264_), .ZN(new_n2247_));
  NAND2_X1   g1984(.A1(new_n2246_), .A2(new_n2247_), .ZN(\result[85] ));
  OAI21_X1   g1985(.A1(new_n1706_), .A2(new_n1709_), .B(\shift[6] ), .ZN(new_n2249_));
  OAI21_X1   g1986(.A1(new_n1713_), .A2(new_n1716_), .B(new_n264_), .ZN(new_n2250_));
  NAND2_X1   g1987(.A1(new_n2249_), .A2(new_n2250_), .ZN(\result[86] ));
  OAI21_X1   g1988(.A1(new_n1726_), .A2(new_n1721_), .B(\shift[6] ), .ZN(new_n2252_));
  OAI21_X1   g1989(.A1(new_n1733_), .A2(new_n1730_), .B(new_n264_), .ZN(new_n2253_));
  NAND2_X1   g1990(.A1(new_n2252_), .A2(new_n2253_), .ZN(\result[87] ));
  OAI21_X1   g1991(.A1(new_n1738_), .A2(new_n1741_), .B(\shift[6] ), .ZN(new_n2255_));
  OAI21_X1   g1992(.A1(new_n1745_), .A2(new_n1748_), .B(new_n264_), .ZN(new_n2256_));
  NAND2_X1   g1993(.A1(new_n2255_), .A2(new_n2256_), .ZN(\result[88] ));
  OAI21_X1   g1994(.A1(new_n1753_), .A2(new_n1756_), .B(\shift[6] ), .ZN(new_n2258_));
  OAI21_X1   g1995(.A1(new_n1760_), .A2(new_n1763_), .B(new_n264_), .ZN(new_n2259_));
  NAND2_X1   g1996(.A1(new_n2259_), .A2(new_n2258_), .ZN(\result[89] ));
  OAI21_X1   g1997(.A1(new_n1768_), .A2(new_n1771_), .B(\shift[6] ), .ZN(new_n2261_));
  OAI21_X1   g1998(.A1(new_n1775_), .A2(new_n1778_), .B(new_n264_), .ZN(new_n2262_));
  NAND2_X1   g1999(.A1(new_n2261_), .A2(new_n2262_), .ZN(\result[90] ));
  OAI21_X1   g2000(.A1(new_n1783_), .A2(new_n1786_), .B(\shift[6] ), .ZN(new_n2264_));
  OAI21_X1   g2001(.A1(new_n1793_), .A2(new_n1790_), .B(new_n264_), .ZN(new_n2265_));
  NAND2_X1   g2002(.A1(new_n2264_), .A2(new_n2265_), .ZN(\result[91] ));
  OAI21_X1   g2003(.A1(new_n1798_), .A2(new_n1801_), .B(\shift[6] ), .ZN(new_n2267_));
  OAI21_X1   g2004(.A1(new_n1805_), .A2(new_n1808_), .B(new_n264_), .ZN(new_n2268_));
  NAND2_X1   g2005(.A1(new_n2267_), .A2(new_n2268_), .ZN(\result[92] ));
  OAI21_X1   g2006(.A1(new_n1816_), .A2(new_n1813_), .B(\shift[6] ), .ZN(new_n2270_));
  OAI21_X1   g2007(.A1(new_n1820_), .A2(new_n1823_), .B(new_n264_), .ZN(new_n2271_));
  NAND2_X1   g2008(.A1(new_n2270_), .A2(new_n2271_), .ZN(\result[93] ));
  OAI21_X1   g2009(.A1(new_n1828_), .A2(new_n1831_), .B(\shift[6] ), .ZN(new_n2273_));
  OAI21_X1   g2010(.A1(new_n1835_), .A2(new_n1838_), .B(new_n264_), .ZN(new_n2274_));
  NAND2_X1   g2011(.A1(new_n2273_), .A2(new_n2274_), .ZN(\result[94] ));
  OAI21_X1   g2012(.A1(new_n1843_), .A2(new_n1846_), .B(\shift[6] ), .ZN(new_n2276_));
  OAI21_X1   g2013(.A1(new_n1850_), .A2(new_n1853_), .B(new_n264_), .ZN(new_n2277_));
  NAND2_X1   g2014(.A1(new_n2276_), .A2(new_n2277_), .ZN(\result[95] ));
  OAI21_X1   g2015(.A1(new_n1856_), .A2(new_n1857_), .B(\shift[6] ), .ZN(new_n2279_));
  OAI21_X1   g2016(.A1(new_n1859_), .A2(new_n1860_), .B(new_n264_), .ZN(new_n2280_));
  NAND2_X1   g2017(.A1(new_n2279_), .A2(new_n2280_), .ZN(\result[96] ));
  OAI21_X1   g2018(.A1(new_n1866_), .A2(new_n1863_), .B(\shift[6] ), .ZN(new_n2282_));
  OAI21_X1   g2019(.A1(new_n1870_), .A2(new_n1873_), .B(new_n264_), .ZN(new_n2283_));
  NAND2_X1   g2020(.A1(new_n2282_), .A2(new_n2283_), .ZN(\result[97] ));
  OAI21_X1   g2021(.A1(new_n1876_), .A2(new_n1879_), .B(\shift[6] ), .ZN(new_n2285_));
  OAI21_X1   g2022(.A1(new_n1882_), .A2(new_n1885_), .B(new_n264_), .ZN(new_n2286_));
  NAND2_X1   g2023(.A1(new_n2285_), .A2(new_n2286_), .ZN(\result[98] ));
  OAI21_X1   g2024(.A1(new_n1890_), .A2(new_n1893_), .B(\shift[6] ), .ZN(new_n2288_));
  OAI21_X1   g2025(.A1(new_n1900_), .A2(new_n1897_), .B(new_n264_), .ZN(new_n2289_));
  NAND2_X1   g2026(.A1(new_n2289_), .A2(new_n2288_), .ZN(\result[99] ));
  OAI21_X1   g2027(.A1(new_n1903_), .A2(new_n1904_), .B(\shift[6] ), .ZN(new_n2291_));
  OAI21_X1   g2028(.A1(new_n1906_), .A2(new_n1907_), .B(new_n264_), .ZN(new_n2292_));
  NAND2_X1   g2029(.A1(new_n2291_), .A2(new_n2292_), .ZN(\result[100] ));
  OAI21_X1   g2030(.A1(new_n1910_), .A2(new_n1911_), .B(\shift[6] ), .ZN(new_n2294_));
  OAI21_X1   g2031(.A1(new_n1913_), .A2(new_n1914_), .B(new_n264_), .ZN(new_n2295_));
  NAND2_X1   g2032(.A1(new_n2294_), .A2(new_n2295_), .ZN(\result[101] ));
  OAI21_X1   g2033(.A1(new_n1917_), .A2(new_n1918_), .B(\shift[6] ), .ZN(new_n2297_));
  OAI21_X1   g2034(.A1(new_n1920_), .A2(new_n1921_), .B(new_n264_), .ZN(new_n2298_));
  NAND2_X1   g2035(.A1(new_n2297_), .A2(new_n2298_), .ZN(\result[102] ));
  OAI21_X1   g2036(.A1(new_n1925_), .A2(new_n1924_), .B(\shift[6] ), .ZN(new_n2300_));
  OAI21_X1   g2037(.A1(new_n1928_), .A2(new_n1927_), .B(new_n264_), .ZN(new_n2301_));
  NAND2_X1   g2038(.A1(new_n2300_), .A2(new_n2301_), .ZN(\result[103] ));
  OAI21_X1   g2039(.A1(new_n1931_), .A2(new_n1932_), .B(\shift[6] ), .ZN(new_n2303_));
  OAI21_X1   g2040(.A1(new_n1934_), .A2(new_n1935_), .B(new_n264_), .ZN(new_n2304_));
  NAND2_X1   g2041(.A1(new_n2303_), .A2(new_n2304_), .ZN(\result[104] ));
  OAI21_X1   g2042(.A1(new_n1939_), .A2(new_n1938_), .B(\shift[6] ), .ZN(new_n2306_));
  OAI21_X1   g2043(.A1(new_n1942_), .A2(new_n1941_), .B(new_n264_), .ZN(new_n2307_));
  NAND2_X1   g2044(.A1(new_n2306_), .A2(new_n2307_), .ZN(\result[105] ));
  OAI21_X1   g2045(.A1(new_n1945_), .A2(new_n1946_), .B(\shift[6] ), .ZN(new_n2309_));
  OAI21_X1   g2046(.A1(new_n1948_), .A2(new_n1949_), .B(new_n264_), .ZN(new_n2310_));
  NAND2_X1   g2047(.A1(new_n2309_), .A2(new_n2310_), .ZN(\result[106] ));
  OAI21_X1   g2048(.A1(new_n1952_), .A2(new_n1953_), .B(\shift[6] ), .ZN(new_n2312_));
  OAI21_X1   g2049(.A1(new_n1956_), .A2(new_n1955_), .B(new_n264_), .ZN(new_n2313_));
  NAND2_X1   g2050(.A1(new_n2312_), .A2(new_n2313_), .ZN(\result[107] ));
  OAI21_X1   g2051(.A1(new_n1959_), .A2(new_n1960_), .B(\shift[6] ), .ZN(new_n2315_));
  OAI21_X1   g2052(.A1(new_n1962_), .A2(new_n1963_), .B(new_n264_), .ZN(new_n2316_));
  NAND2_X1   g2053(.A1(new_n2315_), .A2(new_n2316_), .ZN(\result[108] ));
  OAI21_X1   g2054(.A1(new_n1966_), .A2(new_n1967_), .B(\shift[6] ), .ZN(new_n2318_));
  OAI21_X1   g2055(.A1(new_n1969_), .A2(new_n1970_), .B(new_n264_), .ZN(new_n2319_));
  NAND2_X1   g2056(.A1(new_n2319_), .A2(new_n2318_), .ZN(\result[109] ));
  OAI21_X1   g2057(.A1(new_n1973_), .A2(new_n1974_), .B(\shift[6] ), .ZN(new_n2321_));
  OAI21_X1   g2058(.A1(new_n1976_), .A2(new_n1977_), .B(new_n264_), .ZN(new_n2322_));
  NAND2_X1   g2059(.A1(new_n2321_), .A2(new_n2322_), .ZN(\result[110] ));
  OAI21_X1   g2060(.A1(new_n1980_), .A2(new_n1981_), .B(\shift[6] ), .ZN(new_n2324_));
  OAI21_X1   g2061(.A1(new_n1984_), .A2(new_n1983_), .B(new_n264_), .ZN(new_n2325_));
  NAND2_X1   g2062(.A1(new_n2325_), .A2(new_n2324_), .ZN(\result[111] ));
  OAI21_X1   g2063(.A1(new_n1987_), .A2(new_n1990_), .B(\shift[6] ), .ZN(new_n2327_));
  OAI21_X1   g2064(.A1(new_n1993_), .A2(new_n1996_), .B(new_n264_), .ZN(new_n2328_));
  NAND2_X1   g2065(.A1(new_n2327_), .A2(new_n2328_), .ZN(\result[112] ));
  OAI21_X1   g2066(.A1(new_n1999_), .A2(new_n2000_), .B(\shift[6] ), .ZN(new_n2330_));
  OAI21_X1   g2067(.A1(new_n2002_), .A2(new_n2003_), .B(new_n264_), .ZN(new_n2331_));
  NAND2_X1   g2068(.A1(new_n2331_), .A2(new_n2330_), .ZN(\result[113] ));
  OAI21_X1   g2069(.A1(new_n2006_), .A2(new_n2007_), .B(\shift[6] ), .ZN(new_n2333_));
  OAI21_X1   g2070(.A1(new_n2009_), .A2(new_n2010_), .B(new_n264_), .ZN(new_n2334_));
  NAND2_X1   g2071(.A1(new_n2333_), .A2(new_n2334_), .ZN(\result[114] ));
  OAI21_X1   g2072(.A1(new_n2014_), .A2(new_n2013_), .B(\shift[6] ), .ZN(new_n2336_));
  OAI21_X1   g2073(.A1(new_n2017_), .A2(new_n2016_), .B(new_n264_), .ZN(new_n2337_));
  NAND2_X1   g2074(.A1(new_n2337_), .A2(new_n2336_), .ZN(\result[115] ));
  OAI21_X1   g2075(.A1(new_n2022_), .A2(new_n2025_), .B(\shift[6] ), .ZN(new_n2339_));
  OAI21_X1   g2076(.A1(new_n2029_), .A2(new_n2032_), .B(new_n264_), .ZN(new_n2340_));
  NAND2_X1   g2077(.A1(new_n2339_), .A2(new_n2340_), .ZN(\result[116] ));
  OAI21_X1   g2078(.A1(new_n2040_), .A2(new_n2037_), .B(\shift[6] ), .ZN(new_n2342_));
  OAI21_X1   g2079(.A1(new_n2044_), .A2(new_n2047_), .B(new_n264_), .ZN(new_n2343_));
  NAND2_X1   g2080(.A1(new_n2343_), .A2(new_n2342_), .ZN(\result[117] ));
  OAI21_X1   g2081(.A1(new_n2052_), .A2(new_n2055_), .B(\shift[6] ), .ZN(new_n2345_));
  OAI21_X1   g2082(.A1(new_n2059_), .A2(new_n2062_), .B(new_n264_), .ZN(new_n2346_));
  NAND2_X1   g2083(.A1(new_n2345_), .A2(new_n2346_), .ZN(\result[118] ));
  OAI21_X1   g2084(.A1(new_n2070_), .A2(new_n2067_), .B(\shift[6] ), .ZN(new_n2348_));
  OAI21_X1   g2085(.A1(new_n2077_), .A2(new_n2074_), .B(new_n264_), .ZN(new_n2349_));
  NAND2_X1   g2086(.A1(new_n2349_), .A2(new_n2348_), .ZN(\result[119] ));
  OAI21_X1   g2087(.A1(new_n2082_), .A2(new_n2085_), .B(\shift[6] ), .ZN(new_n2351_));
  OAI21_X1   g2088(.A1(new_n2089_), .A2(new_n2092_), .B(new_n264_), .ZN(new_n2352_));
  NAND2_X1   g2089(.A1(new_n2351_), .A2(new_n2352_), .ZN(\result[120] ));
  OAI21_X1   g2090(.A1(new_n2097_), .A2(new_n2100_), .B(\shift[6] ), .ZN(new_n2354_));
  OAI21_X1   g2091(.A1(new_n2104_), .A2(new_n2107_), .B(new_n264_), .ZN(new_n2355_));
  NAND2_X1   g2092(.A1(new_n2355_), .A2(new_n2354_), .ZN(\result[121] ));
  OAI21_X1   g2093(.A1(new_n2111_), .A2(new_n2114_), .B(\shift[6] ), .ZN(new_n2357_));
  OAI21_X1   g2094(.A1(new_n2118_), .A2(new_n2119_), .B(new_n264_), .ZN(new_n2358_));
  NAND2_X1   g2095(.A1(new_n2358_), .A2(new_n2357_), .ZN(\result[122] ));
  OAI21_X1   g2096(.A1(new_n2126_), .A2(new_n2124_), .B(\shift[6] ), .ZN(new_n2360_));
  OAI21_X1   g2097(.A1(new_n2131_), .A2(new_n2130_), .B(new_n264_), .ZN(new_n2361_));
  NAND2_X1   g2098(.A1(new_n2361_), .A2(new_n2360_), .ZN(\result[123] ));
  OAI21_X1   g2099(.A1(new_n2135_), .A2(new_n2138_), .B(\shift[6] ), .ZN(new_n2363_));
  OAI21_X1   g2100(.A1(new_n2142_), .A2(new_n2143_), .B(new_n264_), .ZN(new_n2364_));
  NAND2_X1   g2101(.A1(new_n2364_), .A2(new_n2363_), .ZN(\result[124] ));
  OAI21_X1   g2102(.A1(new_n2148_), .A2(new_n2151_), .B(\shift[6] ), .ZN(new_n2366_));
  OAI21_X1   g2103(.A1(new_n2155_), .A2(new_n2156_), .B(new_n264_), .ZN(new_n2367_));
  NAND2_X1   g2104(.A1(new_n2367_), .A2(new_n2366_), .ZN(\result[125] ));
  OAI21_X1   g2105(.A1(new_n2160_), .A2(new_n2163_), .B(\shift[6] ), .ZN(new_n2369_));
  OAI21_X1   g2106(.A1(new_n2167_), .A2(new_n2168_), .B(new_n264_), .ZN(new_n2370_));
  NAND2_X1   g2107(.A1(new_n2370_), .A2(new_n2369_), .ZN(\result[126] ));
  OAI21_X1   g2108(.A1(new_n2172_), .A2(new_n2175_), .B(\shift[6] ), .ZN(new_n2372_));
  OAI21_X1   g2109(.A1(new_n2180_), .A2(new_n2179_), .B(new_n264_), .ZN(new_n2373_));
  NAND2_X1   g2110(.A1(new_n2373_), .A2(new_n2372_), .ZN(\result[127] ));
endmodule


