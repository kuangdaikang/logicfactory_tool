// Benchmark "source.pla" written by ABC on Fri Feb 25 15:13:04 2022

module x7dn  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29,
    v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43,
    v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57,
    v58, v59, v60, v61, v62, v63, v64, v65,
    \v66.0 , \v66.1 , \v66.2 , \v66.3 , \v66.4 , \v66.5 , \v66.6 , \v66.7 ,
    \v66.8 , \v66.9 , \v66.10 , \v66.11 , \v66.12 , \v66.13 , \v66.14   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28,
    v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42,
    v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56,
    v57, v58, v59, v60, v61, v62, v63, v64, v65;
  output \v66.0 , \v66.1 , \v66.2 , \v66.3 , \v66.4 , \v66.5 , \v66.6 ,
    \v66.7 , \v66.8 , \v66.9 , \v66.10 , \v66.11 , \v66.12 , \v66.13 ,
    \v66.14 ;
  wire new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_,
    new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_,
    new_n96_, new_n97_, new_n98_, new_n99_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n122_, new_n123_, new_n124_, new_n125_, new_n126_, new_n127_,
    new_n128_, new_n129_, new_n130_, new_n131_, new_n132_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_,
    new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_;
  assign new_n82_ = ~v0 & ~v1;
  assign new_n83_ = v6 & v8;
  assign new_n84_ = v9 & ~v10;
  assign new_n85_ = new_n83_ & new_n84_;
  assign new_n86_ = ~v4 & ~new_n85_;
  assign new_n87_ = v2 & v3;
  assign new_n88_ = ~v3 & v5;
  assign new_n89_ = ~new_n87_ & ~new_n88_;
  assign new_n90_ = ~new_n86_ & ~new_n89_;
  assign new_n91_ = v8 & v9;
  assign new_n92_ = ~v8 & ~v9;
  assign new_n93_ = ~new_n91_ & ~new_n92_;
  assign new_n94_ = ~v7 & ~new_n93_;
  assign new_n95_ = v7 & new_n84_;
  assign new_n96_ = ~new_n94_ & ~new_n95_;
  assign new_n97_ = ~v6 & ~new_n96_;
  assign new_n98_ = v5 & new_n97_;
  assign new_n99_ = ~new_n90_ & ~new_n98_;
  assign \v66.0  = ~new_n82_ & ~new_n99_;
  assign new_n101_ = v3 & v11;
  assign new_n102_ = ~v3 & v12;
  assign new_n103_ = ~new_n101_ & ~new_n102_;
  assign new_n104_ = ~new_n82_ & ~new_n103_;
  assign new_n105_ = v14 & ~v15;
  assign new_n106_ = ~v3 & new_n105_;
  assign new_n107_ = v14 & ~new_n106_;
  assign new_n108_ = v13 & ~new_n107_;
  assign new_n109_ = v3 & v16;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = ~v1 & ~new_n110_;
  assign new_n112_ = ~v0 & new_n111_;
  assign new_n113_ = ~new_n104_ & ~new_n112_;
  assign new_n114_ = ~new_n86_ & ~new_n113_;
  assign new_n115_ = v12 & ~new_n82_;
  assign new_n116_ = ~v1 & v13;
  assign new_n117_ = ~v0 & new_n116_;
  assign new_n118_ = ~new_n115_ & ~new_n117_;
  assign new_n119_ = ~new_n96_ & ~new_n118_;
  assign new_n120_ = ~v6 & new_n119_;
  assign \v66.1  = new_n114_ | new_n120_;
  assign new_n122_ = v3 & v17;
  assign new_n123_ = ~v3 & v18;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = ~new_n82_ & ~new_n124_;
  assign new_n126_ = v3 & v20;
  assign new_n127_ = v19 & ~new_n107_;
  assign new_n128_ = ~new_n126_ & ~new_n127_;
  assign new_n129_ = ~v1 & ~new_n128_;
  assign new_n130_ = ~v0 & new_n129_;
  assign new_n131_ = ~new_n125_ & ~new_n130_;
  assign new_n132_ = ~new_n86_ & ~new_n131_;
  assign new_n133_ = v18 & ~new_n82_;
  assign new_n134_ = ~v1 & v19;
  assign new_n135_ = ~v0 & new_n134_;
  assign new_n136_ = ~new_n133_ & ~new_n135_;
  assign new_n137_ = ~new_n96_ & ~new_n136_;
  assign new_n138_ = ~v6 & new_n137_;
  assign \v66.2  = new_n132_ | new_n138_;
  assign new_n140_ = v3 & v21;
  assign new_n141_ = ~v3 & v22;
  assign new_n142_ = ~new_n140_ & ~new_n141_;
  assign new_n143_ = ~new_n82_ & ~new_n142_;
  assign new_n144_ = v3 & v24;
  assign new_n145_ = v23 & ~new_n107_;
  assign new_n146_ = ~new_n144_ & ~new_n145_;
  assign new_n147_ = ~v1 & ~new_n146_;
  assign new_n148_ = ~v0 & new_n147_;
  assign new_n149_ = ~new_n143_ & ~new_n148_;
  assign new_n150_ = ~new_n86_ & ~new_n149_;
  assign new_n151_ = v22 & ~new_n82_;
  assign new_n152_ = ~v1 & v23;
  assign new_n153_ = ~v0 & new_n152_;
  assign new_n154_ = ~new_n151_ & ~new_n153_;
  assign new_n155_ = ~new_n96_ & ~new_n154_;
  assign new_n156_ = ~v6 & new_n155_;
  assign \v66.3  = new_n150_ | new_n156_;
  assign new_n158_ = v3 & v25;
  assign new_n159_ = ~v3 & v26;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~new_n82_ & ~new_n160_;
  assign new_n162_ = v3 & v28;
  assign new_n163_ = v27 & ~new_n107_;
  assign new_n164_ = ~new_n162_ & ~new_n163_;
  assign new_n165_ = ~v1 & ~new_n164_;
  assign new_n166_ = ~v0 & new_n165_;
  assign new_n167_ = ~new_n161_ & ~new_n166_;
  assign new_n168_ = ~new_n86_ & ~new_n167_;
  assign new_n169_ = v26 & ~new_n82_;
  assign new_n170_ = ~v1 & v27;
  assign new_n171_ = ~v0 & new_n170_;
  assign new_n172_ = ~new_n169_ & ~new_n171_;
  assign new_n173_ = ~new_n96_ & ~new_n172_;
  assign new_n174_ = ~v6 & new_n173_;
  assign \v66.4  = new_n168_ | new_n174_;
  assign new_n176_ = v3 & v29;
  assign new_n177_ = ~v3 & v30;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~new_n82_ & ~new_n178_;
  assign new_n180_ = v3 & v32;
  assign new_n181_ = v31 & ~new_n107_;
  assign new_n182_ = ~new_n180_ & ~new_n181_;
  assign new_n183_ = ~v1 & ~new_n182_;
  assign new_n184_ = ~v0 & new_n183_;
  assign new_n185_ = ~new_n179_ & ~new_n184_;
  assign new_n186_ = ~new_n86_ & ~new_n185_;
  assign new_n187_ = v30 & ~new_n82_;
  assign new_n188_ = ~v1 & v31;
  assign new_n189_ = ~v0 & new_n188_;
  assign new_n190_ = ~new_n187_ & ~new_n189_;
  assign new_n191_ = ~new_n96_ & ~new_n190_;
  assign new_n192_ = ~v6 & new_n191_;
  assign \v66.5  = new_n186_ | new_n192_;
  assign new_n194_ = v3 & v33;
  assign new_n195_ = ~v3 & v34;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = ~new_n82_ & ~new_n196_;
  assign new_n198_ = v3 & v36;
  assign new_n199_ = v35 & ~new_n107_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = ~v1 & ~new_n200_;
  assign new_n202_ = ~v0 & new_n201_;
  assign new_n203_ = ~new_n197_ & ~new_n202_;
  assign new_n204_ = ~new_n86_ & ~new_n203_;
  assign new_n205_ = v34 & ~new_n82_;
  assign new_n206_ = ~v1 & v35;
  assign new_n207_ = ~v0 & new_n206_;
  assign new_n208_ = ~new_n205_ & ~new_n207_;
  assign new_n209_ = ~new_n96_ & ~new_n208_;
  assign new_n210_ = ~v6 & new_n209_;
  assign \v66.6  = new_n204_ | new_n210_;
  assign new_n212_ = v3 & v37;
  assign new_n213_ = ~v3 & v38;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = ~new_n82_ & ~new_n214_;
  assign new_n216_ = ~v1 & ~new_n89_;
  assign new_n217_ = ~v0 & new_n216_;
  assign new_n218_ = ~new_n215_ & ~new_n217_;
  assign new_n219_ = ~new_n86_ & ~new_n218_;
  assign new_n220_ = v38 & ~new_n82_;
  assign new_n221_ = ~v1 & v5;
  assign new_n222_ = ~v0 & new_n221_;
  assign new_n223_ = ~new_n220_ & ~new_n222_;
  assign new_n224_ = ~new_n96_ & ~new_n223_;
  assign new_n225_ = ~v6 & new_n224_;
  assign \v66.7  = new_n219_ | new_n225_;
  assign new_n227_ = ~new_n86_ & ~new_n103_;
  assign new_n228_ = v12 & ~new_n96_;
  assign new_n229_ = ~v6 & new_n228_;
  assign new_n230_ = ~new_n227_ & ~new_n229_;
  assign new_n231_ = ~v1 & ~new_n230_;
  assign new_n232_ = ~v0 & new_n231_;
  assign new_n233_ = v45 & v46;
  assign new_n234_ = v47 & v48;
  assign new_n235_ = new_n233_ & new_n234_;
  assign new_n236_ = v49 & v50;
  assign new_n237_ = v51 & v52;
  assign new_n238_ = new_n236_ & new_n237_;
  assign new_n239_ = new_n235_ & new_n238_;
  assign new_n240_ = ~v45 & ~v46;
  assign new_n241_ = ~v47 & ~v48;
  assign new_n242_ = new_n240_ & new_n241_;
  assign new_n243_ = ~v49 & ~v50;
  assign new_n244_ = ~v52 & v53;
  assign new_n245_ = ~v51 & new_n244_;
  assign new_n246_ = new_n243_ & new_n245_;
  assign new_n247_ = new_n242_ & new_n246_;
  assign new_n248_ = ~new_n239_ & ~new_n247_;
  assign new_n249_ = ~v39 & ~new_n248_;
  assign new_n250_ = v46 & v47;
  assign new_n251_ = v45 & new_n250_;
  assign new_n252_ = v48 & v49;
  assign new_n253_ = v50 & v51;
  assign new_n254_ = new_n252_ & new_n253_;
  assign new_n255_ = new_n251_ & new_n254_;
  assign new_n256_ = v52 & ~new_n255_;
  assign new_n257_ = ~v46 & ~v47;
  assign new_n258_ = ~v45 & new_n257_;
  assign new_n259_ = ~v48 & ~v49;
  assign new_n260_ = ~v50 & ~v51;
  assign new_n261_ = new_n259_ & new_n260_;
  assign new_n262_ = new_n258_ & new_n261_;
  assign new_n263_ = v53 & ~new_n262_;
  assign new_n264_ = v53 & ~new_n263_;
  assign new_n265_ = ~v52 & ~new_n264_;
  assign new_n266_ = ~new_n256_ & ~new_n265_;
  assign new_n267_ = v39 & ~new_n266_;
  assign new_n268_ = ~new_n249_ & ~new_n267_;
  assign new_n269_ = ~v10 & ~new_n268_;
  assign new_n270_ = v7 & new_n269_;
  assign new_n271_ = v8 & v44;
  assign new_n272_ = ~v7 & new_n271_;
  assign new_n273_ = ~new_n270_ & ~new_n272_;
  assign new_n274_ = v9 & ~new_n273_;
  assign new_n275_ = v39 & v42;
  assign new_n276_ = ~v42 & v44;
  assign new_n277_ = ~new_n275_ & ~new_n276_;
  assign new_n278_ = ~v43 & ~new_n277_;
  assign new_n279_ = v41 & new_n278_;
  assign new_n280_ = ~v42 & v43;
  assign new_n281_ = v40 & new_n280_;
  assign new_n282_ = ~new_n279_ & ~new_n281_;
  assign new_n283_ = ~v9 & ~new_n282_;
  assign new_n284_ = ~v8 & new_n283_;
  assign new_n285_ = ~v7 & new_n284_;
  assign new_n286_ = ~new_n274_ & ~new_n285_;
  assign new_n287_ = ~v6 & ~new_n286_;
  assign new_n288_ = v4 & v39;
  assign new_n289_ = ~v7 & ~new_n268_;
  assign new_n290_ = v7 & v39;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = ~v10 & ~new_n291_;
  assign new_n293_ = v9 & new_n292_;
  assign new_n294_ = v8 & new_n293_;
  assign new_n295_ = v6 & new_n294_;
  assign new_n296_ = ~new_n288_ & ~new_n295_;
  assign new_n297_ = ~new_n287_ & new_n296_;
  assign new_n298_ = ~new_n82_ & ~new_n297_;
  assign \v66.8  = new_n232_ | new_n298_;
  assign new_n300_ = ~new_n86_ & ~new_n124_;
  assign new_n301_ = v18 & ~new_n96_;
  assign new_n302_ = ~v6 & new_n301_;
  assign new_n303_ = ~new_n300_ & ~new_n302_;
  assign new_n304_ = ~v1 & ~new_n303_;
  assign new_n305_ = ~v0 & new_n304_;
  assign new_n306_ = v10 & v56;
  assign new_n307_ = v3 & new_n306_;
  assign new_n308_ = ~v55 & ~new_n307_;
  assign new_n309_ = v8 & ~new_n308_;
  assign new_n310_ = ~v7 & new_n309_;
  assign new_n311_ = v46 & new_n234_;
  assign new_n312_ = new_n238_ & new_n311_;
  assign new_n313_ = new_n257_ & new_n259_;
  assign new_n314_ = new_n244_ & new_n260_;
  assign new_n315_ = new_n313_ & new_n314_;
  assign new_n316_ = ~new_n312_ & ~new_n315_;
  assign new_n317_ = ~v45 & ~new_n316_;
  assign new_n318_ = v49 & new_n253_;
  assign new_n319_ = new_n311_ & new_n318_;
  assign new_n320_ = v52 & ~new_n319_;
  assign new_n321_ = ~v46 & new_n241_;
  assign new_n322_ = ~v49 & new_n260_;
  assign new_n323_ = new_n321_ & new_n322_;
  assign new_n324_ = v53 & ~new_n323_;
  assign new_n325_ = v53 & ~new_n324_;
  assign new_n326_ = ~v52 & ~new_n325_;
  assign new_n327_ = ~new_n320_ & ~new_n326_;
  assign new_n328_ = v45 & ~new_n327_;
  assign new_n329_ = ~new_n317_ & ~new_n328_;
  assign new_n330_ = ~v10 & ~new_n329_;
  assign new_n331_ = v7 & new_n330_;
  assign new_n332_ = ~new_n310_ & ~new_n331_;
  assign new_n333_ = v9 & ~new_n332_;
  assign new_n334_ = v42 & v45;
  assign new_n335_ = ~v42 & v55;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = ~v43 & ~new_n336_;
  assign new_n338_ = v41 & new_n337_;
  assign new_n339_ = v43 & v54;
  assign new_n340_ = ~v42 & new_n339_;
  assign new_n341_ = ~new_n338_ & ~new_n340_;
  assign new_n342_ = ~v9 & ~new_n341_;
  assign new_n343_ = ~v8 & new_n342_;
  assign new_n344_ = ~v7 & new_n343_;
  assign new_n345_ = ~new_n333_ & ~new_n344_;
  assign new_n346_ = ~v6 & ~new_n345_;
  assign new_n347_ = ~v7 & ~new_n329_;
  assign new_n348_ = v7 & v45;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_ = ~v10 & ~new_n349_;
  assign new_n351_ = v9 & new_n350_;
  assign new_n352_ = v8 & new_n351_;
  assign new_n353_ = v6 & new_n352_;
  assign new_n354_ = v4 & v45;
  assign new_n355_ = ~new_n353_ & ~new_n354_;
  assign new_n356_ = ~new_n346_ & new_n355_;
  assign new_n357_ = ~new_n82_ & ~new_n356_;
  assign \v66.9  = new_n305_ | new_n357_;
  assign new_n359_ = ~new_n86_ & ~new_n142_;
  assign new_n360_ = v22 & ~new_n96_;
  assign new_n361_ = ~v6 & new_n360_;
  assign new_n362_ = ~new_n359_ & ~new_n361_;
  assign new_n363_ = ~v1 & ~new_n362_;
  assign new_n364_ = ~v0 & new_n363_;
  assign new_n365_ = ~v42 & ~v43;
  assign new_n366_ = v41 & new_n365_;
  assign new_n367_ = new_n92_ & new_n366_;
  assign new_n368_ = ~new_n91_ & ~new_n367_;
  assign new_n369_ = v16 & ~new_n368_;
  assign new_n370_ = v13 & new_n280_;
  assign new_n371_ = v41 & v42;
  assign new_n372_ = ~v43 & v46;
  assign new_n373_ = new_n371_ & new_n372_;
  assign new_n374_ = ~new_n370_ & ~new_n373_;
  assign new_n375_ = ~v9 & ~new_n374_;
  assign new_n376_ = ~v8 & new_n375_;
  assign new_n377_ = ~new_n369_ & ~new_n376_;
  assign new_n378_ = ~v7 & ~new_n377_;
  assign new_n379_ = v47 & new_n252_;
  assign new_n380_ = v50 & new_n237_;
  assign new_n381_ = new_n379_ & new_n380_;
  assign new_n382_ = ~v47 & new_n259_;
  assign new_n383_ = new_n314_ & new_n382_;
  assign new_n384_ = ~new_n381_ & ~new_n383_;
  assign new_n385_ = ~v46 & ~new_n384_;
  assign new_n386_ = new_n234_ & new_n318_;
  assign new_n387_ = v52 & ~new_n386_;
  assign new_n388_ = new_n241_ & new_n322_;
  assign new_n389_ = v53 & ~new_n388_;
  assign new_n390_ = v53 & ~new_n389_;
  assign new_n391_ = ~v52 & ~new_n390_;
  assign new_n392_ = ~new_n387_ & ~new_n391_;
  assign new_n393_ = v46 & ~new_n392_;
  assign new_n394_ = ~new_n385_ & ~new_n393_;
  assign new_n395_ = ~v10 & ~new_n394_;
  assign new_n396_ = v9 & new_n395_;
  assign new_n397_ = v7 & new_n396_;
  assign new_n398_ = ~new_n378_ & ~new_n397_;
  assign new_n399_ = ~v6 & ~new_n398_;
  assign new_n400_ = ~v7 & ~new_n394_;
  assign new_n401_ = v7 & v46;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign new_n403_ = ~v10 & ~new_n402_;
  assign new_n404_ = v9 & new_n403_;
  assign new_n405_ = v8 & new_n404_;
  assign new_n406_ = v6 & new_n405_;
  assign new_n407_ = v4 & v46;
  assign new_n408_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = ~new_n399_ & new_n408_;
  assign new_n410_ = ~new_n82_ & ~new_n409_;
  assign \v66.10  = new_n364_ | new_n410_;
  assign new_n412_ = ~new_n86_ & ~new_n160_;
  assign new_n413_ = v26 & ~new_n96_;
  assign new_n414_ = ~v6 & new_n413_;
  assign new_n415_ = ~new_n412_ & ~new_n414_;
  assign new_n416_ = ~v1 & ~new_n415_;
  assign new_n417_ = ~v0 & new_n416_;
  assign new_n418_ = v20 & ~new_n368_;
  assign new_n419_ = v19 & new_n280_;
  assign new_n420_ = ~v43 & v47;
  assign new_n421_ = new_n371_ & new_n420_;
  assign new_n422_ = ~new_n419_ & ~new_n421_;
  assign new_n423_ = ~v9 & ~new_n422_;
  assign new_n424_ = ~v8 & new_n423_;
  assign new_n425_ = ~new_n418_ & ~new_n424_;
  assign new_n426_ = ~v7 & ~new_n425_;
  assign new_n427_ = new_n252_ & new_n380_;
  assign new_n428_ = ~v48 & new_n243_;
  assign new_n429_ = new_n245_ & new_n428_;
  assign new_n430_ = ~new_n427_ & ~new_n429_;
  assign new_n431_ = ~v47 & ~new_n430_;
  assign new_n432_ = v52 & ~new_n254_;
  assign new_n433_ = v53 & ~new_n261_;
  assign new_n434_ = v53 & ~new_n433_;
  assign new_n435_ = ~v52 & ~new_n434_;
  assign new_n436_ = ~new_n432_ & ~new_n435_;
  assign new_n437_ = v47 & ~new_n436_;
  assign new_n438_ = ~new_n431_ & ~new_n437_;
  assign new_n439_ = ~v10 & ~new_n438_;
  assign new_n440_ = v9 & new_n439_;
  assign new_n441_ = v7 & new_n440_;
  assign new_n442_ = ~new_n426_ & ~new_n441_;
  assign new_n443_ = ~v6 & ~new_n442_;
  assign new_n444_ = v4 & v47;
  assign new_n445_ = v7 & v47;
  assign new_n446_ = ~v7 & ~new_n438_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = ~v10 & ~new_n447_;
  assign new_n449_ = v9 & new_n448_;
  assign new_n450_ = v8 & new_n449_;
  assign new_n451_ = v6 & new_n450_;
  assign new_n452_ = ~new_n444_ & ~new_n451_;
  assign new_n453_ = ~new_n443_ & new_n452_;
  assign new_n454_ = ~new_n82_ & ~new_n453_;
  assign \v66.11  = new_n417_ | new_n454_;
  assign new_n456_ = ~new_n86_ & ~new_n178_;
  assign new_n457_ = v30 & ~new_n96_;
  assign new_n458_ = ~v6 & new_n457_;
  assign new_n459_ = ~new_n456_ & ~new_n458_;
  assign new_n460_ = ~v1 & ~new_n459_;
  assign new_n461_ = ~v0 & new_n460_;
  assign new_n462_ = v24 & ~new_n368_;
  assign new_n463_ = v23 & new_n280_;
  assign new_n464_ = ~v43 & v48;
  assign new_n465_ = new_n371_ & new_n464_;
  assign new_n466_ = ~new_n463_ & ~new_n465_;
  assign new_n467_ = ~v9 & ~new_n466_;
  assign new_n468_ = ~v8 & new_n467_;
  assign new_n469_ = ~new_n462_ & ~new_n468_;
  assign new_n470_ = ~v7 & ~new_n469_;
  assign new_n471_ = ~new_n238_ & ~new_n246_;
  assign new_n472_ = ~v48 & ~new_n471_;
  assign new_n473_ = v52 & ~new_n318_;
  assign new_n474_ = v53 & ~new_n322_;
  assign new_n475_ = v53 & ~new_n474_;
  assign new_n476_ = ~v52 & ~new_n475_;
  assign new_n477_ = ~new_n473_ & ~new_n476_;
  assign new_n478_ = v48 & ~new_n477_;
  assign new_n479_ = ~new_n472_ & ~new_n478_;
  assign new_n480_ = ~v10 & ~new_n479_;
  assign new_n481_ = v9 & new_n480_;
  assign new_n482_ = v7 & new_n481_;
  assign new_n483_ = ~new_n470_ & ~new_n482_;
  assign new_n484_ = ~v6 & ~new_n483_;
  assign new_n485_ = v4 & v48;
  assign new_n486_ = v7 & v48;
  assign new_n487_ = ~v7 & ~new_n479_;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = ~v10 & ~new_n488_;
  assign new_n490_ = v9 & new_n489_;
  assign new_n491_ = v8 & new_n490_;
  assign new_n492_ = v6 & new_n491_;
  assign new_n493_ = ~new_n485_ & ~new_n492_;
  assign new_n494_ = ~new_n484_ & new_n493_;
  assign new_n495_ = ~new_n82_ & ~new_n494_;
  assign \v66.12  = new_n461_ | new_n495_;
  assign new_n497_ = ~new_n86_ & ~new_n196_;
  assign new_n498_ = v34 & ~new_n96_;
  assign new_n499_ = ~v6 & new_n498_;
  assign new_n500_ = ~new_n497_ & ~new_n499_;
  assign new_n501_ = ~v1 & ~new_n500_;
  assign new_n502_ = ~v0 & new_n501_;
  assign new_n503_ = v28 & ~new_n368_;
  assign new_n504_ = v27 & new_n280_;
  assign new_n505_ = ~v43 & v49;
  assign new_n506_ = v43 & v57;
  assign new_n507_ = v58 & ~v59;
  assign new_n508_ = new_n506_ & new_n507_;
  assign new_n509_ = ~v60 & ~v61;
  assign new_n510_ = ~v62 & ~v63;
  assign new_n511_ = new_n509_ & new_n510_;
  assign new_n512_ = new_n508_ & new_n511_;
  assign new_n513_ = ~new_n505_ & ~new_n512_;
  assign new_n514_ = v42 & ~new_n513_;
  assign new_n515_ = v41 & new_n514_;
  assign new_n516_ = ~new_n504_ & ~new_n515_;
  assign new_n517_ = ~v9 & ~new_n516_;
  assign new_n518_ = ~v8 & new_n517_;
  assign new_n519_ = ~new_n503_ & ~new_n518_;
  assign new_n520_ = ~v7 & ~new_n519_;
  assign new_n521_ = ~new_n314_ & ~new_n380_;
  assign new_n522_ = ~v49 & ~new_n521_;
  assign new_n523_ = v52 & ~new_n253_;
  assign new_n524_ = v53 & ~new_n260_;
  assign new_n525_ = v53 & ~new_n524_;
  assign new_n526_ = ~v52 & ~new_n525_;
  assign new_n527_ = ~new_n523_ & ~new_n526_;
  assign new_n528_ = v49 & ~new_n527_;
  assign new_n529_ = ~new_n522_ & ~new_n528_;
  assign new_n530_ = ~v10 & ~new_n529_;
  assign new_n531_ = v9 & new_n530_;
  assign new_n532_ = v7 & new_n531_;
  assign new_n533_ = ~new_n520_ & ~new_n532_;
  assign new_n534_ = ~v6 & ~new_n533_;
  assign new_n535_ = v4 & v49;
  assign new_n536_ = v7 & v49;
  assign new_n537_ = ~v7 & ~new_n529_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~v10 & ~new_n538_;
  assign new_n540_ = v9 & new_n539_;
  assign new_n541_ = v8 & new_n540_;
  assign new_n542_ = v6 & new_n541_;
  assign new_n543_ = ~new_n535_ & ~new_n542_;
  assign new_n544_ = ~new_n534_ & new_n543_;
  assign new_n545_ = ~new_n82_ & ~new_n544_;
  assign \v66.13  = new_n502_ | new_n545_;
  assign new_n547_ = ~new_n86_ & ~new_n214_;
  assign new_n548_ = v38 & ~new_n96_;
  assign new_n549_ = ~v6 & new_n548_;
  assign new_n550_ = ~new_n547_ & ~new_n549_;
  assign new_n551_ = ~v1 & ~new_n550_;
  assign new_n552_ = ~v0 & new_n551_;
  assign new_n553_ = v32 & ~new_n368_;
  assign new_n554_ = v31 & new_n280_;
  assign new_n555_ = ~v43 & v50;
  assign new_n556_ = v63 & v64;
  assign new_n557_ = ~v58 & new_n556_;
  assign new_n558_ = ~v63 & v65;
  assign new_n559_ = v58 & new_n558_;
  assign new_n560_ = ~new_n557_ & ~new_n559_;
  assign new_n561_ = ~v62 & ~new_n560_;
  assign new_n562_ = ~v61 & new_n561_;
  assign new_n563_ = ~v60 & new_n562_;
  assign new_n564_ = ~v59 & new_n563_;
  assign new_n565_ = v43 & new_n564_;
  assign new_n566_ = ~new_n555_ & ~new_n565_;
  assign new_n567_ = v42 & ~new_n566_;
  assign new_n568_ = v41 & new_n567_;
  assign new_n569_ = ~new_n554_ & ~new_n568_;
  assign new_n570_ = ~v9 & ~new_n569_;
  assign new_n571_ = ~v8 & new_n570_;
  assign new_n572_ = ~new_n553_ & ~new_n571_;
  assign new_n573_ = ~v7 & ~new_n572_;
  assign new_n574_ = ~new_n237_ & ~new_n245_;
  assign new_n575_ = ~v50 & ~new_n574_;
  assign new_n576_ = v51 & v53;
  assign new_n577_ = v53 & ~new_n576_;
  assign new_n578_ = ~v52 & ~new_n577_;
  assign new_n579_ = ~v51 & v52;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = v50 & ~new_n580_;
  assign new_n582_ = ~new_n575_ & ~new_n581_;
  assign new_n583_ = ~v10 & ~new_n582_;
  assign new_n584_ = v9 & new_n583_;
  assign new_n585_ = v7 & new_n584_;
  assign new_n586_ = ~new_n573_ & ~new_n585_;
  assign new_n587_ = ~v6 & ~new_n586_;
  assign new_n588_ = v4 & v50;
  assign new_n589_ = v7 & v50;
  assign new_n590_ = ~v7 & ~new_n582_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~v10 & ~new_n591_;
  assign new_n593_ = v9 & new_n592_;
  assign new_n594_ = v8 & new_n593_;
  assign new_n595_ = v6 & new_n594_;
  assign new_n596_ = ~new_n588_ & ~new_n595_;
  assign new_n597_ = ~new_n587_ & new_n596_;
  assign new_n598_ = ~new_n82_ & ~new_n597_;
  assign \v66.14  = new_n552_ | new_n598_;
endmodule


