// Benchmark "c5315.blif" written by ABC on Fri Feb 25 15:12:33 2022

module c5315  ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire new_n310_, new_n311_, new_n312_, new_n314_, new_n315_, new_n316_,
    new_n318_, new_n319_, new_n320_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_,
    new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_,
    new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_,
    new_n1039_, new_n1040_, new_n1042_, new_n1043_, new_n1044_, new_n1045_,
    new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1296_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1308_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1349_, new_n1350_, new_n1351_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_,
    new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_,
    new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_,
    new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_,
    new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_,
    new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_,
    new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_,
    new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_,
    new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_,
    new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_,
    new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_,
    new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_,
    new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_,
    new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_,
    new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_,
    new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_,
    new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_,
    new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_;
  assign G601 = G552 & G562;
  assign G810 = G141 & G145;
  assign G634 = G1 & G373;
  assign G815 = G136 & ~G3173;
  assign G845 = ~G27 | G2824;
  assign G847 = ~G386 | ~G556;
  assign G809 = ~G27 | ~G31;
  assign G656 = ~G140 | G809;
  assign new_n310_ = G87 & G2358;
  assign new_n311_ = G86 & ~G2358;
  assign new_n312_ = ~new_n310_ & ~new_n311_;
  assign G636 = G809 | new_n312_;
  assign new_n314_ = G34 & G2358;
  assign new_n315_ = G88 & ~G2358;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign G704 = G809 | new_n316_;
  assign new_n318_ = G83 & G2358;
  assign new_n319_ = G83 & ~G2358;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign G820 = G809 | new_n320_;
  assign new_n322_ = G24 & ~G2358;
  assign new_n323_ = ~G809 & new_n322_;
  assign new_n324_ = G25 & G2358;
  assign new_n325_ = ~G809 & new_n324_;
  assign new_n326_ = ~G2358 & G809;
  assign new_n327_ = G2358 & G809;
  assign new_n328_ = ~new_n323_ & ~new_n325_;
  assign new_n329_ = ~new_n326_ & ~new_n327_;
  assign new_n330_ = new_n328_ & new_n329_;
  assign G639 = G141 & ~new_n330_;
  assign new_n332_ = G26 & ~G2358;
  assign new_n333_ = ~G809 & new_n332_;
  assign new_n334_ = G81 & G2358;
  assign new_n335_ = ~G809 & new_n334_;
  assign new_n336_ = ~new_n333_ & ~new_n335_;
  assign new_n337_ = new_n329_ & new_n336_;
  assign G673 = G141 & ~new_n337_;
  assign new_n339_ = G79 & ~G2358;
  assign new_n340_ = ~G809 & new_n339_;
  assign new_n341_ = G23 & G2358;
  assign new_n342_ = ~G809 & new_n341_;
  assign new_n343_ = ~new_n340_ & ~new_n342_;
  assign new_n344_ = new_n329_ & new_n343_;
  assign G707 = G141 & ~new_n344_;
  assign new_n346_ = G82 & ~G2358;
  assign new_n347_ = ~G809 & new_n346_;
  assign new_n348_ = G80 & G2358;
  assign new_n349_ = ~G809 & new_n348_;
  assign new_n350_ = ~new_n347_ & ~new_n349_;
  assign new_n351_ = new_n329_ & new_n350_;
  assign G715 = G141 & ~new_n351_;
  assign new_n353_ = G248 & G490;
  assign new_n354_ = G316 & new_n353_;
  assign new_n355_ = G251 & G490;
  assign new_n356_ = ~G316 & new_n355_;
  assign new_n357_ = ~new_n354_ & ~new_n356_;
  assign new_n358_ = G242 & G316;
  assign new_n359_ = G254 & ~G316;
  assign new_n360_ = ~new_n358_ & ~new_n359_;
  assign new_n361_ = ~G490 & new_n360_;
  assign new_n362_ = new_n357_ & ~new_n361_;
  assign new_n363_ = G248 & G479;
  assign new_n364_ = G308 & new_n363_;
  assign new_n365_ = G251 & G479;
  assign new_n366_ = ~G308 & new_n365_;
  assign new_n367_ = ~new_n364_ & ~new_n366_;
  assign new_n368_ = G242 & G308;
  assign new_n369_ = G254 & ~G308;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = ~G479 & new_n370_;
  assign new_n372_ = new_n367_ & ~new_n371_;
  assign new_n373_ = G248 & G302;
  assign new_n374_ = G251 & ~G302;
  assign new_n375_ = ~new_n373_ & ~new_n374_;
  assign new_n376_ = G242 & G293;
  assign new_n377_ = G254 & ~G293;
  assign new_n378_ = ~new_n376_ & ~new_n377_;
  assign new_n379_ = ~new_n362_ & ~new_n372_;
  assign new_n380_ = ~new_n375_ & new_n379_;
  assign new_n381_ = new_n378_ & new_n380_;
  assign new_n382_ = G534 & ~G3552;
  assign new_n383_ = G351 & new_n382_;
  assign new_n384_ = G534 & ~G3550;
  assign new_n385_ = ~G351 & new_n384_;
  assign new_n386_ = ~new_n383_ & ~new_n385_;
  assign new_n387_ = G351 & ~G3546;
  assign new_n388_ = ~G351 & ~G3548;
  assign new_n389_ = ~new_n387_ & ~new_n388_;
  assign new_n390_ = ~G534 & new_n389_;
  assign new_n391_ = new_n386_ & ~new_n390_;
  assign new_n392_ = G523 & ~G3552;
  assign new_n393_ = G341 & new_n392_;
  assign new_n394_ = G523 & ~G3550;
  assign new_n395_ = ~G341 & new_n394_;
  assign new_n396_ = ~new_n393_ & ~new_n395_;
  assign new_n397_ = G341 & ~G3546;
  assign new_n398_ = ~G341 & ~G3548;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = ~G523 & new_n399_;
  assign new_n401_ = new_n396_ & ~new_n400_;
  assign new_n402_ = G514 & ~G3552;
  assign new_n403_ = ~G514 & G3546;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = G503 & ~G3552;
  assign new_n406_ = G324 & new_n405_;
  assign new_n407_ = G503 & ~G3550;
  assign new_n408_ = ~G324 & new_n407_;
  assign new_n409_ = ~new_n406_ & ~new_n408_;
  assign new_n410_ = G324 & ~G3546;
  assign new_n411_ = ~G324 & ~G3548;
  assign new_n412_ = ~new_n410_ & ~new_n411_;
  assign new_n413_ = ~G503 & new_n412_;
  assign new_n414_ = new_n409_ & ~new_n413_;
  assign new_n415_ = ~new_n391_ & ~new_n401_;
  assign new_n416_ = ~new_n404_ & new_n415_;
  assign new_n417_ = ~new_n414_ & new_n416_;
  assign new_n418_ = G248 & G361;
  assign new_n419_ = G251 & ~G361;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = new_n381_ & new_n417_;
  assign G598 = ~new_n420_ & new_n421_;
  assign new_n423_ = G435 & ~G3552;
  assign new_n424_ = G234 & new_n423_;
  assign new_n425_ = G435 & ~G3550;
  assign new_n426_ = ~G234 & new_n425_;
  assign new_n427_ = ~new_n424_ & ~new_n426_;
  assign new_n428_ = G234 & ~G3546;
  assign new_n429_ = ~G234 & ~G3548;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = ~G435 & new_n430_;
  assign new_n432_ = new_n427_ & ~new_n431_;
  assign new_n433_ = G422 & ~G3552;
  assign new_n434_ = G226 & new_n433_;
  assign new_n435_ = G422 & ~G3550;
  assign new_n436_ = ~G226 & new_n435_;
  assign new_n437_ = ~new_n434_ & ~new_n436_;
  assign new_n438_ = G226 & ~G3546;
  assign new_n439_ = ~G226 & ~G3548;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~G422 & new_n440_;
  assign new_n442_ = new_n437_ & ~new_n441_;
  assign new_n443_ = G468 & ~G3552;
  assign new_n444_ = G218 & new_n443_;
  assign new_n445_ = G468 & ~G3550;
  assign new_n446_ = ~G218 & new_n445_;
  assign new_n447_ = ~new_n444_ & ~new_n446_;
  assign new_n448_ = G218 & ~G3546;
  assign new_n449_ = ~G218 & ~G3548;
  assign new_n450_ = ~new_n448_ & ~new_n449_;
  assign new_n451_ = ~G468 & new_n450_;
  assign new_n452_ = new_n447_ & ~new_n451_;
  assign new_n453_ = G457 & ~G3552;
  assign new_n454_ = G210 & new_n453_;
  assign new_n455_ = G457 & ~G3550;
  assign new_n456_ = ~G210 & new_n455_;
  assign new_n457_ = ~new_n454_ & ~new_n456_;
  assign new_n458_ = G210 & ~G3546;
  assign new_n459_ = ~G210 & ~G3548;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~G457 & new_n460_;
  assign new_n462_ = new_n457_ & ~new_n461_;
  assign new_n463_ = ~new_n432_ & ~new_n442_;
  assign new_n464_ = ~new_n452_ & new_n463_;
  assign new_n465_ = ~new_n462_ & new_n464_;
  assign new_n466_ = G374 & ~G3552;
  assign new_n467_ = G281 & new_n466_;
  assign new_n468_ = G374 & ~G3550;
  assign new_n469_ = ~G281 & new_n468_;
  assign new_n470_ = ~new_n467_ & ~new_n469_;
  assign new_n471_ = G281 & ~G3546;
  assign new_n472_ = ~G281 & ~G3548;
  assign new_n473_ = ~new_n471_ & ~new_n472_;
  assign new_n474_ = ~G374 & new_n473_;
  assign new_n475_ = new_n470_ & ~new_n474_;
  assign new_n476_ = G411 & ~G3552;
  assign new_n477_ = G273 & new_n476_;
  assign new_n478_ = G411 & ~G3550;
  assign new_n479_ = ~G273 & new_n478_;
  assign new_n480_ = ~new_n477_ & ~new_n479_;
  assign new_n481_ = G273 & ~G3546;
  assign new_n482_ = ~G273 & ~G3548;
  assign new_n483_ = ~new_n481_ & ~new_n482_;
  assign new_n484_ = ~G411 & new_n483_;
  assign new_n485_ = new_n480_ & ~new_n484_;
  assign new_n486_ = G400 & ~G3552;
  assign new_n487_ = G265 & new_n486_;
  assign new_n488_ = G400 & ~G3550;
  assign new_n489_ = ~G265 & new_n488_;
  assign new_n490_ = ~new_n487_ & ~new_n489_;
  assign new_n491_ = G265 & ~G3546;
  assign new_n492_ = ~G265 & ~G3548;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = ~G400 & new_n493_;
  assign new_n495_ = new_n490_ & ~new_n494_;
  assign new_n496_ = G389 & ~G3552;
  assign new_n497_ = G257 & new_n496_;
  assign new_n498_ = G389 & ~G3550;
  assign new_n499_ = ~G257 & new_n498_;
  assign new_n500_ = ~new_n497_ & ~new_n499_;
  assign new_n501_ = G257 & ~G3546;
  assign new_n502_ = ~G257 & ~G3548;
  assign new_n503_ = ~new_n501_ & ~new_n502_;
  assign new_n504_ = ~G389 & new_n503_;
  assign new_n505_ = new_n500_ & ~new_n504_;
  assign new_n506_ = ~new_n475_ & ~new_n485_;
  assign new_n507_ = ~new_n495_ & new_n506_;
  assign new_n508_ = ~new_n505_ & new_n507_;
  assign new_n509_ = G248 & G446;
  assign new_n510_ = G206 & new_n509_;
  assign new_n511_ = G251 & G446;
  assign new_n512_ = ~G206 & new_n511_;
  assign new_n513_ = ~new_n510_ & ~new_n512_;
  assign new_n514_ = G206 & G242;
  assign new_n515_ = ~G206 & G254;
  assign new_n516_ = ~new_n514_ & ~new_n515_;
  assign new_n517_ = ~G446 & new_n516_;
  assign new_n518_ = new_n513_ & ~new_n517_;
  assign new_n519_ = new_n465_ & new_n508_;
  assign G610 = ~new_n518_ & new_n519_;
  assign new_n521_ = G226 & ~G335;
  assign new_n522_ = G233 & G335;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign new_n524_ = ~G422 & ~new_n523_;
  assign new_n525_ = G422 & new_n523_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = G218 & ~G335;
  assign new_n528_ = G225 & G335;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_ = ~G468 & ~new_n529_;
  assign new_n531_ = G468 & new_n529_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = G210 & ~G335;
  assign new_n534_ = G217 & G335;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~G457 & ~new_n535_;
  assign new_n537_ = G457 & new_n535_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = G206 & ~G335;
  assign new_n540_ = G209 & G335;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = ~G446 & ~new_n541_;
  assign new_n543_ = G446 & new_n541_;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = ~new_n526_ & ~new_n532_;
  assign new_n546_ = ~new_n538_ & new_n545_;
  assign new_n547_ = ~new_n544_ & new_n546_;
  assign new_n548_ = G281 & ~G335;
  assign new_n549_ = G288 & G335;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = ~G374 & ~new_n550_;
  assign new_n552_ = G374 & new_n550_;
  assign new_n553_ = ~new_n551_ & ~new_n552_;
  assign new_n554_ = G273 & ~G335;
  assign new_n555_ = G280 & G335;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = ~G411 & ~new_n556_;
  assign new_n558_ = G411 & new_n556_;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = G265 & ~G335;
  assign new_n561_ = G272 & G335;
  assign new_n562_ = ~new_n560_ & ~new_n561_;
  assign new_n563_ = ~G400 & ~new_n562_;
  assign new_n564_ = G400 & new_n562_;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = G257 & ~G335;
  assign new_n567_ = G264 & G335;
  assign new_n568_ = ~new_n566_ & ~new_n567_;
  assign new_n569_ = ~G389 & ~new_n568_;
  assign new_n570_ = G389 & new_n568_;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign new_n572_ = G234 & ~G335;
  assign new_n573_ = G241 & G335;
  assign new_n574_ = ~new_n572_ & ~new_n573_;
  assign new_n575_ = ~G435 & ~new_n574_;
  assign new_n576_ = G435 & new_n574_;
  assign new_n577_ = ~new_n575_ & ~new_n576_;
  assign new_n578_ = ~new_n553_ & ~new_n559_;
  assign new_n579_ = ~new_n565_ & new_n578_;
  assign new_n580_ = ~new_n571_ & new_n579_;
  assign new_n581_ = ~new_n577_ & new_n580_;
  assign G588 = new_n547_ & new_n581_;
  assign new_n583_ = G302 & ~G332;
  assign new_n584_ = G307 & G332;
  assign new_n585_ = ~new_n583_ & ~new_n584_;
  assign new_n586_ = G316 & ~G332;
  assign new_n587_ = G323 & G332;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = G490 & new_n588_;
  assign new_n590_ = ~G490 & ~new_n588_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = G308 & ~G332;
  assign new_n593_ = G315 & G332;
  assign new_n594_ = ~new_n592_ & ~new_n593_;
  assign new_n595_ = G479 & new_n594_;
  assign new_n596_ = ~G479 & ~new_n594_;
  assign new_n597_ = ~new_n595_ & ~new_n596_;
  assign new_n598_ = G293 & ~G332;
  assign new_n599_ = G299 & G332;
  assign new_n600_ = ~new_n598_ & ~new_n599_;
  assign new_n601_ = new_n585_ & ~new_n591_;
  assign new_n602_ = ~new_n597_ & new_n601_;
  assign new_n603_ = new_n600_ & new_n602_;
  assign new_n604_ = G332 & G338;
  assign new_n605_ = G332 & ~new_n604_;
  assign new_n606_ = G514 & new_n605_;
  assign new_n607_ = ~G514 & ~new_n605_;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = ~G332 & G361;
  assign new_n610_ = G332 & G366;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = ~G332 & G341;
  assign new_n613_ = G332 & G348;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = G523 & new_n614_;
  assign new_n616_ = ~G523 & ~new_n614_;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = G324 & ~G332;
  assign new_n619_ = G331 & G332;
  assign new_n620_ = ~new_n618_ & ~new_n619_;
  assign new_n621_ = G503 & new_n620_;
  assign new_n622_ = ~G503 & ~new_n620_;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_ = ~G332 & G351;
  assign new_n625_ = G332 & G358;
  assign new_n626_ = ~new_n624_ & ~new_n625_;
  assign new_n627_ = G534 & new_n626_;
  assign new_n628_ = ~G534 & ~new_n626_;
  assign new_n629_ = ~new_n627_ & ~new_n628_;
  assign new_n630_ = ~new_n608_ & new_n611_;
  assign new_n631_ = ~new_n617_ & new_n630_;
  assign new_n632_ = ~new_n623_ & new_n631_;
  assign new_n633_ = ~new_n629_ & new_n632_;
  assign G615 = new_n603_ & new_n633_;
  assign new_n635_ = ~new_n591_ & ~new_n597_;
  assign new_n636_ = new_n585_ & new_n635_;
  assign new_n637_ = new_n600_ & new_n636_;
  assign new_n638_ = new_n611_ & ~new_n629_;
  assign new_n639_ = ~new_n617_ & new_n638_;
  assign new_n640_ = ~new_n608_ & new_n639_;
  assign new_n641_ = ~new_n623_ & new_n640_;
  assign G626 = new_n637_ & new_n641_;
  assign new_n643_ = ~new_n526_ & ~new_n538_;
  assign new_n644_ = ~new_n532_ & new_n643_;
  assign new_n645_ = ~new_n544_ & new_n644_;
  assign new_n646_ = ~new_n553_ & ~new_n571_;
  assign new_n647_ = ~new_n565_ & new_n646_;
  assign new_n648_ = ~new_n577_ & new_n647_;
  assign new_n649_ = ~new_n559_ & new_n648_;
  assign G632 = new_n645_ & new_n649_;
  assign new_n651_ = ~G308 & G316;
  assign new_n652_ = G308 & ~G316;
  assign new_n653_ = ~new_n651_ & ~new_n652_;
  assign new_n654_ = ~G293 & G302;
  assign new_n655_ = G293 & ~G302;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = ~new_n653_ & new_n656_;
  assign new_n658_ = new_n653_ & ~new_n656_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~G361 & G369;
  assign new_n661_ = G361 & ~G369;
  assign new_n662_ = ~new_n660_ & ~new_n661_;
  assign new_n663_ = ~G341 & G351;
  assign new_n664_ = G341 & ~G351;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = ~new_n662_ & new_n665_;
  assign new_n667_ = G324 & new_n666_;
  assign new_n668_ = new_n662_ & new_n665_;
  assign new_n669_ = ~G324 & new_n668_;
  assign new_n670_ = ~new_n667_ & ~new_n669_;
  assign new_n671_ = new_n662_ & ~new_n665_;
  assign new_n672_ = G324 & new_n671_;
  assign new_n673_ = ~new_n662_ & ~new_n665_;
  assign new_n674_ = ~G324 & new_n673_;
  assign new_n675_ = ~new_n672_ & ~new_n674_;
  assign new_n676_ = new_n670_ & new_n675_;
  assign new_n677_ = ~new_n659_ & new_n676_;
  assign new_n678_ = new_n659_ & ~new_n676_;
  assign G1002 = new_n677_ | new_n678_;
  assign new_n680_ = ~G218 & G226;
  assign new_n681_ = G218 & ~G226;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~G206 & G210;
  assign new_n684_ = G206 & ~G210;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign new_n686_ = ~new_n682_ & new_n685_;
  assign new_n687_ = new_n682_ & ~new_n685_;
  assign new_n688_ = ~new_n686_ & ~new_n687_;
  assign new_n689_ = ~G281 & G289;
  assign new_n690_ = G281 & ~G289;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = ~G265 & G273;
  assign new_n693_ = G265 & ~G273;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = ~G234 & G257;
  assign new_n696_ = G234 & ~G257;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~new_n691_ & new_n694_;
  assign new_n699_ = new_n697_ & new_n698_;
  assign new_n700_ = new_n691_ & new_n694_;
  assign new_n701_ = ~new_n697_ & new_n700_;
  assign new_n702_ = ~new_n699_ & ~new_n701_;
  assign new_n703_ = new_n691_ & ~new_n694_;
  assign new_n704_ = new_n697_ & new_n703_;
  assign new_n705_ = ~new_n691_ & ~new_n694_;
  assign new_n706_ = ~new_n697_ & new_n705_;
  assign new_n707_ = ~new_n704_ & ~new_n706_;
  assign new_n708_ = new_n702_ & new_n707_;
  assign new_n709_ = ~new_n688_ & new_n708_;
  assign new_n710_ = new_n688_ & ~new_n708_;
  assign G1004 = new_n709_ | new_n710_;
  assign new_n712_ = G446 & ~new_n541_;
  assign new_n713_ = G457 & ~new_n535_;
  assign new_n714_ = ~new_n544_ & new_n713_;
  assign new_n715_ = G468 & ~new_n529_;
  assign new_n716_ = ~new_n538_ & ~new_n544_;
  assign new_n717_ = new_n715_ & new_n716_;
  assign new_n718_ = G422 & ~new_n523_;
  assign new_n719_ = ~new_n532_ & ~new_n544_;
  assign new_n720_ = new_n718_ & new_n719_;
  assign new_n721_ = ~new_n538_ & new_n720_;
  assign new_n722_ = ~new_n712_ & ~new_n714_;
  assign new_n723_ = ~new_n717_ & ~new_n721_;
  assign new_n724_ = new_n722_ & new_n723_;
  assign new_n725_ = G435 & ~new_n574_;
  assign new_n726_ = G389 & ~new_n568_;
  assign new_n727_ = ~new_n577_ & new_n726_;
  assign new_n728_ = G400 & ~new_n562_;
  assign new_n729_ = ~new_n571_ & ~new_n577_;
  assign new_n730_ = new_n728_ & new_n729_;
  assign new_n731_ = G411 & ~new_n556_;
  assign new_n732_ = ~new_n565_ & ~new_n577_;
  assign new_n733_ = new_n731_ & new_n732_;
  assign new_n734_ = ~new_n571_ & new_n733_;
  assign new_n735_ = G374 & ~new_n550_;
  assign new_n736_ = ~new_n559_ & ~new_n565_;
  assign new_n737_ = ~new_n577_ & new_n736_;
  assign new_n738_ = new_n735_ & new_n737_;
  assign new_n739_ = ~new_n571_ & new_n738_;
  assign new_n740_ = ~new_n725_ & ~new_n727_;
  assign new_n741_ = ~new_n730_ & new_n740_;
  assign new_n742_ = ~new_n734_ & ~new_n739_;
  assign new_n743_ = new_n741_ & new_n742_;
  assign new_n744_ = new_n547_ & ~new_n743_;
  assign G591 = ~new_n724_ | new_n744_;
  assign new_n746_ = ~new_n585_ & new_n600_;
  assign new_n747_ = G479 & ~new_n594_;
  assign new_n748_ = new_n585_ & new_n600_;
  assign new_n749_ = new_n747_ & new_n748_;
  assign new_n750_ = G490 & ~new_n588_;
  assign new_n751_ = ~new_n597_ & new_n600_;
  assign new_n752_ = new_n750_ & new_n751_;
  assign new_n753_ = new_n585_ & new_n752_;
  assign new_n754_ = new_n600_ & ~new_n746_;
  assign new_n755_ = ~new_n749_ & ~new_n753_;
  assign new_n756_ = new_n754_ & new_n755_;
  assign new_n757_ = G503 & ~new_n620_;
  assign new_n758_ = G514 & ~new_n605_;
  assign new_n759_ = ~new_n623_ & new_n758_;
  assign new_n760_ = G523 & ~new_n614_;
  assign new_n761_ = ~new_n608_ & ~new_n623_;
  assign new_n762_ = new_n760_ & new_n761_;
  assign new_n763_ = G534 & ~new_n626_;
  assign new_n764_ = ~new_n617_ & ~new_n623_;
  assign new_n765_ = new_n763_ & new_n764_;
  assign new_n766_ = ~new_n608_ & new_n765_;
  assign new_n767_ = ~new_n617_ & ~new_n629_;
  assign new_n768_ = ~new_n623_ & new_n767_;
  assign new_n769_ = ~new_n611_ & new_n768_;
  assign new_n770_ = ~new_n608_ & new_n769_;
  assign new_n771_ = ~new_n757_ & ~new_n759_;
  assign new_n772_ = ~new_n762_ & new_n771_;
  assign new_n773_ = ~new_n766_ & ~new_n770_;
  assign new_n774_ = new_n772_ & new_n773_;
  assign new_n775_ = new_n603_ & ~new_n774_;
  assign G618 = ~new_n756_ | new_n775_;
  assign new_n777_ = new_n645_ & ~new_n743_;
  assign G621 = ~new_n724_ | new_n777_;
  assign new_n779_ = new_n637_ & ~new_n774_;
  assign G629 = ~new_n756_ | new_n779_;
  assign new_n781_ = ~G4091 & new_n420_;
  assign new_n782_ = ~G4092 & new_n781_;
  assign new_n783_ = ~G54 & new_n611_;
  assign new_n784_ = G54 & ~new_n611_;
  assign new_n785_ = ~new_n783_ & ~new_n784_;
  assign new_n786_ = G4091 & ~new_n785_;
  assign new_n787_ = ~G4092 & new_n786_;
  assign new_n788_ = G131 & ~G4091;
  assign new_n789_ = G4092 & new_n788_;
  assign new_n790_ = ~new_n782_ & ~new_n787_;
  assign G822 = ~new_n789_ & new_n790_;
  assign new_n792_ = ~G4091 & new_n391_;
  assign new_n793_ = ~G4092 & new_n792_;
  assign new_n794_ = G54 & new_n611_;
  assign new_n795_ = new_n611_ & ~new_n794_;
  assign new_n796_ = ~new_n629_ & new_n795_;
  assign new_n797_ = new_n629_ & ~new_n795_;
  assign new_n798_ = ~new_n796_ & ~new_n797_;
  assign new_n799_ = G4091 & ~new_n798_;
  assign new_n800_ = ~G4092 & new_n799_;
  assign new_n801_ = G129 & ~G4091;
  assign new_n802_ = G4092 & new_n801_;
  assign new_n803_ = ~new_n793_ & ~new_n800_;
  assign G838 = ~new_n802_ & new_n803_;
  assign new_n805_ = ~G4091 & new_n475_;
  assign new_n806_ = ~G4092 & new_n805_;
  assign new_n807_ = ~G4 & ~new_n553_;
  assign new_n808_ = G4 & new_n553_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = G4091 & ~new_n809_;
  assign new_n811_ = ~G4092 & new_n810_;
  assign new_n812_ = G117 & ~G4091;
  assign new_n813_ = G4092 & new_n812_;
  assign new_n814_ = ~new_n806_ & ~new_n811_;
  assign G861 = ~new_n813_ & new_n814_;
  assign new_n816_ = new_n585_ & new_n747_;
  assign new_n817_ = ~new_n597_ & new_n750_;
  assign new_n818_ = new_n585_ & new_n817_;
  assign new_n819_ = new_n585_ & ~new_n816_;
  assign new_n820_ = ~new_n818_ & new_n819_;
  assign new_n821_ = new_n600_ & ~new_n820_;
  assign new_n822_ = ~new_n600_ & new_n820_;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = G54 & new_n633_;
  assign new_n825_ = new_n774_ & ~new_n824_;
  assign new_n826_ = new_n823_ & new_n825_;
  assign new_n827_ = ~new_n636_ & ~new_n818_;
  assign new_n828_ = new_n819_ & new_n827_;
  assign new_n829_ = new_n600_ & new_n828_;
  assign new_n830_ = ~new_n600_ & ~new_n828_;
  assign new_n831_ = ~new_n829_ & ~new_n830_;
  assign new_n832_ = ~new_n825_ & ~new_n831_;
  assign G623 = ~new_n826_ & ~new_n832_;
  assign new_n834_ = ~G4088 & ~G822;
  assign new_n835_ = ~G4087 & new_n834_;
  assign new_n836_ = G4088 & ~G861;
  assign new_n837_ = ~G4087 & new_n836_;
  assign new_n838_ = G11 & ~G4088;
  assign new_n839_ = G4087 & new_n838_;
  assign new_n840_ = G61 & G4088;
  assign new_n841_ = G4087 & new_n840_;
  assign new_n842_ = ~new_n835_ & ~new_n837_;
  assign new_n843_ = ~new_n839_ & ~new_n841_;
  assign G722 = ~new_n842_ | ~new_n843_;
  assign new_n845_ = ~G4091 & new_n414_;
  assign new_n846_ = ~G4092 & new_n845_;
  assign new_n847_ = ~new_n608_ & new_n760_;
  assign new_n848_ = ~new_n617_ & new_n763_;
  assign new_n849_ = ~new_n608_ & new_n848_;
  assign new_n850_ = ~new_n611_ & new_n767_;
  assign new_n851_ = ~new_n608_ & new_n850_;
  assign new_n852_ = ~new_n617_ & new_n794_;
  assign new_n853_ = ~new_n629_ & new_n852_;
  assign new_n854_ = ~new_n608_ & new_n853_;
  assign new_n855_ = ~new_n758_ & ~new_n847_;
  assign new_n856_ = ~new_n849_ & new_n855_;
  assign new_n857_ = ~new_n851_ & ~new_n854_;
  assign new_n858_ = new_n856_ & new_n857_;
  assign new_n859_ = ~new_n623_ & new_n858_;
  assign new_n860_ = new_n623_ & ~new_n858_;
  assign new_n861_ = ~new_n859_ & ~new_n860_;
  assign new_n862_ = G4091 & ~new_n861_;
  assign new_n863_ = ~G4092 & new_n862_;
  assign new_n864_ = G52 & ~G4091;
  assign new_n865_ = G4092 & new_n864_;
  assign new_n866_ = ~new_n846_ & ~new_n863_;
  assign G832 = ~new_n865_ & new_n866_;
  assign new_n868_ = ~G4091 & new_n404_;
  assign new_n869_ = ~G4092 & new_n868_;
  assign new_n870_ = ~new_n760_ & ~new_n848_;
  assign new_n871_ = ~new_n850_ & ~new_n853_;
  assign new_n872_ = new_n870_ & new_n871_;
  assign new_n873_ = ~new_n608_ & new_n872_;
  assign new_n874_ = new_n608_ & ~new_n872_;
  assign new_n875_ = ~new_n873_ & ~new_n874_;
  assign new_n876_ = G4091 & ~new_n875_;
  assign new_n877_ = ~G4092 & new_n876_;
  assign new_n878_ = G130 & ~G4091;
  assign new_n879_ = G4092 & new_n878_;
  assign new_n880_ = ~new_n869_ & ~new_n877_;
  assign G834 = ~new_n879_ & new_n880_;
  assign new_n882_ = ~G4091 & new_n401_;
  assign new_n883_ = ~G4092 & new_n882_;
  assign new_n884_ = ~new_n611_ & ~new_n629_;
  assign new_n885_ = ~new_n629_ & new_n794_;
  assign new_n886_ = ~new_n763_ & ~new_n884_;
  assign new_n887_ = ~new_n885_ & new_n886_;
  assign new_n888_ = ~new_n617_ & new_n887_;
  assign new_n889_ = new_n617_ & ~new_n887_;
  assign new_n890_ = ~new_n888_ & ~new_n889_;
  assign new_n891_ = G4091 & ~new_n890_;
  assign new_n892_ = ~G4092 & new_n891_;
  assign new_n893_ = G119 & ~G4091;
  assign new_n894_ = G4092 & new_n893_;
  assign new_n895_ = ~new_n883_ & ~new_n892_;
  assign G836 = ~new_n894_ & new_n895_;
  assign new_n897_ = ~G4089 & ~G822;
  assign new_n898_ = ~G4090 & new_n897_;
  assign new_n899_ = G4089 & ~G861;
  assign new_n900_ = ~G4090 & new_n899_;
  assign new_n901_ = G11 & ~G4089;
  assign new_n902_ = G4090 & new_n901_;
  assign new_n903_ = G61 & G4089;
  assign new_n904_ = G4090 & new_n903_;
  assign new_n905_ = ~new_n898_ & ~new_n900_;
  assign new_n906_ = ~new_n902_ & ~new_n904_;
  assign G859 = ~new_n905_ | ~new_n906_;
  assign new_n908_ = ~G4091 & new_n432_;
  assign new_n909_ = ~G4092 & new_n908_;
  assign new_n910_ = ~new_n571_ & new_n728_;
  assign new_n911_ = ~new_n565_ & new_n731_;
  assign new_n912_ = ~new_n571_ & new_n911_;
  assign new_n913_ = new_n735_ & new_n736_;
  assign new_n914_ = ~new_n571_ & new_n913_;
  assign new_n915_ = G4 & ~new_n553_;
  assign new_n916_ = ~new_n565_ & new_n915_;
  assign new_n917_ = ~new_n559_ & new_n916_;
  assign new_n918_ = ~new_n571_ & new_n917_;
  assign new_n919_ = ~new_n726_ & ~new_n910_;
  assign new_n920_ = ~new_n912_ & new_n919_;
  assign new_n921_ = ~new_n914_ & ~new_n918_;
  assign new_n922_ = new_n920_ & new_n921_;
  assign new_n923_ = ~new_n577_ & new_n922_;
  assign new_n924_ = new_n577_ & ~new_n922_;
  assign new_n925_ = ~new_n923_ & ~new_n924_;
  assign new_n926_ = G4091 & ~new_n925_;
  assign new_n927_ = ~G4092 & new_n926_;
  assign new_n928_ = G122 & ~G4091;
  assign new_n929_ = G4092 & new_n928_;
  assign new_n930_ = ~new_n909_ & ~new_n927_;
  assign G871 = ~new_n929_ & new_n930_;
  assign new_n932_ = ~G4091 & new_n505_;
  assign new_n933_ = ~G4092 & new_n932_;
  assign new_n934_ = ~new_n728_ & ~new_n911_;
  assign new_n935_ = ~new_n913_ & ~new_n917_;
  assign new_n936_ = new_n934_ & new_n935_;
  assign new_n937_ = ~new_n571_ & new_n936_;
  assign new_n938_ = new_n571_ & ~new_n936_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = G4091 & ~new_n939_;
  assign new_n941_ = ~G4092 & new_n940_;
  assign new_n942_ = G128 & ~G4091;
  assign new_n943_ = G4092 & new_n942_;
  assign new_n944_ = ~new_n933_ & ~new_n941_;
  assign G873 = ~new_n943_ & new_n944_;
  assign new_n946_ = ~G4091 & new_n495_;
  assign new_n947_ = ~G4092 & new_n946_;
  assign new_n948_ = ~new_n559_ & new_n735_;
  assign new_n949_ = ~new_n559_ & new_n915_;
  assign new_n950_ = ~new_n731_ & ~new_n948_;
  assign new_n951_ = ~new_n949_ & new_n950_;
  assign new_n952_ = ~new_n565_ & new_n951_;
  assign new_n953_ = new_n565_ & ~new_n951_;
  assign new_n954_ = ~new_n952_ & ~new_n953_;
  assign new_n955_ = G4091 & ~new_n954_;
  assign new_n956_ = ~G4092 & new_n955_;
  assign new_n957_ = G127 & ~G4091;
  assign new_n958_ = G4092 & new_n957_;
  assign new_n959_ = ~new_n947_ & ~new_n956_;
  assign G875 = ~new_n958_ & new_n959_;
  assign new_n961_ = ~G4091 & new_n485_;
  assign new_n962_ = ~G4092 & new_n961_;
  assign new_n963_ = ~new_n735_ & ~new_n915_;
  assign new_n964_ = ~new_n559_ & new_n963_;
  assign new_n965_ = new_n559_ & ~new_n963_;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = G4091 & ~new_n966_;
  assign new_n968_ = ~G4092 & new_n967_;
  assign new_n969_ = G126 & ~G4091;
  assign new_n970_ = G4092 & new_n969_;
  assign new_n971_ = ~new_n962_ & ~new_n968_;
  assign G877 = ~new_n970_ & new_n971_;
  assign new_n973_ = ~new_n588_ & new_n594_;
  assign new_n974_ = new_n588_ & ~new_n594_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign new_n976_ = new_n585_ & ~new_n600_;
  assign new_n977_ = ~new_n746_ & ~new_n976_;
  assign new_n978_ = ~new_n975_ & new_n977_;
  assign new_n979_ = new_n975_ & ~new_n977_;
  assign new_n980_ = ~new_n978_ & ~new_n979_;
  assign new_n981_ = ~new_n614_ & new_n626_;
  assign new_n982_ = new_n614_ & ~new_n626_;
  assign new_n983_ = ~new_n981_ & ~new_n982_;
  assign new_n984_ = ~G332 & G369;
  assign new_n985_ = G332 & G372;
  assign new_n986_ = ~new_n984_ & ~new_n985_;
  assign new_n987_ = ~new_n611_ & new_n986_;
  assign new_n988_ = new_n611_ & ~new_n986_;
  assign new_n989_ = ~new_n987_ & ~new_n988_;
  assign new_n990_ = ~new_n605_ & new_n620_;
  assign new_n991_ = new_n605_ & ~new_n620_;
  assign new_n992_ = ~new_n990_ & ~new_n991_;
  assign new_n993_ = ~new_n983_ & new_n989_;
  assign new_n994_ = new_n992_ & new_n993_;
  assign new_n995_ = new_n983_ & new_n989_;
  assign new_n996_ = ~new_n992_ & new_n995_;
  assign new_n997_ = ~new_n994_ & ~new_n996_;
  assign new_n998_ = new_n983_ & ~new_n989_;
  assign new_n999_ = new_n992_ & new_n998_;
  assign new_n1000_ = ~new_n983_ & ~new_n989_;
  assign new_n1001_ = ~new_n992_ & new_n1000_;
  assign new_n1002_ = ~new_n999_ & ~new_n1001_;
  assign new_n1003_ = new_n997_ & new_n1002_;
  assign new_n1004_ = ~new_n980_ & new_n1003_;
  assign new_n1005_ = new_n980_ & ~new_n1003_;
  assign G998 = new_n1004_ | new_n1005_;
  assign new_n1007_ = ~new_n550_ & new_n556_;
  assign new_n1008_ = new_n550_ & ~new_n556_;
  assign new_n1009_ = ~new_n1007_ & ~new_n1008_;
  assign new_n1010_ = ~new_n562_ & new_n568_;
  assign new_n1011_ = new_n562_ & ~new_n568_;
  assign new_n1012_ = ~new_n1010_ & ~new_n1011_;
  assign new_n1013_ = ~new_n1009_ & new_n1012_;
  assign new_n1014_ = new_n1009_ & ~new_n1012_;
  assign new_n1015_ = ~new_n1013_ & ~new_n1014_;
  assign new_n1016_ = new_n523_ & ~new_n574_;
  assign new_n1017_ = ~new_n523_ & new_n574_;
  assign new_n1018_ = ~new_n1016_ & ~new_n1017_;
  assign new_n1019_ = ~new_n529_ & new_n535_;
  assign new_n1020_ = new_n529_ & ~new_n535_;
  assign new_n1021_ = ~new_n1019_ & ~new_n1020_;
  assign new_n1022_ = G289 & ~G335;
  assign new_n1023_ = G292 & G335;
  assign new_n1024_ = ~new_n1022_ & ~new_n1023_;
  assign new_n1025_ = ~new_n541_ & new_n1024_;
  assign new_n1026_ = new_n541_ & ~new_n1024_;
  assign new_n1027_ = ~new_n1025_ & ~new_n1026_;
  assign new_n1028_ = ~new_n1018_ & new_n1021_;
  assign new_n1029_ = new_n1027_ & new_n1028_;
  assign new_n1030_ = new_n1018_ & new_n1021_;
  assign new_n1031_ = ~new_n1027_ & new_n1030_;
  assign new_n1032_ = ~new_n1029_ & ~new_n1031_;
  assign new_n1033_ = new_n1018_ & ~new_n1021_;
  assign new_n1034_ = new_n1027_ & new_n1033_;
  assign new_n1035_ = ~new_n1018_ & ~new_n1021_;
  assign new_n1036_ = ~new_n1027_ & new_n1035_;
  assign new_n1037_ = ~new_n1034_ & ~new_n1036_;
  assign new_n1038_ = new_n1032_ & new_n1037_;
  assign new_n1039_ = ~new_n1015_ & new_n1038_;
  assign new_n1040_ = new_n1015_ & ~new_n1038_;
  assign G1000 = new_n1039_ | new_n1040_;
  assign new_n1042_ = G4 & new_n649_;
  assign new_n1043_ = new_n743_ & ~new_n1042_;
  assign new_n1044_ = ~new_n526_ & new_n1043_;
  assign new_n1045_ = new_n526_ & ~new_n1043_;
  assign new_n1046_ = ~new_n1044_ & ~new_n1045_;
  assign new_n1047_ = ~new_n532_ & ~new_n718_;
  assign new_n1048_ = new_n532_ & new_n718_;
  assign new_n1049_ = ~new_n1047_ & ~new_n1048_;
  assign new_n1050_ = new_n1043_ & ~new_n1049_;
  assign new_n1051_ = ~G422 & new_n523_;
  assign new_n1052_ = ~new_n532_ & ~new_n1051_;
  assign new_n1053_ = new_n532_ & new_n1051_;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = ~new_n1043_ & new_n1054_;
  assign new_n1056_ = ~new_n1050_ & ~new_n1055_;
  assign new_n1057_ = ~new_n532_ & new_n718_;
  assign new_n1058_ = ~new_n715_ & ~new_n1057_;
  assign new_n1059_ = ~new_n538_ & ~new_n1058_;
  assign new_n1060_ = new_n538_ & new_n1058_;
  assign new_n1061_ = ~new_n1059_ & ~new_n1060_;
  assign new_n1062_ = new_n1043_ & new_n1061_;
  assign new_n1063_ = ~new_n545_ & new_n1058_;
  assign new_n1064_ = ~new_n538_ & new_n1063_;
  assign new_n1065_ = new_n538_ & ~new_n1063_;
  assign new_n1066_ = ~new_n1064_ & ~new_n1065_;
  assign new_n1067_ = ~new_n1043_ & ~new_n1066_;
  assign new_n1068_ = ~new_n1062_ & ~new_n1067_;
  assign new_n1069_ = ~new_n538_ & new_n715_;
  assign new_n1070_ = ~new_n538_ & new_n1057_;
  assign new_n1071_ = ~new_n713_ & ~new_n1069_;
  assign new_n1072_ = ~new_n1070_ & new_n1071_;
  assign new_n1073_ = ~new_n544_ & ~new_n1072_;
  assign new_n1074_ = new_n544_ & new_n1072_;
  assign new_n1075_ = ~new_n1073_ & ~new_n1074_;
  assign new_n1076_ = new_n1043_ & new_n1075_;
  assign new_n1077_ = ~new_n546_ & ~new_n1070_;
  assign new_n1078_ = new_n1071_ & new_n1077_;
  assign new_n1079_ = ~new_n544_ & new_n1078_;
  assign new_n1080_ = new_n544_ & ~new_n1078_;
  assign new_n1081_ = ~new_n1079_ & ~new_n1080_;
  assign new_n1082_ = ~new_n1043_ & ~new_n1081_;
  assign new_n1083_ = ~new_n1076_ & ~new_n1082_;
  assign new_n1084_ = new_n809_ & new_n966_;
  assign new_n1085_ = new_n954_ & new_n1084_;
  assign new_n1086_ = new_n939_ & new_n1085_;
  assign new_n1087_ = new_n925_ & new_n1086_;
  assign new_n1088_ = new_n1046_ & new_n1087_;
  assign new_n1089_ = new_n1056_ & new_n1088_;
  assign new_n1090_ = new_n1068_ & new_n1089_;
  assign G575 = new_n1083_ & new_n1090_;
  assign new_n1092_ = ~new_n591_ & new_n825_;
  assign new_n1093_ = new_n591_ & ~new_n825_;
  assign new_n1094_ = ~new_n1092_ & ~new_n1093_;
  assign new_n1095_ = ~new_n597_ & ~new_n750_;
  assign new_n1096_ = new_n597_ & new_n750_;
  assign new_n1097_ = ~new_n1095_ & ~new_n1096_;
  assign new_n1098_ = new_n825_ & ~new_n1097_;
  assign new_n1099_ = ~G490 & new_n588_;
  assign new_n1100_ = ~new_n597_ & ~new_n1099_;
  assign new_n1101_ = new_n597_ & new_n1099_;
  assign new_n1102_ = ~new_n1100_ & ~new_n1101_;
  assign new_n1103_ = ~new_n825_ & new_n1102_;
  assign new_n1104_ = ~new_n1098_ & ~new_n1103_;
  assign new_n1105_ = ~new_n747_ & ~new_n817_;
  assign new_n1106_ = new_n585_ & ~new_n1105_;
  assign new_n1107_ = ~new_n585_ & new_n1105_;
  assign new_n1108_ = ~new_n1106_ & ~new_n1107_;
  assign new_n1109_ = new_n825_ & new_n1108_;
  assign new_n1110_ = ~new_n635_ & new_n1105_;
  assign new_n1111_ = new_n585_ & new_n1110_;
  assign new_n1112_ = ~new_n585_ & ~new_n1110_;
  assign new_n1113_ = ~new_n1111_ & ~new_n1112_;
  assign new_n1114_ = ~new_n825_ & ~new_n1113_;
  assign new_n1115_ = ~new_n1109_ & ~new_n1114_;
  assign new_n1116_ = new_n785_ & new_n798_;
  assign new_n1117_ = new_n890_ & new_n1116_;
  assign new_n1118_ = new_n875_ & new_n1117_;
  assign new_n1119_ = new_n861_ & new_n1118_;
  assign new_n1120_ = new_n1094_ & new_n1119_;
  assign new_n1121_ = new_n1104_ & new_n1120_;
  assign new_n1122_ = new_n1115_ & new_n1121_;
  assign G585 = G623 & new_n1122_;
  assign new_n1124_ = ~G1689 & ~G822;
  assign new_n1125_ = ~G1690 & new_n1124_;
  assign new_n1126_ = G1689 & ~G861;
  assign new_n1127_ = ~G1690 & new_n1126_;
  assign new_n1128_ = G182 & ~G1689;
  assign new_n1129_ = G1690 & new_n1128_;
  assign new_n1130_ = G185 & G1689;
  assign new_n1131_ = G1690 & new_n1130_;
  assign new_n1132_ = ~new_n1125_ & ~new_n1127_;
  assign new_n1133_ = ~new_n1129_ & ~new_n1131_;
  assign new_n1134_ = new_n1132_ & new_n1133_;
  assign G661 = G137 & ~new_n1134_;
  assign new_n1136_ = ~G1691 & ~G822;
  assign new_n1137_ = ~G1694 & new_n1136_;
  assign new_n1138_ = G1691 & ~G861;
  assign new_n1139_ = ~G1694 & new_n1138_;
  assign new_n1140_ = G182 & ~G1691;
  assign new_n1141_ = G1694 & new_n1140_;
  assign new_n1142_ = G185 & G1691;
  assign new_n1143_ = G1694 & new_n1142_;
  assign new_n1144_ = ~new_n1137_ & ~new_n1139_;
  assign new_n1145_ = ~new_n1141_ & ~new_n1143_;
  assign new_n1146_ = new_n1144_ & new_n1145_;
  assign G693 = G137 & ~new_n1146_;
  assign new_n1148_ = ~G4088 & ~G832;
  assign new_n1149_ = ~G4087 & new_n1148_;
  assign new_n1150_ = G4088 & ~G871;
  assign new_n1151_ = ~G4087 & new_n1150_;
  assign new_n1152_ = G43 & ~G4088;
  assign new_n1153_ = G4087 & new_n1152_;
  assign new_n1154_ = G37 & G4088;
  assign new_n1155_ = G4087 & new_n1154_;
  assign new_n1156_ = ~new_n1149_ & ~new_n1151_;
  assign new_n1157_ = ~new_n1153_ & ~new_n1155_;
  assign G747 = ~new_n1156_ | ~new_n1157_;
  assign new_n1159_ = ~G4088 & ~G834;
  assign new_n1160_ = ~G4087 & new_n1159_;
  assign new_n1161_ = G4088 & ~G873;
  assign new_n1162_ = ~G4087 & new_n1161_;
  assign new_n1163_ = G76 & ~G4088;
  assign new_n1164_ = G4087 & new_n1163_;
  assign new_n1165_ = G20 & G4088;
  assign new_n1166_ = G4087 & new_n1165_;
  assign new_n1167_ = ~new_n1160_ & ~new_n1162_;
  assign new_n1168_ = ~new_n1164_ & ~new_n1166_;
  assign G752 = ~new_n1167_ | ~new_n1168_;
  assign new_n1170_ = ~G4088 & ~G836;
  assign new_n1171_ = ~G4087 & new_n1170_;
  assign new_n1172_ = G4088 & ~G875;
  assign new_n1173_ = ~G4087 & new_n1172_;
  assign new_n1174_ = G73 & ~G4088;
  assign new_n1175_ = G4087 & new_n1174_;
  assign new_n1176_ = G17 & G4088;
  assign new_n1177_ = G4087 & new_n1176_;
  assign new_n1178_ = ~new_n1171_ & ~new_n1173_;
  assign new_n1179_ = ~new_n1175_ & ~new_n1177_;
  assign G757 = ~new_n1178_ | ~new_n1179_;
  assign new_n1181_ = ~G4088 & ~G838;
  assign new_n1182_ = ~G4087 & new_n1181_;
  assign new_n1183_ = G4088 & ~G877;
  assign new_n1184_ = ~G4087 & new_n1183_;
  assign new_n1185_ = G67 & ~G4088;
  assign new_n1186_ = G4087 & new_n1185_;
  assign new_n1187_ = G70 & G4088;
  assign new_n1188_ = G4087 & new_n1187_;
  assign new_n1189_ = ~new_n1182_ & ~new_n1184_;
  assign new_n1190_ = ~new_n1186_ & ~new_n1188_;
  assign G762 = ~new_n1189_ | ~new_n1190_;
  assign new_n1192_ = ~G4089 & ~G832;
  assign new_n1193_ = ~G4090 & new_n1192_;
  assign new_n1194_ = G4089 & ~G871;
  assign new_n1195_ = ~G4090 & new_n1194_;
  assign new_n1196_ = G43 & ~G4089;
  assign new_n1197_ = G4090 & new_n1196_;
  assign new_n1198_ = G37 & G4089;
  assign new_n1199_ = G4090 & new_n1198_;
  assign new_n1200_ = ~new_n1193_ & ~new_n1195_;
  assign new_n1201_ = ~new_n1197_ & ~new_n1199_;
  assign G787 = ~new_n1200_ | ~new_n1201_;
  assign new_n1203_ = ~G4089 & ~G834;
  assign new_n1204_ = ~G4090 & new_n1203_;
  assign new_n1205_ = G4089 & ~G873;
  assign new_n1206_ = ~G4090 & new_n1205_;
  assign new_n1207_ = G76 & ~G4089;
  assign new_n1208_ = G4090 & new_n1207_;
  assign new_n1209_ = G20 & G4089;
  assign new_n1210_ = G4090 & new_n1209_;
  assign new_n1211_ = ~new_n1204_ & ~new_n1206_;
  assign new_n1212_ = ~new_n1208_ & ~new_n1210_;
  assign G792 = ~new_n1211_ | ~new_n1212_;
  assign new_n1214_ = ~G4089 & ~G836;
  assign new_n1215_ = ~G4090 & new_n1214_;
  assign new_n1216_ = G4089 & ~G875;
  assign new_n1217_ = ~G4090 & new_n1216_;
  assign new_n1218_ = G73 & ~G4089;
  assign new_n1219_ = G4090 & new_n1218_;
  assign new_n1220_ = G17 & G4089;
  assign new_n1221_ = G4090 & new_n1220_;
  assign new_n1222_ = ~new_n1215_ & ~new_n1217_;
  assign new_n1223_ = ~new_n1219_ & ~new_n1221_;
  assign G797 = ~new_n1222_ | ~new_n1223_;
  assign new_n1225_ = ~G4089 & ~G838;
  assign new_n1226_ = ~G4090 & new_n1225_;
  assign new_n1227_ = G4089 & ~G877;
  assign new_n1228_ = ~G4090 & new_n1227_;
  assign new_n1229_ = G67 & ~G4089;
  assign new_n1230_ = G4090 & new_n1229_;
  assign new_n1231_ = G70 & G4089;
  assign new_n1232_ = G4090 & new_n1231_;
  assign new_n1233_ = ~new_n1226_ & ~new_n1228_;
  assign new_n1234_ = ~new_n1230_ & ~new_n1232_;
  assign G802 = ~new_n1233_ | ~new_n1234_;
  assign new_n1236_ = ~G1689 & ~G832;
  assign new_n1237_ = ~G1690 & new_n1236_;
  assign new_n1238_ = G1689 & ~G871;
  assign new_n1239_ = ~G1690 & new_n1238_;
  assign new_n1240_ = G200 & ~G1689;
  assign new_n1241_ = G1690 & new_n1240_;
  assign new_n1242_ = G170 & G1689;
  assign new_n1243_ = G1690 & new_n1242_;
  assign new_n1244_ = ~new_n1237_ & ~new_n1239_;
  assign new_n1245_ = ~new_n1241_ & ~new_n1243_;
  assign new_n1246_ = new_n1244_ & new_n1245_;
  assign G642 = G137 & ~new_n1246_;
  assign new_n1248_ = ~G1689 & ~G838;
  assign new_n1249_ = ~G1690 & new_n1248_;
  assign new_n1250_ = G1689 & ~G877;
  assign new_n1251_ = ~G1690 & new_n1250_;
  assign new_n1252_ = G188 & ~G1689;
  assign new_n1253_ = G1690 & new_n1252_;
  assign new_n1254_ = G158 & G1689;
  assign new_n1255_ = G1690 & new_n1254_;
  assign new_n1256_ = ~new_n1249_ & ~new_n1251_;
  assign new_n1257_ = ~new_n1253_ & ~new_n1255_;
  assign new_n1258_ = new_n1256_ & new_n1257_;
  assign G664 = G137 & ~new_n1258_;
  assign new_n1260_ = ~G1689 & ~G836;
  assign new_n1261_ = ~G1690 & new_n1260_;
  assign new_n1262_ = G1689 & ~G875;
  assign new_n1263_ = ~G1690 & new_n1262_;
  assign new_n1264_ = G155 & ~G1689;
  assign new_n1265_ = G1690 & new_n1264_;
  assign new_n1266_ = G152 & G1689;
  assign new_n1267_ = G1690 & new_n1266_;
  assign new_n1268_ = ~new_n1261_ & ~new_n1263_;
  assign new_n1269_ = ~new_n1265_ & ~new_n1267_;
  assign new_n1270_ = new_n1268_ & new_n1269_;
  assign G667 = G137 & ~new_n1270_;
  assign new_n1272_ = ~G1689 & ~G834;
  assign new_n1273_ = ~G1690 & new_n1272_;
  assign new_n1274_ = G1689 & ~G873;
  assign new_n1275_ = ~G1690 & new_n1274_;
  assign new_n1276_ = G149 & ~G1689;
  assign new_n1277_ = G1690 & new_n1276_;
  assign new_n1278_ = G146 & G1689;
  assign new_n1279_ = G1690 & new_n1278_;
  assign new_n1280_ = ~new_n1273_ & ~new_n1275_;
  assign new_n1281_ = ~new_n1277_ & ~new_n1279_;
  assign new_n1282_ = new_n1280_ & new_n1281_;
  assign G670 = G137 & ~new_n1282_;
  assign new_n1284_ = ~G1691 & ~G832;
  assign new_n1285_ = ~G1694 & new_n1284_;
  assign new_n1286_ = G1691 & ~G871;
  assign new_n1287_ = ~G1694 & new_n1286_;
  assign new_n1288_ = G200 & ~G1691;
  assign new_n1289_ = G1694 & new_n1288_;
  assign new_n1290_ = G170 & G1691;
  assign new_n1291_ = G1694 & new_n1290_;
  assign new_n1292_ = ~new_n1285_ & ~new_n1287_;
  assign new_n1293_ = ~new_n1289_ & ~new_n1291_;
  assign new_n1294_ = new_n1292_ & new_n1293_;
  assign G676 = G137 & ~new_n1294_;
  assign new_n1296_ = ~G1691 & ~G838;
  assign new_n1297_ = ~G1694 & new_n1296_;
  assign new_n1298_ = G1691 & ~G877;
  assign new_n1299_ = ~G1694 & new_n1298_;
  assign new_n1300_ = G188 & ~G1691;
  assign new_n1301_ = G1694 & new_n1300_;
  assign new_n1302_ = G158 & G1691;
  assign new_n1303_ = G1694 & new_n1302_;
  assign new_n1304_ = ~new_n1297_ & ~new_n1299_;
  assign new_n1305_ = ~new_n1301_ & ~new_n1303_;
  assign new_n1306_ = new_n1304_ & new_n1305_;
  assign G696 = G137 & ~new_n1306_;
  assign new_n1308_ = ~G1691 & ~G836;
  assign new_n1309_ = ~G1694 & new_n1308_;
  assign new_n1310_ = G1691 & ~G875;
  assign new_n1311_ = ~G1694 & new_n1310_;
  assign new_n1312_ = G155 & ~G1691;
  assign new_n1313_ = G1694 & new_n1312_;
  assign new_n1314_ = G152 & G1691;
  assign new_n1315_ = G1694 & new_n1314_;
  assign new_n1316_ = ~new_n1309_ & ~new_n1311_;
  assign new_n1317_ = ~new_n1313_ & ~new_n1315_;
  assign new_n1318_ = new_n1316_ & new_n1317_;
  assign G699 = G137 & ~new_n1318_;
  assign new_n1320_ = ~G1691 & ~G834;
  assign new_n1321_ = ~G1694 & new_n1320_;
  assign new_n1322_ = G1691 & ~G873;
  assign new_n1323_ = ~G1694 & new_n1322_;
  assign new_n1324_ = G149 & ~G1691;
  assign new_n1325_ = G1694 & new_n1324_;
  assign new_n1326_ = G146 & G1691;
  assign new_n1327_ = G1694 & new_n1326_;
  assign new_n1328_ = ~new_n1321_ & ~new_n1323_;
  assign new_n1329_ = ~new_n1325_ & ~new_n1327_;
  assign new_n1330_ = new_n1328_ & new_n1329_;
  assign G702 = G137 & ~new_n1330_;
  assign new_n1332_ = G135 & G4115;
  assign new_n1333_ = ~G3724 & ~new_n378_;
  assign new_n1334_ = ~G3717 & new_n1333_;
  assign new_n1335_ = G132 & new_n600_;
  assign new_n1336_ = new_n600_ & ~new_n1335_;
  assign new_n1337_ = G132 & ~new_n1335_;
  assign new_n1338_ = ~new_n1336_ & ~new_n1337_;
  assign new_n1339_ = G3724 & ~new_n1338_;
  assign new_n1340_ = ~G3717 & new_n1339_;
  assign new_n1341_ = G123 & ~G3724;
  assign new_n1342_ = G3717 & new_n1341_;
  assign new_n1343_ = G3724 & ~G623;
  assign new_n1344_ = G3717 & new_n1343_;
  assign new_n1345_ = ~new_n1334_ & ~new_n1340_;
  assign new_n1346_ = ~new_n1342_ & ~new_n1344_;
  assign new_n1347_ = new_n1345_ & new_n1346_;
  assign G818 = ~new_n1332_ & ~new_n1347_;
  assign new_n1349_ = ~G623 & ~new_n1338_;
  assign new_n1350_ = ~new_n1338_ & ~new_n1349_;
  assign new_n1351_ = ~G623 & ~new_n1349_;
  assign G813 = new_n1350_ | new_n1351_;
  assign new_n1353_ = ~G4091 & ~new_n378_;
  assign new_n1354_ = ~G4092 & new_n1353_;
  assign new_n1355_ = G4091 & ~G623;
  assign new_n1356_ = ~G4092 & new_n1355_;
  assign new_n1357_ = G123 & ~G4091;
  assign new_n1358_ = G4092 & new_n1357_;
  assign new_n1359_ = ~new_n1354_ & ~new_n1356_;
  assign G824 = ~new_n1358_ & new_n1359_;
  assign new_n1361_ = ~G4091 & new_n375_;
  assign new_n1362_ = ~G4092 & new_n1361_;
  assign new_n1363_ = G4091 & ~new_n1115_;
  assign new_n1364_ = ~G4092 & new_n1363_;
  assign new_n1365_ = G121 & ~G4091;
  assign new_n1366_ = G4092 & new_n1365_;
  assign new_n1367_ = ~new_n1362_ & ~new_n1364_;
  assign G826 = ~new_n1366_ & new_n1367_;
  assign new_n1369_ = ~G4091 & new_n372_;
  assign new_n1370_ = ~G4092 & new_n1369_;
  assign new_n1371_ = G4091 & ~new_n1104_;
  assign new_n1372_ = ~G4092 & new_n1371_;
  assign new_n1373_ = G116 & ~G4091;
  assign new_n1374_ = G4092 & new_n1373_;
  assign new_n1375_ = ~new_n1370_ & ~new_n1372_;
  assign G828 = ~new_n1374_ & new_n1375_;
  assign new_n1377_ = ~G4091 & new_n362_;
  assign new_n1378_ = ~G4092 & new_n1377_;
  assign new_n1379_ = G4091 & ~new_n1094_;
  assign new_n1380_ = ~G4092 & new_n1379_;
  assign new_n1381_ = G112 & ~G4091;
  assign new_n1382_ = G4092 & new_n1381_;
  assign new_n1383_ = ~new_n1378_ & ~new_n1380_;
  assign G830 = ~new_n1382_ & new_n1383_;
  assign new_n1385_ = G386 & G559;
  assign new_n1386_ = G556 & new_n1385_;
  assign new_n1387_ = G552 & new_n1386_;
  assign new_n1388_ = G562 & ~G998;
  assign new_n1389_ = ~G1000 & new_n1388_;
  assign new_n1390_ = ~G1002 & new_n1389_;
  assign new_n1391_ = ~G1004 & new_n1390_;
  assign new_n1392_ = new_n1387_ & new_n1391_;
  assign G854 = G245 & new_n1392_;
  assign new_n1394_ = ~G4091 & new_n518_;
  assign new_n1395_ = ~G4092 & new_n1394_;
  assign new_n1396_ = G4091 & ~new_n1083_;
  assign new_n1397_ = ~G4092 & new_n1396_;
  assign new_n1398_ = G115 & ~G4091;
  assign new_n1399_ = G4092 & new_n1398_;
  assign new_n1400_ = ~new_n1395_ & ~new_n1397_;
  assign G863 = ~new_n1399_ & new_n1400_;
  assign new_n1402_ = ~G4091 & new_n462_;
  assign new_n1403_ = ~G4092 & new_n1402_;
  assign new_n1404_ = G4091 & ~new_n1068_;
  assign new_n1405_ = ~G4092 & new_n1404_;
  assign new_n1406_ = G114 & ~G4091;
  assign new_n1407_ = G4092 & new_n1406_;
  assign new_n1408_ = ~new_n1403_ & ~new_n1405_;
  assign G865 = ~new_n1407_ & new_n1408_;
  assign new_n1410_ = ~G4091 & new_n452_;
  assign new_n1411_ = ~G4092 & new_n1410_;
  assign new_n1412_ = G4091 & ~new_n1056_;
  assign new_n1413_ = ~G4092 & new_n1412_;
  assign new_n1414_ = G53 & ~G4091;
  assign new_n1415_ = G4092 & new_n1414_;
  assign new_n1416_ = ~new_n1411_ & ~new_n1413_;
  assign G867 = ~new_n1415_ & new_n1416_;
  assign new_n1418_ = ~G4091 & new_n442_;
  assign new_n1419_ = ~G4092 & new_n1418_;
  assign new_n1420_ = G4091 & ~new_n1046_;
  assign new_n1421_ = ~G4092 & new_n1420_;
  assign new_n1422_ = G113 & ~G4091;
  assign new_n1423_ = G4092 & new_n1422_;
  assign new_n1424_ = ~new_n1419_ & ~new_n1421_;
  assign G869 = ~new_n1423_ & new_n1424_;
  assign new_n1426_ = ~G4089 & ~G824;
  assign new_n1427_ = ~G4090 & new_n1426_;
  assign new_n1428_ = G4089 & ~G863;
  assign new_n1429_ = ~G4090 & new_n1428_;
  assign new_n1430_ = G109 & ~G4089;
  assign new_n1431_ = G4090 & new_n1430_;
  assign new_n1432_ = G106 & G4089;
  assign new_n1433_ = G4090 & new_n1432_;
  assign new_n1434_ = ~new_n1427_ & ~new_n1429_;
  assign new_n1435_ = ~new_n1431_ & ~new_n1433_;
  assign G712 = ~new_n1434_ | ~new_n1435_;
  assign new_n1437_ = ~G4088 & ~G824;
  assign new_n1438_ = ~G4087 & new_n1437_;
  assign new_n1439_ = G4088 & ~G863;
  assign new_n1440_ = ~G4087 & new_n1439_;
  assign new_n1441_ = G109 & ~G4088;
  assign new_n1442_ = G4087 & new_n1441_;
  assign new_n1443_ = G106 & G4088;
  assign new_n1444_ = G4087 & new_n1443_;
  assign new_n1445_ = ~new_n1438_ & ~new_n1440_;
  assign new_n1446_ = ~new_n1442_ & ~new_n1444_;
  assign G727 = ~new_n1445_ | ~new_n1446_;
  assign new_n1448_ = ~G4088 & ~G826;
  assign new_n1449_ = ~G4087 & new_n1448_;
  assign new_n1450_ = G4088 & ~G865;
  assign new_n1451_ = ~G4087 & new_n1450_;
  assign new_n1452_ = G46 & ~G4088;
  assign new_n1453_ = G4087 & new_n1452_;
  assign new_n1454_ = G49 & G4088;
  assign new_n1455_ = G4087 & new_n1454_;
  assign new_n1456_ = ~new_n1449_ & ~new_n1451_;
  assign new_n1457_ = ~new_n1453_ & ~new_n1455_;
  assign G732 = ~new_n1456_ | ~new_n1457_;
  assign new_n1459_ = ~G4088 & ~G828;
  assign new_n1460_ = ~G4087 & new_n1459_;
  assign new_n1461_ = G4088 & ~G867;
  assign new_n1462_ = ~G4087 & new_n1461_;
  assign new_n1463_ = G100 & ~G4088;
  assign new_n1464_ = G4087 & new_n1463_;
  assign new_n1465_ = G103 & G4088;
  assign new_n1466_ = G4087 & new_n1465_;
  assign new_n1467_ = ~new_n1460_ & ~new_n1462_;
  assign new_n1468_ = ~new_n1464_ & ~new_n1466_;
  assign G737 = ~new_n1467_ | ~new_n1468_;
  assign new_n1470_ = ~G4088 & ~G830;
  assign new_n1471_ = ~G4087 & new_n1470_;
  assign new_n1472_ = G4088 & ~G869;
  assign new_n1473_ = ~G4087 & new_n1472_;
  assign new_n1474_ = G91 & ~G4088;
  assign new_n1475_ = G4087 & new_n1474_;
  assign new_n1476_ = G40 & G4088;
  assign new_n1477_ = G4087 & new_n1476_;
  assign new_n1478_ = ~new_n1471_ & ~new_n1473_;
  assign new_n1479_ = ~new_n1475_ & ~new_n1477_;
  assign G742 = ~new_n1478_ | ~new_n1479_;
  assign new_n1481_ = ~G4089 & ~G826;
  assign new_n1482_ = ~G4090 & new_n1481_;
  assign new_n1483_ = G4089 & ~G865;
  assign new_n1484_ = ~G4090 & new_n1483_;
  assign new_n1485_ = G46 & ~G4089;
  assign new_n1486_ = G4090 & new_n1485_;
  assign new_n1487_ = G49 & G4089;
  assign new_n1488_ = G4090 & new_n1487_;
  assign new_n1489_ = ~new_n1482_ & ~new_n1484_;
  assign new_n1490_ = ~new_n1486_ & ~new_n1488_;
  assign G772 = ~new_n1489_ | ~new_n1490_;
  assign new_n1492_ = ~G4089 & ~G828;
  assign new_n1493_ = ~G4090 & new_n1492_;
  assign new_n1494_ = G4089 & ~G867;
  assign new_n1495_ = ~G4090 & new_n1494_;
  assign new_n1496_ = G100 & ~G4089;
  assign new_n1497_ = G4090 & new_n1496_;
  assign new_n1498_ = G103 & G4089;
  assign new_n1499_ = G4090 & new_n1498_;
  assign new_n1500_ = ~new_n1493_ & ~new_n1495_;
  assign new_n1501_ = ~new_n1497_ & ~new_n1499_;
  assign G777 = ~new_n1500_ | ~new_n1501_;
  assign new_n1503_ = ~G4089 & ~G830;
  assign new_n1504_ = ~G4090 & new_n1503_;
  assign new_n1505_ = G4089 & ~G869;
  assign new_n1506_ = ~G4090 & new_n1505_;
  assign new_n1507_ = G91 & ~G4089;
  assign new_n1508_ = G4090 & new_n1507_;
  assign new_n1509_ = G40 & G4089;
  assign new_n1510_ = G4090 & new_n1509_;
  assign new_n1511_ = ~new_n1504_ & ~new_n1506_;
  assign new_n1512_ = ~new_n1508_ & ~new_n1510_;
  assign G782 = ~new_n1511_ | ~new_n1512_;
  assign new_n1514_ = ~G1689 & ~G830;
  assign new_n1515_ = ~G1690 & new_n1514_;
  assign new_n1516_ = G1689 & ~G869;
  assign new_n1517_ = ~G1690 & new_n1516_;
  assign new_n1518_ = G203 & ~G1689;
  assign new_n1519_ = G1690 & new_n1518_;
  assign new_n1520_ = G173 & G1689;
  assign new_n1521_ = G1690 & new_n1520_;
  assign new_n1522_ = ~new_n1515_ & ~new_n1517_;
  assign new_n1523_ = ~new_n1519_ & ~new_n1521_;
  assign new_n1524_ = new_n1522_ & new_n1523_;
  assign G645 = G137 & ~new_n1524_;
  assign new_n1526_ = ~G1689 & ~G828;
  assign new_n1527_ = ~G1690 & new_n1526_;
  assign new_n1528_ = G1689 & ~G867;
  assign new_n1529_ = ~G1690 & new_n1528_;
  assign new_n1530_ = G197 & ~G1689;
  assign new_n1531_ = G1690 & new_n1530_;
  assign new_n1532_ = G167 & G1689;
  assign new_n1533_ = G1690 & new_n1532_;
  assign new_n1534_ = ~new_n1527_ & ~new_n1529_;
  assign new_n1535_ = ~new_n1531_ & ~new_n1533_;
  assign new_n1536_ = new_n1534_ & new_n1535_;
  assign G648 = G137 & ~new_n1536_;
  assign new_n1538_ = ~G1689 & ~G826;
  assign new_n1539_ = ~G1690 & new_n1538_;
  assign new_n1540_ = G1689 & ~G865;
  assign new_n1541_ = ~G1690 & new_n1540_;
  assign new_n1542_ = G194 & ~G1689;
  assign new_n1543_ = G1690 & new_n1542_;
  assign new_n1544_ = G164 & G1689;
  assign new_n1545_ = G1690 & new_n1544_;
  assign new_n1546_ = ~new_n1539_ & ~new_n1541_;
  assign new_n1547_ = ~new_n1543_ & ~new_n1545_;
  assign new_n1548_ = new_n1546_ & new_n1547_;
  assign G651 = G137 & ~new_n1548_;
  assign new_n1550_ = ~G1689 & ~G824;
  assign new_n1551_ = ~G1690 & new_n1550_;
  assign new_n1552_ = G1689 & ~G863;
  assign new_n1553_ = ~G1690 & new_n1552_;
  assign new_n1554_ = G191 & ~G1689;
  assign new_n1555_ = G1690 & new_n1554_;
  assign new_n1556_ = G161 & G1689;
  assign new_n1557_ = G1690 & new_n1556_;
  assign new_n1558_ = ~new_n1551_ & ~new_n1553_;
  assign new_n1559_ = ~new_n1555_ & ~new_n1557_;
  assign new_n1560_ = new_n1558_ & new_n1559_;
  assign G654 = G137 & ~new_n1560_;
  assign new_n1562_ = ~G1691 & ~G830;
  assign new_n1563_ = ~G1694 & new_n1562_;
  assign new_n1564_ = G1691 & ~G869;
  assign new_n1565_ = ~G1694 & new_n1564_;
  assign new_n1566_ = G203 & ~G1691;
  assign new_n1567_ = G1694 & new_n1566_;
  assign new_n1568_ = G173 & G1691;
  assign new_n1569_ = G1694 & new_n1568_;
  assign new_n1570_ = ~new_n1563_ & ~new_n1565_;
  assign new_n1571_ = ~new_n1567_ & ~new_n1569_;
  assign new_n1572_ = new_n1570_ & new_n1571_;
  assign G679 = G137 & ~new_n1572_;
  assign new_n1574_ = ~G1691 & ~G828;
  assign new_n1575_ = ~G1694 & new_n1574_;
  assign new_n1576_ = G1691 & ~G867;
  assign new_n1577_ = ~G1694 & new_n1576_;
  assign new_n1578_ = G197 & ~G1691;
  assign new_n1579_ = G1694 & new_n1578_;
  assign new_n1580_ = G167 & G1691;
  assign new_n1581_ = G1694 & new_n1580_;
  assign new_n1582_ = ~new_n1575_ & ~new_n1577_;
  assign new_n1583_ = ~new_n1579_ & ~new_n1581_;
  assign new_n1584_ = new_n1582_ & new_n1583_;
  assign G682 = G137 & ~new_n1584_;
  assign new_n1586_ = ~G1691 & ~G826;
  assign new_n1587_ = ~G1694 & new_n1586_;
  assign new_n1588_ = G1691 & ~G865;
  assign new_n1589_ = ~G1694 & new_n1588_;
  assign new_n1590_ = G194 & ~G1691;
  assign new_n1591_ = G1694 & new_n1590_;
  assign new_n1592_ = G164 & G1691;
  assign new_n1593_ = G1694 & new_n1592_;
  assign new_n1594_ = ~new_n1587_ & ~new_n1589_;
  assign new_n1595_ = ~new_n1591_ & ~new_n1593_;
  assign new_n1596_ = new_n1594_ & new_n1595_;
  assign G685 = G137 & ~new_n1596_;
  assign new_n1598_ = ~G1691 & ~G824;
  assign new_n1599_ = ~G1694 & new_n1598_;
  assign new_n1600_ = G1691 & ~G863;
  assign new_n1601_ = ~G1694 & new_n1600_;
  assign new_n1602_ = G191 & ~G1691;
  assign new_n1603_ = G1694 & new_n1602_;
  assign new_n1604_ = G161 & G1691;
  assign new_n1605_ = G1694 & new_n1604_;
  assign new_n1606_ = ~new_n1599_ & ~new_n1601_;
  assign new_n1607_ = ~new_n1603_ & ~new_n1605_;
  assign new_n1608_ = new_n1606_ & new_n1607_;
  assign G688 = G137 & ~new_n1608_;
  assign new_n1610_ = new_n362_ & ~new_n372_;
  assign new_n1611_ = ~new_n362_ & new_n372_;
  assign new_n1612_ = ~new_n1610_ & ~new_n1611_;
  assign new_n1613_ = new_n375_ & new_n378_;
  assign new_n1614_ = ~new_n375_ & ~new_n378_;
  assign new_n1615_ = ~new_n1613_ & ~new_n1614_;
  assign new_n1616_ = ~new_n1612_ & new_n1615_;
  assign new_n1617_ = new_n1612_ & ~new_n1615_;
  assign new_n1618_ = ~new_n1616_ & ~new_n1617_;
  assign new_n1619_ = G248 & G534;
  assign new_n1620_ = G351 & new_n1619_;
  assign new_n1621_ = G251 & G534;
  assign new_n1622_ = ~G351 & new_n1621_;
  assign new_n1623_ = ~new_n1620_ & ~new_n1622_;
  assign new_n1624_ = G242 & G351;
  assign new_n1625_ = G254 & ~G351;
  assign new_n1626_ = ~new_n1624_ & ~new_n1625_;
  assign new_n1627_ = ~G534 & new_n1626_;
  assign new_n1628_ = new_n1623_ & ~new_n1627_;
  assign new_n1629_ = G248 & G523;
  assign new_n1630_ = G341 & new_n1629_;
  assign new_n1631_ = G251 & G523;
  assign new_n1632_ = ~G341 & new_n1631_;
  assign new_n1633_ = ~new_n1630_ & ~new_n1632_;
  assign new_n1634_ = G242 & G341;
  assign new_n1635_ = G254 & ~G341;
  assign new_n1636_ = ~new_n1634_ & ~new_n1635_;
  assign new_n1637_ = ~G523 & new_n1636_;
  assign new_n1638_ = new_n1633_ & ~new_n1637_;
  assign new_n1639_ = new_n1628_ & ~new_n1638_;
  assign new_n1640_ = ~new_n1628_ & new_n1638_;
  assign new_n1641_ = ~new_n1639_ & ~new_n1640_;
  assign new_n1642_ = G248 & G514;
  assign new_n1643_ = ~G242 & ~G514;
  assign new_n1644_ = ~new_n1642_ & ~new_n1643_;
  assign new_n1645_ = G248 & G503;
  assign new_n1646_ = G324 & new_n1645_;
  assign new_n1647_ = G251 & G503;
  assign new_n1648_ = ~G324 & new_n1647_;
  assign new_n1649_ = ~new_n1646_ & ~new_n1648_;
  assign new_n1650_ = G242 & G324;
  assign new_n1651_ = G254 & ~G324;
  assign new_n1652_ = ~new_n1650_ & ~new_n1651_;
  assign new_n1653_ = ~G503 & new_n1652_;
  assign new_n1654_ = new_n1649_ & ~new_n1653_;
  assign new_n1655_ = new_n1644_ & ~new_n1654_;
  assign new_n1656_ = ~new_n1644_ & new_n1654_;
  assign new_n1657_ = ~new_n1655_ & ~new_n1656_;
  assign new_n1658_ = ~new_n420_ & new_n1641_;
  assign new_n1659_ = new_n1657_ & new_n1658_;
  assign new_n1660_ = new_n420_ & new_n1641_;
  assign new_n1661_ = ~new_n1657_ & new_n1660_;
  assign new_n1662_ = ~new_n1659_ & ~new_n1661_;
  assign new_n1663_ = new_n420_ & ~new_n1641_;
  assign new_n1664_ = new_n1657_ & new_n1663_;
  assign new_n1665_ = ~new_n420_ & ~new_n1641_;
  assign new_n1666_ = ~new_n1657_ & new_n1665_;
  assign new_n1667_ = ~new_n1664_ & ~new_n1666_;
  assign new_n1668_ = new_n1662_ & new_n1667_;
  assign new_n1669_ = ~new_n1618_ & new_n1668_;
  assign new_n1670_ = new_n1618_ & ~new_n1668_;
  assign new_n1671_ = ~new_n1669_ & ~new_n1670_;
  assign new_n1672_ = ~G4091 & new_n1671_;
  assign new_n1673_ = ~G4092 & new_n1672_;
  assign new_n1674_ = ~new_n851_ & new_n856_;
  assign new_n1675_ = ~new_n850_ & new_n870_;
  assign new_n1676_ = new_n611_ & new_n1675_;
  assign new_n1677_ = ~new_n611_ & ~new_n1675_;
  assign new_n1678_ = ~new_n1676_ & ~new_n1677_;
  assign new_n1679_ = new_n886_ & new_n1678_;
  assign new_n1680_ = ~new_n886_ & ~new_n1678_;
  assign new_n1681_ = ~new_n1679_ & ~new_n1680_;
  assign new_n1682_ = new_n1674_ & new_n1681_;
  assign new_n1683_ = ~new_n1674_ & ~new_n1681_;
  assign new_n1684_ = ~new_n1682_ & ~new_n1683_;
  assign new_n1685_ = new_n611_ & new_n1684_;
  assign new_n1686_ = ~new_n611_ & ~new_n1684_;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = ~new_n629_ & new_n1687_;
  assign new_n1689_ = new_n629_ & ~new_n1687_;
  assign new_n1690_ = ~new_n1688_ & ~new_n1689_;
  assign new_n1691_ = ~new_n623_ & new_n1690_;
  assign new_n1692_ = new_n623_ & ~new_n1690_;
  assign new_n1693_ = ~new_n1691_ & ~new_n1692_;
  assign new_n1694_ = ~new_n617_ & new_n1693_;
  assign new_n1695_ = new_n617_ & ~new_n1693_;
  assign new_n1696_ = ~new_n1694_ & ~new_n1695_;
  assign new_n1697_ = ~new_n608_ & new_n1696_;
  assign new_n1698_ = new_n608_ & ~new_n1696_;
  assign new_n1699_ = ~new_n1697_ & ~new_n1698_;
  assign new_n1700_ = ~G2174 & new_n1699_;
  assign new_n1701_ = new_n611_ & ~new_n617_;
  assign new_n1702_ = ~new_n608_ & new_n1701_;
  assign new_n1703_ = ~new_n629_ & new_n1702_;
  assign new_n1704_ = ~new_n851_ & ~new_n1703_;
  assign new_n1705_ = new_n856_ & new_n1704_;
  assign new_n1706_ = ~new_n638_ & new_n886_;
  assign new_n1707_ = ~new_n629_ & new_n1701_;
  assign new_n1708_ = ~new_n850_ & ~new_n1707_;
  assign new_n1709_ = new_n870_ & new_n1708_;
  assign new_n1710_ = ~new_n1706_ & new_n1709_;
  assign new_n1711_ = new_n1706_ & ~new_n1709_;
  assign new_n1712_ = ~new_n1710_ & ~new_n1711_;
  assign new_n1713_ = ~new_n1705_ & new_n1712_;
  assign new_n1714_ = new_n1705_ & ~new_n1712_;
  assign new_n1715_ = ~new_n1713_ & ~new_n1714_;
  assign new_n1716_ = new_n611_ & new_n1715_;
  assign new_n1717_ = ~new_n611_ & ~new_n1715_;
  assign new_n1718_ = ~new_n1716_ & ~new_n1717_;
  assign new_n1719_ = ~new_n629_ & new_n1718_;
  assign new_n1720_ = new_n629_ & ~new_n1718_;
  assign new_n1721_ = ~new_n1719_ & ~new_n1720_;
  assign new_n1722_ = ~new_n623_ & new_n1721_;
  assign new_n1723_ = new_n623_ & ~new_n1721_;
  assign new_n1724_ = ~new_n1722_ & ~new_n1723_;
  assign new_n1725_ = ~new_n617_ & new_n1724_;
  assign new_n1726_ = new_n617_ & ~new_n1724_;
  assign new_n1727_ = ~new_n1725_ & ~new_n1726_;
  assign new_n1728_ = ~new_n608_ & new_n1727_;
  assign new_n1729_ = new_n608_ & ~new_n1727_;
  assign new_n1730_ = ~new_n1728_ & ~new_n1729_;
  assign new_n1731_ = G2174 & ~new_n1730_;
  assign new_n1732_ = ~new_n1700_ & ~new_n1731_;
  assign new_n1733_ = ~new_n750_ & new_n1105_;
  assign new_n1734_ = new_n750_ & ~new_n1105_;
  assign new_n1735_ = ~new_n1733_ & ~new_n1734_;
  assign new_n1736_ = new_n820_ & new_n1735_;
  assign new_n1737_ = ~new_n820_ & ~new_n1735_;
  assign new_n1738_ = ~new_n1736_ & ~new_n1737_;
  assign new_n1739_ = ~new_n591_ & new_n1738_;
  assign new_n1740_ = new_n591_ & ~new_n1738_;
  assign new_n1741_ = ~new_n1739_ & ~new_n1740_;
  assign new_n1742_ = ~new_n597_ & new_n1741_;
  assign new_n1743_ = new_n597_ & ~new_n1741_;
  assign new_n1744_ = ~new_n1742_ & ~new_n1743_;
  assign new_n1745_ = new_n600_ & new_n1744_;
  assign new_n1746_ = ~new_n600_ & ~new_n1744_;
  assign new_n1747_ = ~new_n1745_ & ~new_n1746_;
  assign new_n1748_ = new_n585_ & new_n1747_;
  assign new_n1749_ = ~new_n585_ & ~new_n1747_;
  assign new_n1750_ = ~new_n1748_ & ~new_n1749_;
  assign new_n1751_ = new_n774_ & ~new_n1750_;
  assign new_n1752_ = ~G2174 & new_n1751_;
  assign new_n1753_ = ~new_n1099_ & ~new_n1110_;
  assign new_n1754_ = new_n1099_ & new_n1110_;
  assign new_n1755_ = ~new_n1753_ & ~new_n1754_;
  assign new_n1756_ = ~new_n828_ & new_n1755_;
  assign new_n1757_ = new_n828_ & ~new_n1755_;
  assign new_n1758_ = ~new_n1756_ & ~new_n1757_;
  assign new_n1759_ = ~new_n591_ & new_n1758_;
  assign new_n1760_ = new_n591_ & ~new_n1758_;
  assign new_n1761_ = ~new_n1759_ & ~new_n1760_;
  assign new_n1762_ = ~new_n597_ & new_n1761_;
  assign new_n1763_ = new_n597_ & ~new_n1761_;
  assign new_n1764_ = ~new_n1762_ & ~new_n1763_;
  assign new_n1765_ = new_n600_ & new_n1764_;
  assign new_n1766_ = ~new_n600_ & ~new_n1764_;
  assign new_n1767_ = ~new_n1765_ & ~new_n1766_;
  assign new_n1768_ = new_n585_ & new_n1767_;
  assign new_n1769_ = ~new_n585_ & ~new_n1767_;
  assign new_n1770_ = ~new_n1768_ & ~new_n1769_;
  assign new_n1771_ = ~new_n774_ & ~new_n1770_;
  assign new_n1772_ = ~G2174 & new_n1771_;
  assign new_n1773_ = ~new_n641_ & new_n774_;
  assign new_n1774_ = ~new_n1750_ & new_n1773_;
  assign new_n1775_ = G2174 & new_n1774_;
  assign new_n1776_ = ~new_n1770_ & ~new_n1773_;
  assign new_n1777_ = G2174 & new_n1776_;
  assign new_n1778_ = ~new_n1752_ & ~new_n1772_;
  assign new_n1779_ = ~new_n1775_ & ~new_n1777_;
  assign new_n1780_ = new_n1778_ & new_n1779_;
  assign new_n1781_ = ~new_n1732_ & new_n1780_;
  assign new_n1782_ = new_n1732_ & ~new_n1780_;
  assign new_n1783_ = ~new_n1781_ & ~new_n1782_;
  assign new_n1784_ = G4091 & ~new_n1783_;
  assign new_n1785_ = ~G4092 & new_n1784_;
  assign new_n1786_ = G120 & ~G4091;
  assign new_n1787_ = G4092 & new_n1786_;
  assign new_n1788_ = G4091 & G4092;
  assign new_n1789_ = ~new_n1673_ & ~new_n1785_;
  assign new_n1790_ = ~new_n1787_ & ~new_n1788_;
  assign G843 = ~new_n1789_ | ~new_n1790_;
  assign new_n1792_ = G248 & G422;
  assign new_n1793_ = G226 & new_n1792_;
  assign new_n1794_ = G251 & G422;
  assign new_n1795_ = ~G226 & new_n1794_;
  assign new_n1796_ = ~new_n1793_ & ~new_n1795_;
  assign new_n1797_ = G226 & G242;
  assign new_n1798_ = ~G226 & G254;
  assign new_n1799_ = ~new_n1797_ & ~new_n1798_;
  assign new_n1800_ = ~G422 & new_n1799_;
  assign new_n1801_ = new_n1796_ & ~new_n1800_;
  assign new_n1802_ = G248 & G468;
  assign new_n1803_ = G218 & new_n1802_;
  assign new_n1804_ = G251 & G468;
  assign new_n1805_ = ~G218 & new_n1804_;
  assign new_n1806_ = ~new_n1803_ & ~new_n1805_;
  assign new_n1807_ = G218 & G242;
  assign new_n1808_ = ~G218 & G254;
  assign new_n1809_ = ~new_n1807_ & ~new_n1808_;
  assign new_n1810_ = ~G468 & new_n1809_;
  assign new_n1811_ = new_n1806_ & ~new_n1810_;
  assign new_n1812_ = new_n1801_ & ~new_n1811_;
  assign new_n1813_ = ~new_n1801_ & new_n1811_;
  assign new_n1814_ = ~new_n1812_ & ~new_n1813_;
  assign new_n1815_ = G248 & G457;
  assign new_n1816_ = G210 & new_n1815_;
  assign new_n1817_ = G251 & G457;
  assign new_n1818_ = ~G210 & new_n1817_;
  assign new_n1819_ = ~new_n1816_ & ~new_n1818_;
  assign new_n1820_ = G210 & G242;
  assign new_n1821_ = ~G210 & G254;
  assign new_n1822_ = ~new_n1820_ & ~new_n1821_;
  assign new_n1823_ = ~G457 & new_n1822_;
  assign new_n1824_ = new_n1819_ & ~new_n1823_;
  assign new_n1825_ = ~new_n518_ & new_n1824_;
  assign new_n1826_ = new_n518_ & ~new_n1824_;
  assign new_n1827_ = ~new_n1825_ & ~new_n1826_;
  assign new_n1828_ = ~new_n1814_ & new_n1827_;
  assign new_n1829_ = new_n1814_ & ~new_n1827_;
  assign new_n1830_ = ~new_n1828_ & ~new_n1829_;
  assign new_n1831_ = G248 & G374;
  assign new_n1832_ = G281 & new_n1831_;
  assign new_n1833_ = G251 & G374;
  assign new_n1834_ = ~G281 & new_n1833_;
  assign new_n1835_ = ~new_n1832_ & ~new_n1834_;
  assign new_n1836_ = G242 & G281;
  assign new_n1837_ = G254 & ~G281;
  assign new_n1838_ = ~new_n1836_ & ~new_n1837_;
  assign new_n1839_ = ~G374 & new_n1838_;
  assign new_n1840_ = new_n1835_ & ~new_n1839_;
  assign new_n1841_ = G248 & G411;
  assign new_n1842_ = G273 & new_n1841_;
  assign new_n1843_ = G251 & G411;
  assign new_n1844_ = ~G273 & new_n1843_;
  assign new_n1845_ = ~new_n1842_ & ~new_n1844_;
  assign new_n1846_ = G242 & G273;
  assign new_n1847_ = G254 & ~G273;
  assign new_n1848_ = ~new_n1846_ & ~new_n1847_;
  assign new_n1849_ = ~G411 & new_n1848_;
  assign new_n1850_ = new_n1845_ & ~new_n1849_;
  assign new_n1851_ = G248 & G400;
  assign new_n1852_ = G265 & new_n1851_;
  assign new_n1853_ = G251 & G400;
  assign new_n1854_ = ~G265 & new_n1853_;
  assign new_n1855_ = ~new_n1852_ & ~new_n1854_;
  assign new_n1856_ = G242 & G265;
  assign new_n1857_ = G254 & ~G265;
  assign new_n1858_ = ~new_n1856_ & ~new_n1857_;
  assign new_n1859_ = ~G400 & new_n1858_;
  assign new_n1860_ = new_n1855_ & ~new_n1859_;
  assign new_n1861_ = new_n1850_ & ~new_n1860_;
  assign new_n1862_ = ~new_n1850_ & new_n1860_;
  assign new_n1863_ = ~new_n1861_ & ~new_n1862_;
  assign new_n1864_ = G248 & G389;
  assign new_n1865_ = G257 & new_n1864_;
  assign new_n1866_ = G251 & G389;
  assign new_n1867_ = ~G257 & new_n1866_;
  assign new_n1868_ = ~new_n1865_ & ~new_n1867_;
  assign new_n1869_ = G242 & G257;
  assign new_n1870_ = G254 & ~G257;
  assign new_n1871_ = ~new_n1869_ & ~new_n1870_;
  assign new_n1872_ = ~G389 & new_n1871_;
  assign new_n1873_ = new_n1868_ & ~new_n1872_;
  assign new_n1874_ = G248 & G435;
  assign new_n1875_ = G234 & new_n1874_;
  assign new_n1876_ = G251 & G435;
  assign new_n1877_ = ~G234 & new_n1876_;
  assign new_n1878_ = ~new_n1875_ & ~new_n1877_;
  assign new_n1879_ = G234 & G242;
  assign new_n1880_ = ~G234 & G254;
  assign new_n1881_ = ~new_n1879_ & ~new_n1880_;
  assign new_n1882_ = ~G435 & new_n1881_;
  assign new_n1883_ = new_n1878_ & ~new_n1882_;
  assign new_n1884_ = new_n1873_ & ~new_n1883_;
  assign new_n1885_ = ~new_n1873_ & new_n1883_;
  assign new_n1886_ = ~new_n1884_ & ~new_n1885_;
  assign new_n1887_ = ~new_n1840_ & new_n1863_;
  assign new_n1888_ = new_n1886_ & new_n1887_;
  assign new_n1889_ = new_n1840_ & new_n1863_;
  assign new_n1890_ = ~new_n1886_ & new_n1889_;
  assign new_n1891_ = ~new_n1888_ & ~new_n1890_;
  assign new_n1892_ = new_n1840_ & ~new_n1863_;
  assign new_n1893_ = new_n1886_ & new_n1892_;
  assign new_n1894_ = ~new_n1840_ & ~new_n1863_;
  assign new_n1895_ = ~new_n1886_ & new_n1894_;
  assign new_n1896_ = ~new_n1893_ & ~new_n1895_;
  assign new_n1897_ = new_n1891_ & new_n1896_;
  assign new_n1898_ = ~new_n1830_ & new_n1897_;
  assign new_n1899_ = new_n1830_ & ~new_n1897_;
  assign new_n1900_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1901_ = ~G4091 & new_n1900_;
  assign new_n1902_ = ~G4092 & new_n1901_;
  assign new_n1903_ = ~new_n914_ & new_n920_;
  assign new_n1904_ = ~new_n913_ & new_n934_;
  assign new_n1905_ = ~new_n735_ & new_n1904_;
  assign new_n1906_ = new_n735_ & ~new_n1904_;
  assign new_n1907_ = ~new_n1905_ & ~new_n1906_;
  assign new_n1908_ = new_n950_ & new_n1907_;
  assign new_n1909_ = ~new_n950_ & ~new_n1907_;
  assign new_n1910_ = ~new_n1908_ & ~new_n1909_;
  assign new_n1911_ = new_n1903_ & new_n1910_;
  assign new_n1912_ = ~new_n1903_ & ~new_n1910_;
  assign new_n1913_ = ~new_n1911_ & ~new_n1912_;
  assign new_n1914_ = ~new_n553_ & new_n1913_;
  assign new_n1915_ = new_n553_ & ~new_n1913_;
  assign new_n1916_ = ~new_n1914_ & ~new_n1915_;
  assign new_n1917_ = ~new_n559_ & new_n1916_;
  assign new_n1918_ = new_n559_ & ~new_n1916_;
  assign new_n1919_ = ~new_n1917_ & ~new_n1918_;
  assign new_n1920_ = ~new_n577_ & new_n1919_;
  assign new_n1921_ = new_n577_ & ~new_n1919_;
  assign new_n1922_ = ~new_n1920_ & ~new_n1921_;
  assign new_n1923_ = ~new_n565_ & new_n1922_;
  assign new_n1924_ = new_n565_ & ~new_n1922_;
  assign new_n1925_ = ~new_n1923_ & ~new_n1924_;
  assign new_n1926_ = ~new_n571_ & new_n1925_;
  assign new_n1927_ = new_n571_ & ~new_n1925_;
  assign new_n1928_ = ~new_n1926_ & ~new_n1927_;
  assign new_n1929_ = ~G1497 & new_n1928_;
  assign new_n1930_ = ~new_n553_ & ~new_n565_;
  assign new_n1931_ = ~new_n571_ & new_n1930_;
  assign new_n1932_ = ~new_n559_ & new_n1931_;
  assign new_n1933_ = ~new_n914_ & ~new_n1932_;
  assign new_n1934_ = new_n920_ & new_n1933_;
  assign new_n1935_ = ~new_n578_ & new_n950_;
  assign new_n1936_ = ~new_n559_ & new_n1930_;
  assign new_n1937_ = ~new_n913_ & ~new_n1936_;
  assign new_n1938_ = new_n934_ & new_n1937_;
  assign new_n1939_ = ~G374 & new_n550_;
  assign new_n1940_ = ~new_n1938_ & ~new_n1939_;
  assign new_n1941_ = new_n1938_ & new_n1939_;
  assign new_n1942_ = ~new_n1940_ & ~new_n1941_;
  assign new_n1943_ = ~new_n1935_ & new_n1942_;
  assign new_n1944_ = new_n1935_ & ~new_n1942_;
  assign new_n1945_ = ~new_n1943_ & ~new_n1944_;
  assign new_n1946_ = ~new_n1934_ & new_n1945_;
  assign new_n1947_ = new_n1934_ & ~new_n1945_;
  assign new_n1948_ = ~new_n1946_ & ~new_n1947_;
  assign new_n1949_ = ~new_n553_ & new_n1948_;
  assign new_n1950_ = new_n553_ & ~new_n1948_;
  assign new_n1951_ = ~new_n1949_ & ~new_n1950_;
  assign new_n1952_ = ~new_n559_ & new_n1951_;
  assign new_n1953_ = new_n559_ & ~new_n1951_;
  assign new_n1954_ = ~new_n1952_ & ~new_n1953_;
  assign new_n1955_ = ~new_n577_ & new_n1954_;
  assign new_n1956_ = new_n577_ & ~new_n1954_;
  assign new_n1957_ = ~new_n1955_ & ~new_n1956_;
  assign new_n1958_ = ~new_n565_ & new_n1957_;
  assign new_n1959_ = new_n565_ & ~new_n1957_;
  assign new_n1960_ = ~new_n1958_ & ~new_n1959_;
  assign new_n1961_ = ~new_n571_ & new_n1960_;
  assign new_n1962_ = new_n571_ & ~new_n1960_;
  assign new_n1963_ = ~new_n1961_ & ~new_n1962_;
  assign new_n1964_ = G1497 & ~new_n1963_;
  assign new_n1965_ = ~new_n1929_ & ~new_n1964_;
  assign new_n1966_ = ~new_n718_ & new_n1058_;
  assign new_n1967_ = new_n718_ & ~new_n1058_;
  assign new_n1968_ = ~new_n1966_ & ~new_n1967_;
  assign new_n1969_ = new_n1072_ & new_n1968_;
  assign new_n1970_ = ~new_n1072_ & ~new_n1968_;
  assign new_n1971_ = ~new_n1969_ & ~new_n1970_;
  assign new_n1972_ = ~new_n526_ & new_n1971_;
  assign new_n1973_ = new_n526_ & ~new_n1971_;
  assign new_n1974_ = ~new_n1972_ & ~new_n1973_;
  assign new_n1975_ = ~new_n532_ & new_n1974_;
  assign new_n1976_ = new_n532_ & ~new_n1974_;
  assign new_n1977_ = ~new_n1975_ & ~new_n1976_;
  assign new_n1978_ = ~new_n544_ & new_n1977_;
  assign new_n1979_ = new_n544_ & ~new_n1977_;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = ~new_n538_ & new_n1980_;
  assign new_n1982_ = new_n538_ & ~new_n1980_;
  assign new_n1983_ = ~new_n1981_ & ~new_n1982_;
  assign new_n1984_ = new_n743_ & ~new_n1983_;
  assign new_n1985_ = ~G1497 & new_n1984_;
  assign new_n1986_ = ~new_n1051_ & ~new_n1063_;
  assign new_n1987_ = new_n1051_ & new_n1063_;
  assign new_n1988_ = ~new_n1986_ & ~new_n1987_;
  assign new_n1989_ = ~new_n1078_ & new_n1988_;
  assign new_n1990_ = new_n1078_ & ~new_n1988_;
  assign new_n1991_ = ~new_n1989_ & ~new_n1990_;
  assign new_n1992_ = ~new_n526_ & new_n1991_;
  assign new_n1993_ = new_n526_ & ~new_n1991_;
  assign new_n1994_ = ~new_n1992_ & ~new_n1993_;
  assign new_n1995_ = ~new_n532_ & new_n1994_;
  assign new_n1996_ = new_n532_ & ~new_n1994_;
  assign new_n1997_ = ~new_n1995_ & ~new_n1996_;
  assign new_n1998_ = ~new_n544_ & new_n1997_;
  assign new_n1999_ = new_n544_ & ~new_n1997_;
  assign new_n2000_ = ~new_n1998_ & ~new_n1999_;
  assign new_n2001_ = ~new_n538_ & new_n2000_;
  assign new_n2002_ = new_n538_ & ~new_n2000_;
  assign new_n2003_ = ~new_n2001_ & ~new_n2002_;
  assign new_n2004_ = ~new_n743_ & ~new_n2003_;
  assign new_n2005_ = ~G1497 & new_n2004_;
  assign new_n2006_ = ~new_n581_ & new_n743_;
  assign new_n2007_ = ~new_n1983_ & new_n2006_;
  assign new_n2008_ = G1497 & new_n2007_;
  assign new_n2009_ = ~new_n2003_ & ~new_n2006_;
  assign new_n2010_ = G1497 & new_n2009_;
  assign new_n2011_ = ~new_n1985_ & ~new_n2005_;
  assign new_n2012_ = ~new_n2008_ & ~new_n2010_;
  assign new_n2013_ = new_n2011_ & new_n2012_;
  assign new_n2014_ = ~new_n1965_ & new_n2013_;
  assign new_n2015_ = new_n1965_ & ~new_n2013_;
  assign new_n2016_ = ~new_n2014_ & ~new_n2015_;
  assign new_n2017_ = G4091 & ~new_n2016_;
  assign new_n2018_ = ~G4092 & new_n2017_;
  assign new_n2019_ = G118 & ~G4091;
  assign new_n2020_ = G4092 & new_n2019_;
  assign new_n2021_ = ~new_n1902_ & ~new_n2018_;
  assign new_n2022_ = ~new_n1788_ & ~new_n2020_;
  assign G882 = ~new_n2021_ | ~new_n2022_;
  assign new_n2024_ = ~G4091 & ~new_n1671_;
  assign new_n2025_ = G4091 & new_n1783_;
  assign new_n2026_ = ~new_n2024_ & ~new_n2025_;
  assign new_n2027_ = ~G4092 & ~new_n2026_;
  assign new_n2028_ = G94 & G4092;
  assign new_n2029_ = ~new_n2027_ & ~new_n2028_;
  assign new_n2030_ = ~G4088 & ~new_n2029_;
  assign new_n2031_ = ~G4087 & new_n2030_;
  assign new_n2032_ = ~G4091 & ~new_n1900_;
  assign new_n2033_ = G4091 & new_n2016_;
  assign new_n2034_ = ~new_n2032_ & ~new_n2033_;
  assign new_n2035_ = ~G4092 & ~new_n2034_;
  assign new_n2036_ = G97 & G4092;
  assign new_n2037_ = ~new_n2035_ & ~new_n2036_;
  assign new_n2038_ = G4088 & ~new_n2037_;
  assign new_n2039_ = ~G4087 & new_n2038_;
  assign new_n2040_ = G14 & ~G4088;
  assign new_n2041_ = G4087 & new_n2040_;
  assign new_n2042_ = G64 & G4088;
  assign new_n2043_ = G4087 & new_n2042_;
  assign new_n2044_ = ~new_n2031_ & ~new_n2039_;
  assign new_n2045_ = ~new_n2041_ & ~new_n2043_;
  assign G767 = ~new_n2044_ | ~new_n2045_;
  assign new_n2047_ = ~G4089 & ~new_n2029_;
  assign new_n2048_ = ~G4090 & new_n2047_;
  assign new_n2049_ = G4089 & ~new_n2037_;
  assign new_n2050_ = ~G4090 & new_n2049_;
  assign new_n2051_ = G14 & ~G4089;
  assign new_n2052_ = G4090 & new_n2051_;
  assign new_n2053_ = G64 & G4089;
  assign new_n2054_ = G4090 & new_n2053_;
  assign new_n2055_ = ~new_n2048_ & ~new_n2050_;
  assign new_n2056_ = ~new_n2052_ & ~new_n2054_;
  assign G807 = ~new_n2055_ | ~new_n2056_;
  assign new_n2058_ = ~G1689 & ~new_n2029_;
  assign new_n2059_ = ~G1690 & new_n2058_;
  assign new_n2060_ = G1689 & ~new_n2037_;
  assign new_n2061_ = ~G1690 & new_n2060_;
  assign new_n2062_ = G176 & ~G1689;
  assign new_n2063_ = G1690 & new_n2062_;
  assign new_n2064_ = G179 & G1689;
  assign new_n2065_ = G1690 & new_n2064_;
  assign new_n2066_ = ~new_n2059_ & ~new_n2061_;
  assign new_n2067_ = ~new_n2063_ & ~new_n2065_;
  assign new_n2068_ = new_n2066_ & new_n2067_;
  assign G658 = ~G137 | new_n2068_;
  assign new_n2070_ = ~G1691 & ~new_n2029_;
  assign new_n2071_ = ~G1694 & new_n2070_;
  assign new_n2072_ = G1691 & ~new_n2037_;
  assign new_n2073_ = ~G1694 & new_n2072_;
  assign new_n2074_ = G176 & ~G1691;
  assign new_n2075_ = G1694 & new_n2074_;
  assign new_n2076_ = G179 & G1691;
  assign new_n2077_ = G1694 & new_n2076_;
  assign new_n2078_ = ~new_n2071_ & ~new_n2073_;
  assign new_n2079_ = ~new_n2075_ & ~new_n2077_;
  assign new_n2080_ = new_n2078_ & new_n2079_;
  assign G690 = ~G137 | new_n2080_;
  assign G594 = ~G545;
  assign G599 = ~G348;
  assign G600 = ~G366;
  assign G602 = ~G549;
  assign G611 = ~G338;
  assign G612 = ~G358;
  assign G848 = ~G245;
  assign G849 = ~G552;
  assign G850 = ~G562;
  assign G851 = ~G559;
  assign G593 = ~G299;
  assign G144 = G141;
  assign G298 = G293;
  assign G973 = G3173;
  assign G603 = G594;
  assign G604 = G594;
  assign G926 = G137;
  assign G923 = G141;
  assign G921 = G1;
  assign G892 = G549;
  assign G887 = G299;
  assign G606 = G602;
  assign G993 = G1;
  assign G978 = G1;
  assign G949 = G1;
  assign G939 = G1;
  assign G889 = G299;
  assign G717 = G704;
endmodule


