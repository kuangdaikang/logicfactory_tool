// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:38 2022

module e64  ( 
    i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_, i_10_,
    i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_, i_20_,
    i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_, i_30_,
    i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_, i_40_,
    i_41_, i_42_, i_43_, i_44_, i_45_, i_46_, i_47_, i_48_, i_49_, i_50_,
    i_51_, i_52_, i_53_, i_54_, i_55_, i_56_, i_57_, i_58_, i_59_, i_60_,
    i_61_, i_62_, i_63_, i_64_,
    o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_,
    o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_,
    o_61_, o_62_, o_63_, o_64_  );
  input  i_0_, i_1_, i_2_, i_3_, i_4_, i_5_, i_6_, i_7_, i_8_, i_9_,
    i_10_, i_11_, i_12_, i_13_, i_14_, i_15_, i_16_, i_17_, i_18_, i_19_,
    i_20_, i_21_, i_22_, i_23_, i_24_, i_25_, i_26_, i_27_, i_28_, i_29_,
    i_30_, i_31_, i_32_, i_33_, i_34_, i_35_, i_36_, i_37_, i_38_, i_39_,
    i_40_, i_41_, i_42_, i_43_, i_44_, i_45_, i_46_, i_47_, i_48_, i_49_,
    i_50_, i_51_, i_52_, i_53_, i_54_, i_55_, i_56_, i_57_, i_58_, i_59_,
    i_60_, i_61_, i_62_, i_63_, i_64_;
  output o_0_, o_1_, o_2_, o_3_, o_4_, o_5_, o_6_, o_7_, o_8_, o_9_, o_10_,
    o_11_, o_12_, o_13_, o_14_, o_15_, o_16_, o_17_, o_18_, o_19_, o_20_,
    o_21_, o_22_, o_23_, o_24_, o_25_, o_26_, o_27_, o_28_, o_29_, o_30_,
    o_31_, o_32_, o_33_, o_34_, o_35_, o_36_, o_37_, o_38_, o_39_, o_40_,
    o_41_, o_42_, o_43_, o_44_, o_45_, o_46_, o_47_, o_48_, o_49_, o_50_,
    o_51_, o_52_, o_53_, o_54_, o_55_, o_56_, o_57_, o_58_, o_59_, o_60_,
    o_61_, o_62_, o_63_, o_64_;
  wire new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_,
    new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_,
    new_n314_, new_n315_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n323_, new_n324_, new_n325_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n392_, new_n393_, new_n395_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_,
    new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1342_, new_n1343_, new_n1344_, new_n1345_,
    new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_,
    new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_,
    new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_,
    new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_,
    new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_,
    new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_,
    new_n1383_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1474_, new_n1475_, new_n1476_, new_n1477_,
    new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_,
    new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_,
    new_n1490_, new_n1491_, new_n1493_, new_n1494_, new_n1495_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1554_,
    new_n1555_, new_n1556_, new_n1558_, new_n1559_, new_n1560_, new_n1561_,
    new_n1562_, new_n1563_, new_n1564_, new_n1565_;
  assign new_n131_ = ~i_0_ & ~i_3_;
  assign new_n132_ = ~i_4_ & new_n131_;
  assign new_n133_ = ~i_5_ & new_n132_;
  assign new_n134_ = ~i_6_ & new_n133_;
  assign new_n135_ = ~i_7_ & new_n134_;
  assign new_n136_ = ~i_8_ & new_n135_;
  assign new_n137_ = ~i_9_ & new_n136_;
  assign new_n138_ = ~i_10_ & new_n137_;
  assign new_n139_ = ~i_11_ & new_n138_;
  assign new_n140_ = ~i_14_ & new_n139_;
  assign new_n141_ = ~i_15_ & new_n140_;
  assign new_n142_ = ~i_17_ & new_n141_;
  assign new_n143_ = ~i_18_ & new_n142_;
  assign new_n144_ = ~i_22_ & new_n143_;
  assign new_n145_ = ~i_24_ & new_n144_;
  assign new_n146_ = ~i_25_ & new_n145_;
  assign new_n147_ = ~i_26_ & new_n146_;
  assign new_n148_ = ~i_28_ & new_n147_;
  assign new_n149_ = i_29_ & new_n148_;
  assign new_n150_ = ~i_30_ & new_n149_;
  assign new_n151_ = ~i_31_ & new_n150_;
  assign new_n152_ = ~i_33_ & new_n151_;
  assign new_n153_ = ~i_34_ & new_n152_;
  assign new_n154_ = ~i_35_ & new_n153_;
  assign new_n155_ = ~i_37_ & new_n154_;
  assign new_n156_ = ~i_39_ & new_n155_;
  assign new_n157_ = ~i_40_ & new_n156_;
  assign new_n158_ = ~i_41_ & new_n157_;
  assign new_n159_ = ~i_42_ & new_n158_;
  assign new_n160_ = ~i_43_ & new_n159_;
  assign new_n161_ = i_45_ & new_n160_;
  assign new_n162_ = ~i_46_ & new_n161_;
  assign new_n163_ = ~i_47_ & new_n162_;
  assign new_n164_ = ~i_50_ & new_n163_;
  assign new_n165_ = ~i_51_ & new_n164_;
  assign new_n166_ = ~i_53_ & new_n165_;
  assign new_n167_ = ~i_54_ & new_n166_;
  assign new_n168_ = ~i_55_ & new_n167_;
  assign new_n169_ = ~i_56_ & new_n168_;
  assign new_n170_ = ~i_58_ & new_n169_;
  assign new_n171_ = ~i_59_ & new_n170_;
  assign new_n172_ = ~i_60_ & new_n171_;
  assign new_n173_ = ~i_61_ & new_n172_;
  assign o_0_ = ~i_62_ & new_n173_;
  assign new_n175_ = i_5_ & new_n132_;
  assign new_n176_ = ~i_6_ & new_n175_;
  assign new_n177_ = ~i_7_ & new_n176_;
  assign new_n178_ = ~i_8_ & new_n177_;
  assign new_n179_ = ~i_9_ & new_n178_;
  assign new_n180_ = ~i_10_ & new_n179_;
  assign new_n181_ = ~i_11_ & new_n180_;
  assign new_n182_ = ~i_14_ & new_n181_;
  assign new_n183_ = ~i_15_ & new_n182_;
  assign new_n184_ = ~i_17_ & new_n183_;
  assign new_n185_ = ~i_18_ & new_n184_;
  assign new_n186_ = ~i_22_ & new_n185_;
  assign new_n187_ = ~i_24_ & new_n186_;
  assign new_n188_ = ~i_25_ & new_n187_;
  assign new_n189_ = ~i_26_ & new_n188_;
  assign new_n190_ = ~i_28_ & new_n189_;
  assign new_n191_ = i_29_ & new_n190_;
  assign new_n192_ = ~i_30_ & new_n191_;
  assign new_n193_ = ~i_31_ & new_n192_;
  assign new_n194_ = ~i_33_ & new_n193_;
  assign new_n195_ = ~i_34_ & new_n194_;
  assign new_n196_ = ~i_35_ & new_n195_;
  assign new_n197_ = ~i_37_ & new_n196_;
  assign new_n198_ = ~i_39_ & new_n197_;
  assign new_n199_ = ~i_40_ & new_n198_;
  assign new_n200_ = ~i_41_ & new_n199_;
  assign new_n201_ = ~i_42_ & new_n200_;
  assign new_n202_ = ~i_43_ & new_n201_;
  assign new_n203_ = ~i_46_ & new_n202_;
  assign new_n204_ = ~i_47_ & new_n203_;
  assign new_n205_ = ~i_50_ & new_n204_;
  assign new_n206_ = ~i_51_ & new_n205_;
  assign new_n207_ = ~i_53_ & new_n206_;
  assign new_n208_ = ~i_54_ & new_n207_;
  assign new_n209_ = ~i_55_ & new_n208_;
  assign new_n210_ = ~i_56_ & new_n209_;
  assign new_n211_ = ~i_58_ & new_n210_;
  assign new_n212_ = ~i_59_ & new_n211_;
  assign new_n213_ = ~i_60_ & new_n212_;
  assign new_n214_ = ~i_61_ & new_n213_;
  assign o_1_ = ~i_62_ & new_n214_;
  assign new_n216_ = ~i_0_ & ~i_1_;
  assign new_n217_ = ~i_2_ & new_n216_;
  assign new_n218_ = ~i_3_ & new_n217_;
  assign new_n219_ = ~i_4_ & new_n218_;
  assign new_n220_ = ~i_5_ & new_n219_;
  assign new_n221_ = ~i_6_ & new_n220_;
  assign new_n222_ = ~i_7_ & new_n221_;
  assign new_n223_ = ~i_8_ & new_n222_;
  assign new_n224_ = ~i_9_ & new_n223_;
  assign new_n225_ = ~i_10_ & new_n224_;
  assign new_n226_ = ~i_11_ & new_n225_;
  assign new_n227_ = ~i_12_ & new_n226_;
  assign new_n228_ = ~i_13_ & new_n227_;
  assign new_n229_ = ~i_14_ & new_n228_;
  assign new_n230_ = ~i_15_ & new_n229_;
  assign new_n231_ = ~i_16_ & new_n230_;
  assign new_n232_ = ~i_17_ & new_n231_;
  assign new_n233_ = ~i_18_ & new_n232_;
  assign new_n234_ = ~i_19_ & new_n233_;
  assign new_n235_ = ~i_20_ & new_n234_;
  assign new_n236_ = ~i_21_ & new_n235_;
  assign new_n237_ = ~i_22_ & new_n236_;
  assign new_n238_ = ~i_23_ & new_n237_;
  assign new_n239_ = ~i_24_ & new_n238_;
  assign new_n240_ = ~i_25_ & new_n239_;
  assign new_n241_ = ~i_26_ & new_n240_;
  assign new_n242_ = i_27_ & new_n241_;
  assign new_n243_ = ~i_28_ & new_n242_;
  assign new_n244_ = i_29_ & new_n243_;
  assign new_n245_ = ~i_30_ & new_n244_;
  assign new_n246_ = ~i_31_ & new_n245_;
  assign new_n247_ = ~i_32_ & new_n246_;
  assign new_n248_ = ~i_33_ & new_n247_;
  assign new_n249_ = ~i_34_ & new_n248_;
  assign new_n250_ = ~i_35_ & new_n249_;
  assign new_n251_ = ~i_36_ & new_n250_;
  assign new_n252_ = ~i_37_ & new_n251_;
  assign new_n253_ = ~i_38_ & new_n252_;
  assign new_n254_ = ~i_39_ & new_n253_;
  assign new_n255_ = ~i_40_ & new_n254_;
  assign new_n256_ = ~i_41_ & new_n255_;
  assign new_n257_ = ~i_42_ & new_n256_;
  assign new_n258_ = ~i_43_ & new_n257_;
  assign new_n259_ = ~i_44_ & new_n258_;
  assign new_n260_ = ~i_45_ & new_n259_;
  assign new_n261_ = ~i_46_ & new_n260_;
  assign new_n262_ = ~i_47_ & new_n261_;
  assign new_n263_ = ~i_48_ & new_n262_;
  assign new_n264_ = ~i_49_ & new_n263_;
  assign new_n265_ = ~i_50_ & new_n264_;
  assign new_n266_ = ~i_51_ & new_n265_;
  assign new_n267_ = ~i_52_ & new_n266_;
  assign new_n268_ = ~i_53_ & new_n267_;
  assign new_n269_ = ~i_54_ & new_n268_;
  assign new_n270_ = ~i_55_ & new_n269_;
  assign new_n271_ = ~i_56_ & new_n270_;
  assign new_n272_ = ~i_57_ & new_n271_;
  assign new_n273_ = ~i_58_ & new_n272_;
  assign new_n274_ = ~i_59_ & new_n273_;
  assign new_n275_ = ~i_60_ & new_n274_;
  assign new_n276_ = ~i_61_ & new_n275_;
  assign new_n277_ = ~i_62_ & new_n276_;
  assign new_n278_ = ~i_63_ & new_n277_;
  assign o_2_ = ~i_64_ & new_n278_;
  assign new_n280_ = ~i_28_ & new_n241_;
  assign new_n281_ = i_29_ & new_n280_;
  assign new_n282_ = ~i_30_ & new_n281_;
  assign new_n283_ = ~i_31_ & new_n282_;
  assign new_n284_ = ~i_32_ & new_n283_;
  assign new_n285_ = ~i_33_ & new_n284_;
  assign new_n286_ = ~i_34_ & new_n285_;
  assign new_n287_ = ~i_35_ & new_n286_;
  assign new_n288_ = ~i_36_ & new_n287_;
  assign new_n289_ = ~i_37_ & new_n288_;
  assign new_n290_ = ~i_38_ & new_n289_;
  assign new_n291_ = ~i_39_ & new_n290_;
  assign new_n292_ = ~i_40_ & new_n291_;
  assign new_n293_ = ~i_41_ & new_n292_;
  assign new_n294_ = ~i_42_ & new_n293_;
  assign new_n295_ = ~i_43_ & new_n294_;
  assign new_n296_ = i_44_ & new_n295_;
  assign new_n297_ = ~i_45_ & new_n296_;
  assign new_n298_ = ~i_46_ & new_n297_;
  assign new_n299_ = ~i_47_ & new_n298_;
  assign new_n300_ = ~i_48_ & new_n299_;
  assign new_n301_ = ~i_49_ & new_n300_;
  assign new_n302_ = ~i_50_ & new_n301_;
  assign new_n303_ = ~i_51_ & new_n302_;
  assign new_n304_ = ~i_52_ & new_n303_;
  assign new_n305_ = ~i_53_ & new_n304_;
  assign new_n306_ = ~i_54_ & new_n305_;
  assign new_n307_ = ~i_55_ & new_n306_;
  assign new_n308_ = ~i_56_ & new_n307_;
  assign new_n309_ = ~i_57_ & new_n308_;
  assign new_n310_ = ~i_58_ & new_n309_;
  assign new_n311_ = ~i_59_ & new_n310_;
  assign new_n312_ = ~i_60_ & new_n311_;
  assign new_n313_ = ~i_61_ & new_n312_;
  assign new_n314_ = ~i_62_ & new_n313_;
  assign new_n315_ = ~i_63_ & new_n314_;
  assign o_3_ = ~i_64_ & new_n315_;
  assign o_4_ = i_15_ & i_29_;
  assign new_n318_ = i_14_ & ~i_15_;
  assign new_n319_ = ~i_28_ & new_n318_;
  assign new_n320_ = i_29_ & new_n319_;
  assign new_n321_ = ~i_37_ & new_n320_;
  assign o_6_ = ~i_43_ & new_n321_;
  assign new_n323_ = ~i_15_ & ~i_28_;
  assign new_n324_ = i_29_ & new_n323_;
  assign new_n325_ = ~i_37_ & new_n324_;
  assign o_7_ = i_43_ & new_n325_;
  assign new_n327_ = i_38_ & new_n289_;
  assign new_n328_ = ~i_39_ & new_n327_;
  assign new_n329_ = ~i_40_ & new_n328_;
  assign new_n330_ = ~i_41_ & new_n329_;
  assign new_n331_ = ~i_42_ & new_n330_;
  assign new_n332_ = ~i_43_ & new_n331_;
  assign new_n333_ = ~i_45_ & new_n332_;
  assign new_n334_ = ~i_46_ & new_n333_;
  assign new_n335_ = ~i_47_ & new_n334_;
  assign new_n336_ = ~i_48_ & new_n335_;
  assign new_n337_ = ~i_49_ & new_n336_;
  assign new_n338_ = ~i_50_ & new_n337_;
  assign new_n339_ = ~i_51_ & new_n338_;
  assign new_n340_ = ~i_52_ & new_n339_;
  assign new_n341_ = ~i_53_ & new_n340_;
  assign new_n342_ = ~i_54_ & new_n341_;
  assign new_n343_ = ~i_55_ & new_n342_;
  assign new_n344_ = ~i_56_ & new_n343_;
  assign new_n345_ = ~i_57_ & new_n344_;
  assign new_n346_ = ~i_58_ & new_n345_;
  assign new_n347_ = ~i_59_ & new_n346_;
  assign new_n348_ = ~i_60_ & new_n347_;
  assign new_n349_ = ~i_61_ & new_n348_;
  assign new_n350_ = ~i_62_ & new_n349_;
  assign new_n351_ = ~i_63_ & new_n350_;
  assign o_8_ = ~i_64_ & new_n351_;
  assign new_n353_ = i_23_ & new_n237_;
  assign new_n354_ = ~i_24_ & new_n353_;
  assign new_n355_ = ~i_25_ & new_n354_;
  assign new_n356_ = ~i_26_ & new_n355_;
  assign new_n357_ = ~i_28_ & new_n356_;
  assign new_n358_ = i_29_ & new_n357_;
  assign new_n359_ = ~i_30_ & new_n358_;
  assign new_n360_ = ~i_31_ & new_n359_;
  assign new_n361_ = ~i_32_ & new_n360_;
  assign new_n362_ = ~i_33_ & new_n361_;
  assign new_n363_ = ~i_34_ & new_n362_;
  assign new_n364_ = ~i_35_ & new_n363_;
  assign new_n365_ = ~i_36_ & new_n364_;
  assign new_n366_ = ~i_37_ & new_n365_;
  assign new_n367_ = ~i_39_ & new_n366_;
  assign new_n368_ = ~i_40_ & new_n367_;
  assign new_n369_ = ~i_41_ & new_n368_;
  assign new_n370_ = ~i_42_ & new_n369_;
  assign new_n371_ = ~i_43_ & new_n370_;
  assign new_n372_ = ~i_45_ & new_n371_;
  assign new_n373_ = ~i_46_ & new_n372_;
  assign new_n374_ = ~i_47_ & new_n373_;
  assign new_n375_ = ~i_48_ & new_n374_;
  assign new_n376_ = ~i_49_ & new_n375_;
  assign new_n377_ = ~i_50_ & new_n376_;
  assign new_n378_ = ~i_51_ & new_n377_;
  assign new_n379_ = ~i_52_ & new_n378_;
  assign new_n380_ = ~i_53_ & new_n379_;
  assign new_n381_ = ~i_54_ & new_n380_;
  assign new_n382_ = ~i_55_ & new_n381_;
  assign new_n383_ = ~i_56_ & new_n382_;
  assign new_n384_ = ~i_57_ & new_n383_;
  assign new_n385_ = ~i_58_ & new_n384_;
  assign new_n386_ = ~i_59_ & new_n385_;
  assign new_n387_ = ~i_60_ & new_n386_;
  assign new_n388_ = ~i_61_ & new_n387_;
  assign new_n389_ = ~i_62_ & new_n388_;
  assign new_n390_ = ~i_63_ & new_n389_;
  assign o_9_ = ~i_64_ & new_n390_;
  assign new_n392_ = ~i_15_ & i_28_;
  assign new_n393_ = i_29_ & new_n392_;
  assign o_10_ = ~i_37_ & new_n393_;
  assign new_n395_ = ~i_15_ & i_29_;
  assign o_11_ = i_37_ & new_n395_;
  assign new_n397_ = ~i_3_ & i_6_;
  assign new_n398_ = ~i_7_ & new_n397_;
  assign new_n399_ = ~i_8_ & new_n398_;
  assign new_n400_ = ~i_10_ & new_n399_;
  assign new_n401_ = ~i_11_ & new_n400_;
  assign new_n402_ = ~i_14_ & new_n401_;
  assign new_n403_ = ~i_15_ & new_n402_;
  assign new_n404_ = ~i_24_ & new_n403_;
  assign new_n405_ = ~i_25_ & new_n404_;
  assign new_n406_ = ~i_26_ & new_n405_;
  assign new_n407_ = ~i_28_ & new_n406_;
  assign new_n408_ = i_29_ & new_n407_;
  assign new_n409_ = ~i_30_ & new_n408_;
  assign new_n410_ = ~i_37_ & new_n409_;
  assign new_n411_ = ~i_39_ & new_n410_;
  assign new_n412_ = ~i_40_ & new_n411_;
  assign new_n413_ = ~i_41_ & new_n412_;
  assign new_n414_ = ~i_43_ & new_n413_;
  assign new_n415_ = ~i_46_ & new_n414_;
  assign new_n416_ = ~i_47_ & new_n415_;
  assign new_n417_ = ~i_50_ & new_n416_;
  assign new_n418_ = ~i_56_ & new_n417_;
  assign new_n419_ = ~i_58_ & new_n418_;
  assign new_n420_ = ~i_60_ & new_n419_;
  assign o_12_ = ~i_62_ & new_n420_;
  assign new_n422_ = ~i_3_ & ~i_7_;
  assign new_n423_ = ~i_8_ & new_n422_;
  assign new_n424_ = ~i_10_ & new_n423_;
  assign new_n425_ = ~i_11_ & new_n424_;
  assign new_n426_ = ~i_14_ & new_n425_;
  assign new_n427_ = ~i_15_ & new_n426_;
  assign new_n428_ = ~i_24_ & new_n427_;
  assign new_n429_ = ~i_25_ & new_n428_;
  assign new_n430_ = ~i_26_ & new_n429_;
  assign new_n431_ = ~i_28_ & new_n430_;
  assign new_n432_ = i_29_ & new_n431_;
  assign new_n433_ = ~i_30_ & new_n432_;
  assign new_n434_ = ~i_37_ & new_n433_;
  assign new_n435_ = ~i_39_ & new_n434_;
  assign new_n436_ = ~i_40_ & new_n435_;
  assign new_n437_ = i_41_ & new_n436_;
  assign new_n438_ = ~i_43_ & new_n437_;
  assign new_n439_ = ~i_46_ & new_n438_;
  assign new_n440_ = ~i_47_ & new_n439_;
  assign new_n441_ = ~i_50_ & new_n440_;
  assign new_n442_ = ~i_56_ & new_n441_;
  assign new_n443_ = ~i_58_ & new_n442_;
  assign new_n444_ = ~i_60_ & new_n443_;
  assign o_13_ = ~i_62_ & new_n444_;
  assign new_n446_ = ~i_10_ & ~i_14_;
  assign new_n447_ = ~i_15_ & new_n446_;
  assign new_n448_ = ~i_28_ & new_n447_;
  assign new_n449_ = i_29_ & new_n448_;
  assign new_n450_ = ~i_37_ & new_n449_;
  assign new_n451_ = ~i_43_ & new_n450_;
  assign new_n452_ = i_50_ & new_n451_;
  assign o_14_ = ~i_58_ & new_n452_;
  assign new_n454_ = i_10_ & ~i_14_;
  assign new_n455_ = ~i_15_ & new_n454_;
  assign new_n456_ = ~i_28_ & new_n455_;
  assign new_n457_ = i_29_ & new_n456_;
  assign new_n458_ = ~i_37_ & new_n457_;
  assign new_n459_ = ~i_43_ & new_n458_;
  assign o_15_ = ~i_58_ & new_n459_;
  assign new_n461_ = i_26_ & new_n429_;
  assign new_n462_ = ~i_28_ & new_n461_;
  assign new_n463_ = i_29_ & new_n462_;
  assign new_n464_ = ~i_30_ & new_n463_;
  assign new_n465_ = ~i_37_ & new_n464_;
  assign new_n466_ = ~i_39_ & new_n465_;
  assign new_n467_ = ~i_40_ & new_n466_;
  assign new_n468_ = ~i_43_ & new_n467_;
  assign new_n469_ = ~i_46_ & new_n468_;
  assign new_n470_ = ~i_47_ & new_n469_;
  assign new_n471_ = ~i_50_ & new_n470_;
  assign new_n472_ = ~i_56_ & new_n471_;
  assign new_n473_ = ~i_58_ & new_n472_;
  assign new_n474_ = ~i_60_ & new_n473_;
  assign o_16_ = ~i_62_ & new_n474_;
  assign new_n476_ = i_3_ & ~i_7_;
  assign new_n477_ = ~i_8_ & new_n476_;
  assign new_n478_ = ~i_10_ & new_n477_;
  assign new_n479_ = ~i_11_ & new_n478_;
  assign new_n480_ = ~i_14_ & new_n479_;
  assign new_n481_ = ~i_15_ & new_n480_;
  assign new_n482_ = ~i_24_ & new_n481_;
  assign new_n483_ = ~i_25_ & new_n482_;
  assign new_n484_ = ~i_28_ & new_n483_;
  assign new_n485_ = i_29_ & new_n484_;
  assign new_n486_ = ~i_30_ & new_n485_;
  assign new_n487_ = ~i_37_ & new_n486_;
  assign new_n488_ = ~i_39_ & new_n487_;
  assign new_n489_ = ~i_40_ & new_n488_;
  assign new_n490_ = ~i_43_ & new_n489_;
  assign new_n491_ = ~i_46_ & new_n490_;
  assign new_n492_ = ~i_47_ & new_n491_;
  assign new_n493_ = ~i_50_ & new_n492_;
  assign new_n494_ = ~i_56_ & new_n493_;
  assign new_n495_ = ~i_58_ & new_n494_;
  assign new_n496_ = ~i_60_ & new_n495_;
  assign o_17_ = ~i_62_ & new_n496_;
  assign new_n498_ = ~i_7_ & ~i_8_;
  assign new_n499_ = ~i_10_ & new_n498_;
  assign new_n500_ = ~i_11_ & new_n499_;
  assign new_n501_ = ~i_14_ & new_n500_;
  assign new_n502_ = ~i_15_ & new_n501_;
  assign new_n503_ = ~i_24_ & new_n502_;
  assign new_n504_ = ~i_25_ & new_n503_;
  assign new_n505_ = ~i_28_ & new_n504_;
  assign new_n506_ = i_29_ & new_n505_;
  assign new_n507_ = ~i_30_ & new_n506_;
  assign new_n508_ = ~i_37_ & new_n507_;
  assign new_n509_ = ~i_39_ & new_n508_;
  assign new_n510_ = ~i_40_ & new_n509_;
  assign new_n511_ = ~i_43_ & new_n510_;
  assign new_n512_ = ~i_46_ & new_n511_;
  assign new_n513_ = ~i_47_ & new_n512_;
  assign new_n514_ = ~i_50_ & new_n513_;
  assign new_n515_ = ~i_56_ & new_n514_;
  assign new_n516_ = ~i_58_ & new_n515_;
  assign new_n517_ = ~i_60_ & new_n516_;
  assign o_18_ = i_62_ & new_n517_;
  assign new_n519_ = ~i_14_ & new_n226_;
  assign new_n520_ = ~i_15_ & new_n519_;
  assign new_n521_ = ~i_17_ & new_n520_;
  assign new_n522_ = ~i_18_ & new_n521_;
  assign new_n523_ = ~i_22_ & new_n522_;
  assign new_n524_ = ~i_24_ & new_n523_;
  assign new_n525_ = ~i_25_ & new_n524_;
  assign new_n526_ = ~i_26_ & new_n525_;
  assign new_n527_ = ~i_28_ & new_n526_;
  assign new_n528_ = i_29_ & new_n527_;
  assign new_n529_ = ~i_30_ & new_n528_;
  assign new_n530_ = ~i_31_ & new_n529_;
  assign new_n531_ = ~i_33_ & new_n530_;
  assign new_n532_ = ~i_34_ & new_n531_;
  assign new_n533_ = ~i_35_ & new_n532_;
  assign new_n534_ = ~i_37_ & new_n533_;
  assign new_n535_ = ~i_39_ & new_n534_;
  assign new_n536_ = ~i_40_ & new_n535_;
  assign new_n537_ = ~i_41_ & new_n536_;
  assign new_n538_ = ~i_42_ & new_n537_;
  assign new_n539_ = ~i_43_ & new_n538_;
  assign new_n540_ = ~i_45_ & new_n539_;
  assign new_n541_ = ~i_46_ & new_n540_;
  assign new_n542_ = ~i_47_ & new_n541_;
  assign new_n543_ = ~i_48_ & new_n542_;
  assign new_n544_ = ~i_49_ & new_n543_;
  assign new_n545_ = ~i_50_ & new_n544_;
  assign new_n546_ = ~i_51_ & new_n545_;
  assign new_n547_ = ~i_53_ & new_n546_;
  assign new_n548_ = ~i_54_ & new_n547_;
  assign new_n549_ = ~i_55_ & new_n548_;
  assign new_n550_ = ~i_56_ & new_n549_;
  assign new_n551_ = ~i_57_ & new_n550_;
  assign new_n552_ = ~i_58_ & new_n551_;
  assign new_n553_ = ~i_59_ & new_n552_;
  assign new_n554_ = ~i_60_ & new_n553_;
  assign new_n555_ = ~i_61_ & new_n554_;
  assign new_n556_ = ~i_62_ & new_n555_;
  assign o_19_ = i_64_ & new_n556_;
  assign new_n558_ = ~i_6_ & new_n131_;
  assign new_n559_ = ~i_7_ & new_n558_;
  assign new_n560_ = ~i_8_ & new_n559_;
  assign new_n561_ = ~i_10_ & new_n560_;
  assign new_n562_ = ~i_11_ & new_n561_;
  assign new_n563_ = ~i_14_ & new_n562_;
  assign new_n564_ = ~i_15_ & new_n563_;
  assign new_n565_ = ~i_18_ & new_n564_;
  assign new_n566_ = ~i_22_ & new_n565_;
  assign new_n567_ = ~i_24_ & new_n566_;
  assign new_n568_ = ~i_25_ & new_n567_;
  assign new_n569_ = ~i_26_ & new_n568_;
  assign new_n570_ = ~i_28_ & new_n569_;
  assign new_n571_ = i_29_ & new_n570_;
  assign new_n572_ = ~i_30_ & new_n571_;
  assign new_n573_ = ~i_37_ & new_n572_;
  assign new_n574_ = ~i_39_ & new_n573_;
  assign new_n575_ = ~i_40_ & new_n574_;
  assign new_n576_ = ~i_41_ & new_n575_;
  assign new_n577_ = ~i_43_ & new_n576_;
  assign new_n578_ = ~i_46_ & new_n577_;
  assign new_n579_ = ~i_47_ & new_n578_;
  assign new_n580_ = ~i_50_ & new_n579_;
  assign new_n581_ = i_51_ & new_n580_;
  assign new_n582_ = ~i_56_ & new_n581_;
  assign new_n583_ = ~i_58_ & new_n582_;
  assign new_n584_ = ~i_60_ & new_n583_;
  assign o_20_ = ~i_62_ & new_n584_;
  assign new_n586_ = i_0_ & ~i_3_;
  assign new_n587_ = ~i_6_ & new_n586_;
  assign new_n588_ = ~i_7_ & new_n587_;
  assign new_n589_ = ~i_8_ & new_n588_;
  assign new_n590_ = ~i_10_ & new_n589_;
  assign new_n591_ = ~i_11_ & new_n590_;
  assign new_n592_ = ~i_14_ & new_n591_;
  assign new_n593_ = ~i_15_ & new_n592_;
  assign new_n594_ = ~i_18_ & new_n593_;
  assign new_n595_ = ~i_22_ & new_n594_;
  assign new_n596_ = ~i_24_ & new_n595_;
  assign new_n597_ = ~i_25_ & new_n596_;
  assign new_n598_ = ~i_26_ & new_n597_;
  assign new_n599_ = ~i_28_ & new_n598_;
  assign new_n600_ = i_29_ & new_n599_;
  assign new_n601_ = ~i_30_ & new_n600_;
  assign new_n602_ = ~i_37_ & new_n601_;
  assign new_n603_ = ~i_39_ & new_n602_;
  assign new_n604_ = ~i_40_ & new_n603_;
  assign new_n605_ = ~i_41_ & new_n604_;
  assign new_n606_ = ~i_43_ & new_n605_;
  assign new_n607_ = ~i_46_ & new_n606_;
  assign new_n608_ = ~i_47_ & new_n607_;
  assign new_n609_ = ~i_50_ & new_n608_;
  assign new_n610_ = ~i_56_ & new_n609_;
  assign new_n611_ = ~i_58_ & new_n610_;
  assign new_n612_ = ~i_60_ & new_n611_;
  assign o_21_ = ~i_62_ & new_n612_;
  assign new_n614_ = ~i_14_ & new_n227_;
  assign new_n615_ = ~i_15_ & new_n614_;
  assign new_n616_ = ~i_17_ & new_n615_;
  assign new_n617_ = ~i_18_ & new_n616_;
  assign new_n618_ = ~i_22_ & new_n617_;
  assign new_n619_ = ~i_24_ & new_n618_;
  assign new_n620_ = ~i_25_ & new_n619_;
  assign new_n621_ = ~i_26_ & new_n620_;
  assign new_n622_ = ~i_28_ & new_n621_;
  assign new_n623_ = i_29_ & new_n622_;
  assign new_n624_ = ~i_30_ & new_n623_;
  assign new_n625_ = ~i_31_ & new_n624_;
  assign new_n626_ = ~i_33_ & new_n625_;
  assign new_n627_ = ~i_34_ & new_n626_;
  assign new_n628_ = ~i_35_ & new_n627_;
  assign new_n629_ = i_36_ & new_n628_;
  assign new_n630_ = ~i_37_ & new_n629_;
  assign new_n631_ = ~i_39_ & new_n630_;
  assign new_n632_ = ~i_40_ & new_n631_;
  assign new_n633_ = ~i_41_ & new_n632_;
  assign new_n634_ = ~i_42_ & new_n633_;
  assign new_n635_ = ~i_43_ & new_n634_;
  assign new_n636_ = ~i_45_ & new_n635_;
  assign new_n637_ = ~i_46_ & new_n636_;
  assign new_n638_ = ~i_47_ & new_n637_;
  assign new_n639_ = ~i_48_ & new_n638_;
  assign new_n640_ = ~i_49_ & new_n639_;
  assign new_n641_ = ~i_50_ & new_n640_;
  assign new_n642_ = ~i_51_ & new_n641_;
  assign new_n643_ = ~i_53_ & new_n642_;
  assign new_n644_ = ~i_54_ & new_n643_;
  assign new_n645_ = ~i_55_ & new_n644_;
  assign new_n646_ = ~i_56_ & new_n645_;
  assign new_n647_ = ~i_57_ & new_n646_;
  assign new_n648_ = ~i_58_ & new_n647_;
  assign new_n649_ = ~i_59_ & new_n648_;
  assign new_n650_ = ~i_60_ & new_n649_;
  assign new_n651_ = ~i_61_ & new_n650_;
  assign new_n652_ = ~i_62_ & new_n651_;
  assign new_n653_ = ~i_63_ & new_n652_;
  assign o_22_ = ~i_64_ & new_n653_;
  assign new_n655_ = i_16_ & new_n615_;
  assign new_n656_ = ~i_17_ & new_n655_;
  assign new_n657_ = ~i_18_ & new_n656_;
  assign new_n658_ = ~i_21_ & new_n657_;
  assign new_n659_ = ~i_22_ & new_n658_;
  assign new_n660_ = ~i_24_ & new_n659_;
  assign new_n661_ = ~i_25_ & new_n660_;
  assign new_n662_ = ~i_26_ & new_n661_;
  assign new_n663_ = ~i_28_ & new_n662_;
  assign new_n664_ = i_29_ & new_n663_;
  assign new_n665_ = ~i_30_ & new_n664_;
  assign new_n666_ = ~i_31_ & new_n665_;
  assign new_n667_ = ~i_33_ & new_n666_;
  assign new_n668_ = ~i_34_ & new_n667_;
  assign new_n669_ = ~i_35_ & new_n668_;
  assign new_n670_ = ~i_36_ & new_n669_;
  assign new_n671_ = ~i_37_ & new_n670_;
  assign new_n672_ = ~i_39_ & new_n671_;
  assign new_n673_ = ~i_40_ & new_n672_;
  assign new_n674_ = ~i_41_ & new_n673_;
  assign new_n675_ = ~i_42_ & new_n674_;
  assign new_n676_ = ~i_43_ & new_n675_;
  assign new_n677_ = ~i_45_ & new_n676_;
  assign new_n678_ = ~i_46_ & new_n677_;
  assign new_n679_ = ~i_47_ & new_n678_;
  assign new_n680_ = ~i_48_ & new_n679_;
  assign new_n681_ = ~i_49_ & new_n680_;
  assign new_n682_ = ~i_50_ & new_n681_;
  assign new_n683_ = ~i_51_ & new_n682_;
  assign new_n684_ = ~i_52_ & new_n683_;
  assign new_n685_ = ~i_53_ & new_n684_;
  assign new_n686_ = ~i_54_ & new_n685_;
  assign new_n687_ = ~i_55_ & new_n686_;
  assign new_n688_ = ~i_56_ & new_n687_;
  assign new_n689_ = ~i_57_ & new_n688_;
  assign new_n690_ = ~i_58_ & new_n689_;
  assign new_n691_ = ~i_59_ & new_n690_;
  assign new_n692_ = ~i_60_ & new_n691_;
  assign new_n693_ = ~i_61_ & new_n692_;
  assign new_n694_ = ~i_62_ & new_n693_;
  assign new_n695_ = ~i_63_ & new_n694_;
  assign o_23_ = ~i_64_ & new_n695_;
  assign new_n697_ = ~i_10_ & i_11_;
  assign new_n698_ = ~i_14_ & new_n697_;
  assign new_n699_ = ~i_15_ & new_n698_;
  assign new_n700_ = ~i_24_ & new_n699_;
  assign new_n701_ = ~i_25_ & new_n700_;
  assign new_n702_ = ~i_28_ & new_n701_;
  assign new_n703_ = i_29_ & new_n702_;
  assign new_n704_ = ~i_37_ & new_n703_;
  assign new_n705_ = ~i_39_ & new_n704_;
  assign new_n706_ = ~i_40_ & new_n705_;
  assign new_n707_ = ~i_43_ & new_n706_;
  assign new_n708_ = ~i_46_ & new_n707_;
  assign new_n709_ = ~i_50_ & new_n708_;
  assign new_n710_ = ~i_58_ & new_n709_;
  assign o_24_ = ~i_60_ & new_n710_;
  assign new_n712_ = i_24_ & new_n447_;
  assign new_n713_ = ~i_25_ & new_n712_;
  assign new_n714_ = ~i_28_ & new_n713_;
  assign new_n715_ = i_29_ & new_n714_;
  assign new_n716_ = ~i_37_ & new_n715_;
  assign new_n717_ = ~i_39_ & new_n716_;
  assign new_n718_ = ~i_40_ & new_n717_;
  assign new_n719_ = ~i_43_ & new_n718_;
  assign new_n720_ = ~i_46_ & new_n719_;
  assign new_n721_ = ~i_50_ & new_n720_;
  assign new_n722_ = ~i_58_ & new_n721_;
  assign o_25_ = ~i_60_ & new_n722_;
  assign new_n724_ = ~i_20_ & new_n233_;
  assign new_n725_ = ~i_21_ & new_n724_;
  assign new_n726_ = ~i_22_ & new_n725_;
  assign new_n727_ = ~i_24_ & new_n726_;
  assign new_n728_ = ~i_25_ & new_n727_;
  assign new_n729_ = ~i_26_ & new_n728_;
  assign new_n730_ = ~i_28_ & new_n729_;
  assign new_n731_ = i_29_ & new_n730_;
  assign new_n732_ = ~i_30_ & new_n731_;
  assign new_n733_ = ~i_31_ & new_n732_;
  assign new_n734_ = i_32_ & new_n733_;
  assign new_n735_ = ~i_33_ & new_n734_;
  assign new_n736_ = ~i_34_ & new_n735_;
  assign new_n737_ = ~i_35_ & new_n736_;
  assign new_n738_ = ~i_36_ & new_n737_;
  assign new_n739_ = ~i_37_ & new_n738_;
  assign new_n740_ = ~i_39_ & new_n739_;
  assign new_n741_ = ~i_40_ & new_n740_;
  assign new_n742_ = ~i_41_ & new_n741_;
  assign new_n743_ = ~i_42_ & new_n742_;
  assign new_n744_ = ~i_43_ & new_n743_;
  assign new_n745_ = ~i_45_ & new_n744_;
  assign new_n746_ = ~i_46_ & new_n745_;
  assign new_n747_ = ~i_47_ & new_n746_;
  assign new_n748_ = ~i_48_ & new_n747_;
  assign new_n749_ = ~i_49_ & new_n748_;
  assign new_n750_ = ~i_50_ & new_n749_;
  assign new_n751_ = ~i_51_ & new_n750_;
  assign new_n752_ = ~i_52_ & new_n751_;
  assign new_n753_ = ~i_53_ & new_n752_;
  assign new_n754_ = ~i_54_ & new_n753_;
  assign new_n755_ = ~i_55_ & new_n754_;
  assign new_n756_ = ~i_56_ & new_n755_;
  assign new_n757_ = ~i_57_ & new_n756_;
  assign new_n758_ = ~i_58_ & new_n757_;
  assign new_n759_ = ~i_59_ & new_n758_;
  assign new_n760_ = ~i_60_ & new_n759_;
  assign new_n761_ = ~i_61_ & new_n760_;
  assign new_n762_ = ~i_62_ & new_n761_;
  assign new_n763_ = ~i_63_ & new_n762_;
  assign o_26_ = ~i_64_ & new_n763_;
  assign new_n765_ = i_13_ & new_n227_;
  assign new_n766_ = ~i_14_ & new_n765_;
  assign new_n767_ = ~i_15_ & new_n766_;
  assign new_n768_ = ~i_16_ & new_n767_;
  assign new_n769_ = ~i_17_ & new_n768_;
  assign new_n770_ = ~i_18_ & new_n769_;
  assign new_n771_ = ~i_20_ & new_n770_;
  assign new_n772_ = ~i_21_ & new_n771_;
  assign new_n773_ = ~i_22_ & new_n772_;
  assign new_n774_ = ~i_24_ & new_n773_;
  assign new_n775_ = ~i_25_ & new_n774_;
  assign new_n776_ = ~i_26_ & new_n775_;
  assign new_n777_ = ~i_28_ & new_n776_;
  assign new_n778_ = i_29_ & new_n777_;
  assign new_n779_ = ~i_30_ & new_n778_;
  assign new_n780_ = ~i_31_ & new_n779_;
  assign new_n781_ = ~i_33_ & new_n780_;
  assign new_n782_ = ~i_34_ & new_n781_;
  assign new_n783_ = ~i_35_ & new_n782_;
  assign new_n784_ = ~i_36_ & new_n783_;
  assign new_n785_ = ~i_37_ & new_n784_;
  assign new_n786_ = ~i_39_ & new_n785_;
  assign new_n787_ = ~i_40_ & new_n786_;
  assign new_n788_ = ~i_41_ & new_n787_;
  assign new_n789_ = ~i_42_ & new_n788_;
  assign new_n790_ = ~i_43_ & new_n789_;
  assign new_n791_ = ~i_45_ & new_n790_;
  assign new_n792_ = ~i_46_ & new_n791_;
  assign new_n793_ = ~i_47_ & new_n792_;
  assign new_n794_ = ~i_48_ & new_n793_;
  assign new_n795_ = ~i_49_ & new_n794_;
  assign new_n796_ = ~i_50_ & new_n795_;
  assign new_n797_ = ~i_51_ & new_n796_;
  assign new_n798_ = ~i_52_ & new_n797_;
  assign new_n799_ = ~i_53_ & new_n798_;
  assign new_n800_ = ~i_54_ & new_n799_;
  assign new_n801_ = ~i_55_ & new_n800_;
  assign new_n802_ = ~i_56_ & new_n801_;
  assign new_n803_ = ~i_57_ & new_n802_;
  assign new_n804_ = ~i_58_ & new_n803_;
  assign new_n805_ = ~i_59_ & new_n804_;
  assign new_n806_ = ~i_60_ & new_n805_;
  assign new_n807_ = ~i_61_ & new_n806_;
  assign new_n808_ = ~i_62_ & new_n807_;
  assign new_n809_ = ~i_63_ & new_n808_;
  assign o_27_ = ~i_64_ & new_n809_;
  assign new_n811_ = i_25_ & new_n447_;
  assign new_n812_ = ~i_28_ & new_n811_;
  assign new_n813_ = i_29_ & new_n812_;
  assign new_n814_ = ~i_37_ & new_n813_;
  assign new_n815_ = ~i_39_ & new_n814_;
  assign new_n816_ = ~i_40_ & new_n815_;
  assign new_n817_ = ~i_43_ & new_n816_;
  assign new_n818_ = ~i_46_ & new_n817_;
  assign new_n819_ = ~i_50_ & new_n818_;
  assign new_n820_ = ~i_58_ & new_n819_;
  assign o_28_ = ~i_60_ & new_n820_;
  assign new_n822_ = ~i_39_ & new_n450_;
  assign new_n823_ = ~i_40_ & new_n822_;
  assign new_n824_ = ~i_43_ & new_n823_;
  assign new_n825_ = ~i_46_ & new_n824_;
  assign new_n826_ = ~i_50_ & new_n825_;
  assign new_n827_ = ~i_58_ & new_n826_;
  assign o_29_ = i_60_ & new_n827_;
  assign new_n829_ = ~i_21_ & new_n617_;
  assign new_n830_ = ~i_22_ & new_n829_;
  assign new_n831_ = ~i_24_ & new_n830_;
  assign new_n832_ = ~i_25_ & new_n831_;
  assign new_n833_ = ~i_26_ & new_n832_;
  assign new_n834_ = ~i_28_ & new_n833_;
  assign new_n835_ = i_29_ & new_n834_;
  assign new_n836_ = ~i_30_ & new_n835_;
  assign new_n837_ = ~i_31_ & new_n836_;
  assign new_n838_ = ~i_33_ & new_n837_;
  assign new_n839_ = ~i_34_ & new_n838_;
  assign new_n840_ = ~i_35_ & new_n839_;
  assign new_n841_ = ~i_36_ & new_n840_;
  assign new_n842_ = ~i_37_ & new_n841_;
  assign new_n843_ = ~i_39_ & new_n842_;
  assign new_n844_ = ~i_40_ & new_n843_;
  assign new_n845_ = ~i_41_ & new_n844_;
  assign new_n846_ = ~i_42_ & new_n845_;
  assign new_n847_ = ~i_43_ & new_n846_;
  assign new_n848_ = ~i_45_ & new_n847_;
  assign new_n849_ = ~i_46_ & new_n848_;
  assign new_n850_ = ~i_47_ & new_n849_;
  assign new_n851_ = ~i_48_ & new_n850_;
  assign new_n852_ = ~i_49_ & new_n851_;
  assign new_n853_ = ~i_50_ & new_n852_;
  assign new_n854_ = ~i_51_ & new_n853_;
  assign new_n855_ = i_52_ & new_n854_;
  assign new_n856_ = ~i_53_ & new_n855_;
  assign new_n857_ = ~i_54_ & new_n856_;
  assign new_n858_ = ~i_55_ & new_n857_;
  assign new_n859_ = ~i_56_ & new_n858_;
  assign new_n860_ = ~i_57_ & new_n859_;
  assign new_n861_ = ~i_58_ & new_n860_;
  assign new_n862_ = ~i_59_ & new_n861_;
  assign new_n863_ = ~i_60_ & new_n862_;
  assign new_n864_ = ~i_61_ & new_n863_;
  assign new_n865_ = ~i_62_ & new_n864_;
  assign new_n866_ = ~i_63_ & new_n865_;
  assign o_30_ = ~i_64_ & new_n866_;
  assign new_n868_ = i_21_ & new_n617_;
  assign new_n869_ = ~i_22_ & new_n868_;
  assign new_n870_ = ~i_24_ & new_n869_;
  assign new_n871_ = ~i_25_ & new_n870_;
  assign new_n872_ = ~i_26_ & new_n871_;
  assign new_n873_ = ~i_28_ & new_n872_;
  assign new_n874_ = i_29_ & new_n873_;
  assign new_n875_ = ~i_30_ & new_n874_;
  assign new_n876_ = ~i_31_ & new_n875_;
  assign new_n877_ = ~i_33_ & new_n876_;
  assign new_n878_ = ~i_34_ & new_n877_;
  assign new_n879_ = ~i_35_ & new_n878_;
  assign new_n880_ = ~i_36_ & new_n879_;
  assign new_n881_ = ~i_37_ & new_n880_;
  assign new_n882_ = ~i_39_ & new_n881_;
  assign new_n883_ = ~i_40_ & new_n882_;
  assign new_n884_ = ~i_41_ & new_n883_;
  assign new_n885_ = ~i_42_ & new_n884_;
  assign new_n886_ = ~i_43_ & new_n885_;
  assign new_n887_ = ~i_45_ & new_n886_;
  assign new_n888_ = ~i_46_ & new_n887_;
  assign new_n889_ = ~i_47_ & new_n888_;
  assign new_n890_ = ~i_48_ & new_n889_;
  assign new_n891_ = ~i_49_ & new_n890_;
  assign new_n892_ = ~i_50_ & new_n891_;
  assign new_n893_ = ~i_51_ & new_n892_;
  assign new_n894_ = ~i_53_ & new_n893_;
  assign new_n895_ = ~i_54_ & new_n894_;
  assign new_n896_ = ~i_55_ & new_n895_;
  assign new_n897_ = ~i_56_ & new_n896_;
  assign new_n898_ = ~i_57_ & new_n897_;
  assign new_n899_ = ~i_58_ & new_n898_;
  assign new_n900_ = ~i_59_ & new_n899_;
  assign new_n901_ = ~i_60_ & new_n900_;
  assign new_n902_ = ~i_61_ & new_n901_;
  assign new_n903_ = ~i_62_ & new_n902_;
  assign new_n904_ = ~i_63_ & new_n903_;
  assign o_31_ = ~i_64_ & new_n904_;
  assign new_n906_ = i_46_ & new_n824_;
  assign new_n907_ = ~i_50_ & new_n906_;
  assign o_32_ = ~i_58_ & new_n907_;
  assign new_n909_ = i_39_ & new_n450_;
  assign new_n910_ = ~i_40_ & new_n909_;
  assign new_n911_ = ~i_43_ & new_n910_;
  assign new_n912_ = ~i_50_ & new_n911_;
  assign o_33_ = ~i_58_ & new_n912_;
  assign new_n914_ = ~i_14_ & ~i_15_;
  assign new_n915_ = ~i_28_ & new_n914_;
  assign new_n916_ = i_29_ & new_n915_;
  assign new_n917_ = ~i_37_ & new_n916_;
  assign new_n918_ = ~i_43_ & new_n917_;
  assign o_34_ = i_58_ & new_n918_;
  assign new_n920_ = i_4_ & new_n131_;
  assign new_n921_ = ~i_6_ & new_n920_;
  assign new_n922_ = ~i_7_ & new_n921_;
  assign new_n923_ = ~i_8_ & new_n922_;
  assign new_n924_ = ~i_10_ & new_n923_;
  assign new_n925_ = ~i_11_ & new_n924_;
  assign new_n926_ = ~i_14_ & new_n925_;
  assign new_n927_ = ~i_15_ & new_n926_;
  assign new_n928_ = ~i_18_ & new_n927_;
  assign new_n929_ = ~i_22_ & new_n928_;
  assign new_n930_ = ~i_24_ & new_n929_;
  assign new_n931_ = ~i_25_ & new_n930_;
  assign new_n932_ = ~i_26_ & new_n931_;
  assign new_n933_ = ~i_28_ & new_n932_;
  assign new_n934_ = i_29_ & new_n933_;
  assign new_n935_ = ~i_30_ & new_n934_;
  assign new_n936_ = ~i_35_ & new_n935_;
  assign new_n937_ = ~i_37_ & new_n936_;
  assign new_n938_ = ~i_39_ & new_n937_;
  assign new_n939_ = ~i_40_ & new_n938_;
  assign new_n940_ = ~i_41_ & new_n939_;
  assign new_n941_ = ~i_43_ & new_n940_;
  assign new_n942_ = ~i_46_ & new_n941_;
  assign new_n943_ = ~i_47_ & new_n942_;
  assign new_n944_ = ~i_50_ & new_n943_;
  assign new_n945_ = ~i_51_ & new_n944_;
  assign new_n946_ = ~i_55_ & new_n945_;
  assign new_n947_ = ~i_56_ & new_n946_;
  assign new_n948_ = ~i_58_ & new_n947_;
  assign new_n949_ = ~i_60_ & new_n948_;
  assign new_n950_ = ~i_61_ & new_n949_;
  assign o_35_ = ~i_62_ & new_n950_;
  assign new_n952_ = ~i_35_ & new_n572_;
  assign new_n953_ = ~i_37_ & new_n952_;
  assign new_n954_ = ~i_39_ & new_n953_;
  assign new_n955_ = ~i_40_ & new_n954_;
  assign new_n956_ = ~i_41_ & new_n955_;
  assign new_n957_ = ~i_43_ & new_n956_;
  assign new_n958_ = ~i_46_ & new_n957_;
  assign new_n959_ = ~i_47_ & new_n958_;
  assign new_n960_ = ~i_50_ & new_n959_;
  assign new_n961_ = ~i_51_ & new_n960_;
  assign new_n962_ = ~i_55_ & new_n961_;
  assign new_n963_ = ~i_56_ & new_n962_;
  assign new_n964_ = ~i_58_ & new_n963_;
  assign new_n965_ = ~i_60_ & new_n964_;
  assign new_n966_ = i_61_ & new_n965_;
  assign o_36_ = ~i_62_ & new_n966_;
  assign new_n968_ = i_19_ & new_n233_;
  assign new_n969_ = ~i_20_ & new_n968_;
  assign new_n970_ = ~i_21_ & new_n969_;
  assign new_n971_ = ~i_22_ & new_n970_;
  assign new_n972_ = ~i_24_ & new_n971_;
  assign new_n973_ = ~i_25_ & new_n972_;
  assign new_n974_ = ~i_26_ & new_n973_;
  assign new_n975_ = ~i_28_ & new_n974_;
  assign new_n976_ = i_29_ & new_n975_;
  assign new_n977_ = ~i_30_ & new_n976_;
  assign new_n978_ = ~i_31_ & new_n977_;
  assign new_n979_ = ~i_32_ & new_n978_;
  assign new_n980_ = ~i_33_ & new_n979_;
  assign new_n981_ = ~i_34_ & new_n980_;
  assign new_n982_ = ~i_35_ & new_n981_;
  assign new_n983_ = ~i_36_ & new_n982_;
  assign new_n984_ = ~i_37_ & new_n983_;
  assign new_n985_ = ~i_39_ & new_n984_;
  assign new_n986_ = ~i_40_ & new_n985_;
  assign new_n987_ = ~i_41_ & new_n986_;
  assign new_n988_ = ~i_42_ & new_n987_;
  assign new_n989_ = ~i_43_ & new_n988_;
  assign new_n990_ = ~i_45_ & new_n989_;
  assign new_n991_ = ~i_46_ & new_n990_;
  assign new_n992_ = ~i_47_ & new_n991_;
  assign new_n993_ = ~i_48_ & new_n992_;
  assign new_n994_ = ~i_49_ & new_n993_;
  assign new_n995_ = ~i_50_ & new_n994_;
  assign new_n996_ = ~i_51_ & new_n995_;
  assign new_n997_ = ~i_52_ & new_n996_;
  assign new_n998_ = ~i_53_ & new_n997_;
  assign new_n999_ = ~i_54_ & new_n998_;
  assign new_n1000_ = ~i_55_ & new_n999_;
  assign new_n1001_ = ~i_56_ & new_n1000_;
  assign new_n1002_ = ~i_57_ & new_n1001_;
  assign new_n1003_ = ~i_58_ & new_n1002_;
  assign new_n1004_ = ~i_59_ & new_n1003_;
  assign new_n1005_ = ~i_60_ & new_n1004_;
  assign new_n1006_ = ~i_61_ & new_n1005_;
  assign new_n1007_ = ~i_62_ & new_n1006_;
  assign new_n1008_ = ~i_63_ & new_n1007_;
  assign o_37_ = ~i_64_ & new_n1008_;
  assign new_n1010_ = ~i_6_ & new_n132_;
  assign new_n1011_ = ~i_7_ & new_n1010_;
  assign new_n1012_ = ~i_8_ & new_n1011_;
  assign new_n1013_ = ~i_10_ & new_n1012_;
  assign new_n1014_ = ~i_11_ & new_n1013_;
  assign new_n1015_ = ~i_14_ & new_n1014_;
  assign new_n1016_ = ~i_15_ & new_n1015_;
  assign new_n1017_ = ~i_18_ & new_n1016_;
  assign new_n1018_ = ~i_22_ & new_n1017_;
  assign new_n1019_ = ~i_24_ & new_n1018_;
  assign new_n1020_ = ~i_25_ & new_n1019_;
  assign new_n1021_ = ~i_26_ & new_n1020_;
  assign new_n1022_ = ~i_28_ & new_n1021_;
  assign new_n1023_ = i_29_ & new_n1022_;
  assign new_n1024_ = ~i_30_ & new_n1023_;
  assign new_n1025_ = ~i_35_ & new_n1024_;
  assign new_n1026_ = ~i_37_ & new_n1025_;
  assign new_n1027_ = ~i_39_ & new_n1026_;
  assign new_n1028_ = ~i_40_ & new_n1027_;
  assign new_n1029_ = ~i_41_ & new_n1028_;
  assign new_n1030_ = ~i_42_ & new_n1029_;
  assign new_n1031_ = ~i_43_ & new_n1030_;
  assign new_n1032_ = ~i_46_ & new_n1031_;
  assign new_n1033_ = ~i_47_ & new_n1032_;
  assign new_n1034_ = ~i_50_ & new_n1033_;
  assign new_n1035_ = ~i_51_ & new_n1034_;
  assign new_n1036_ = ~i_55_ & new_n1035_;
  assign new_n1037_ = ~i_56_ & new_n1036_;
  assign new_n1038_ = ~i_58_ & new_n1037_;
  assign new_n1039_ = i_59_ & new_n1038_;
  assign new_n1040_ = ~i_60_ & new_n1039_;
  assign new_n1041_ = ~i_61_ & new_n1040_;
  assign o_38_ = ~i_62_ & new_n1041_;
  assign new_n1043_ = i_42_ & new_n1029_;
  assign new_n1044_ = ~i_43_ & new_n1043_;
  assign new_n1045_ = ~i_46_ & new_n1044_;
  assign new_n1046_ = ~i_47_ & new_n1045_;
  assign new_n1047_ = ~i_50_ & new_n1046_;
  assign new_n1048_ = ~i_51_ & new_n1047_;
  assign new_n1049_ = ~i_55_ & new_n1048_;
  assign new_n1050_ = ~i_56_ & new_n1049_;
  assign new_n1051_ = ~i_58_ & new_n1050_;
  assign new_n1052_ = ~i_60_ & new_n1051_;
  assign new_n1053_ = ~i_61_ & new_n1052_;
  assign o_39_ = ~i_62_ & new_n1053_;
  assign new_n1055_ = ~i_9_ & new_n1012_;
  assign new_n1056_ = ~i_10_ & new_n1055_;
  assign new_n1057_ = ~i_11_ & new_n1056_;
  assign new_n1058_ = ~i_14_ & new_n1057_;
  assign new_n1059_ = ~i_15_ & new_n1058_;
  assign new_n1060_ = ~i_17_ & new_n1059_;
  assign new_n1061_ = ~i_18_ & new_n1060_;
  assign new_n1062_ = ~i_22_ & new_n1061_;
  assign new_n1063_ = ~i_24_ & new_n1062_;
  assign new_n1064_ = ~i_25_ & new_n1063_;
  assign new_n1065_ = ~i_26_ & new_n1064_;
  assign new_n1066_ = ~i_28_ & new_n1065_;
  assign new_n1067_ = i_29_ & new_n1066_;
  assign new_n1068_ = ~i_30_ & new_n1067_;
  assign new_n1069_ = ~i_33_ & new_n1068_;
  assign new_n1070_ = ~i_34_ & new_n1069_;
  assign new_n1071_ = ~i_35_ & new_n1070_;
  assign new_n1072_ = ~i_37_ & new_n1071_;
  assign new_n1073_ = ~i_39_ & new_n1072_;
  assign new_n1074_ = ~i_40_ & new_n1073_;
  assign new_n1075_ = ~i_41_ & new_n1074_;
  assign new_n1076_ = ~i_42_ & new_n1075_;
  assign new_n1077_ = ~i_43_ & new_n1076_;
  assign new_n1078_ = ~i_46_ & new_n1077_;
  assign new_n1079_ = ~i_47_ & new_n1078_;
  assign new_n1080_ = ~i_50_ & new_n1079_;
  assign new_n1081_ = ~i_51_ & new_n1080_;
  assign new_n1082_ = i_54_ & new_n1081_;
  assign new_n1083_ = ~i_55_ & new_n1082_;
  assign new_n1084_ = ~i_56_ & new_n1083_;
  assign new_n1085_ = ~i_58_ & new_n1084_;
  assign new_n1086_ = ~i_59_ & new_n1085_;
  assign new_n1087_ = ~i_60_ & new_n1086_;
  assign new_n1088_ = ~i_61_ & new_n1087_;
  assign o_40_ = ~i_62_ & new_n1088_;
  assign new_n1090_ = i_33_ & new_n1068_;
  assign new_n1091_ = ~i_34_ & new_n1090_;
  assign new_n1092_ = ~i_35_ & new_n1091_;
  assign new_n1093_ = ~i_37_ & new_n1092_;
  assign new_n1094_ = ~i_39_ & new_n1093_;
  assign new_n1095_ = ~i_40_ & new_n1094_;
  assign new_n1096_ = ~i_41_ & new_n1095_;
  assign new_n1097_ = ~i_42_ & new_n1096_;
  assign new_n1098_ = ~i_43_ & new_n1097_;
  assign new_n1099_ = ~i_46_ & new_n1098_;
  assign new_n1100_ = ~i_47_ & new_n1099_;
  assign new_n1101_ = ~i_50_ & new_n1100_;
  assign new_n1102_ = ~i_51_ & new_n1101_;
  assign new_n1103_ = ~i_55_ & new_n1102_;
  assign new_n1104_ = ~i_56_ & new_n1103_;
  assign new_n1105_ = ~i_58_ & new_n1104_;
  assign new_n1106_ = ~i_59_ & new_n1105_;
  assign new_n1107_ = ~i_60_ & new_n1106_;
  assign new_n1108_ = ~i_61_ & new_n1107_;
  assign o_41_ = ~i_62_ & new_n1108_;
  assign new_n1110_ = i_49_ & new_n542_;
  assign new_n1111_ = ~i_50_ & new_n1110_;
  assign new_n1112_ = ~i_51_ & new_n1111_;
  assign new_n1113_ = ~i_53_ & new_n1112_;
  assign new_n1114_ = ~i_54_ & new_n1113_;
  assign new_n1115_ = ~i_55_ & new_n1114_;
  assign new_n1116_ = ~i_56_ & new_n1115_;
  assign new_n1117_ = ~i_58_ & new_n1116_;
  assign new_n1118_ = ~i_59_ & new_n1117_;
  assign new_n1119_ = ~i_60_ & new_n1118_;
  assign new_n1120_ = ~i_61_ & new_n1119_;
  assign o_42_ = ~i_62_ & new_n1120_;
  assign new_n1122_ = ~i_0_ & i_1_;
  assign new_n1123_ = ~i_2_ & new_n1122_;
  assign new_n1124_ = ~i_3_ & new_n1123_;
  assign new_n1125_ = ~i_4_ & new_n1124_;
  assign new_n1126_ = ~i_5_ & new_n1125_;
  assign new_n1127_ = ~i_6_ & new_n1126_;
  assign new_n1128_ = ~i_7_ & new_n1127_;
  assign new_n1129_ = ~i_8_ & new_n1128_;
  assign new_n1130_ = ~i_9_ & new_n1129_;
  assign new_n1131_ = ~i_10_ & new_n1130_;
  assign new_n1132_ = ~i_11_ & new_n1131_;
  assign new_n1133_ = ~i_14_ & new_n1132_;
  assign new_n1134_ = ~i_15_ & new_n1133_;
  assign new_n1135_ = ~i_17_ & new_n1134_;
  assign new_n1136_ = ~i_18_ & new_n1135_;
  assign new_n1137_ = ~i_22_ & new_n1136_;
  assign new_n1138_ = ~i_24_ & new_n1137_;
  assign new_n1139_ = ~i_25_ & new_n1138_;
  assign new_n1140_ = ~i_26_ & new_n1139_;
  assign new_n1141_ = ~i_28_ & new_n1140_;
  assign new_n1142_ = i_29_ & new_n1141_;
  assign new_n1143_ = ~i_30_ & new_n1142_;
  assign new_n1144_ = ~i_31_ & new_n1143_;
  assign new_n1145_ = ~i_33_ & new_n1144_;
  assign new_n1146_ = ~i_34_ & new_n1145_;
  assign new_n1147_ = ~i_35_ & new_n1146_;
  assign new_n1148_ = ~i_37_ & new_n1147_;
  assign new_n1149_ = ~i_39_ & new_n1148_;
  assign new_n1150_ = ~i_40_ & new_n1149_;
  assign new_n1151_ = ~i_41_ & new_n1150_;
  assign new_n1152_ = ~i_42_ & new_n1151_;
  assign new_n1153_ = ~i_43_ & new_n1152_;
  assign new_n1154_ = ~i_45_ & new_n1153_;
  assign new_n1155_ = ~i_46_ & new_n1154_;
  assign new_n1156_ = ~i_47_ & new_n1155_;
  assign new_n1157_ = ~i_50_ & new_n1156_;
  assign new_n1158_ = ~i_51_ & new_n1157_;
  assign new_n1159_ = ~i_53_ & new_n1158_;
  assign new_n1160_ = ~i_54_ & new_n1159_;
  assign new_n1161_ = ~i_55_ & new_n1160_;
  assign new_n1162_ = ~i_56_ & new_n1161_;
  assign new_n1163_ = ~i_58_ & new_n1162_;
  assign new_n1164_ = ~i_59_ & new_n1163_;
  assign new_n1165_ = ~i_60_ & new_n1164_;
  assign new_n1166_ = ~i_61_ & new_n1165_;
  assign o_43_ = ~i_62_ & new_n1166_;
  assign new_n1168_ = ~i_0_ & i_2_;
  assign new_n1169_ = ~i_3_ & new_n1168_;
  assign new_n1170_ = ~i_4_ & new_n1169_;
  assign new_n1171_ = ~i_5_ & new_n1170_;
  assign new_n1172_ = ~i_6_ & new_n1171_;
  assign new_n1173_ = ~i_7_ & new_n1172_;
  assign new_n1174_ = ~i_8_ & new_n1173_;
  assign new_n1175_ = ~i_9_ & new_n1174_;
  assign new_n1176_ = ~i_10_ & new_n1175_;
  assign new_n1177_ = ~i_11_ & new_n1176_;
  assign new_n1178_ = ~i_14_ & new_n1177_;
  assign new_n1179_ = ~i_15_ & new_n1178_;
  assign new_n1180_ = ~i_17_ & new_n1179_;
  assign new_n1181_ = ~i_18_ & new_n1180_;
  assign new_n1182_ = ~i_22_ & new_n1181_;
  assign new_n1183_ = ~i_24_ & new_n1182_;
  assign new_n1184_ = ~i_25_ & new_n1183_;
  assign new_n1185_ = ~i_26_ & new_n1184_;
  assign new_n1186_ = ~i_28_ & new_n1185_;
  assign new_n1187_ = i_29_ & new_n1186_;
  assign new_n1188_ = ~i_30_ & new_n1187_;
  assign new_n1189_ = ~i_31_ & new_n1188_;
  assign new_n1190_ = ~i_33_ & new_n1189_;
  assign new_n1191_ = ~i_34_ & new_n1190_;
  assign new_n1192_ = ~i_35_ & new_n1191_;
  assign new_n1193_ = ~i_37_ & new_n1192_;
  assign new_n1194_ = ~i_39_ & new_n1193_;
  assign new_n1195_ = ~i_40_ & new_n1194_;
  assign new_n1196_ = ~i_41_ & new_n1195_;
  assign new_n1197_ = ~i_42_ & new_n1196_;
  assign new_n1198_ = ~i_43_ & new_n1197_;
  assign new_n1199_ = ~i_45_ & new_n1198_;
  assign new_n1200_ = ~i_46_ & new_n1199_;
  assign new_n1201_ = ~i_47_ & new_n1200_;
  assign new_n1202_ = ~i_50_ & new_n1201_;
  assign new_n1203_ = ~i_51_ & new_n1202_;
  assign new_n1204_ = ~i_53_ & new_n1203_;
  assign new_n1205_ = ~i_54_ & new_n1204_;
  assign new_n1206_ = ~i_55_ & new_n1205_;
  assign new_n1207_ = ~i_56_ & new_n1206_;
  assign new_n1208_ = ~i_58_ & new_n1207_;
  assign new_n1209_ = ~i_59_ & new_n1208_;
  assign new_n1210_ = ~i_60_ & new_n1209_;
  assign new_n1211_ = ~i_61_ & new_n1210_;
  assign o_44_ = ~i_62_ & new_n1211_;
  assign new_n1213_ = i_34_ & new_n1068_;
  assign new_n1214_ = ~i_35_ & new_n1213_;
  assign new_n1215_ = ~i_37_ & new_n1214_;
  assign new_n1216_ = ~i_39_ & new_n1215_;
  assign new_n1217_ = ~i_40_ & new_n1216_;
  assign new_n1218_ = ~i_41_ & new_n1217_;
  assign new_n1219_ = ~i_42_ & new_n1218_;
  assign new_n1220_ = ~i_43_ & new_n1219_;
  assign new_n1221_ = ~i_46_ & new_n1220_;
  assign new_n1222_ = ~i_47_ & new_n1221_;
  assign new_n1223_ = ~i_50_ & new_n1222_;
  assign new_n1224_ = ~i_51_ & new_n1223_;
  assign new_n1225_ = ~i_55_ & new_n1224_;
  assign new_n1226_ = ~i_56_ & new_n1225_;
  assign new_n1227_ = ~i_58_ & new_n1226_;
  assign new_n1228_ = ~i_59_ & new_n1227_;
  assign new_n1229_ = ~i_60_ & new_n1228_;
  assign new_n1230_ = ~i_61_ & new_n1229_;
  assign o_45_ = ~i_62_ & new_n1230_;
  assign new_n1232_ = i_9_ & new_n1012_;
  assign new_n1233_ = ~i_10_ & new_n1232_;
  assign new_n1234_ = ~i_11_ & new_n1233_;
  assign new_n1235_ = ~i_14_ & new_n1234_;
  assign new_n1236_ = ~i_15_ & new_n1235_;
  assign new_n1237_ = ~i_17_ & new_n1236_;
  assign new_n1238_ = ~i_18_ & new_n1237_;
  assign new_n1239_ = ~i_22_ & new_n1238_;
  assign new_n1240_ = ~i_24_ & new_n1239_;
  assign new_n1241_ = ~i_25_ & new_n1240_;
  assign new_n1242_ = ~i_26_ & new_n1241_;
  assign new_n1243_ = ~i_28_ & new_n1242_;
  assign new_n1244_ = i_29_ & new_n1243_;
  assign new_n1245_ = ~i_30_ & new_n1244_;
  assign new_n1246_ = ~i_35_ & new_n1245_;
  assign new_n1247_ = ~i_37_ & new_n1246_;
  assign new_n1248_ = ~i_39_ & new_n1247_;
  assign new_n1249_ = ~i_40_ & new_n1248_;
  assign new_n1250_ = ~i_41_ & new_n1249_;
  assign new_n1251_ = ~i_42_ & new_n1250_;
  assign new_n1252_ = ~i_43_ & new_n1251_;
  assign new_n1253_ = ~i_46_ & new_n1252_;
  assign new_n1254_ = ~i_47_ & new_n1253_;
  assign new_n1255_ = ~i_50_ & new_n1254_;
  assign new_n1256_ = ~i_51_ & new_n1255_;
  assign new_n1257_ = ~i_55_ & new_n1256_;
  assign new_n1258_ = ~i_56_ & new_n1257_;
  assign new_n1259_ = ~i_58_ & new_n1258_;
  assign new_n1260_ = ~i_59_ & new_n1259_;
  assign new_n1261_ = ~i_60_ & new_n1260_;
  assign new_n1262_ = ~i_61_ & new_n1261_;
  assign o_46_ = ~i_62_ & new_n1262_;
  assign new_n1264_ = i_17_ & new_n1016_;
  assign new_n1265_ = ~i_18_ & new_n1264_;
  assign new_n1266_ = ~i_22_ & new_n1265_;
  assign new_n1267_ = ~i_24_ & new_n1266_;
  assign new_n1268_ = ~i_25_ & new_n1267_;
  assign new_n1269_ = ~i_26_ & new_n1268_;
  assign new_n1270_ = ~i_28_ & new_n1269_;
  assign new_n1271_ = i_29_ & new_n1270_;
  assign new_n1272_ = ~i_30_ & new_n1271_;
  assign new_n1273_ = ~i_35_ & new_n1272_;
  assign new_n1274_ = ~i_37_ & new_n1273_;
  assign new_n1275_ = ~i_39_ & new_n1274_;
  assign new_n1276_ = ~i_40_ & new_n1275_;
  assign new_n1277_ = ~i_41_ & new_n1276_;
  assign new_n1278_ = ~i_42_ & new_n1277_;
  assign new_n1279_ = ~i_43_ & new_n1278_;
  assign new_n1280_ = ~i_46_ & new_n1279_;
  assign new_n1281_ = ~i_47_ & new_n1280_;
  assign new_n1282_ = ~i_50_ & new_n1281_;
  assign new_n1283_ = ~i_51_ & new_n1282_;
  assign new_n1284_ = ~i_55_ & new_n1283_;
  assign new_n1285_ = ~i_56_ & new_n1284_;
  assign new_n1286_ = ~i_58_ & new_n1285_;
  assign new_n1287_ = ~i_59_ & new_n1286_;
  assign new_n1288_ = ~i_60_ & new_n1287_;
  assign new_n1289_ = ~i_61_ & new_n1288_;
  assign o_47_ = ~i_62_ & new_n1289_;
  assign new_n1291_ = i_31_ & new_n1068_;
  assign new_n1292_ = ~i_33_ & new_n1291_;
  assign new_n1293_ = ~i_34_ & new_n1292_;
  assign new_n1294_ = ~i_35_ & new_n1293_;
  assign new_n1295_ = ~i_37_ & new_n1294_;
  assign new_n1296_ = ~i_39_ & new_n1295_;
  assign new_n1297_ = ~i_40_ & new_n1296_;
  assign new_n1298_ = ~i_41_ & new_n1297_;
  assign new_n1299_ = ~i_42_ & new_n1298_;
  assign new_n1300_ = ~i_43_ & new_n1299_;
  assign new_n1301_ = ~i_46_ & new_n1300_;
  assign new_n1302_ = ~i_47_ & new_n1301_;
  assign new_n1303_ = ~i_50_ & new_n1302_;
  assign new_n1304_ = ~i_51_ & new_n1303_;
  assign new_n1305_ = ~i_53_ & new_n1304_;
  assign new_n1306_ = ~i_54_ & new_n1305_;
  assign new_n1307_ = ~i_55_ & new_n1306_;
  assign new_n1308_ = ~i_56_ & new_n1307_;
  assign new_n1309_ = ~i_58_ & new_n1308_;
  assign new_n1310_ = ~i_59_ & new_n1309_;
  assign new_n1311_ = ~i_60_ & new_n1310_;
  assign new_n1312_ = ~i_61_ & new_n1311_;
  assign o_48_ = ~i_62_ & new_n1312_;
  assign new_n1314_ = i_53_ & new_n1081_;
  assign new_n1315_ = ~i_54_ & new_n1314_;
  assign new_n1316_ = ~i_55_ & new_n1315_;
  assign new_n1317_ = ~i_56_ & new_n1316_;
  assign new_n1318_ = ~i_58_ & new_n1317_;
  assign new_n1319_ = ~i_59_ & new_n1318_;
  assign new_n1320_ = ~i_60_ & new_n1319_;
  assign new_n1321_ = ~i_61_ & new_n1320_;
  assign o_49_ = ~i_62_ & new_n1321_;
  assign new_n1323_ = i_57_ & new_n550_;
  assign new_n1324_ = ~i_58_ & new_n1323_;
  assign new_n1325_ = ~i_59_ & new_n1324_;
  assign new_n1326_ = ~i_60_ & new_n1325_;
  assign new_n1327_ = ~i_61_ & new_n1326_;
  assign o_50_ = ~i_62_ & new_n1327_;
  assign new_n1329_ = i_48_ & new_n542_;
  assign new_n1330_ = ~i_49_ & new_n1329_;
  assign new_n1331_ = ~i_50_ & new_n1330_;
  assign new_n1332_ = ~i_51_ & new_n1331_;
  assign new_n1333_ = ~i_53_ & new_n1332_;
  assign new_n1334_ = ~i_54_ & new_n1333_;
  assign new_n1335_ = ~i_55_ & new_n1334_;
  assign new_n1336_ = ~i_56_ & new_n1335_;
  assign new_n1337_ = ~i_58_ & new_n1336_;
  assign new_n1338_ = ~i_59_ & new_n1337_;
  assign new_n1339_ = ~i_60_ & new_n1338_;
  assign new_n1340_ = ~i_61_ & new_n1339_;
  assign o_51_ = ~i_62_ & new_n1340_;
  assign new_n1342_ = i_12_ & new_n226_;
  assign new_n1343_ = ~i_14_ & new_n1342_;
  assign new_n1344_ = ~i_15_ & new_n1343_;
  assign new_n1345_ = ~i_17_ & new_n1344_;
  assign new_n1346_ = ~i_18_ & new_n1345_;
  assign new_n1347_ = ~i_22_ & new_n1346_;
  assign new_n1348_ = ~i_24_ & new_n1347_;
  assign new_n1349_ = ~i_25_ & new_n1348_;
  assign new_n1350_ = ~i_26_ & new_n1349_;
  assign new_n1351_ = ~i_28_ & new_n1350_;
  assign new_n1352_ = i_29_ & new_n1351_;
  assign new_n1353_ = ~i_30_ & new_n1352_;
  assign new_n1354_ = ~i_31_ & new_n1353_;
  assign new_n1355_ = ~i_33_ & new_n1354_;
  assign new_n1356_ = ~i_34_ & new_n1355_;
  assign new_n1357_ = ~i_35_ & new_n1356_;
  assign new_n1358_ = ~i_37_ & new_n1357_;
  assign new_n1359_ = ~i_39_ & new_n1358_;
  assign new_n1360_ = ~i_40_ & new_n1359_;
  assign new_n1361_ = ~i_41_ & new_n1360_;
  assign new_n1362_ = ~i_42_ & new_n1361_;
  assign new_n1363_ = ~i_43_ & new_n1362_;
  assign new_n1364_ = ~i_45_ & new_n1363_;
  assign new_n1365_ = ~i_46_ & new_n1364_;
  assign new_n1366_ = ~i_47_ & new_n1365_;
  assign new_n1367_ = ~i_48_ & new_n1366_;
  assign new_n1368_ = ~i_49_ & new_n1367_;
  assign new_n1369_ = ~i_50_ & new_n1368_;
  assign new_n1370_ = ~i_51_ & new_n1369_;
  assign new_n1371_ = ~i_53_ & new_n1370_;
  assign new_n1372_ = ~i_54_ & new_n1371_;
  assign new_n1373_ = ~i_55_ & new_n1372_;
  assign new_n1374_ = ~i_56_ & new_n1373_;
  assign new_n1375_ = ~i_57_ & new_n1374_;
  assign new_n1376_ = ~i_58_ & new_n1375_;
  assign new_n1377_ = ~i_59_ & new_n1376_;
  assign new_n1378_ = ~i_60_ & new_n1377_;
  assign new_n1379_ = ~i_61_ & new_n1378_;
  assign new_n1380_ = ~i_62_ & new_n1379_;
  assign new_n1381_ = ~i_63_ & new_n1380_;
  assign o_52_ = ~i_64_ & new_n1381_;
  assign new_n1383_ = i_63_ & new_n556_;
  assign o_53_ = ~i_64_ & new_n1383_;
  assign new_n1385_ = i_55_ & new_n961_;
  assign new_n1386_ = ~i_56_ & new_n1385_;
  assign new_n1387_ = ~i_58_ & new_n1386_;
  assign new_n1388_ = ~i_60_ & new_n1387_;
  assign o_54_ = ~i_62_ & new_n1388_;
  assign new_n1390_ = i_35_ & new_n572_;
  assign new_n1391_ = ~i_37_ & new_n1390_;
  assign new_n1392_ = ~i_39_ & new_n1391_;
  assign new_n1393_ = ~i_40_ & new_n1392_;
  assign new_n1394_ = ~i_41_ & new_n1393_;
  assign new_n1395_ = ~i_43_ & new_n1394_;
  assign new_n1396_ = ~i_46_ & new_n1395_;
  assign new_n1397_ = ~i_47_ & new_n1396_;
  assign new_n1398_ = ~i_50_ & new_n1397_;
  assign new_n1399_ = ~i_51_ & new_n1398_;
  assign new_n1400_ = ~i_56_ & new_n1399_;
  assign new_n1401_ = ~i_58_ & new_n1400_;
  assign new_n1402_ = ~i_60_ & new_n1401_;
  assign o_55_ = ~i_62_ & new_n1402_;
  assign new_n1404_ = ~i_16_ & new_n615_;
  assign new_n1405_ = ~i_17_ & new_n1404_;
  assign new_n1406_ = ~i_18_ & new_n1405_;
  assign new_n1407_ = i_20_ & new_n1406_;
  assign new_n1408_ = ~i_21_ & new_n1407_;
  assign new_n1409_ = ~i_22_ & new_n1408_;
  assign new_n1410_ = ~i_24_ & new_n1409_;
  assign new_n1411_ = ~i_25_ & new_n1410_;
  assign new_n1412_ = ~i_26_ & new_n1411_;
  assign new_n1413_ = ~i_28_ & new_n1412_;
  assign new_n1414_ = i_29_ & new_n1413_;
  assign new_n1415_ = ~i_30_ & new_n1414_;
  assign new_n1416_ = ~i_31_ & new_n1415_;
  assign new_n1417_ = ~i_33_ & new_n1416_;
  assign new_n1418_ = ~i_34_ & new_n1417_;
  assign new_n1419_ = ~i_35_ & new_n1418_;
  assign new_n1420_ = ~i_36_ & new_n1419_;
  assign new_n1421_ = ~i_37_ & new_n1420_;
  assign new_n1422_ = ~i_39_ & new_n1421_;
  assign new_n1423_ = ~i_40_ & new_n1422_;
  assign new_n1424_ = ~i_41_ & new_n1423_;
  assign new_n1425_ = ~i_42_ & new_n1424_;
  assign new_n1426_ = ~i_43_ & new_n1425_;
  assign new_n1427_ = ~i_45_ & new_n1426_;
  assign new_n1428_ = ~i_46_ & new_n1427_;
  assign new_n1429_ = ~i_47_ & new_n1428_;
  assign new_n1430_ = ~i_48_ & new_n1429_;
  assign new_n1431_ = ~i_49_ & new_n1430_;
  assign new_n1432_ = ~i_50_ & new_n1431_;
  assign new_n1433_ = ~i_51_ & new_n1432_;
  assign new_n1434_ = ~i_52_ & new_n1433_;
  assign new_n1435_ = ~i_53_ & new_n1434_;
  assign new_n1436_ = ~i_54_ & new_n1435_;
  assign new_n1437_ = ~i_55_ & new_n1436_;
  assign new_n1438_ = ~i_56_ & new_n1437_;
  assign new_n1439_ = ~i_57_ & new_n1438_;
  assign new_n1440_ = ~i_58_ & new_n1439_;
  assign new_n1441_ = ~i_59_ & new_n1440_;
  assign new_n1442_ = ~i_60_ & new_n1441_;
  assign new_n1443_ = ~i_61_ & new_n1442_;
  assign new_n1444_ = ~i_62_ & new_n1443_;
  assign new_n1445_ = ~i_63_ & new_n1444_;
  assign o_56_ = ~i_64_ & new_n1445_;
  assign new_n1447_ = ~i_3_ & ~i_6_;
  assign new_n1448_ = ~i_7_ & new_n1447_;
  assign new_n1449_ = ~i_8_ & new_n1448_;
  assign new_n1450_ = ~i_10_ & new_n1449_;
  assign new_n1451_ = ~i_11_ & new_n1450_;
  assign new_n1452_ = ~i_14_ & new_n1451_;
  assign new_n1453_ = ~i_15_ & new_n1452_;
  assign new_n1454_ = i_18_ & new_n1453_;
  assign new_n1455_ = ~i_22_ & new_n1454_;
  assign new_n1456_ = ~i_24_ & new_n1455_;
  assign new_n1457_ = ~i_25_ & new_n1456_;
  assign new_n1458_ = ~i_26_ & new_n1457_;
  assign new_n1459_ = ~i_28_ & new_n1458_;
  assign new_n1460_ = i_29_ & new_n1459_;
  assign new_n1461_ = ~i_30_ & new_n1460_;
  assign new_n1462_ = ~i_37_ & new_n1461_;
  assign new_n1463_ = ~i_39_ & new_n1462_;
  assign new_n1464_ = ~i_40_ & new_n1463_;
  assign new_n1465_ = ~i_41_ & new_n1464_;
  assign new_n1466_ = ~i_43_ & new_n1465_;
  assign new_n1467_ = ~i_46_ & new_n1466_;
  assign new_n1468_ = ~i_47_ & new_n1467_;
  assign new_n1469_ = ~i_50_ & new_n1468_;
  assign new_n1470_ = ~i_56_ & new_n1469_;
  assign new_n1471_ = ~i_58_ & new_n1470_;
  assign new_n1472_ = ~i_60_ & new_n1471_;
  assign o_57_ = ~i_62_ & new_n1472_;
  assign new_n1474_ = i_22_ & new_n1453_;
  assign new_n1475_ = ~i_24_ & new_n1474_;
  assign new_n1476_ = ~i_25_ & new_n1475_;
  assign new_n1477_ = ~i_26_ & new_n1476_;
  assign new_n1478_ = ~i_28_ & new_n1477_;
  assign new_n1479_ = i_29_ & new_n1478_;
  assign new_n1480_ = ~i_30_ & new_n1479_;
  assign new_n1481_ = ~i_37_ & new_n1480_;
  assign new_n1482_ = ~i_39_ & new_n1481_;
  assign new_n1483_ = ~i_40_ & new_n1482_;
  assign new_n1484_ = ~i_41_ & new_n1483_;
  assign new_n1485_ = ~i_43_ & new_n1484_;
  assign new_n1486_ = ~i_46_ & new_n1485_;
  assign new_n1487_ = ~i_47_ & new_n1486_;
  assign new_n1488_ = ~i_50_ & new_n1487_;
  assign new_n1489_ = ~i_56_ & new_n1488_;
  assign new_n1490_ = ~i_58_ & new_n1489_;
  assign new_n1491_ = ~i_60_ & new_n1490_;
  assign o_58_ = ~i_62_ & new_n1491_;
  assign new_n1493_ = i_40_ & new_n450_;
  assign new_n1494_ = ~i_43_ & new_n1493_;
  assign new_n1495_ = ~i_50_ & new_n1494_;
  assign o_59_ = ~i_58_ & new_n1495_;
  assign new_n1497_ = i_7_ & ~i_8_;
  assign new_n1498_ = ~i_10_ & new_n1497_;
  assign new_n1499_ = ~i_11_ & new_n1498_;
  assign new_n1500_ = ~i_14_ & new_n1499_;
  assign new_n1501_ = ~i_15_ & new_n1500_;
  assign new_n1502_ = ~i_24_ & new_n1501_;
  assign new_n1503_ = ~i_25_ & new_n1502_;
  assign new_n1504_ = ~i_28_ & new_n1503_;
  assign new_n1505_ = i_29_ & new_n1504_;
  assign new_n1506_ = ~i_30_ & new_n1505_;
  assign new_n1507_ = ~i_37_ & new_n1506_;
  assign new_n1508_ = ~i_39_ & new_n1507_;
  assign new_n1509_ = ~i_40_ & new_n1508_;
  assign new_n1510_ = ~i_43_ & new_n1509_;
  assign new_n1511_ = ~i_46_ & new_n1510_;
  assign new_n1512_ = ~i_47_ & new_n1511_;
  assign new_n1513_ = ~i_50_ & new_n1512_;
  assign new_n1514_ = ~i_56_ & new_n1513_;
  assign new_n1515_ = ~i_58_ & new_n1514_;
  assign o_60_ = ~i_60_ & new_n1515_;
  assign new_n1517_ = i_8_ & ~i_10_;
  assign new_n1518_ = ~i_11_ & new_n1517_;
  assign new_n1519_ = ~i_14_ & new_n1518_;
  assign new_n1520_ = ~i_15_ & new_n1519_;
  assign new_n1521_ = ~i_24_ & new_n1520_;
  assign new_n1522_ = ~i_25_ & new_n1521_;
  assign new_n1523_ = ~i_28_ & new_n1522_;
  assign new_n1524_ = i_29_ & new_n1523_;
  assign new_n1525_ = ~i_30_ & new_n1524_;
  assign new_n1526_ = ~i_37_ & new_n1525_;
  assign new_n1527_ = ~i_39_ & new_n1526_;
  assign new_n1528_ = ~i_40_ & new_n1527_;
  assign new_n1529_ = ~i_43_ & new_n1528_;
  assign new_n1530_ = ~i_46_ & new_n1529_;
  assign new_n1531_ = ~i_47_ & new_n1530_;
  assign new_n1532_ = ~i_50_ & new_n1531_;
  assign new_n1533_ = ~i_56_ & new_n1532_;
  assign new_n1534_ = ~i_58_ & new_n1533_;
  assign o_61_ = ~i_60_ & new_n1534_;
  assign new_n1536_ = ~i_10_ & ~i_11_;
  assign new_n1537_ = ~i_14_ & new_n1536_;
  assign new_n1538_ = ~i_15_ & new_n1537_;
  assign new_n1539_ = ~i_24_ & new_n1538_;
  assign new_n1540_ = ~i_25_ & new_n1539_;
  assign new_n1541_ = ~i_28_ & new_n1540_;
  assign new_n1542_ = i_29_ & new_n1541_;
  assign new_n1543_ = ~i_30_ & new_n1542_;
  assign new_n1544_ = ~i_37_ & new_n1543_;
  assign new_n1545_ = ~i_39_ & new_n1544_;
  assign new_n1546_ = ~i_40_ & new_n1545_;
  assign new_n1547_ = ~i_43_ & new_n1546_;
  assign new_n1548_ = ~i_46_ & new_n1547_;
  assign new_n1549_ = i_47_ & new_n1548_;
  assign new_n1550_ = ~i_50_ & new_n1549_;
  assign new_n1551_ = ~i_56_ & new_n1550_;
  assign new_n1552_ = ~i_58_ & new_n1551_;
  assign o_62_ = ~i_60_ & new_n1552_;
  assign new_n1554_ = ~i_50_ & new_n1548_;
  assign new_n1555_ = i_56_ & new_n1554_;
  assign new_n1556_ = ~i_58_ & new_n1555_;
  assign o_63_ = ~i_60_ & new_n1556_;
  assign new_n1558_ = i_30_ & new_n1542_;
  assign new_n1559_ = ~i_37_ & new_n1558_;
  assign new_n1560_ = ~i_39_ & new_n1559_;
  assign new_n1561_ = ~i_40_ & new_n1560_;
  assign new_n1562_ = ~i_43_ & new_n1561_;
  assign new_n1563_ = ~i_46_ & new_n1562_;
  assign new_n1564_ = ~i_50_ & new_n1563_;
  assign new_n1565_ = ~i_58_ & new_n1564_;
  assign o_64_ = ~i_60_ & new_n1565_;
  assign o_5_ = i_29_;
endmodule


