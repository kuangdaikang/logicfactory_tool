// Benchmark "testing" written by ABC on Fri Feb 25 15:13:09 2022

module 25_13 ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A74  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A74;
  wire new_n27_, new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_,
    new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_;
  assign new_n27_ = A302 & A299;
  assign new_n28_ = ~A298 & new_n27_;
  assign new_n29_ = A203 & ~A200;
  assign new_n30_ = new_n28_ & new_n29_;
  assign new_n31_ = A199 & A166;
  assign new_n32_ = A167 & new_n31_;
  assign new_n33_ = ~A168 & ~A169;
  assign new_n34_ = new_n32_ & new_n33_;
  assign new_n35_ = new_n30_ & new_n34_;
  assign new_n36_ = A302 & ~A299;
  assign new_n37_ = A298 & new_n36_;
  assign new_n38_ = new_n29_ & new_n37_;
  assign new_n39_ = new_n34_ & new_n38_;
  assign new_n40_ = ~new_n35_ & ~new_n39_;
  assign new_n41_ = A203 & A200;
  assign new_n42_ = new_n28_ & new_n41_;
  assign new_n43_ = ~A199 & A166;
  assign new_n44_ = A167 & new_n43_;
  assign new_n45_ = new_n33_ & new_n44_;
  assign new_n46_ = new_n42_ & new_n45_;
  assign new_n47_ = new_n37_ & new_n41_;
  assign new_n48_ = new_n45_ & new_n47_;
  assign new_n49_ = ~new_n46_ & ~new_n48_;
  assign new_n50_ = new_n40_ & new_n49_;
  assign new_n51_ = ~A202 & ~A201;
  assign new_n52_ = new_n28_ & new_n51_;
  assign new_n53_ = A200 & A199;
  assign new_n54_ = ~A166 & new_n53_;
  assign new_n55_ = A167 & A170;
  assign new_n56_ = new_n54_ & new_n55_;
  assign new_n57_ = new_n52_ & new_n56_;
  assign new_n58_ = A166 & new_n53_;
  assign new_n59_ = ~A167 & A170;
  assign new_n60_ = new_n58_ & new_n59_;
  assign new_n61_ = new_n52_ & new_n60_;
  assign new_n62_ = new_n37_ & new_n51_;
  assign new_n63_ = new_n60_ & new_n62_;
  assign new_n64_ = ~new_n61_ & ~new_n63_;
  assign new_n65_ = ~new_n57_ & new_n64_;
  assign new_n66_ = new_n50_ & new_n65_;
  assign new_n67_ = A199 & ~A168;
  assign new_n68_ = ~A169 & ~A170;
  assign new_n69_ = new_n67_ & new_n68_;
  assign new_n70_ = new_n38_ & new_n69_;
  assign new_n71_ = new_n56_ & new_n62_;
  assign new_n72_ = new_n30_ & new_n69_;
  assign new_n73_ = ~new_n71_ & ~new_n72_;
  assign new_n74_ = ~new_n70_ & new_n73_;
  assign new_n75_ = A300 & A298;
  assign new_n76_ = A203 & new_n75_;
  assign new_n77_ = ~A200 & A199;
  assign new_n78_ = new_n76_ & new_n77_;
  assign new_n79_ = A166 & A167;
  assign new_n80_ = new_n33_ & new_n79_;
  assign new_n81_ = new_n78_ & new_n80_;
  assign new_n82_ = ~A199 & ~A168;
  assign new_n83_ = new_n68_ & new_n82_;
  assign new_n84_ = new_n42_ & new_n83_;
  assign new_n85_ = new_n47_ & new_n83_;
  assign new_n86_ = ~new_n84_ & ~new_n85_;
  assign new_n87_ = ~new_n81_ & new_n86_;
  assign new_n88_ = new_n74_ & new_n87_;
  assign new_n89_ = new_n66_ & new_n88_;
  assign new_n90_ = A300 & A299;
  assign new_n91_ = A203 & new_n90_;
  assign new_n92_ = new_n77_ & new_n91_;
  assign new_n93_ = new_n80_ & new_n92_;
  assign new_n94_ = A200 & ~A199;
  assign new_n95_ = new_n76_ & new_n94_;
  assign new_n96_ = new_n80_ & new_n95_;
  assign new_n97_ = ~new_n93_ & ~new_n96_;
  assign new_n98_ = new_n91_ & new_n94_;
  assign new_n99_ = new_n80_ & new_n98_;
  assign new_n100_ = A201 & A200;
  assign new_n101_ = new_n28_ & new_n100_;
  assign new_n102_ = new_n80_ & new_n101_;
  assign new_n103_ = ~new_n99_ & ~new_n102_;
  assign new_n104_ = new_n97_ & new_n103_;
  assign new_n105_ = A201 & A199;
  assign new_n106_ = new_n37_ & new_n105_;
  assign new_n107_ = new_n80_ & new_n106_;
  assign new_n108_ = new_n37_ & new_n100_;
  assign new_n109_ = new_n80_ & new_n108_;
  assign new_n110_ = new_n28_ & new_n105_;
  assign new_n111_ = new_n80_ & new_n110_;
  assign new_n112_ = ~new_n109_ & ~new_n111_;
  assign new_n113_ = ~new_n107_ & new_n112_;
  assign new_n114_ = new_n104_ & new_n113_;
  assign new_n115_ = ~A199 & ~A166;
  assign new_n116_ = ~A167 & ~A169;
  assign new_n117_ = new_n115_ & new_n116_;
  assign new_n118_ = new_n42_ & new_n117_;
  assign new_n119_ = A199 & ~A166;
  assign new_n120_ = new_n116_ & new_n119_;
  assign new_n121_ = new_n30_ & new_n120_;
  assign new_n122_ = new_n38_ & new_n120_;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = ~new_n118_ & new_n123_;
  assign new_n125_ = ~A202 & ~A200;
  assign new_n126_ = new_n37_ & new_n125_;
  assign new_n127_ = new_n43_ & new_n59_;
  assign new_n128_ = new_n126_ & new_n127_;
  assign new_n129_ = new_n47_ & new_n117_;
  assign new_n130_ = new_n28_ & new_n125_;
  assign new_n131_ = new_n127_ & new_n130_;
  assign new_n132_ = ~new_n129_ & ~new_n131_;
  assign new_n133_ = ~new_n128_ & new_n132_;
  assign new_n134_ = new_n124_ & new_n133_;
  assign new_n135_ = new_n114_ & new_n134_;
  assign new_n136_ = new_n89_ & new_n135_;
  assign new_n137_ = ~A202 & new_n75_;
  assign new_n138_ = ~A201 & A200;
  assign new_n139_ = new_n137_ & new_n138_;
  assign new_n140_ = new_n31_ & new_n59_;
  assign new_n141_ = new_n139_ & new_n140_;
  assign new_n142_ = ~A202 & new_n90_;
  assign new_n143_ = new_n138_ & new_n142_;
  assign new_n144_ = new_n140_ & new_n143_;
  assign new_n145_ = ~new_n141_ & ~new_n144_;
  assign new_n146_ = ~A203 & ~A202;
  assign new_n147_ = new_n28_ & new_n146_;
  assign new_n148_ = ~A201 & A166;
  assign new_n149_ = new_n59_ & new_n148_;
  assign new_n150_ = new_n147_ & new_n149_;
  assign new_n151_ = new_n37_ & new_n146_;
  assign new_n152_ = new_n149_ & new_n151_;
  assign new_n153_ = ~new_n150_ & ~new_n152_;
  assign new_n154_ = new_n145_ & new_n153_;
  assign new_n155_ = new_n55_ & new_n119_;
  assign new_n156_ = new_n139_ & new_n155_;
  assign new_n157_ = new_n55_ & new_n115_;
  assign new_n158_ = new_n130_ & new_n157_;
  assign new_n159_ = new_n126_ & new_n157_;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_ = ~new_n156_ & new_n160_;
  assign new_n162_ = new_n154_ & new_n161_;
  assign new_n163_ = ~A201 & ~A166;
  assign new_n164_ = new_n55_ & new_n163_;
  assign new_n165_ = new_n151_ & new_n164_;
  assign new_n166_ = new_n143_ & new_n155_;
  assign new_n167_ = new_n147_ & new_n164_;
  assign new_n168_ = ~new_n166_ & ~new_n167_;
  assign new_n169_ = ~new_n165_ & new_n168_;
  assign new_n170_ = A166 & A168;
  assign new_n171_ = new_n53_ & new_n170_;
  assign new_n172_ = new_n52_ & new_n171_;
  assign new_n173_ = A167 & A168;
  assign new_n174_ = new_n53_ & new_n173_;
  assign new_n175_ = new_n52_ & new_n174_;
  assign new_n176_ = new_n62_ & new_n174_;
  assign new_n177_ = ~new_n175_ & ~new_n176_;
  assign new_n178_ = ~new_n172_ & new_n177_;
  assign new_n179_ = new_n169_ & new_n178_;
  assign new_n180_ = new_n162_ & new_n179_;
  assign new_n181_ = new_n62_ & new_n171_;
  assign new_n182_ = new_n29_ & new_n75_;
  assign new_n183_ = new_n69_ & new_n182_;
  assign new_n184_ = ~new_n181_ & ~new_n183_;
  assign new_n185_ = new_n29_ & new_n90_;
  assign new_n186_ = new_n69_ & new_n185_;
  assign new_n187_ = new_n41_ & new_n75_;
  assign new_n188_ = new_n83_ & new_n187_;
  assign new_n189_ = ~new_n186_ & ~new_n188_;
  assign new_n190_ = new_n184_ & new_n189_;
  assign new_n191_ = A298 & A201;
  assign new_n192_ = new_n36_ & new_n191_;
  assign new_n193_ = A200 & ~A168;
  assign new_n194_ = new_n68_ & new_n193_;
  assign new_n195_ = new_n192_ & new_n194_;
  assign new_n196_ = new_n41_ & new_n90_;
  assign new_n197_ = new_n83_ & new_n196_;
  assign new_n198_ = ~A298 & A201;
  assign new_n199_ = new_n27_ & new_n198_;
  assign new_n200_ = new_n194_ & new_n199_;
  assign new_n201_ = ~new_n197_ & ~new_n200_;
  assign new_n202_ = ~new_n195_ & new_n201_;
  assign new_n203_ = new_n190_ & new_n202_;
  assign new_n204_ = A301 & A203;
  assign new_n205_ = new_n77_ & new_n204_;
  assign new_n206_ = new_n80_ & new_n205_;
  assign new_n207_ = new_n69_ & new_n199_;
  assign new_n208_ = new_n69_ & new_n192_;
  assign new_n209_ = ~new_n207_ & ~new_n208_;
  assign new_n210_ = ~new_n206_ & new_n209_;
  assign new_n211_ = new_n90_ & new_n100_;
  assign new_n212_ = new_n80_ & new_n211_;
  assign new_n213_ = new_n94_ & new_n204_;
  assign new_n214_ = new_n80_ & new_n213_;
  assign new_n215_ = new_n75_ & new_n100_;
  assign new_n216_ = new_n80_ & new_n215_;
  assign new_n217_ = ~new_n214_ & ~new_n216_;
  assign new_n218_ = ~new_n212_ & new_n217_;
  assign new_n219_ = new_n210_ & new_n218_;
  assign new_n220_ = new_n203_ & new_n219_;
  assign new_n221_ = new_n180_ & new_n220_;
  assign new_n222_ = new_n136_ & new_n221_;
  assign new_n223_ = new_n75_ & new_n105_;
  assign new_n224_ = new_n80_ & new_n223_;
  assign new_n225_ = new_n90_ & new_n105_;
  assign new_n226_ = new_n80_ & new_n225_;
  assign new_n227_ = ~new_n224_ & ~new_n226_;
  assign new_n228_ = ~A298 & A202;
  assign new_n229_ = new_n27_ & new_n228_;
  assign new_n230_ = new_n80_ & new_n229_;
  assign new_n231_ = A298 & A202;
  assign new_n232_ = new_n36_ & new_n231_;
  assign new_n233_ = new_n80_ & new_n232_;
  assign new_n234_ = ~new_n230_ & ~new_n233_;
  assign new_n235_ = new_n227_ & new_n234_;
  assign new_n236_ = new_n117_ & new_n187_;
  assign new_n237_ = new_n120_ & new_n182_;
  assign new_n238_ = new_n120_ & new_n185_;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign new_n240_ = ~new_n236_ & new_n239_;
  assign new_n241_ = new_n235_ & new_n240_;
  assign new_n242_ = A200 & ~A166;
  assign new_n243_ = new_n116_ & new_n242_;
  assign new_n244_ = new_n192_ & new_n243_;
  assign new_n245_ = new_n117_ & new_n196_;
  assign new_n246_ = new_n199_ & new_n243_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = ~new_n244_ & new_n247_;
  assign new_n249_ = ~A298 & ~A202;
  assign new_n250_ = new_n27_ & new_n249_;
  assign new_n251_ = A199 & A169;
  assign new_n252_ = new_n138_ & new_n251_;
  assign new_n253_ = new_n250_ & new_n252_;
  assign new_n254_ = new_n120_ & new_n199_;
  assign new_n255_ = new_n120_ & new_n192_;
  assign new_n256_ = ~new_n254_ & ~new_n255_;
  assign new_n257_ = ~new_n253_ & new_n256_;
  assign new_n258_ = new_n248_ & new_n257_;
  assign new_n259_ = new_n241_ & new_n258_;
  assign new_n260_ = A298 & ~A202;
  assign new_n261_ = new_n36_ & new_n260_;
  assign new_n262_ = new_n252_ & new_n261_;
  assign new_n263_ = new_n75_ & new_n125_;
  assign new_n264_ = new_n127_ & new_n263_;
  assign new_n265_ = ~new_n262_ & ~new_n264_;
  assign new_n266_ = new_n90_ & new_n125_;
  assign new_n267_ = new_n127_ & new_n266_;
  assign new_n268_ = A301 & ~A202;
  assign new_n269_ = new_n138_ & new_n268_;
  assign new_n270_ = new_n140_ & new_n269_;
  assign new_n271_ = ~new_n267_ & ~new_n270_;
  assign new_n272_ = new_n265_ & new_n271_;
  assign new_n273_ = new_n157_ & new_n263_;
  assign new_n274_ = new_n75_ & new_n146_;
  assign new_n275_ = new_n149_ & new_n274_;
  assign new_n276_ = new_n90_ & new_n146_;
  assign new_n277_ = new_n149_ & new_n276_;
  assign new_n278_ = ~new_n275_ & ~new_n277_;
  assign new_n279_ = ~new_n273_ & new_n278_;
  assign new_n280_ = new_n272_ & new_n279_;
  assign new_n281_ = new_n164_ & new_n274_;
  assign new_n282_ = new_n157_ & new_n266_;
  assign new_n283_ = new_n155_ & new_n269_;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = ~new_n281_ & new_n284_;
  assign new_n286_ = ~A200 & ~A199;
  assign new_n287_ = new_n173_ & new_n286_;
  assign new_n288_ = new_n261_ & new_n287_;
  assign new_n289_ = new_n164_ & new_n276_;
  assign new_n290_ = new_n250_ & new_n287_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = ~new_n288_ & new_n291_;
  assign new_n293_ = new_n285_ & new_n292_;
  assign new_n294_ = new_n280_ & new_n293_;
  assign new_n295_ = new_n259_ & new_n294_;
  assign new_n296_ = new_n51_ & new_n75_;
  assign new_n297_ = new_n174_ & new_n296_;
  assign new_n298_ = new_n51_ & new_n90_;
  assign new_n299_ = new_n174_ & new_n298_;
  assign new_n300_ = ~new_n297_ & ~new_n299_;
  assign new_n301_ = ~A298 & ~A203;
  assign new_n302_ = new_n27_ & new_n301_;
  assign new_n303_ = new_n51_ & new_n173_;
  assign new_n304_ = new_n302_ & new_n303_;
  assign new_n305_ = A298 & ~A203;
  assign new_n306_ = new_n36_ & new_n305_;
  assign new_n307_ = new_n303_ & new_n306_;
  assign new_n308_ = ~new_n304_ & ~new_n307_;
  assign new_n309_ = new_n300_ & new_n308_;
  assign new_n310_ = new_n171_ & new_n296_;
  assign new_n311_ = new_n170_ & new_n286_;
  assign new_n312_ = new_n250_ & new_n311_;
  assign new_n313_ = new_n261_ & new_n311_;
  assign new_n314_ = ~new_n312_ & ~new_n313_;
  assign new_n315_ = ~new_n310_ & new_n314_;
  assign new_n316_ = new_n309_ & new_n315_;
  assign new_n317_ = new_n51_ & new_n170_;
  assign new_n318_ = new_n306_ & new_n317_;
  assign new_n319_ = new_n171_ & new_n298_;
  assign new_n320_ = new_n302_ & new_n317_;
  assign new_n321_ = ~new_n319_ & ~new_n320_;
  assign new_n322_ = ~new_n318_ & new_n321_;
  assign new_n323_ = ~A170 & new_n33_;
  assign new_n324_ = new_n215_ & new_n323_;
  assign new_n325_ = new_n205_ & new_n323_;
  assign new_n326_ = new_n213_ & new_n323_;
  assign new_n327_ = ~new_n325_ & ~new_n326_;
  assign new_n328_ = ~new_n324_ & new_n327_;
  assign new_n329_ = new_n322_ & new_n328_;
  assign new_n330_ = new_n316_ & new_n329_;
  assign new_n331_ = new_n225_ & new_n323_;
  assign new_n332_ = new_n211_ & new_n323_;
  assign new_n333_ = new_n223_ & new_n323_;
  assign new_n334_ = ~new_n332_ & ~new_n333_;
  assign new_n335_ = ~new_n331_ & new_n334_;
  assign new_n336_ = A301 & A201;
  assign new_n337_ = A200 & A166;
  assign new_n338_ = new_n336_ & new_n337_;
  assign new_n339_ = A167 & ~A168;
  assign new_n340_ = ~A169 & new_n339_;
  assign new_n341_ = new_n338_ & new_n340_;
  assign new_n342_ = new_n229_ & new_n323_;
  assign new_n343_ = new_n232_ & new_n323_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign new_n345_ = ~new_n341_ & new_n344_;
  assign new_n346_ = new_n335_ & new_n345_;
  assign new_n347_ = A202 & A166;
  assign new_n348_ = new_n90_ & new_n347_;
  assign new_n349_ = new_n340_ & new_n348_;
  assign new_n350_ = new_n31_ & new_n336_;
  assign new_n351_ = new_n340_ & new_n350_;
  assign new_n352_ = new_n75_ & new_n347_;
  assign new_n353_ = new_n340_ & new_n352_;
  assign new_n354_ = ~new_n351_ & ~new_n353_;
  assign new_n355_ = ~new_n349_ & new_n354_;
  assign new_n356_ = ~A166 & ~A167;
  assign new_n357_ = ~A169 & new_n356_;
  assign new_n358_ = new_n215_ & new_n357_;
  assign new_n359_ = new_n205_ & new_n357_;
  assign new_n360_ = new_n213_ & new_n357_;
  assign new_n361_ = ~new_n359_ & ~new_n360_;
  assign new_n362_ = ~new_n358_ & new_n361_;
  assign new_n363_ = new_n355_ & new_n362_;
  assign new_n364_ = new_n346_ & new_n363_;
  assign new_n365_ = new_n330_ & new_n364_;
  assign new_n366_ = new_n295_ & new_n365_;
  assign new_n367_ = new_n222_ & new_n366_;
  assign new_n368_ = new_n211_ & new_n357_;
  assign new_n369_ = new_n223_ & new_n357_;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = new_n225_ & new_n357_;
  assign new_n372_ = new_n229_ & new_n357_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = new_n370_ & new_n373_;
  assign new_n375_ = A169 & new_n286_;
  assign new_n376_ = new_n261_ & new_n375_;
  assign new_n377_ = new_n232_ & new_n357_;
  assign new_n378_ = new_n250_ & new_n375_;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_ = ~new_n376_ & new_n379_;
  assign new_n381_ = new_n374_ & new_n380_;
  assign new_n382_ = A169 & new_n51_;
  assign new_n383_ = new_n302_ & new_n382_;
  assign new_n384_ = A169 & new_n53_;
  assign new_n385_ = new_n296_ & new_n384_;
  assign new_n386_ = new_n298_ & new_n384_;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign new_n388_ = ~new_n383_ & new_n387_;
  assign new_n389_ = A301 & ~A203;
  assign new_n390_ = new_n51_ & new_n389_;
  assign new_n391_ = A166 & ~A167;
  assign new_n392_ = A170 & new_n391_;
  assign new_n393_ = new_n390_ & new_n392_;
  assign new_n394_ = new_n306_ & new_n382_;
  assign new_n395_ = new_n268_ & new_n286_;
  assign new_n396_ = new_n392_ & new_n395_;
  assign new_n397_ = ~new_n394_ & ~new_n396_;
  assign new_n398_ = ~new_n393_ & new_n397_;
  assign new_n399_ = new_n388_ & new_n398_;
  assign new_n400_ = new_n381_ & new_n399_;
  assign new_n401_ = ~A166 & A167;
  assign new_n402_ = A170 & new_n401_;
  assign new_n403_ = new_n395_ & new_n402_;
  assign new_n404_ = new_n390_ & new_n402_;
  assign new_n405_ = ~new_n403_ & ~new_n404_;
  assign new_n406_ = ~A199 & A167;
  assign new_n407_ = A168 & new_n406_;
  assign new_n408_ = new_n263_ & new_n407_;
  assign new_n409_ = new_n266_ & new_n407_;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = new_n405_ & new_n410_;
  assign new_n412_ = ~A201 & A167;
  assign new_n413_ = A168 & new_n412_;
  assign new_n414_ = new_n276_ & new_n413_;
  assign new_n415_ = A199 & A167;
  assign new_n416_ = A168 & new_n415_;
  assign new_n417_ = new_n269_ & new_n416_;
  assign new_n418_ = new_n274_ & new_n413_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = ~new_n414_ & new_n419_;
  assign new_n421_ = new_n411_ & new_n420_;
  assign new_n422_ = A168 & new_n31_;
  assign new_n423_ = new_n269_ & new_n422_;
  assign new_n424_ = A168 & new_n43_;
  assign new_n425_ = new_n263_ & new_n424_;
  assign new_n426_ = new_n266_ & new_n424_;
  assign new_n427_ = ~new_n425_ & ~new_n426_;
  assign new_n428_ = ~new_n423_ & new_n427_;
  assign new_n429_ = A200 & new_n336_;
  assign new_n430_ = new_n323_ & new_n429_;
  assign new_n431_ = A168 & new_n148_;
  assign new_n432_ = new_n274_ & new_n431_;
  assign new_n433_ = new_n276_ & new_n431_;
  assign new_n434_ = ~new_n432_ & ~new_n433_;
  assign new_n435_ = ~new_n430_ & new_n434_;
  assign new_n436_ = new_n428_ & new_n435_;
  assign new_n437_ = new_n421_ & new_n436_;
  assign new_n438_ = new_n400_ & new_n437_;
  assign new_n439_ = A199 & new_n336_;
  assign new_n440_ = new_n323_ & new_n439_;
  assign new_n441_ = A202 & new_n75_;
  assign new_n442_ = new_n323_ & new_n441_;
  assign new_n443_ = ~new_n440_ & ~new_n442_;
  assign new_n444_ = A202 & new_n90_;
  assign new_n445_ = new_n323_ & new_n444_;
  assign new_n446_ = A301 & A202;
  assign new_n447_ = A166 & new_n446_;
  assign new_n448_ = new_n340_ & new_n447_;
  assign new_n449_ = ~new_n445_ & ~new_n448_;
  assign new_n450_ = new_n443_ & new_n449_;
  assign new_n451_ = new_n357_ & new_n441_;
  assign new_n452_ = new_n357_ & new_n429_;
  assign new_n453_ = new_n357_ & new_n439_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~new_n451_ & new_n454_;
  assign new_n456_ = new_n450_ & new_n455_;
  assign new_n457_ = new_n142_ & new_n375_;
  assign new_n458_ = new_n357_ & new_n444_;
  assign new_n459_ = new_n137_ & new_n375_;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~new_n457_ & new_n460_;
  assign new_n462_ = ~A203 & new_n90_;
  assign new_n463_ = new_n382_ & new_n462_;
  assign new_n464_ = ~A201 & new_n268_;
  assign new_n465_ = new_n384_ & new_n464_;
  assign new_n466_ = ~A203 & new_n75_;
  assign new_n467_ = new_n382_ & new_n466_;
  assign new_n468_ = ~new_n465_ & ~new_n467_;
  assign new_n469_ = ~new_n463_ & new_n468_;
  assign new_n470_ = new_n461_ & new_n469_;
  assign new_n471_ = new_n456_ & new_n470_;
  assign new_n472_ = A236 & ~A233;
  assign new_n473_ = A232 & new_n472_;
  assign new_n474_ = new_n402_ & new_n473_;
  assign new_n475_ = new_n392_ & new_n473_;
  assign new_n476_ = A236 & A233;
  assign new_n477_ = ~A232 & new_n476_;
  assign new_n478_ = new_n392_ & new_n477_;
  assign new_n479_ = ~new_n475_ & ~new_n478_;
  assign new_n480_ = ~new_n474_ & new_n479_;
  assign new_n481_ = ~A202 & new_n389_;
  assign new_n482_ = new_n413_ & new_n481_;
  assign new_n483_ = new_n402_ & new_n477_;
  assign new_n484_ = ~A200 & new_n268_;
  assign new_n485_ = new_n407_ & new_n484_;
  assign new_n486_ = ~new_n483_ & ~new_n485_;
  assign new_n487_ = ~new_n482_ & new_n486_;
  assign new_n488_ = new_n480_ & new_n487_;
  assign new_n489_ = A199 & new_n29_;
  assign new_n490_ = new_n473_ & new_n489_;
  assign new_n491_ = new_n424_ & new_n484_;
  assign new_n492_ = new_n431_ & new_n481_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = ~new_n490_ & new_n493_;
  assign new_n495_ = ~A199 & new_n41_;
  assign new_n496_ = new_n477_ & new_n495_;
  assign new_n497_ = new_n477_ & new_n489_;
  assign new_n498_ = new_n473_ & new_n495_;
  assign new_n499_ = ~new_n497_ & ~new_n498_;
  assign new_n500_ = ~new_n496_ & new_n499_;
  assign new_n501_ = new_n494_ & new_n500_;
  assign new_n502_ = new_n488_ & new_n501_;
  assign new_n503_ = new_n471_ & new_n502_;
  assign new_n504_ = new_n438_ & new_n503_;
  assign new_n505_ = ~A168 & new_n446_;
  assign new_n506_ = new_n68_ & new_n505_;
  assign new_n507_ = ~A166 & new_n446_;
  assign new_n508_ = new_n116_ & new_n507_;
  assign new_n509_ = ~new_n506_ & ~new_n508_;
  assign new_n510_ = ~A199 & A169;
  assign new_n511_ = new_n484_ & new_n510_;
  assign new_n512_ = ~A201 & A169;
  assign new_n513_ = new_n481_ & new_n512_;
  assign new_n514_ = ~new_n511_ & ~new_n513_;
  assign new_n515_ = new_n509_ & new_n514_;
  assign new_n516_ = A234 & A233;
  assign new_n517_ = ~A166 & new_n516_;
  assign new_n518_ = new_n55_ & new_n517_;
  assign new_n519_ = A166 & new_n516_;
  assign new_n520_ = new_n59_ & new_n519_;
  assign new_n521_ = A234 & A232;
  assign new_n522_ = A166 & new_n521_;
  assign new_n523_ = new_n59_ & new_n522_;
  assign new_n524_ = ~new_n520_ & ~new_n523_;
  assign new_n525_ = ~new_n518_ & new_n524_;
  assign new_n526_ = new_n515_ & new_n525_;
  assign new_n527_ = new_n173_ & new_n477_;
  assign new_n528_ = ~A166 & new_n521_;
  assign new_n529_ = new_n55_ & new_n528_;
  assign new_n530_ = new_n173_ & new_n473_;
  assign new_n531_ = ~new_n529_ & ~new_n530_;
  assign new_n532_ = ~new_n527_ & new_n531_;
  assign new_n533_ = A203 & new_n516_;
  assign new_n534_ = new_n77_ & new_n533_;
  assign new_n535_ = new_n170_ & new_n473_;
  assign new_n536_ = new_n170_ & new_n477_;
  assign new_n537_ = ~new_n535_ & ~new_n536_;
  assign new_n538_ = ~new_n534_ & new_n537_;
  assign new_n539_ = new_n532_ & new_n538_;
  assign new_n540_ = new_n526_ & new_n539_;
  assign new_n541_ = A203 & new_n521_;
  assign new_n542_ = new_n77_ & new_n541_;
  assign new_n543_ = new_n94_ & new_n533_;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = new_n94_ & new_n541_;
  assign new_n546_ = new_n100_ & new_n473_;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = new_n544_ & new_n547_;
  assign new_n549_ = new_n105_ & new_n477_;
  assign new_n550_ = new_n100_ & new_n477_;
  assign new_n551_ = new_n105_ & new_n473_;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = ~new_n549_ & new_n552_;
  assign new_n554_ = new_n548_ & new_n553_;
  assign new_n555_ = A235 & A166;
  assign new_n556_ = new_n59_ & new_n555_;
  assign new_n557_ = A232 & A169;
  assign new_n558_ = new_n472_ & new_n557_;
  assign new_n559_ = ~A232 & A169;
  assign new_n560_ = new_n476_ & new_n559_;
  assign new_n561_ = ~new_n558_ & ~new_n560_;
  assign new_n562_ = ~new_n556_ & new_n561_;
  assign new_n563_ = new_n173_ & new_n521_;
  assign new_n564_ = A235 & ~A166;
  assign new_n565_ = new_n55_ & new_n564_;
  assign new_n566_ = new_n173_ & new_n516_;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = ~new_n563_ & new_n567_;
  assign new_n569_ = new_n562_ & new_n568_;
  assign new_n570_ = new_n554_ & new_n569_;
  assign new_n571_ = new_n540_ & new_n570_;
  assign new_n572_ = new_n170_ & new_n516_;
  assign new_n573_ = new_n170_ & new_n521_;
  assign new_n574_ = ~new_n572_ & ~new_n573_;
  assign new_n575_ = A235 & A203;
  assign new_n576_ = new_n77_ & new_n575_;
  assign new_n577_ = new_n94_ & new_n575_;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = new_n574_ & new_n578_;
  assign new_n580_ = new_n105_ & new_n516_;
  assign new_n581_ = new_n100_ & new_n516_;
  assign new_n582_ = new_n100_ & new_n521_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = ~new_n580_ & new_n583_;
  assign new_n585_ = new_n579_ & new_n584_;
  assign new_n586_ = ~A232 & A202;
  assign new_n587_ = new_n476_ & new_n586_;
  assign new_n588_ = new_n105_ & new_n521_;
  assign new_n589_ = A232 & A202;
  assign new_n590_ = new_n472_ & new_n589_;
  assign new_n591_ = ~new_n588_ & ~new_n590_;
  assign new_n592_ = ~new_n587_ & new_n591_;
  assign new_n593_ = A235 & A167;
  assign new_n594_ = A168 & new_n593_;
  assign new_n595_ = A169 & new_n516_;
  assign new_n596_ = A169 & new_n521_;
  assign new_n597_ = ~new_n595_ & ~new_n596_;
  assign new_n598_ = ~new_n594_ & new_n597_;
  assign new_n599_ = new_n592_ & new_n598_;
  assign new_n600_ = new_n585_ & new_n599_;
  assign new_n601_ = A235 & A201;
  assign new_n602_ = A199 & new_n601_;
  assign new_n603_ = A168 & new_n555_;
  assign new_n604_ = A200 & new_n601_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n602_ & new_n605_;
  assign new_n607_ = A269 & ~A266;
  assign new_n608_ = A265 & new_n607_;
  assign new_n609_ = A202 & new_n516_;
  assign new_n610_ = A202 & new_n521_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = ~new_n608_ & new_n611_;
  assign new_n613_ = new_n606_ & new_n612_;
  assign new_n614_ = A235 & A202;
  assign new_n615_ = A269 & A266;
  assign new_n616_ = ~A265 & new_n615_;
  assign new_n617_ = A235 & A169;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = ~new_n614_ & new_n618_;
  assign new_n620_ = A267 & A266;
  assign new_n621_ = A267 & A265;
  assign new_n622_ = ~new_n620_ & ~new_n621_;
  assign new_n623_ = ~A268 & new_n622_;
  assign new_n624_ = new_n619_ & new_n623_;
  assign new_n625_ = new_n613_ & new_n624_;
  assign new_n626_ = new_n600_ & new_n625_;
  assign new_n627_ = new_n571_ & new_n626_;
  assign new_n628_ = new_n504_ & new_n627_;
  assign A74 = ~new_n367_ | ~new_n628_;
endmodule


