// Benchmark "adder" written by ABC on Tue Sep  5 17:43:40 2023

module adder ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387_, new_n388_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n410_, new_n411_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_,
    new_n552_, new_n553_, new_n554_, new_n555_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_,
    new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1309_,
    new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_,
    new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_,
    new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1457_, new_n1458_, new_n1459_,
    new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_,
    new_n1466_, new_n1467_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1753_,
    new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1901_, new_n1902_, new_n1903_,
    new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_,
    new_n1910_, new_n1911_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1937_, new_n1938_, new_n1939_;
  XOR2_X1    g0000(.A1(\a[0] ), .A2(\b[0] ), .Z(\f[0] ));
  NAND2_X1   g0001(.A1(\a[0] ), .A2(\b[0] ), .ZN(new_n387_));
  XNOR2_X1   g0002(.A1(new_n387_), .A2(\b[1] ), .ZN(new_n388_));
  XOR2_X1    g0003(.A1(new_n388_), .A2(\a[1] ), .Z(\f[1] ));
  NAND2_X1   g0004(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n390_));
  NOR2_X1    g0005(.A1(\a[1] ), .A2(\b[1] ), .ZN(new_n391_));
  OAI21_X1   g0006(.A1(new_n387_), .A2(new_n391_), .B(new_n390_), .ZN(new_n392_));
  INV_X1     g0007(.I(\b[2] ), .ZN(new_n393_));
  NOR2_X1    g0008(.A1(new_n393_), .A2(\a[2] ), .ZN(new_n394_));
  INV_X1     g0009(.I(\a[2] ), .ZN(new_n395_));
  NOR2_X1    g0010(.A1(new_n395_), .A2(\b[2] ), .ZN(new_n396_));
  OAI21_X1   g0011(.A1(new_n394_), .A2(new_n396_), .B(new_n392_), .ZN(new_n397_));
  NAND2_X1   g0012(.A1(\a[2] ), .A2(\b[2] ), .ZN(new_n398_));
  INV_X1     g0013(.I(new_n398_), .ZN(new_n399_));
  NOR2_X1    g0014(.A1(\a[2] ), .A2(\b[2] ), .ZN(new_n400_));
  NOR2_X1    g0015(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1   g0016(.A1(new_n392_), .A2(new_n401_), .B(new_n397_), .ZN(\f[2] ));
  AOI21_X1   g0017(.A1(new_n392_), .A2(new_n398_), .B(new_n400_), .ZN(new_n403_));
  XNOR2_X1   g0018(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n404_));
  NAND2_X1   g0019(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n405_));
  INV_X1     g0020(.I(new_n405_), .ZN(new_n406_));
  NOR2_X1    g0021(.A1(\a[3] ), .A2(\b[3] ), .ZN(new_n407_));
  OAI21_X1   g0022(.A1(new_n406_), .A2(new_n407_), .B(new_n403_), .ZN(new_n408_));
  OAI21_X1   g0023(.A1(new_n403_), .A2(new_n404_), .B(new_n408_), .ZN(\f[3] ));
  INV_X1     g0024(.I(\a[4] ), .ZN(new_n410_));
  INV_X1     g0025(.I(\b[4] ), .ZN(new_n411_));
  NOR4_X1    g0026(.A1(\a[2] ), .A2(\a[3] ), .A3(\b[2] ), .A4(\b[3] ), .ZN(new_n413_));
  OAI21_X1   g0027(.A1(new_n406_), .A2(new_n413_), .B(new_n411_), .ZN(new_n414_));
  INV_X1     g0028(.I(new_n414_), .ZN(new_n415_));
  NOR3_X1    g0029(.A1(new_n406_), .A2(new_n413_), .A3(new_n411_), .ZN(new_n416_));
  OAI21_X1   g0030(.A1(new_n415_), .A2(new_n416_), .B(new_n410_), .ZN(new_n417_));
  INV_X1     g0031(.I(new_n416_), .ZN(new_n418_));
  NAND3_X1   g0032(.A1(new_n418_), .A2(\a[4] ), .A3(new_n414_), .ZN(new_n419_));
  NAND2_X1   g0033(.A1(new_n417_), .A2(new_n419_), .ZN(\f[4] ));
  NOR2_X1    g0034(.A1(\a[4] ), .A2(\b[4] ), .ZN(new_n421_));
  AND2_X2    g0035(.A1(\a[4] ), .A2(\b[4] ), .Z(new_n422_));
  NOR3_X1    g0036(.A1(new_n406_), .A2(new_n422_), .A3(new_n413_), .ZN(new_n423_));
  NOR2_X1    g0037(.A1(new_n423_), .A2(new_n421_), .ZN(new_n424_));
  XOR2_X1    g0038(.A1(\a[5] ), .A2(\b[5] ), .Z(new_n425_));
  NAND2_X1   g0039(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1     g0040(.I(\a[5] ), .ZN(new_n427_));
  INV_X1     g0041(.I(\b[5] ), .ZN(new_n428_));
  NOR2_X1    g0042(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1    g0043(.A1(\a[5] ), .A2(\b[5] ), .ZN(new_n430_));
  NOR2_X1    g0044(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1   g0045(.A1(new_n424_), .A2(new_n431_), .B(new_n426_), .ZN(\f[5] ));
  NOR3_X1    g0046(.A1(new_n423_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n433_));
  XOR2_X1    g0047(.A1(\a[6] ), .A2(\b[6] ), .Z(new_n434_));
  OAI21_X1   g0048(.A1(new_n433_), .A2(new_n430_), .B(new_n434_), .ZN(new_n435_));
  INV_X1     g0049(.I(new_n430_), .ZN(new_n436_));
  INV_X1     g0050(.I(new_n421_), .ZN(new_n437_));
  OR4_X2     g0051(.A1(\a[2] ), .A2(\a[3] ), .A3(\b[2] ), .A4(\b[3] ), .Z(new_n438_));
  NAND2_X1   g0052(.A1(\a[4] ), .A2(\b[4] ), .ZN(new_n439_));
  NAND3_X1   g0053(.A1(new_n438_), .A2(new_n405_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1     g0054(.I(new_n429_), .ZN(new_n441_));
  NAND3_X1   g0055(.A1(new_n440_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1   g0056(.A1(\a[6] ), .A2(\b[6] ), .ZN(new_n443_));
  NAND3_X1   g0057(.A1(new_n442_), .A2(new_n436_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1   g0058(.A1(new_n444_), .A2(new_n435_), .ZN(\f[6] ));
  INV_X1     g0059(.I(\a[7] ), .ZN(new_n446_));
  INV_X1     g0060(.I(\b[7] ), .ZN(new_n447_));
  NAND2_X1   g0061(.A1(\a[6] ), .A2(\b[6] ), .ZN(new_n448_));
  INV_X1     g0062(.I(new_n448_), .ZN(new_n449_));
  NOR4_X1    g0063(.A1(\a[5] ), .A2(\a[6] ), .A3(\b[5] ), .A4(\b[6] ), .ZN(new_n450_));
  OAI21_X1   g0064(.A1(new_n449_), .A2(new_n450_), .B(new_n447_), .ZN(new_n451_));
  INV_X1     g0065(.I(new_n451_), .ZN(new_n452_));
  NOR3_X1    g0066(.A1(new_n449_), .A2(new_n450_), .A3(new_n447_), .ZN(new_n453_));
  OAI21_X1   g0067(.A1(new_n452_), .A2(new_n453_), .B(new_n446_), .ZN(new_n454_));
  INV_X1     g0068(.I(new_n453_), .ZN(new_n455_));
  NAND3_X1   g0069(.A1(new_n455_), .A2(\a[7] ), .A3(new_n451_), .ZN(new_n456_));
  NAND2_X1   g0070(.A1(new_n454_), .A2(new_n456_), .ZN(\f[7] ));
  NOR2_X1    g0071(.A1(\a[7] ), .A2(\b[7] ), .ZN(new_n458_));
  AND2_X2    g0072(.A1(\a[7] ), .A2(\b[7] ), .Z(new_n459_));
  NOR3_X1    g0073(.A1(new_n449_), .A2(new_n459_), .A3(new_n450_), .ZN(new_n460_));
  NOR2_X1    g0074(.A1(new_n460_), .A2(new_n458_), .ZN(new_n461_));
  XOR2_X1    g0075(.A1(\a[8] ), .A2(\b[8] ), .Z(new_n462_));
  NAND2_X1   g0076(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1     g0077(.I(\a[8] ), .ZN(new_n464_));
  INV_X1     g0078(.I(\b[8] ), .ZN(new_n465_));
  NOR2_X1    g0079(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1    g0080(.A1(\a[8] ), .A2(\b[8] ), .ZN(new_n467_));
  NOR2_X1    g0081(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1   g0082(.A1(new_n461_), .A2(new_n468_), .B(new_n463_), .ZN(\f[8] ));
  NOR3_X1    g0083(.A1(new_n460_), .A2(new_n458_), .A3(new_n466_), .ZN(new_n470_));
  XOR2_X1    g0084(.A1(\a[9] ), .A2(\b[9] ), .Z(new_n471_));
  OAI21_X1   g0085(.A1(new_n470_), .A2(new_n467_), .B(new_n471_), .ZN(new_n472_));
  INV_X1     g0086(.I(new_n467_), .ZN(new_n473_));
  INV_X1     g0087(.I(new_n458_), .ZN(new_n474_));
  OR4_X2     g0088(.A1(\a[5] ), .A2(\a[6] ), .A3(\b[5] ), .A4(\b[6] ), .Z(new_n475_));
  NAND2_X1   g0089(.A1(\a[7] ), .A2(\b[7] ), .ZN(new_n476_));
  NAND3_X1   g0090(.A1(new_n475_), .A2(new_n448_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1     g0091(.I(new_n466_), .ZN(new_n478_));
  NAND3_X1   g0092(.A1(new_n477_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1   g0093(.A1(\a[9] ), .A2(\b[9] ), .ZN(new_n480_));
  NAND3_X1   g0094(.A1(new_n479_), .A2(new_n473_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1   g0095(.A1(new_n481_), .A2(new_n472_), .ZN(\f[9] ));
  INV_X1     g0096(.I(\a[10] ), .ZN(new_n483_));
  INV_X1     g0097(.I(\b[10] ), .ZN(new_n484_));
  NAND2_X1   g0098(.A1(\a[9] ), .A2(\b[9] ), .ZN(new_n485_));
  INV_X1     g0099(.I(new_n485_), .ZN(new_n486_));
  NOR4_X1    g0100(.A1(\a[8] ), .A2(\a[9] ), .A3(\b[8] ), .A4(\b[9] ), .ZN(new_n487_));
  OAI21_X1   g0101(.A1(new_n486_), .A2(new_n487_), .B(new_n484_), .ZN(new_n488_));
  INV_X1     g0102(.I(new_n488_), .ZN(new_n489_));
  NOR3_X1    g0103(.A1(new_n486_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n490_));
  OAI21_X1   g0104(.A1(new_n489_), .A2(new_n490_), .B(new_n483_), .ZN(new_n491_));
  INV_X1     g0105(.I(new_n490_), .ZN(new_n492_));
  NAND3_X1   g0106(.A1(new_n492_), .A2(\a[10] ), .A3(new_n488_), .ZN(new_n493_));
  NAND2_X1   g0107(.A1(new_n491_), .A2(new_n493_), .ZN(\f[10] ));
  NOR2_X1    g0108(.A1(\a[10] ), .A2(\b[10] ), .ZN(new_n495_));
  AND2_X2    g0109(.A1(\a[10] ), .A2(\b[10] ), .Z(new_n496_));
  NOR3_X1    g0110(.A1(new_n486_), .A2(new_n496_), .A3(new_n487_), .ZN(new_n497_));
  NOR2_X1    g0111(.A1(new_n497_), .A2(new_n495_), .ZN(new_n498_));
  XOR2_X1    g0112(.A1(\a[11] ), .A2(\b[11] ), .Z(new_n499_));
  NAND2_X1   g0113(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1     g0114(.I(\a[11] ), .ZN(new_n501_));
  INV_X1     g0115(.I(\b[11] ), .ZN(new_n502_));
  NOR2_X1    g0116(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1    g0117(.A1(\a[11] ), .A2(\b[11] ), .ZN(new_n504_));
  NOR2_X1    g0118(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  OAI21_X1   g0119(.A1(new_n498_), .A2(new_n505_), .B(new_n500_), .ZN(\f[11] ));
  NOR3_X1    g0120(.A1(new_n497_), .A2(new_n495_), .A3(new_n503_), .ZN(new_n507_));
  XOR2_X1    g0121(.A1(\a[12] ), .A2(\b[12] ), .Z(new_n508_));
  OAI21_X1   g0122(.A1(new_n507_), .A2(new_n504_), .B(new_n508_), .ZN(new_n509_));
  INV_X1     g0123(.I(new_n504_), .ZN(new_n510_));
  INV_X1     g0124(.I(new_n495_), .ZN(new_n511_));
  OR4_X2     g0125(.A1(\a[8] ), .A2(\a[9] ), .A3(\b[8] ), .A4(\b[9] ), .Z(new_n512_));
  NAND2_X1   g0126(.A1(\a[10] ), .A2(\b[10] ), .ZN(new_n513_));
  NAND3_X1   g0127(.A1(new_n512_), .A2(new_n485_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1     g0128(.I(new_n503_), .ZN(new_n515_));
  NAND3_X1   g0129(.A1(new_n514_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1   g0130(.A1(\a[12] ), .A2(\b[12] ), .ZN(new_n517_));
  NAND3_X1   g0131(.A1(new_n516_), .A2(new_n510_), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1   g0132(.A1(new_n518_), .A2(new_n509_), .ZN(\f[12] ));
  INV_X1     g0133(.I(\a[13] ), .ZN(new_n520_));
  INV_X1     g0134(.I(\b[13] ), .ZN(new_n521_));
  NAND2_X1   g0135(.A1(\a[12] ), .A2(\b[12] ), .ZN(new_n522_));
  INV_X1     g0136(.I(new_n522_), .ZN(new_n523_));
  NOR4_X1    g0137(.A1(\a[11] ), .A2(\a[12] ), .A3(\b[11] ), .A4(\b[12] ), .ZN(new_n524_));
  OAI21_X1   g0138(.A1(new_n523_), .A2(new_n524_), .B(new_n521_), .ZN(new_n525_));
  INV_X1     g0139(.I(new_n525_), .ZN(new_n526_));
  NOR3_X1    g0140(.A1(new_n523_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n527_));
  OAI21_X1   g0141(.A1(new_n526_), .A2(new_n527_), .B(new_n520_), .ZN(new_n528_));
  INV_X1     g0142(.I(new_n527_), .ZN(new_n529_));
  NAND3_X1   g0143(.A1(new_n529_), .A2(\a[13] ), .A3(new_n525_), .ZN(new_n530_));
  NAND2_X1   g0144(.A1(new_n528_), .A2(new_n530_), .ZN(\f[13] ));
  NOR2_X1    g0145(.A1(\a[13] ), .A2(\b[13] ), .ZN(new_n532_));
  AND2_X2    g0146(.A1(\a[13] ), .A2(\b[13] ), .Z(new_n533_));
  NOR3_X1    g0147(.A1(new_n523_), .A2(new_n533_), .A3(new_n524_), .ZN(new_n534_));
  NOR2_X1    g0148(.A1(new_n534_), .A2(new_n532_), .ZN(new_n535_));
  XOR2_X1    g0149(.A1(\a[14] ), .A2(\b[14] ), .Z(new_n536_));
  NAND2_X1   g0150(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1     g0151(.I(\a[14] ), .ZN(new_n538_));
  INV_X1     g0152(.I(\b[14] ), .ZN(new_n539_));
  NOR2_X1    g0153(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1    g0154(.A1(\a[14] ), .A2(\b[14] ), .ZN(new_n541_));
  NOR2_X1    g0155(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1   g0156(.A1(new_n535_), .A2(new_n542_), .B(new_n537_), .ZN(\f[14] ));
  NOR3_X1    g0157(.A1(new_n534_), .A2(new_n532_), .A3(new_n540_), .ZN(new_n544_));
  XOR2_X1    g0158(.A1(\a[15] ), .A2(\b[15] ), .Z(new_n545_));
  OAI21_X1   g0159(.A1(new_n544_), .A2(new_n541_), .B(new_n545_), .ZN(new_n546_));
  INV_X1     g0160(.I(new_n541_), .ZN(new_n547_));
  INV_X1     g0161(.I(new_n532_), .ZN(new_n548_));
  OR4_X2     g0162(.A1(\a[11] ), .A2(\a[12] ), .A3(\b[11] ), .A4(\b[12] ), .Z(new_n549_));
  NAND2_X1   g0163(.A1(\a[13] ), .A2(\b[13] ), .ZN(new_n550_));
  NAND3_X1   g0164(.A1(new_n549_), .A2(new_n522_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1     g0165(.I(new_n540_), .ZN(new_n552_));
  NAND3_X1   g0166(.A1(new_n551_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1   g0167(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n554_));
  NAND3_X1   g0168(.A1(new_n553_), .A2(new_n547_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1   g0169(.A1(new_n555_), .A2(new_n546_), .ZN(\f[15] ));
  INV_X1     g0170(.I(\a[16] ), .ZN(new_n557_));
  INV_X1     g0171(.I(\b[16] ), .ZN(new_n558_));
  NAND2_X1   g0172(.A1(\a[15] ), .A2(\b[15] ), .ZN(new_n559_));
  INV_X1     g0173(.I(new_n559_), .ZN(new_n560_));
  NOR4_X1    g0174(.A1(\a[14] ), .A2(\a[15] ), .A3(\b[14] ), .A4(\b[15] ), .ZN(new_n561_));
  OAI21_X1   g0175(.A1(new_n560_), .A2(new_n561_), .B(new_n558_), .ZN(new_n562_));
  INV_X1     g0176(.I(new_n562_), .ZN(new_n563_));
  NOR3_X1    g0177(.A1(new_n560_), .A2(new_n561_), .A3(new_n558_), .ZN(new_n564_));
  OAI21_X1   g0178(.A1(new_n563_), .A2(new_n564_), .B(new_n557_), .ZN(new_n565_));
  INV_X1     g0179(.I(new_n564_), .ZN(new_n566_));
  NAND3_X1   g0180(.A1(new_n566_), .A2(\a[16] ), .A3(new_n562_), .ZN(new_n567_));
  NAND2_X1   g0181(.A1(new_n565_), .A2(new_n567_), .ZN(\f[16] ));
  NOR2_X1    g0182(.A1(\a[16] ), .A2(\b[16] ), .ZN(new_n569_));
  AND2_X2    g0183(.A1(\a[16] ), .A2(\b[16] ), .Z(new_n570_));
  NOR3_X1    g0184(.A1(new_n560_), .A2(new_n570_), .A3(new_n561_), .ZN(new_n571_));
  NOR2_X1    g0185(.A1(new_n571_), .A2(new_n569_), .ZN(new_n572_));
  XOR2_X1    g0186(.A1(\a[17] ), .A2(\b[17] ), .Z(new_n573_));
  NAND2_X1   g0187(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1     g0188(.I(\a[17] ), .ZN(new_n575_));
  INV_X1     g0189(.I(\b[17] ), .ZN(new_n576_));
  NOR2_X1    g0190(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1    g0191(.A1(\a[17] ), .A2(\b[17] ), .ZN(new_n578_));
  NOR2_X1    g0192(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1   g0193(.A1(new_n572_), .A2(new_n579_), .B(new_n574_), .ZN(\f[17] ));
  NOR3_X1    g0194(.A1(new_n571_), .A2(new_n569_), .A3(new_n577_), .ZN(new_n581_));
  XOR2_X1    g0195(.A1(\a[18] ), .A2(\b[18] ), .Z(new_n582_));
  OAI21_X1   g0196(.A1(new_n581_), .A2(new_n578_), .B(new_n582_), .ZN(new_n583_));
  INV_X1     g0197(.I(new_n578_), .ZN(new_n584_));
  INV_X1     g0198(.I(new_n569_), .ZN(new_n585_));
  OR4_X2     g0199(.A1(\a[14] ), .A2(\a[15] ), .A3(\b[14] ), .A4(\b[15] ), .Z(new_n586_));
  NAND2_X1   g0200(.A1(\a[16] ), .A2(\b[16] ), .ZN(new_n587_));
  NAND3_X1   g0201(.A1(new_n586_), .A2(new_n559_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1     g0202(.I(new_n577_), .ZN(new_n589_));
  NAND3_X1   g0203(.A1(new_n588_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  XNOR2_X1   g0204(.A1(\a[18] ), .A2(\b[18] ), .ZN(new_n591_));
  NAND3_X1   g0205(.A1(new_n590_), .A2(new_n584_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1   g0206(.A1(new_n592_), .A2(new_n583_), .ZN(\f[18] ));
  INV_X1     g0207(.I(\a[19] ), .ZN(new_n594_));
  INV_X1     g0208(.I(\b[19] ), .ZN(new_n595_));
  NAND2_X1   g0209(.A1(\a[18] ), .A2(\b[18] ), .ZN(new_n596_));
  INV_X1     g0210(.I(new_n596_), .ZN(new_n597_));
  NOR4_X1    g0211(.A1(\a[17] ), .A2(\a[18] ), .A3(\b[17] ), .A4(\b[18] ), .ZN(new_n598_));
  OAI21_X1   g0212(.A1(new_n597_), .A2(new_n598_), .B(new_n595_), .ZN(new_n599_));
  INV_X1     g0213(.I(new_n599_), .ZN(new_n600_));
  NOR3_X1    g0214(.A1(new_n597_), .A2(new_n598_), .A3(new_n595_), .ZN(new_n601_));
  OAI21_X1   g0215(.A1(new_n600_), .A2(new_n601_), .B(new_n594_), .ZN(new_n602_));
  INV_X1     g0216(.I(new_n601_), .ZN(new_n603_));
  NAND3_X1   g0217(.A1(new_n603_), .A2(\a[19] ), .A3(new_n599_), .ZN(new_n604_));
  NAND2_X1   g0218(.A1(new_n602_), .A2(new_n604_), .ZN(\f[19] ));
  NOR2_X1    g0219(.A1(\a[19] ), .A2(\b[19] ), .ZN(new_n606_));
  AND2_X2    g0220(.A1(\a[19] ), .A2(\b[19] ), .Z(new_n607_));
  NOR3_X1    g0221(.A1(new_n597_), .A2(new_n607_), .A3(new_n598_), .ZN(new_n608_));
  NOR2_X1    g0222(.A1(new_n608_), .A2(new_n606_), .ZN(new_n609_));
  XOR2_X1    g0223(.A1(\a[20] ), .A2(\b[20] ), .Z(new_n610_));
  NAND2_X1   g0224(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1     g0225(.I(\a[20] ), .ZN(new_n612_));
  INV_X1     g0226(.I(\b[20] ), .ZN(new_n613_));
  NOR2_X1    g0227(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1    g0228(.A1(\a[20] ), .A2(\b[20] ), .ZN(new_n615_));
  NOR2_X1    g0229(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1   g0230(.A1(new_n609_), .A2(new_n616_), .B(new_n611_), .ZN(\f[20] ));
  NOR3_X1    g0231(.A1(new_n608_), .A2(new_n606_), .A3(new_n614_), .ZN(new_n618_));
  XOR2_X1    g0232(.A1(\a[21] ), .A2(\b[21] ), .Z(new_n619_));
  OAI21_X1   g0233(.A1(new_n618_), .A2(new_n615_), .B(new_n619_), .ZN(new_n620_));
  INV_X1     g0234(.I(new_n615_), .ZN(new_n621_));
  INV_X1     g0235(.I(new_n606_), .ZN(new_n622_));
  OR4_X2     g0236(.A1(\a[17] ), .A2(\a[18] ), .A3(\b[17] ), .A4(\b[18] ), .Z(new_n623_));
  NAND2_X1   g0237(.A1(\a[19] ), .A2(\b[19] ), .ZN(new_n624_));
  NAND3_X1   g0238(.A1(new_n623_), .A2(new_n596_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1     g0239(.I(new_n614_), .ZN(new_n626_));
  NAND3_X1   g0240(.A1(new_n625_), .A2(new_n622_), .A3(new_n626_), .ZN(new_n627_));
  XNOR2_X1   g0241(.A1(\a[21] ), .A2(\b[21] ), .ZN(new_n628_));
  NAND3_X1   g0242(.A1(new_n627_), .A2(new_n621_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1   g0243(.A1(new_n629_), .A2(new_n620_), .ZN(\f[21] ));
  INV_X1     g0244(.I(\a[22] ), .ZN(new_n631_));
  INV_X1     g0245(.I(\b[22] ), .ZN(new_n632_));
  NAND2_X1   g0246(.A1(\a[21] ), .A2(\b[21] ), .ZN(new_n633_));
  INV_X1     g0247(.I(new_n633_), .ZN(new_n634_));
  NOR4_X1    g0248(.A1(\a[20] ), .A2(\a[21] ), .A3(\b[20] ), .A4(\b[21] ), .ZN(new_n635_));
  OAI21_X1   g0249(.A1(new_n634_), .A2(new_n635_), .B(new_n632_), .ZN(new_n636_));
  INV_X1     g0250(.I(new_n636_), .ZN(new_n637_));
  NOR3_X1    g0251(.A1(new_n634_), .A2(new_n635_), .A3(new_n632_), .ZN(new_n638_));
  OAI21_X1   g0252(.A1(new_n637_), .A2(new_n638_), .B(new_n631_), .ZN(new_n639_));
  INV_X1     g0253(.I(new_n638_), .ZN(new_n640_));
  NAND3_X1   g0254(.A1(new_n640_), .A2(\a[22] ), .A3(new_n636_), .ZN(new_n641_));
  NAND2_X1   g0255(.A1(new_n639_), .A2(new_n641_), .ZN(\f[22] ));
  NOR2_X1    g0256(.A1(\a[22] ), .A2(\b[22] ), .ZN(new_n643_));
  AND2_X2    g0257(.A1(\a[22] ), .A2(\b[22] ), .Z(new_n644_));
  NOR3_X1    g0258(.A1(new_n634_), .A2(new_n644_), .A3(new_n635_), .ZN(new_n645_));
  NOR2_X1    g0259(.A1(new_n645_), .A2(new_n643_), .ZN(new_n646_));
  XOR2_X1    g0260(.A1(\a[23] ), .A2(\b[23] ), .Z(new_n647_));
  NAND2_X1   g0261(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1     g0262(.I(\a[23] ), .ZN(new_n649_));
  INV_X1     g0263(.I(\b[23] ), .ZN(new_n650_));
  NOR2_X1    g0264(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1    g0265(.A1(\a[23] ), .A2(\b[23] ), .ZN(new_n652_));
  NOR2_X1    g0266(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1   g0267(.A1(new_n646_), .A2(new_n653_), .B(new_n648_), .ZN(\f[23] ));
  NOR3_X1    g0268(.A1(new_n645_), .A2(new_n643_), .A3(new_n651_), .ZN(new_n655_));
  XOR2_X1    g0269(.A1(\a[24] ), .A2(\b[24] ), .Z(new_n656_));
  OAI21_X1   g0270(.A1(new_n655_), .A2(new_n652_), .B(new_n656_), .ZN(new_n657_));
  INV_X1     g0271(.I(new_n652_), .ZN(new_n658_));
  INV_X1     g0272(.I(new_n643_), .ZN(new_n659_));
  OR4_X2     g0273(.A1(\a[20] ), .A2(\a[21] ), .A3(\b[20] ), .A4(\b[21] ), .Z(new_n660_));
  NAND2_X1   g0274(.A1(\a[22] ), .A2(\b[22] ), .ZN(new_n661_));
  NAND3_X1   g0275(.A1(new_n660_), .A2(new_n633_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1     g0276(.I(new_n651_), .ZN(new_n663_));
  NAND3_X1   g0277(.A1(new_n662_), .A2(new_n659_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1   g0278(.A1(\a[24] ), .A2(\b[24] ), .ZN(new_n665_));
  NAND3_X1   g0279(.A1(new_n664_), .A2(new_n658_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1   g0280(.A1(new_n666_), .A2(new_n657_), .ZN(\f[24] ));
  INV_X1     g0281(.I(\a[25] ), .ZN(new_n668_));
  INV_X1     g0282(.I(\b[25] ), .ZN(new_n669_));
  NAND2_X1   g0283(.A1(\a[24] ), .A2(\b[24] ), .ZN(new_n670_));
  INV_X1     g0284(.I(new_n670_), .ZN(new_n671_));
  NOR4_X1    g0285(.A1(\a[23] ), .A2(\a[24] ), .A3(\b[23] ), .A4(\b[24] ), .ZN(new_n672_));
  OAI21_X1   g0286(.A1(new_n671_), .A2(new_n672_), .B(new_n669_), .ZN(new_n673_));
  INV_X1     g0287(.I(new_n673_), .ZN(new_n674_));
  NOR3_X1    g0288(.A1(new_n671_), .A2(new_n672_), .A3(new_n669_), .ZN(new_n675_));
  OAI21_X1   g0289(.A1(new_n674_), .A2(new_n675_), .B(new_n668_), .ZN(new_n676_));
  INV_X1     g0290(.I(new_n675_), .ZN(new_n677_));
  NAND3_X1   g0291(.A1(new_n677_), .A2(\a[25] ), .A3(new_n673_), .ZN(new_n678_));
  NAND2_X1   g0292(.A1(new_n676_), .A2(new_n678_), .ZN(\f[25] ));
  NOR2_X1    g0293(.A1(\a[25] ), .A2(\b[25] ), .ZN(new_n680_));
  AND2_X2    g0294(.A1(\a[25] ), .A2(\b[25] ), .Z(new_n681_));
  NOR3_X1    g0295(.A1(new_n671_), .A2(new_n681_), .A3(new_n672_), .ZN(new_n682_));
  NOR2_X1    g0296(.A1(new_n682_), .A2(new_n680_), .ZN(new_n683_));
  XOR2_X1    g0297(.A1(\a[26] ), .A2(\b[26] ), .Z(new_n684_));
  NAND2_X1   g0298(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1     g0299(.I(\a[26] ), .ZN(new_n686_));
  INV_X1     g0300(.I(\b[26] ), .ZN(new_n687_));
  NOR2_X1    g0301(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1    g0302(.A1(\a[26] ), .A2(\b[26] ), .ZN(new_n689_));
  NOR2_X1    g0303(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1   g0304(.A1(new_n683_), .A2(new_n690_), .B(new_n685_), .ZN(\f[26] ));
  NOR3_X1    g0305(.A1(new_n682_), .A2(new_n680_), .A3(new_n688_), .ZN(new_n692_));
  XOR2_X1    g0306(.A1(\a[27] ), .A2(\b[27] ), .Z(new_n693_));
  OAI21_X1   g0307(.A1(new_n692_), .A2(new_n689_), .B(new_n693_), .ZN(new_n694_));
  INV_X1     g0308(.I(new_n689_), .ZN(new_n695_));
  INV_X1     g0309(.I(new_n680_), .ZN(new_n696_));
  OR4_X2     g0310(.A1(\a[23] ), .A2(\a[24] ), .A3(\b[23] ), .A4(\b[24] ), .Z(new_n697_));
  NAND2_X1   g0311(.A1(\a[25] ), .A2(\b[25] ), .ZN(new_n698_));
  NAND3_X1   g0312(.A1(new_n697_), .A2(new_n670_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1     g0313(.I(new_n688_), .ZN(new_n700_));
  NAND3_X1   g0314(.A1(new_n699_), .A2(new_n696_), .A3(new_n700_), .ZN(new_n701_));
  XNOR2_X1   g0315(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n702_));
  NAND3_X1   g0316(.A1(new_n701_), .A2(new_n695_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1   g0317(.A1(new_n703_), .A2(new_n694_), .ZN(\f[27] ));
  INV_X1     g0318(.I(\a[28] ), .ZN(new_n705_));
  INV_X1     g0319(.I(\b[28] ), .ZN(new_n706_));
  NAND2_X1   g0320(.A1(\a[27] ), .A2(\b[27] ), .ZN(new_n707_));
  INV_X1     g0321(.I(new_n707_), .ZN(new_n708_));
  NOR4_X1    g0322(.A1(\a[26] ), .A2(\a[27] ), .A3(\b[26] ), .A4(\b[27] ), .ZN(new_n709_));
  OAI21_X1   g0323(.A1(new_n708_), .A2(new_n709_), .B(new_n706_), .ZN(new_n710_));
  INV_X1     g0324(.I(new_n710_), .ZN(new_n711_));
  NOR3_X1    g0325(.A1(new_n708_), .A2(new_n709_), .A3(new_n706_), .ZN(new_n712_));
  OAI21_X1   g0326(.A1(new_n711_), .A2(new_n712_), .B(new_n705_), .ZN(new_n713_));
  INV_X1     g0327(.I(new_n712_), .ZN(new_n714_));
  NAND3_X1   g0328(.A1(new_n714_), .A2(\a[28] ), .A3(new_n710_), .ZN(new_n715_));
  NAND2_X1   g0329(.A1(new_n713_), .A2(new_n715_), .ZN(\f[28] ));
  NOR2_X1    g0330(.A1(\a[28] ), .A2(\b[28] ), .ZN(new_n717_));
  AND2_X2    g0331(.A1(\a[28] ), .A2(\b[28] ), .Z(new_n718_));
  NOR3_X1    g0332(.A1(new_n708_), .A2(new_n718_), .A3(new_n709_), .ZN(new_n719_));
  NOR2_X1    g0333(.A1(new_n719_), .A2(new_n717_), .ZN(new_n720_));
  XOR2_X1    g0334(.A1(\a[29] ), .A2(\b[29] ), .Z(new_n721_));
  NAND2_X1   g0335(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1     g0336(.I(\a[29] ), .ZN(new_n723_));
  INV_X1     g0337(.I(\b[29] ), .ZN(new_n724_));
  NOR2_X1    g0338(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1    g0339(.A1(\a[29] ), .A2(\b[29] ), .ZN(new_n726_));
  NOR2_X1    g0340(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1   g0341(.A1(new_n720_), .A2(new_n727_), .B(new_n722_), .ZN(\f[29] ));
  NOR3_X1    g0342(.A1(new_n719_), .A2(new_n717_), .A3(new_n725_), .ZN(new_n729_));
  XOR2_X1    g0343(.A1(\a[30] ), .A2(\b[30] ), .Z(new_n730_));
  OAI21_X1   g0344(.A1(new_n729_), .A2(new_n726_), .B(new_n730_), .ZN(new_n731_));
  INV_X1     g0345(.I(new_n726_), .ZN(new_n732_));
  INV_X1     g0346(.I(new_n717_), .ZN(new_n733_));
  OR4_X2     g0347(.A1(\a[26] ), .A2(\a[27] ), .A3(\b[26] ), .A4(\b[27] ), .Z(new_n734_));
  NAND2_X1   g0348(.A1(\a[28] ), .A2(\b[28] ), .ZN(new_n735_));
  NAND3_X1   g0349(.A1(new_n734_), .A2(new_n707_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1     g0350(.I(new_n725_), .ZN(new_n737_));
  NAND3_X1   g0351(.A1(new_n736_), .A2(new_n733_), .A3(new_n737_), .ZN(new_n738_));
  XNOR2_X1   g0352(.A1(\a[30] ), .A2(\b[30] ), .ZN(new_n739_));
  NAND3_X1   g0353(.A1(new_n738_), .A2(new_n732_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1   g0354(.A1(new_n740_), .A2(new_n731_), .ZN(\f[30] ));
  INV_X1     g0355(.I(\a[31] ), .ZN(new_n742_));
  INV_X1     g0356(.I(\b[31] ), .ZN(new_n743_));
  NAND2_X1   g0357(.A1(\a[30] ), .A2(\b[30] ), .ZN(new_n744_));
  INV_X1     g0358(.I(new_n744_), .ZN(new_n745_));
  NOR4_X1    g0359(.A1(\a[29] ), .A2(\a[30] ), .A3(\b[29] ), .A4(\b[30] ), .ZN(new_n746_));
  OAI21_X1   g0360(.A1(new_n745_), .A2(new_n746_), .B(new_n743_), .ZN(new_n747_));
  INV_X1     g0361(.I(new_n747_), .ZN(new_n748_));
  NOR3_X1    g0362(.A1(new_n745_), .A2(new_n746_), .A3(new_n743_), .ZN(new_n749_));
  OAI21_X1   g0363(.A1(new_n748_), .A2(new_n749_), .B(new_n742_), .ZN(new_n750_));
  INV_X1     g0364(.I(new_n749_), .ZN(new_n751_));
  NAND3_X1   g0365(.A1(new_n751_), .A2(\a[31] ), .A3(new_n747_), .ZN(new_n752_));
  NAND2_X1   g0366(.A1(new_n750_), .A2(new_n752_), .ZN(\f[31] ));
  NOR2_X1    g0367(.A1(\a[31] ), .A2(\b[31] ), .ZN(new_n754_));
  AND2_X2    g0368(.A1(\a[31] ), .A2(\b[31] ), .Z(new_n755_));
  NOR3_X1    g0369(.A1(new_n745_), .A2(new_n755_), .A3(new_n746_), .ZN(new_n756_));
  NOR2_X1    g0370(.A1(new_n756_), .A2(new_n754_), .ZN(new_n757_));
  XOR2_X1    g0371(.A1(\a[32] ), .A2(\b[32] ), .Z(new_n758_));
  NAND2_X1   g0372(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1     g0373(.I(\a[32] ), .ZN(new_n760_));
  INV_X1     g0374(.I(\b[32] ), .ZN(new_n761_));
  NOR2_X1    g0375(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1    g0376(.A1(\a[32] ), .A2(\b[32] ), .ZN(new_n763_));
  NOR2_X1    g0377(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1   g0378(.A1(new_n757_), .A2(new_n764_), .B(new_n759_), .ZN(\f[32] ));
  NOR3_X1    g0379(.A1(new_n756_), .A2(new_n754_), .A3(new_n762_), .ZN(new_n766_));
  XOR2_X1    g0380(.A1(\a[33] ), .A2(\b[33] ), .Z(new_n767_));
  OAI21_X1   g0381(.A1(new_n766_), .A2(new_n763_), .B(new_n767_), .ZN(new_n768_));
  INV_X1     g0382(.I(new_n763_), .ZN(new_n769_));
  INV_X1     g0383(.I(new_n754_), .ZN(new_n770_));
  OR4_X2     g0384(.A1(\a[29] ), .A2(\a[30] ), .A3(\b[29] ), .A4(\b[30] ), .Z(new_n771_));
  NAND2_X1   g0385(.A1(\a[31] ), .A2(\b[31] ), .ZN(new_n772_));
  NAND3_X1   g0386(.A1(new_n771_), .A2(new_n744_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1     g0387(.I(new_n762_), .ZN(new_n774_));
  NAND3_X1   g0388(.A1(new_n773_), .A2(new_n770_), .A3(new_n774_), .ZN(new_n775_));
  XNOR2_X1   g0389(.A1(\a[33] ), .A2(\b[33] ), .ZN(new_n776_));
  NAND3_X1   g0390(.A1(new_n775_), .A2(new_n769_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1   g0391(.A1(new_n777_), .A2(new_n768_), .ZN(\f[33] ));
  INV_X1     g0392(.I(\a[34] ), .ZN(new_n779_));
  INV_X1     g0393(.I(\b[34] ), .ZN(new_n780_));
  NAND2_X1   g0394(.A1(\a[33] ), .A2(\b[33] ), .ZN(new_n781_));
  INV_X1     g0395(.I(new_n781_), .ZN(new_n782_));
  NOR4_X1    g0396(.A1(\a[32] ), .A2(\a[33] ), .A3(\b[32] ), .A4(\b[33] ), .ZN(new_n783_));
  OAI21_X1   g0397(.A1(new_n782_), .A2(new_n783_), .B(new_n780_), .ZN(new_n784_));
  INV_X1     g0398(.I(new_n784_), .ZN(new_n785_));
  NOR3_X1    g0399(.A1(new_n782_), .A2(new_n783_), .A3(new_n780_), .ZN(new_n786_));
  OAI21_X1   g0400(.A1(new_n785_), .A2(new_n786_), .B(new_n779_), .ZN(new_n787_));
  INV_X1     g0401(.I(new_n786_), .ZN(new_n788_));
  NAND3_X1   g0402(.A1(new_n788_), .A2(\a[34] ), .A3(new_n784_), .ZN(new_n789_));
  NAND2_X1   g0403(.A1(new_n787_), .A2(new_n789_), .ZN(\f[34] ));
  NOR2_X1    g0404(.A1(\a[34] ), .A2(\b[34] ), .ZN(new_n791_));
  AND2_X2    g0405(.A1(\a[34] ), .A2(\b[34] ), .Z(new_n792_));
  NOR3_X1    g0406(.A1(new_n782_), .A2(new_n792_), .A3(new_n783_), .ZN(new_n793_));
  NOR2_X1    g0407(.A1(new_n793_), .A2(new_n791_), .ZN(new_n794_));
  XOR2_X1    g0408(.A1(\a[35] ), .A2(\b[35] ), .Z(new_n795_));
  NAND2_X1   g0409(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1     g0410(.I(\a[35] ), .ZN(new_n797_));
  INV_X1     g0411(.I(\b[35] ), .ZN(new_n798_));
  NOR2_X1    g0412(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1    g0413(.A1(\a[35] ), .A2(\b[35] ), .ZN(new_n800_));
  NOR2_X1    g0414(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1   g0415(.A1(new_n794_), .A2(new_n801_), .B(new_n796_), .ZN(\f[35] ));
  NOR3_X1    g0416(.A1(new_n793_), .A2(new_n791_), .A3(new_n799_), .ZN(new_n803_));
  XOR2_X1    g0417(.A1(\a[36] ), .A2(\b[36] ), .Z(new_n804_));
  OAI21_X1   g0418(.A1(new_n803_), .A2(new_n800_), .B(new_n804_), .ZN(new_n805_));
  INV_X1     g0419(.I(new_n800_), .ZN(new_n806_));
  INV_X1     g0420(.I(new_n791_), .ZN(new_n807_));
  OR4_X2     g0421(.A1(\a[32] ), .A2(\a[33] ), .A3(\b[32] ), .A4(\b[33] ), .Z(new_n808_));
  NAND2_X1   g0422(.A1(\a[34] ), .A2(\b[34] ), .ZN(new_n809_));
  NAND3_X1   g0423(.A1(new_n808_), .A2(new_n781_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1     g0424(.I(new_n799_), .ZN(new_n811_));
  NAND3_X1   g0425(.A1(new_n810_), .A2(new_n807_), .A3(new_n811_), .ZN(new_n812_));
  XNOR2_X1   g0426(.A1(\a[36] ), .A2(\b[36] ), .ZN(new_n813_));
  NAND3_X1   g0427(.A1(new_n812_), .A2(new_n806_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1   g0428(.A1(new_n814_), .A2(new_n805_), .ZN(\f[36] ));
  INV_X1     g0429(.I(\a[37] ), .ZN(new_n816_));
  INV_X1     g0430(.I(\b[37] ), .ZN(new_n817_));
  NAND2_X1   g0431(.A1(\a[36] ), .A2(\b[36] ), .ZN(new_n818_));
  INV_X1     g0432(.I(new_n818_), .ZN(new_n819_));
  NOR4_X1    g0433(.A1(\a[35] ), .A2(\a[36] ), .A3(\b[35] ), .A4(\b[36] ), .ZN(new_n820_));
  OAI21_X1   g0434(.A1(new_n819_), .A2(new_n820_), .B(new_n817_), .ZN(new_n821_));
  INV_X1     g0435(.I(new_n821_), .ZN(new_n822_));
  NOR3_X1    g0436(.A1(new_n819_), .A2(new_n820_), .A3(new_n817_), .ZN(new_n823_));
  OAI21_X1   g0437(.A1(new_n822_), .A2(new_n823_), .B(new_n816_), .ZN(new_n824_));
  INV_X1     g0438(.I(new_n823_), .ZN(new_n825_));
  NAND3_X1   g0439(.A1(new_n825_), .A2(\a[37] ), .A3(new_n821_), .ZN(new_n826_));
  NAND2_X1   g0440(.A1(new_n824_), .A2(new_n826_), .ZN(\f[37] ));
  NOR2_X1    g0441(.A1(\a[37] ), .A2(\b[37] ), .ZN(new_n828_));
  AND2_X2    g0442(.A1(\a[37] ), .A2(\b[37] ), .Z(new_n829_));
  NOR3_X1    g0443(.A1(new_n819_), .A2(new_n829_), .A3(new_n820_), .ZN(new_n830_));
  NOR2_X1    g0444(.A1(new_n830_), .A2(new_n828_), .ZN(new_n831_));
  XOR2_X1    g0445(.A1(\a[38] ), .A2(\b[38] ), .Z(new_n832_));
  NAND2_X1   g0446(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1     g0447(.I(\a[38] ), .ZN(new_n834_));
  INV_X1     g0448(.I(\b[38] ), .ZN(new_n835_));
  NOR2_X1    g0449(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1    g0450(.A1(\a[38] ), .A2(\b[38] ), .ZN(new_n837_));
  NOR2_X1    g0451(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1   g0452(.A1(new_n831_), .A2(new_n838_), .B(new_n833_), .ZN(\f[38] ));
  NOR3_X1    g0453(.A1(new_n830_), .A2(new_n828_), .A3(new_n836_), .ZN(new_n840_));
  XOR2_X1    g0454(.A1(\a[39] ), .A2(\b[39] ), .Z(new_n841_));
  OAI21_X1   g0455(.A1(new_n840_), .A2(new_n837_), .B(new_n841_), .ZN(new_n842_));
  INV_X1     g0456(.I(new_n837_), .ZN(new_n843_));
  INV_X1     g0457(.I(new_n828_), .ZN(new_n844_));
  OR4_X2     g0458(.A1(\a[35] ), .A2(\a[36] ), .A3(\b[35] ), .A4(\b[36] ), .Z(new_n845_));
  NAND2_X1   g0459(.A1(\a[37] ), .A2(\b[37] ), .ZN(new_n846_));
  NAND3_X1   g0460(.A1(new_n845_), .A2(new_n818_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1     g0461(.I(new_n836_), .ZN(new_n848_));
  NAND3_X1   g0462(.A1(new_n847_), .A2(new_n844_), .A3(new_n848_), .ZN(new_n849_));
  XNOR2_X1   g0463(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n850_));
  NAND3_X1   g0464(.A1(new_n849_), .A2(new_n843_), .A3(new_n850_), .ZN(new_n851_));
  NAND2_X1   g0465(.A1(new_n851_), .A2(new_n842_), .ZN(\f[39] ));
  INV_X1     g0466(.I(\a[40] ), .ZN(new_n853_));
  INV_X1     g0467(.I(\b[40] ), .ZN(new_n854_));
  NAND2_X1   g0468(.A1(\a[39] ), .A2(\b[39] ), .ZN(new_n855_));
  INV_X1     g0469(.I(new_n855_), .ZN(new_n856_));
  NOR4_X1    g0470(.A1(\a[38] ), .A2(\a[39] ), .A3(\b[38] ), .A4(\b[39] ), .ZN(new_n857_));
  OAI21_X1   g0471(.A1(new_n856_), .A2(new_n857_), .B(new_n854_), .ZN(new_n858_));
  INV_X1     g0472(.I(new_n858_), .ZN(new_n859_));
  NOR3_X1    g0473(.A1(new_n856_), .A2(new_n857_), .A3(new_n854_), .ZN(new_n860_));
  OAI21_X1   g0474(.A1(new_n859_), .A2(new_n860_), .B(new_n853_), .ZN(new_n861_));
  INV_X1     g0475(.I(new_n860_), .ZN(new_n862_));
  NAND3_X1   g0476(.A1(new_n862_), .A2(\a[40] ), .A3(new_n858_), .ZN(new_n863_));
  NAND2_X1   g0477(.A1(new_n861_), .A2(new_n863_), .ZN(\f[40] ));
  NOR2_X1    g0478(.A1(\a[40] ), .A2(\b[40] ), .ZN(new_n865_));
  AND2_X2    g0479(.A1(\a[40] ), .A2(\b[40] ), .Z(new_n866_));
  NOR3_X1    g0480(.A1(new_n856_), .A2(new_n866_), .A3(new_n857_), .ZN(new_n867_));
  NOR2_X1    g0481(.A1(new_n867_), .A2(new_n865_), .ZN(new_n868_));
  XOR2_X1    g0482(.A1(\a[41] ), .A2(\b[41] ), .Z(new_n869_));
  NAND2_X1   g0483(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1     g0484(.I(\a[41] ), .ZN(new_n871_));
  INV_X1     g0485(.I(\b[41] ), .ZN(new_n872_));
  NOR2_X1    g0486(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NOR2_X1    g0487(.A1(\a[41] ), .A2(\b[41] ), .ZN(new_n874_));
  NOR2_X1    g0488(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1   g0489(.A1(new_n868_), .A2(new_n875_), .B(new_n870_), .ZN(\f[41] ));
  NOR3_X1    g0490(.A1(new_n867_), .A2(new_n865_), .A3(new_n873_), .ZN(new_n877_));
  XOR2_X1    g0491(.A1(\a[42] ), .A2(\b[42] ), .Z(new_n878_));
  OAI21_X1   g0492(.A1(new_n877_), .A2(new_n874_), .B(new_n878_), .ZN(new_n879_));
  INV_X1     g0493(.I(new_n874_), .ZN(new_n880_));
  INV_X1     g0494(.I(new_n865_), .ZN(new_n881_));
  OR4_X2     g0495(.A1(\a[38] ), .A2(\a[39] ), .A3(\b[38] ), .A4(\b[39] ), .Z(new_n882_));
  NAND2_X1   g0496(.A1(\a[40] ), .A2(\b[40] ), .ZN(new_n883_));
  NAND3_X1   g0497(.A1(new_n882_), .A2(new_n855_), .A3(new_n883_), .ZN(new_n884_));
  INV_X1     g0498(.I(new_n873_), .ZN(new_n885_));
  NAND3_X1   g0499(.A1(new_n884_), .A2(new_n881_), .A3(new_n885_), .ZN(new_n886_));
  XNOR2_X1   g0500(.A1(\a[42] ), .A2(\b[42] ), .ZN(new_n887_));
  NAND3_X1   g0501(.A1(new_n886_), .A2(new_n880_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1   g0502(.A1(new_n888_), .A2(new_n879_), .ZN(\f[42] ));
  INV_X1     g0503(.I(\a[43] ), .ZN(new_n890_));
  INV_X1     g0504(.I(\b[43] ), .ZN(new_n891_));
  NAND2_X1   g0505(.A1(\a[42] ), .A2(\b[42] ), .ZN(new_n892_));
  INV_X1     g0506(.I(new_n892_), .ZN(new_n893_));
  NOR4_X1    g0507(.A1(\a[41] ), .A2(\a[42] ), .A3(\b[41] ), .A4(\b[42] ), .ZN(new_n894_));
  OAI21_X1   g0508(.A1(new_n893_), .A2(new_n894_), .B(new_n891_), .ZN(new_n895_));
  INV_X1     g0509(.I(new_n895_), .ZN(new_n896_));
  NOR3_X1    g0510(.A1(new_n893_), .A2(new_n894_), .A3(new_n891_), .ZN(new_n897_));
  OAI21_X1   g0511(.A1(new_n896_), .A2(new_n897_), .B(new_n890_), .ZN(new_n898_));
  INV_X1     g0512(.I(new_n897_), .ZN(new_n899_));
  NAND3_X1   g0513(.A1(new_n899_), .A2(\a[43] ), .A3(new_n895_), .ZN(new_n900_));
  NAND2_X1   g0514(.A1(new_n898_), .A2(new_n900_), .ZN(\f[43] ));
  NOR2_X1    g0515(.A1(\a[43] ), .A2(\b[43] ), .ZN(new_n902_));
  AND2_X2    g0516(.A1(\a[43] ), .A2(\b[43] ), .Z(new_n903_));
  NOR3_X1    g0517(.A1(new_n893_), .A2(new_n903_), .A3(new_n894_), .ZN(new_n904_));
  NOR2_X1    g0518(.A1(new_n904_), .A2(new_n902_), .ZN(new_n905_));
  XOR2_X1    g0519(.A1(\a[44] ), .A2(\b[44] ), .Z(new_n906_));
  NAND2_X1   g0520(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1     g0521(.I(\a[44] ), .ZN(new_n908_));
  INV_X1     g0522(.I(\b[44] ), .ZN(new_n909_));
  NOR2_X1    g0523(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1    g0524(.A1(\a[44] ), .A2(\b[44] ), .ZN(new_n911_));
  NOR2_X1    g0525(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1   g0526(.A1(new_n905_), .A2(new_n912_), .B(new_n907_), .ZN(\f[44] ));
  NOR3_X1    g0527(.A1(new_n904_), .A2(new_n902_), .A3(new_n910_), .ZN(new_n914_));
  XOR2_X1    g0528(.A1(\a[45] ), .A2(\b[45] ), .Z(new_n915_));
  OAI21_X1   g0529(.A1(new_n914_), .A2(new_n911_), .B(new_n915_), .ZN(new_n916_));
  INV_X1     g0530(.I(new_n911_), .ZN(new_n917_));
  INV_X1     g0531(.I(new_n902_), .ZN(new_n918_));
  OR4_X2     g0532(.A1(\a[41] ), .A2(\a[42] ), .A3(\b[41] ), .A4(\b[42] ), .Z(new_n919_));
  NAND2_X1   g0533(.A1(\a[43] ), .A2(\b[43] ), .ZN(new_n920_));
  NAND3_X1   g0534(.A1(new_n919_), .A2(new_n892_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1     g0535(.I(new_n910_), .ZN(new_n922_));
  NAND3_X1   g0536(.A1(new_n921_), .A2(new_n918_), .A3(new_n922_), .ZN(new_n923_));
  XNOR2_X1   g0537(.A1(\a[45] ), .A2(\b[45] ), .ZN(new_n924_));
  NAND3_X1   g0538(.A1(new_n923_), .A2(new_n917_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1   g0539(.A1(new_n925_), .A2(new_n916_), .ZN(\f[45] ));
  INV_X1     g0540(.I(\a[46] ), .ZN(new_n927_));
  INV_X1     g0541(.I(\b[46] ), .ZN(new_n928_));
  NAND2_X1   g0542(.A1(\a[45] ), .A2(\b[45] ), .ZN(new_n929_));
  INV_X1     g0543(.I(new_n929_), .ZN(new_n930_));
  NOR4_X1    g0544(.A1(\a[44] ), .A2(\a[45] ), .A3(\b[44] ), .A4(\b[45] ), .ZN(new_n931_));
  OAI21_X1   g0545(.A1(new_n930_), .A2(new_n931_), .B(new_n928_), .ZN(new_n932_));
  INV_X1     g0546(.I(new_n932_), .ZN(new_n933_));
  NOR3_X1    g0547(.A1(new_n930_), .A2(new_n931_), .A3(new_n928_), .ZN(new_n934_));
  OAI21_X1   g0548(.A1(new_n933_), .A2(new_n934_), .B(new_n927_), .ZN(new_n935_));
  INV_X1     g0549(.I(new_n934_), .ZN(new_n936_));
  NAND3_X1   g0550(.A1(new_n936_), .A2(\a[46] ), .A3(new_n932_), .ZN(new_n937_));
  NAND2_X1   g0551(.A1(new_n935_), .A2(new_n937_), .ZN(\f[46] ));
  NOR2_X1    g0552(.A1(\a[46] ), .A2(\b[46] ), .ZN(new_n939_));
  AND2_X2    g0553(.A1(\a[46] ), .A2(\b[46] ), .Z(new_n940_));
  NOR3_X1    g0554(.A1(new_n930_), .A2(new_n940_), .A3(new_n931_), .ZN(new_n941_));
  NOR2_X1    g0555(.A1(new_n941_), .A2(new_n939_), .ZN(new_n942_));
  XOR2_X1    g0556(.A1(\a[47] ), .A2(\b[47] ), .Z(new_n943_));
  NAND2_X1   g0557(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1     g0558(.I(\a[47] ), .ZN(new_n945_));
  INV_X1     g0559(.I(\b[47] ), .ZN(new_n946_));
  NOR2_X1    g0560(.A1(new_n945_), .A2(new_n946_), .ZN(new_n947_));
  NOR2_X1    g0561(.A1(\a[47] ), .A2(\b[47] ), .ZN(new_n948_));
  NOR2_X1    g0562(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  OAI21_X1   g0563(.A1(new_n942_), .A2(new_n949_), .B(new_n944_), .ZN(\f[47] ));
  NOR3_X1    g0564(.A1(new_n941_), .A2(new_n939_), .A3(new_n947_), .ZN(new_n951_));
  XOR2_X1    g0565(.A1(\a[48] ), .A2(\b[48] ), .Z(new_n952_));
  OAI21_X1   g0566(.A1(new_n951_), .A2(new_n948_), .B(new_n952_), .ZN(new_n953_));
  INV_X1     g0567(.I(new_n948_), .ZN(new_n954_));
  INV_X1     g0568(.I(new_n939_), .ZN(new_n955_));
  OR4_X2     g0569(.A1(\a[44] ), .A2(\a[45] ), .A3(\b[44] ), .A4(\b[45] ), .Z(new_n956_));
  NAND2_X1   g0570(.A1(\a[46] ), .A2(\b[46] ), .ZN(new_n957_));
  NAND3_X1   g0571(.A1(new_n956_), .A2(new_n929_), .A3(new_n957_), .ZN(new_n958_));
  INV_X1     g0572(.I(new_n947_), .ZN(new_n959_));
  NAND3_X1   g0573(.A1(new_n958_), .A2(new_n955_), .A3(new_n959_), .ZN(new_n960_));
  XNOR2_X1   g0574(.A1(\a[48] ), .A2(\b[48] ), .ZN(new_n961_));
  NAND3_X1   g0575(.A1(new_n960_), .A2(new_n954_), .A3(new_n961_), .ZN(new_n962_));
  NAND2_X1   g0576(.A1(new_n962_), .A2(new_n953_), .ZN(\f[48] ));
  INV_X1     g0577(.I(\a[49] ), .ZN(new_n964_));
  INV_X1     g0578(.I(\b[49] ), .ZN(new_n965_));
  NAND2_X1   g0579(.A1(\a[48] ), .A2(\b[48] ), .ZN(new_n966_));
  INV_X1     g0580(.I(new_n966_), .ZN(new_n967_));
  NOR4_X1    g0581(.A1(\a[47] ), .A2(\a[48] ), .A3(\b[47] ), .A4(\b[48] ), .ZN(new_n968_));
  OAI21_X1   g0582(.A1(new_n967_), .A2(new_n968_), .B(new_n965_), .ZN(new_n969_));
  INV_X1     g0583(.I(new_n969_), .ZN(new_n970_));
  NOR3_X1    g0584(.A1(new_n967_), .A2(new_n968_), .A3(new_n965_), .ZN(new_n971_));
  OAI21_X1   g0585(.A1(new_n970_), .A2(new_n971_), .B(new_n964_), .ZN(new_n972_));
  INV_X1     g0586(.I(new_n971_), .ZN(new_n973_));
  NAND3_X1   g0587(.A1(new_n973_), .A2(\a[49] ), .A3(new_n969_), .ZN(new_n974_));
  NAND2_X1   g0588(.A1(new_n972_), .A2(new_n974_), .ZN(\f[49] ));
  NOR2_X1    g0589(.A1(\a[49] ), .A2(\b[49] ), .ZN(new_n976_));
  AND2_X2    g0590(.A1(\a[49] ), .A2(\b[49] ), .Z(new_n977_));
  NOR3_X1    g0591(.A1(new_n967_), .A2(new_n977_), .A3(new_n968_), .ZN(new_n978_));
  NOR2_X1    g0592(.A1(new_n978_), .A2(new_n976_), .ZN(new_n979_));
  XOR2_X1    g0593(.A1(\a[50] ), .A2(\b[50] ), .Z(new_n980_));
  NAND2_X1   g0594(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1     g0595(.I(\a[50] ), .ZN(new_n982_));
  INV_X1     g0596(.I(\b[50] ), .ZN(new_n983_));
  NOR2_X1    g0597(.A1(new_n982_), .A2(new_n983_), .ZN(new_n984_));
  NOR2_X1    g0598(.A1(\a[50] ), .A2(\b[50] ), .ZN(new_n985_));
  NOR2_X1    g0599(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  OAI21_X1   g0600(.A1(new_n979_), .A2(new_n986_), .B(new_n981_), .ZN(\f[50] ));
  NOR3_X1    g0601(.A1(new_n978_), .A2(new_n976_), .A3(new_n984_), .ZN(new_n988_));
  XOR2_X1    g0602(.A1(\a[51] ), .A2(\b[51] ), .Z(new_n989_));
  OAI21_X1   g0603(.A1(new_n988_), .A2(new_n985_), .B(new_n989_), .ZN(new_n990_));
  INV_X1     g0604(.I(new_n985_), .ZN(new_n991_));
  INV_X1     g0605(.I(new_n976_), .ZN(new_n992_));
  OR4_X2     g0606(.A1(\a[47] ), .A2(\a[48] ), .A3(\b[47] ), .A4(\b[48] ), .Z(new_n993_));
  NAND2_X1   g0607(.A1(\a[49] ), .A2(\b[49] ), .ZN(new_n994_));
  NAND3_X1   g0608(.A1(new_n993_), .A2(new_n966_), .A3(new_n994_), .ZN(new_n995_));
  INV_X1     g0609(.I(new_n984_), .ZN(new_n996_));
  NAND3_X1   g0610(.A1(new_n995_), .A2(new_n992_), .A3(new_n996_), .ZN(new_n997_));
  XNOR2_X1   g0611(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n998_));
  NAND3_X1   g0612(.A1(new_n997_), .A2(new_n991_), .A3(new_n998_), .ZN(new_n999_));
  NAND2_X1   g0613(.A1(new_n999_), .A2(new_n990_), .ZN(\f[51] ));
  INV_X1     g0614(.I(\a[52] ), .ZN(new_n1001_));
  INV_X1     g0615(.I(\b[52] ), .ZN(new_n1002_));
  NAND2_X1   g0616(.A1(\a[51] ), .A2(\b[51] ), .ZN(new_n1003_));
  INV_X1     g0617(.I(new_n1003_), .ZN(new_n1004_));
  NOR4_X1    g0618(.A1(\a[50] ), .A2(\a[51] ), .A3(\b[50] ), .A4(\b[51] ), .ZN(new_n1005_));
  OAI21_X1   g0619(.A1(new_n1004_), .A2(new_n1005_), .B(new_n1002_), .ZN(new_n1006_));
  INV_X1     g0620(.I(new_n1006_), .ZN(new_n1007_));
  NOR3_X1    g0621(.A1(new_n1004_), .A2(new_n1005_), .A3(new_n1002_), .ZN(new_n1008_));
  OAI21_X1   g0622(.A1(new_n1007_), .A2(new_n1008_), .B(new_n1001_), .ZN(new_n1009_));
  INV_X1     g0623(.I(new_n1008_), .ZN(new_n1010_));
  NAND3_X1   g0624(.A1(new_n1010_), .A2(\a[52] ), .A3(new_n1006_), .ZN(new_n1011_));
  NAND2_X1   g0625(.A1(new_n1009_), .A2(new_n1011_), .ZN(\f[52] ));
  NOR2_X1    g0626(.A1(\a[52] ), .A2(\b[52] ), .ZN(new_n1013_));
  AND2_X2    g0627(.A1(\a[52] ), .A2(\b[52] ), .Z(new_n1014_));
  NOR3_X1    g0628(.A1(new_n1004_), .A2(new_n1014_), .A3(new_n1005_), .ZN(new_n1015_));
  NOR2_X1    g0629(.A1(new_n1015_), .A2(new_n1013_), .ZN(new_n1016_));
  XOR2_X1    g0630(.A1(\a[53] ), .A2(\b[53] ), .Z(new_n1017_));
  NAND2_X1   g0631(.A1(new_n1016_), .A2(new_n1017_), .ZN(new_n1018_));
  INV_X1     g0632(.I(\a[53] ), .ZN(new_n1019_));
  INV_X1     g0633(.I(\b[53] ), .ZN(new_n1020_));
  NOR2_X1    g0634(.A1(new_n1019_), .A2(new_n1020_), .ZN(new_n1021_));
  NOR2_X1    g0635(.A1(\a[53] ), .A2(\b[53] ), .ZN(new_n1022_));
  NOR2_X1    g0636(.A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1023_));
  OAI21_X1   g0637(.A1(new_n1016_), .A2(new_n1023_), .B(new_n1018_), .ZN(\f[53] ));
  NOR3_X1    g0638(.A1(new_n1015_), .A2(new_n1013_), .A3(new_n1021_), .ZN(new_n1025_));
  XOR2_X1    g0639(.A1(\a[54] ), .A2(\b[54] ), .Z(new_n1026_));
  OAI21_X1   g0640(.A1(new_n1025_), .A2(new_n1022_), .B(new_n1026_), .ZN(new_n1027_));
  INV_X1     g0641(.I(new_n1022_), .ZN(new_n1028_));
  INV_X1     g0642(.I(new_n1013_), .ZN(new_n1029_));
  OR4_X2     g0643(.A1(\a[50] ), .A2(\a[51] ), .A3(\b[50] ), .A4(\b[51] ), .Z(new_n1030_));
  NAND2_X1   g0644(.A1(\a[52] ), .A2(\b[52] ), .ZN(new_n1031_));
  NAND3_X1   g0645(.A1(new_n1030_), .A2(new_n1003_), .A3(new_n1031_), .ZN(new_n1032_));
  INV_X1     g0646(.I(new_n1021_), .ZN(new_n1033_));
  NAND3_X1   g0647(.A1(new_n1032_), .A2(new_n1029_), .A3(new_n1033_), .ZN(new_n1034_));
  XNOR2_X1   g0648(.A1(\a[54] ), .A2(\b[54] ), .ZN(new_n1035_));
  NAND3_X1   g0649(.A1(new_n1034_), .A2(new_n1028_), .A3(new_n1035_), .ZN(new_n1036_));
  NAND2_X1   g0650(.A1(new_n1036_), .A2(new_n1027_), .ZN(\f[54] ));
  INV_X1     g0651(.I(\a[55] ), .ZN(new_n1038_));
  INV_X1     g0652(.I(\b[55] ), .ZN(new_n1039_));
  NAND2_X1   g0653(.A1(\a[54] ), .A2(\b[54] ), .ZN(new_n1040_));
  INV_X1     g0654(.I(new_n1040_), .ZN(new_n1041_));
  NOR4_X1    g0655(.A1(\a[53] ), .A2(\a[54] ), .A3(\b[53] ), .A4(\b[54] ), .ZN(new_n1042_));
  OAI21_X1   g0656(.A1(new_n1041_), .A2(new_n1042_), .B(new_n1039_), .ZN(new_n1043_));
  INV_X1     g0657(.I(new_n1043_), .ZN(new_n1044_));
  NOR3_X1    g0658(.A1(new_n1041_), .A2(new_n1042_), .A3(new_n1039_), .ZN(new_n1045_));
  OAI21_X1   g0659(.A1(new_n1044_), .A2(new_n1045_), .B(new_n1038_), .ZN(new_n1046_));
  INV_X1     g0660(.I(new_n1045_), .ZN(new_n1047_));
  NAND3_X1   g0661(.A1(new_n1047_), .A2(\a[55] ), .A3(new_n1043_), .ZN(new_n1048_));
  NAND2_X1   g0662(.A1(new_n1046_), .A2(new_n1048_), .ZN(\f[55] ));
  NOR2_X1    g0663(.A1(\a[55] ), .A2(\b[55] ), .ZN(new_n1050_));
  AND2_X2    g0664(.A1(\a[55] ), .A2(\b[55] ), .Z(new_n1051_));
  NOR3_X1    g0665(.A1(new_n1041_), .A2(new_n1051_), .A3(new_n1042_), .ZN(new_n1052_));
  NOR2_X1    g0666(.A1(new_n1052_), .A2(new_n1050_), .ZN(new_n1053_));
  XOR2_X1    g0667(.A1(\a[56] ), .A2(\b[56] ), .Z(new_n1054_));
  NAND2_X1   g0668(.A1(new_n1053_), .A2(new_n1054_), .ZN(new_n1055_));
  INV_X1     g0669(.I(\a[56] ), .ZN(new_n1056_));
  INV_X1     g0670(.I(\b[56] ), .ZN(new_n1057_));
  NOR2_X1    g0671(.A1(new_n1056_), .A2(new_n1057_), .ZN(new_n1058_));
  NOR2_X1    g0672(.A1(\a[56] ), .A2(\b[56] ), .ZN(new_n1059_));
  NOR2_X1    g0673(.A1(new_n1058_), .A2(new_n1059_), .ZN(new_n1060_));
  OAI21_X1   g0674(.A1(new_n1053_), .A2(new_n1060_), .B(new_n1055_), .ZN(\f[56] ));
  NOR3_X1    g0675(.A1(new_n1052_), .A2(new_n1050_), .A3(new_n1058_), .ZN(new_n1062_));
  XOR2_X1    g0676(.A1(\a[57] ), .A2(\b[57] ), .Z(new_n1063_));
  OAI21_X1   g0677(.A1(new_n1062_), .A2(new_n1059_), .B(new_n1063_), .ZN(new_n1064_));
  INV_X1     g0678(.I(new_n1059_), .ZN(new_n1065_));
  INV_X1     g0679(.I(new_n1050_), .ZN(new_n1066_));
  OR4_X2     g0680(.A1(\a[53] ), .A2(\a[54] ), .A3(\b[53] ), .A4(\b[54] ), .Z(new_n1067_));
  NAND2_X1   g0681(.A1(\a[55] ), .A2(\b[55] ), .ZN(new_n1068_));
  NAND3_X1   g0682(.A1(new_n1067_), .A2(new_n1040_), .A3(new_n1068_), .ZN(new_n1069_));
  INV_X1     g0683(.I(new_n1058_), .ZN(new_n1070_));
  NAND3_X1   g0684(.A1(new_n1069_), .A2(new_n1066_), .A3(new_n1070_), .ZN(new_n1071_));
  XNOR2_X1   g0685(.A1(\a[57] ), .A2(\b[57] ), .ZN(new_n1072_));
  NAND3_X1   g0686(.A1(new_n1071_), .A2(new_n1065_), .A3(new_n1072_), .ZN(new_n1073_));
  NAND2_X1   g0687(.A1(new_n1073_), .A2(new_n1064_), .ZN(\f[57] ));
  INV_X1     g0688(.I(\a[58] ), .ZN(new_n1075_));
  INV_X1     g0689(.I(\b[58] ), .ZN(new_n1076_));
  NAND2_X1   g0690(.A1(\a[57] ), .A2(\b[57] ), .ZN(new_n1077_));
  INV_X1     g0691(.I(new_n1077_), .ZN(new_n1078_));
  NOR4_X1    g0692(.A1(\a[56] ), .A2(\a[57] ), .A3(\b[56] ), .A4(\b[57] ), .ZN(new_n1079_));
  OAI21_X1   g0693(.A1(new_n1078_), .A2(new_n1079_), .B(new_n1076_), .ZN(new_n1080_));
  INV_X1     g0694(.I(new_n1080_), .ZN(new_n1081_));
  NOR3_X1    g0695(.A1(new_n1078_), .A2(new_n1079_), .A3(new_n1076_), .ZN(new_n1082_));
  OAI21_X1   g0696(.A1(new_n1081_), .A2(new_n1082_), .B(new_n1075_), .ZN(new_n1083_));
  INV_X1     g0697(.I(new_n1082_), .ZN(new_n1084_));
  NAND3_X1   g0698(.A1(new_n1084_), .A2(\a[58] ), .A3(new_n1080_), .ZN(new_n1085_));
  NAND2_X1   g0699(.A1(new_n1083_), .A2(new_n1085_), .ZN(\f[58] ));
  NOR2_X1    g0700(.A1(\a[58] ), .A2(\b[58] ), .ZN(new_n1087_));
  AND2_X2    g0701(.A1(\a[58] ), .A2(\b[58] ), .Z(new_n1088_));
  NOR3_X1    g0702(.A1(new_n1078_), .A2(new_n1088_), .A3(new_n1079_), .ZN(new_n1089_));
  NOR2_X1    g0703(.A1(new_n1089_), .A2(new_n1087_), .ZN(new_n1090_));
  XOR2_X1    g0704(.A1(\a[59] ), .A2(\b[59] ), .Z(new_n1091_));
  NAND2_X1   g0705(.A1(new_n1090_), .A2(new_n1091_), .ZN(new_n1092_));
  INV_X1     g0706(.I(\a[59] ), .ZN(new_n1093_));
  INV_X1     g0707(.I(\b[59] ), .ZN(new_n1094_));
  NOR2_X1    g0708(.A1(new_n1093_), .A2(new_n1094_), .ZN(new_n1095_));
  NOR2_X1    g0709(.A1(\a[59] ), .A2(\b[59] ), .ZN(new_n1096_));
  NOR2_X1    g0710(.A1(new_n1095_), .A2(new_n1096_), .ZN(new_n1097_));
  OAI21_X1   g0711(.A1(new_n1090_), .A2(new_n1097_), .B(new_n1092_), .ZN(\f[59] ));
  NOR3_X1    g0712(.A1(new_n1089_), .A2(new_n1087_), .A3(new_n1095_), .ZN(new_n1099_));
  XOR2_X1    g0713(.A1(\a[60] ), .A2(\b[60] ), .Z(new_n1100_));
  OAI21_X1   g0714(.A1(new_n1099_), .A2(new_n1096_), .B(new_n1100_), .ZN(new_n1101_));
  INV_X1     g0715(.I(new_n1096_), .ZN(new_n1102_));
  INV_X1     g0716(.I(new_n1087_), .ZN(new_n1103_));
  OR4_X2     g0717(.A1(\a[56] ), .A2(\a[57] ), .A3(\b[56] ), .A4(\b[57] ), .Z(new_n1104_));
  NAND2_X1   g0718(.A1(\a[58] ), .A2(\b[58] ), .ZN(new_n1105_));
  NAND3_X1   g0719(.A1(new_n1104_), .A2(new_n1077_), .A3(new_n1105_), .ZN(new_n1106_));
  INV_X1     g0720(.I(new_n1095_), .ZN(new_n1107_));
  NAND3_X1   g0721(.A1(new_n1106_), .A2(new_n1103_), .A3(new_n1107_), .ZN(new_n1108_));
  XNOR2_X1   g0722(.A1(\a[60] ), .A2(\b[60] ), .ZN(new_n1109_));
  NAND3_X1   g0723(.A1(new_n1108_), .A2(new_n1102_), .A3(new_n1109_), .ZN(new_n1110_));
  NAND2_X1   g0724(.A1(new_n1110_), .A2(new_n1101_), .ZN(\f[60] ));
  INV_X1     g0725(.I(\a[61] ), .ZN(new_n1112_));
  INV_X1     g0726(.I(\b[61] ), .ZN(new_n1113_));
  NAND2_X1   g0727(.A1(\a[60] ), .A2(\b[60] ), .ZN(new_n1114_));
  INV_X1     g0728(.I(new_n1114_), .ZN(new_n1115_));
  NOR4_X1    g0729(.A1(\a[59] ), .A2(\a[60] ), .A3(\b[59] ), .A4(\b[60] ), .ZN(new_n1116_));
  OAI21_X1   g0730(.A1(new_n1115_), .A2(new_n1116_), .B(new_n1113_), .ZN(new_n1117_));
  INV_X1     g0731(.I(new_n1117_), .ZN(new_n1118_));
  NOR3_X1    g0732(.A1(new_n1115_), .A2(new_n1116_), .A3(new_n1113_), .ZN(new_n1119_));
  OAI21_X1   g0733(.A1(new_n1118_), .A2(new_n1119_), .B(new_n1112_), .ZN(new_n1120_));
  INV_X1     g0734(.I(new_n1119_), .ZN(new_n1121_));
  NAND3_X1   g0735(.A1(new_n1121_), .A2(\a[61] ), .A3(new_n1117_), .ZN(new_n1122_));
  NAND2_X1   g0736(.A1(new_n1120_), .A2(new_n1122_), .ZN(\f[61] ));
  NOR2_X1    g0737(.A1(\a[61] ), .A2(\b[61] ), .ZN(new_n1124_));
  AND2_X2    g0738(.A1(\a[61] ), .A2(\b[61] ), .Z(new_n1125_));
  NOR3_X1    g0739(.A1(new_n1115_), .A2(new_n1125_), .A3(new_n1116_), .ZN(new_n1126_));
  NOR2_X1    g0740(.A1(new_n1126_), .A2(new_n1124_), .ZN(new_n1127_));
  XOR2_X1    g0741(.A1(\a[62] ), .A2(\b[62] ), .Z(new_n1128_));
  NAND2_X1   g0742(.A1(new_n1127_), .A2(new_n1128_), .ZN(new_n1129_));
  INV_X1     g0743(.I(\a[62] ), .ZN(new_n1130_));
  INV_X1     g0744(.I(\b[62] ), .ZN(new_n1131_));
  NOR2_X1    g0745(.A1(new_n1130_), .A2(new_n1131_), .ZN(new_n1132_));
  NOR2_X1    g0746(.A1(\a[62] ), .A2(\b[62] ), .ZN(new_n1133_));
  NOR2_X1    g0747(.A1(new_n1132_), .A2(new_n1133_), .ZN(new_n1134_));
  OAI21_X1   g0748(.A1(new_n1127_), .A2(new_n1134_), .B(new_n1129_), .ZN(\f[62] ));
  NOR3_X1    g0749(.A1(new_n1126_), .A2(new_n1124_), .A3(new_n1132_), .ZN(new_n1136_));
  XOR2_X1    g0750(.A1(\a[63] ), .A2(\b[63] ), .Z(new_n1137_));
  OAI21_X1   g0751(.A1(new_n1136_), .A2(new_n1133_), .B(new_n1137_), .ZN(new_n1138_));
  INV_X1     g0752(.I(new_n1133_), .ZN(new_n1139_));
  INV_X1     g0753(.I(new_n1124_), .ZN(new_n1140_));
  OR4_X2     g0754(.A1(\a[59] ), .A2(\a[60] ), .A3(\b[59] ), .A4(\b[60] ), .Z(new_n1141_));
  NAND2_X1   g0755(.A1(\a[61] ), .A2(\b[61] ), .ZN(new_n1142_));
  NAND3_X1   g0756(.A1(new_n1141_), .A2(new_n1114_), .A3(new_n1142_), .ZN(new_n1143_));
  INV_X1     g0757(.I(new_n1132_), .ZN(new_n1144_));
  NAND3_X1   g0758(.A1(new_n1143_), .A2(new_n1140_), .A3(new_n1144_), .ZN(new_n1145_));
  XNOR2_X1   g0759(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n1146_));
  NAND3_X1   g0760(.A1(new_n1145_), .A2(new_n1139_), .A3(new_n1146_), .ZN(new_n1147_));
  NAND2_X1   g0761(.A1(new_n1147_), .A2(new_n1138_), .ZN(\f[63] ));
  INV_X1     g0762(.I(\a[64] ), .ZN(new_n1149_));
  INV_X1     g0763(.I(\b[64] ), .ZN(new_n1150_));
  NAND2_X1   g0764(.A1(\a[63] ), .A2(\b[63] ), .ZN(new_n1151_));
  INV_X1     g0765(.I(new_n1151_), .ZN(new_n1152_));
  NOR4_X1    g0766(.A1(\a[62] ), .A2(\a[63] ), .A3(\b[62] ), .A4(\b[63] ), .ZN(new_n1153_));
  OAI21_X1   g0767(.A1(new_n1152_), .A2(new_n1153_), .B(new_n1150_), .ZN(new_n1154_));
  INV_X1     g0768(.I(new_n1154_), .ZN(new_n1155_));
  NOR3_X1    g0769(.A1(new_n1152_), .A2(new_n1153_), .A3(new_n1150_), .ZN(new_n1156_));
  OAI21_X1   g0770(.A1(new_n1155_), .A2(new_n1156_), .B(new_n1149_), .ZN(new_n1157_));
  INV_X1     g0771(.I(new_n1156_), .ZN(new_n1158_));
  NAND3_X1   g0772(.A1(new_n1158_), .A2(\a[64] ), .A3(new_n1154_), .ZN(new_n1159_));
  NAND2_X1   g0773(.A1(new_n1157_), .A2(new_n1159_), .ZN(\f[64] ));
  NOR2_X1    g0774(.A1(\a[64] ), .A2(\b[64] ), .ZN(new_n1161_));
  AND2_X2    g0775(.A1(\a[64] ), .A2(\b[64] ), .Z(new_n1162_));
  NOR3_X1    g0776(.A1(new_n1152_), .A2(new_n1162_), .A3(new_n1153_), .ZN(new_n1163_));
  NOR2_X1    g0777(.A1(new_n1163_), .A2(new_n1161_), .ZN(new_n1164_));
  XOR2_X1    g0778(.A1(\a[65] ), .A2(\b[65] ), .Z(new_n1165_));
  NAND2_X1   g0779(.A1(new_n1164_), .A2(new_n1165_), .ZN(new_n1166_));
  INV_X1     g0780(.I(\a[65] ), .ZN(new_n1167_));
  INV_X1     g0781(.I(\b[65] ), .ZN(new_n1168_));
  NOR2_X1    g0782(.A1(new_n1167_), .A2(new_n1168_), .ZN(new_n1169_));
  NOR2_X1    g0783(.A1(\a[65] ), .A2(\b[65] ), .ZN(new_n1170_));
  NOR2_X1    g0784(.A1(new_n1169_), .A2(new_n1170_), .ZN(new_n1171_));
  OAI21_X1   g0785(.A1(new_n1164_), .A2(new_n1171_), .B(new_n1166_), .ZN(\f[65] ));
  NOR3_X1    g0786(.A1(new_n1163_), .A2(new_n1161_), .A3(new_n1169_), .ZN(new_n1173_));
  XOR2_X1    g0787(.A1(\a[66] ), .A2(\b[66] ), .Z(new_n1174_));
  OAI21_X1   g0788(.A1(new_n1173_), .A2(new_n1170_), .B(new_n1174_), .ZN(new_n1175_));
  INV_X1     g0789(.I(new_n1170_), .ZN(new_n1176_));
  INV_X1     g0790(.I(new_n1161_), .ZN(new_n1177_));
  OR4_X2     g0791(.A1(\a[62] ), .A2(\a[63] ), .A3(\b[62] ), .A4(\b[63] ), .Z(new_n1178_));
  NAND2_X1   g0792(.A1(\a[64] ), .A2(\b[64] ), .ZN(new_n1179_));
  NAND3_X1   g0793(.A1(new_n1178_), .A2(new_n1151_), .A3(new_n1179_), .ZN(new_n1180_));
  INV_X1     g0794(.I(new_n1169_), .ZN(new_n1181_));
  NAND3_X1   g0795(.A1(new_n1180_), .A2(new_n1177_), .A3(new_n1181_), .ZN(new_n1182_));
  XNOR2_X1   g0796(.A1(\a[66] ), .A2(\b[66] ), .ZN(new_n1183_));
  NAND3_X1   g0797(.A1(new_n1182_), .A2(new_n1176_), .A3(new_n1183_), .ZN(new_n1184_));
  NAND2_X1   g0798(.A1(new_n1184_), .A2(new_n1175_), .ZN(\f[66] ));
  INV_X1     g0799(.I(\a[67] ), .ZN(new_n1186_));
  INV_X1     g0800(.I(\b[67] ), .ZN(new_n1187_));
  NAND2_X1   g0801(.A1(\a[66] ), .A2(\b[66] ), .ZN(new_n1188_));
  INV_X1     g0802(.I(new_n1188_), .ZN(new_n1189_));
  NOR4_X1    g0803(.A1(\a[65] ), .A2(\a[66] ), .A3(\b[65] ), .A4(\b[66] ), .ZN(new_n1190_));
  OAI21_X1   g0804(.A1(new_n1189_), .A2(new_n1190_), .B(new_n1187_), .ZN(new_n1191_));
  INV_X1     g0805(.I(new_n1191_), .ZN(new_n1192_));
  NOR3_X1    g0806(.A1(new_n1189_), .A2(new_n1190_), .A3(new_n1187_), .ZN(new_n1193_));
  OAI21_X1   g0807(.A1(new_n1192_), .A2(new_n1193_), .B(new_n1186_), .ZN(new_n1194_));
  INV_X1     g0808(.I(new_n1193_), .ZN(new_n1195_));
  NAND3_X1   g0809(.A1(new_n1195_), .A2(\a[67] ), .A3(new_n1191_), .ZN(new_n1196_));
  NAND2_X1   g0810(.A1(new_n1194_), .A2(new_n1196_), .ZN(\f[67] ));
  NOR2_X1    g0811(.A1(\a[67] ), .A2(\b[67] ), .ZN(new_n1198_));
  AND2_X2    g0812(.A1(\a[67] ), .A2(\b[67] ), .Z(new_n1199_));
  NOR3_X1    g0813(.A1(new_n1189_), .A2(new_n1199_), .A3(new_n1190_), .ZN(new_n1200_));
  NOR2_X1    g0814(.A1(new_n1200_), .A2(new_n1198_), .ZN(new_n1201_));
  XOR2_X1    g0815(.A1(\a[68] ), .A2(\b[68] ), .Z(new_n1202_));
  NAND2_X1   g0816(.A1(new_n1201_), .A2(new_n1202_), .ZN(new_n1203_));
  INV_X1     g0817(.I(\a[68] ), .ZN(new_n1204_));
  INV_X1     g0818(.I(\b[68] ), .ZN(new_n1205_));
  NOR2_X1    g0819(.A1(new_n1204_), .A2(new_n1205_), .ZN(new_n1206_));
  NOR2_X1    g0820(.A1(\a[68] ), .A2(\b[68] ), .ZN(new_n1207_));
  NOR2_X1    g0821(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1208_));
  OAI21_X1   g0822(.A1(new_n1201_), .A2(new_n1208_), .B(new_n1203_), .ZN(\f[68] ));
  NOR3_X1    g0823(.A1(new_n1200_), .A2(new_n1198_), .A3(new_n1206_), .ZN(new_n1210_));
  XOR2_X1    g0824(.A1(\a[69] ), .A2(\b[69] ), .Z(new_n1211_));
  OAI21_X1   g0825(.A1(new_n1210_), .A2(new_n1207_), .B(new_n1211_), .ZN(new_n1212_));
  INV_X1     g0826(.I(new_n1207_), .ZN(new_n1213_));
  INV_X1     g0827(.I(new_n1198_), .ZN(new_n1214_));
  OR4_X2     g0828(.A1(\a[65] ), .A2(\a[66] ), .A3(\b[65] ), .A4(\b[66] ), .Z(new_n1215_));
  NAND2_X1   g0829(.A1(\a[67] ), .A2(\b[67] ), .ZN(new_n1216_));
  NAND3_X1   g0830(.A1(new_n1215_), .A2(new_n1188_), .A3(new_n1216_), .ZN(new_n1217_));
  INV_X1     g0831(.I(new_n1206_), .ZN(new_n1218_));
  NAND3_X1   g0832(.A1(new_n1217_), .A2(new_n1214_), .A3(new_n1218_), .ZN(new_n1219_));
  XNOR2_X1   g0833(.A1(\a[69] ), .A2(\b[69] ), .ZN(new_n1220_));
  NAND3_X1   g0834(.A1(new_n1219_), .A2(new_n1213_), .A3(new_n1220_), .ZN(new_n1221_));
  NAND2_X1   g0835(.A1(new_n1221_), .A2(new_n1212_), .ZN(\f[69] ));
  INV_X1     g0836(.I(\a[70] ), .ZN(new_n1223_));
  INV_X1     g0837(.I(\b[70] ), .ZN(new_n1224_));
  NAND2_X1   g0838(.A1(\a[69] ), .A2(\b[69] ), .ZN(new_n1225_));
  INV_X1     g0839(.I(new_n1225_), .ZN(new_n1226_));
  NOR4_X1    g0840(.A1(\a[68] ), .A2(\a[69] ), .A3(\b[68] ), .A4(\b[69] ), .ZN(new_n1227_));
  OAI21_X1   g0841(.A1(new_n1226_), .A2(new_n1227_), .B(new_n1224_), .ZN(new_n1228_));
  INV_X1     g0842(.I(new_n1228_), .ZN(new_n1229_));
  NOR3_X1    g0843(.A1(new_n1226_), .A2(new_n1227_), .A3(new_n1224_), .ZN(new_n1230_));
  OAI21_X1   g0844(.A1(new_n1229_), .A2(new_n1230_), .B(new_n1223_), .ZN(new_n1231_));
  INV_X1     g0845(.I(new_n1230_), .ZN(new_n1232_));
  NAND3_X1   g0846(.A1(new_n1232_), .A2(\a[70] ), .A3(new_n1228_), .ZN(new_n1233_));
  NAND2_X1   g0847(.A1(new_n1231_), .A2(new_n1233_), .ZN(\f[70] ));
  NOR2_X1    g0848(.A1(\a[70] ), .A2(\b[70] ), .ZN(new_n1235_));
  AND2_X2    g0849(.A1(\a[70] ), .A2(\b[70] ), .Z(new_n1236_));
  NOR3_X1    g0850(.A1(new_n1226_), .A2(new_n1236_), .A3(new_n1227_), .ZN(new_n1237_));
  NOR2_X1    g0851(.A1(new_n1237_), .A2(new_n1235_), .ZN(new_n1238_));
  XOR2_X1    g0852(.A1(\a[71] ), .A2(\b[71] ), .Z(new_n1239_));
  NAND2_X1   g0853(.A1(new_n1238_), .A2(new_n1239_), .ZN(new_n1240_));
  INV_X1     g0854(.I(\a[71] ), .ZN(new_n1241_));
  INV_X1     g0855(.I(\b[71] ), .ZN(new_n1242_));
  NOR2_X1    g0856(.A1(new_n1241_), .A2(new_n1242_), .ZN(new_n1243_));
  NOR2_X1    g0857(.A1(\a[71] ), .A2(\b[71] ), .ZN(new_n1244_));
  NOR2_X1    g0858(.A1(new_n1243_), .A2(new_n1244_), .ZN(new_n1245_));
  OAI21_X1   g0859(.A1(new_n1238_), .A2(new_n1245_), .B(new_n1240_), .ZN(\f[71] ));
  NOR3_X1    g0860(.A1(new_n1237_), .A2(new_n1235_), .A3(new_n1243_), .ZN(new_n1247_));
  XOR2_X1    g0861(.A1(\a[72] ), .A2(\b[72] ), .Z(new_n1248_));
  OAI21_X1   g0862(.A1(new_n1247_), .A2(new_n1244_), .B(new_n1248_), .ZN(new_n1249_));
  INV_X1     g0863(.I(new_n1244_), .ZN(new_n1250_));
  INV_X1     g0864(.I(new_n1235_), .ZN(new_n1251_));
  OR4_X2     g0865(.A1(\a[68] ), .A2(\a[69] ), .A3(\b[68] ), .A4(\b[69] ), .Z(new_n1252_));
  NAND2_X1   g0866(.A1(\a[70] ), .A2(\b[70] ), .ZN(new_n1253_));
  NAND3_X1   g0867(.A1(new_n1252_), .A2(new_n1225_), .A3(new_n1253_), .ZN(new_n1254_));
  INV_X1     g0868(.I(new_n1243_), .ZN(new_n1255_));
  NAND3_X1   g0869(.A1(new_n1254_), .A2(new_n1251_), .A3(new_n1255_), .ZN(new_n1256_));
  XNOR2_X1   g0870(.A1(\a[72] ), .A2(\b[72] ), .ZN(new_n1257_));
  NAND3_X1   g0871(.A1(new_n1256_), .A2(new_n1250_), .A3(new_n1257_), .ZN(new_n1258_));
  NAND2_X1   g0872(.A1(new_n1258_), .A2(new_n1249_), .ZN(\f[72] ));
  INV_X1     g0873(.I(\a[73] ), .ZN(new_n1260_));
  INV_X1     g0874(.I(\b[73] ), .ZN(new_n1261_));
  NAND2_X1   g0875(.A1(\a[72] ), .A2(\b[72] ), .ZN(new_n1262_));
  INV_X1     g0876(.I(new_n1262_), .ZN(new_n1263_));
  NOR4_X1    g0877(.A1(\a[71] ), .A2(\a[72] ), .A3(\b[71] ), .A4(\b[72] ), .ZN(new_n1264_));
  OAI21_X1   g0878(.A1(new_n1263_), .A2(new_n1264_), .B(new_n1261_), .ZN(new_n1265_));
  INV_X1     g0879(.I(new_n1265_), .ZN(new_n1266_));
  NOR3_X1    g0880(.A1(new_n1263_), .A2(new_n1264_), .A3(new_n1261_), .ZN(new_n1267_));
  OAI21_X1   g0881(.A1(new_n1266_), .A2(new_n1267_), .B(new_n1260_), .ZN(new_n1268_));
  INV_X1     g0882(.I(new_n1267_), .ZN(new_n1269_));
  NAND3_X1   g0883(.A1(new_n1269_), .A2(\a[73] ), .A3(new_n1265_), .ZN(new_n1270_));
  NAND2_X1   g0884(.A1(new_n1268_), .A2(new_n1270_), .ZN(\f[73] ));
  NOR2_X1    g0885(.A1(\a[73] ), .A2(\b[73] ), .ZN(new_n1272_));
  AND2_X2    g0886(.A1(\a[73] ), .A2(\b[73] ), .Z(new_n1273_));
  NOR3_X1    g0887(.A1(new_n1263_), .A2(new_n1273_), .A3(new_n1264_), .ZN(new_n1274_));
  NOR2_X1    g0888(.A1(new_n1274_), .A2(new_n1272_), .ZN(new_n1275_));
  XOR2_X1    g0889(.A1(\a[74] ), .A2(\b[74] ), .Z(new_n1276_));
  NAND2_X1   g0890(.A1(new_n1275_), .A2(new_n1276_), .ZN(new_n1277_));
  INV_X1     g0891(.I(\a[74] ), .ZN(new_n1278_));
  INV_X1     g0892(.I(\b[74] ), .ZN(new_n1279_));
  NOR2_X1    g0893(.A1(new_n1278_), .A2(new_n1279_), .ZN(new_n1280_));
  NOR2_X1    g0894(.A1(\a[74] ), .A2(\b[74] ), .ZN(new_n1281_));
  NOR2_X1    g0895(.A1(new_n1280_), .A2(new_n1281_), .ZN(new_n1282_));
  OAI21_X1   g0896(.A1(new_n1275_), .A2(new_n1282_), .B(new_n1277_), .ZN(\f[74] ));
  NOR3_X1    g0897(.A1(new_n1274_), .A2(new_n1272_), .A3(new_n1280_), .ZN(new_n1284_));
  XOR2_X1    g0898(.A1(\a[75] ), .A2(\b[75] ), .Z(new_n1285_));
  OAI21_X1   g0899(.A1(new_n1284_), .A2(new_n1281_), .B(new_n1285_), .ZN(new_n1286_));
  INV_X1     g0900(.I(new_n1281_), .ZN(new_n1287_));
  INV_X1     g0901(.I(new_n1272_), .ZN(new_n1288_));
  OR4_X2     g0902(.A1(\a[71] ), .A2(\a[72] ), .A3(\b[71] ), .A4(\b[72] ), .Z(new_n1289_));
  NAND2_X1   g0903(.A1(\a[73] ), .A2(\b[73] ), .ZN(new_n1290_));
  NAND3_X1   g0904(.A1(new_n1289_), .A2(new_n1262_), .A3(new_n1290_), .ZN(new_n1291_));
  INV_X1     g0905(.I(new_n1280_), .ZN(new_n1292_));
  NAND3_X1   g0906(.A1(new_n1291_), .A2(new_n1288_), .A3(new_n1292_), .ZN(new_n1293_));
  XNOR2_X1   g0907(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n1294_));
  NAND3_X1   g0908(.A1(new_n1293_), .A2(new_n1287_), .A3(new_n1294_), .ZN(new_n1295_));
  NAND2_X1   g0909(.A1(new_n1295_), .A2(new_n1286_), .ZN(\f[75] ));
  INV_X1     g0910(.I(\a[76] ), .ZN(new_n1297_));
  INV_X1     g0911(.I(\b[76] ), .ZN(new_n1298_));
  NAND2_X1   g0912(.A1(\a[75] ), .A2(\b[75] ), .ZN(new_n1299_));
  INV_X1     g0913(.I(new_n1299_), .ZN(new_n1300_));
  NOR4_X1    g0914(.A1(\a[74] ), .A2(\a[75] ), .A3(\b[74] ), .A4(\b[75] ), .ZN(new_n1301_));
  OAI21_X1   g0915(.A1(new_n1300_), .A2(new_n1301_), .B(new_n1298_), .ZN(new_n1302_));
  INV_X1     g0916(.I(new_n1302_), .ZN(new_n1303_));
  NOR3_X1    g0917(.A1(new_n1300_), .A2(new_n1301_), .A3(new_n1298_), .ZN(new_n1304_));
  OAI21_X1   g0918(.A1(new_n1303_), .A2(new_n1304_), .B(new_n1297_), .ZN(new_n1305_));
  INV_X1     g0919(.I(new_n1304_), .ZN(new_n1306_));
  NAND3_X1   g0920(.A1(new_n1306_), .A2(\a[76] ), .A3(new_n1302_), .ZN(new_n1307_));
  NAND2_X1   g0921(.A1(new_n1305_), .A2(new_n1307_), .ZN(\f[76] ));
  NOR2_X1    g0922(.A1(\a[76] ), .A2(\b[76] ), .ZN(new_n1309_));
  AND2_X2    g0923(.A1(\a[76] ), .A2(\b[76] ), .Z(new_n1310_));
  NOR3_X1    g0924(.A1(new_n1300_), .A2(new_n1310_), .A3(new_n1301_), .ZN(new_n1311_));
  NOR2_X1    g0925(.A1(new_n1311_), .A2(new_n1309_), .ZN(new_n1312_));
  XOR2_X1    g0926(.A1(\a[77] ), .A2(\b[77] ), .Z(new_n1313_));
  NAND2_X1   g0927(.A1(new_n1312_), .A2(new_n1313_), .ZN(new_n1314_));
  INV_X1     g0928(.I(\a[77] ), .ZN(new_n1315_));
  INV_X1     g0929(.I(\b[77] ), .ZN(new_n1316_));
  NOR2_X1    g0930(.A1(new_n1315_), .A2(new_n1316_), .ZN(new_n1317_));
  NOR2_X1    g0931(.A1(\a[77] ), .A2(\b[77] ), .ZN(new_n1318_));
  NOR2_X1    g0932(.A1(new_n1317_), .A2(new_n1318_), .ZN(new_n1319_));
  OAI21_X1   g0933(.A1(new_n1312_), .A2(new_n1319_), .B(new_n1314_), .ZN(\f[77] ));
  NOR3_X1    g0934(.A1(new_n1311_), .A2(new_n1309_), .A3(new_n1317_), .ZN(new_n1321_));
  XOR2_X1    g0935(.A1(\a[78] ), .A2(\b[78] ), .Z(new_n1322_));
  OAI21_X1   g0936(.A1(new_n1321_), .A2(new_n1318_), .B(new_n1322_), .ZN(new_n1323_));
  INV_X1     g0937(.I(new_n1318_), .ZN(new_n1324_));
  INV_X1     g0938(.I(new_n1309_), .ZN(new_n1325_));
  OR4_X2     g0939(.A1(\a[74] ), .A2(\a[75] ), .A3(\b[74] ), .A4(\b[75] ), .Z(new_n1326_));
  NAND2_X1   g0940(.A1(\a[76] ), .A2(\b[76] ), .ZN(new_n1327_));
  NAND3_X1   g0941(.A1(new_n1326_), .A2(new_n1299_), .A3(new_n1327_), .ZN(new_n1328_));
  INV_X1     g0942(.I(new_n1317_), .ZN(new_n1329_));
  NAND3_X1   g0943(.A1(new_n1328_), .A2(new_n1325_), .A3(new_n1329_), .ZN(new_n1330_));
  XNOR2_X1   g0944(.A1(\a[78] ), .A2(\b[78] ), .ZN(new_n1331_));
  NAND3_X1   g0945(.A1(new_n1330_), .A2(new_n1324_), .A3(new_n1331_), .ZN(new_n1332_));
  NAND2_X1   g0946(.A1(new_n1332_), .A2(new_n1323_), .ZN(\f[78] ));
  INV_X1     g0947(.I(\a[79] ), .ZN(new_n1334_));
  INV_X1     g0948(.I(\b[79] ), .ZN(new_n1335_));
  NAND2_X1   g0949(.A1(\a[78] ), .A2(\b[78] ), .ZN(new_n1336_));
  INV_X1     g0950(.I(new_n1336_), .ZN(new_n1337_));
  NOR4_X1    g0951(.A1(\a[77] ), .A2(\a[78] ), .A3(\b[77] ), .A4(\b[78] ), .ZN(new_n1338_));
  OAI21_X1   g0952(.A1(new_n1337_), .A2(new_n1338_), .B(new_n1335_), .ZN(new_n1339_));
  INV_X1     g0953(.I(new_n1339_), .ZN(new_n1340_));
  NOR3_X1    g0954(.A1(new_n1337_), .A2(new_n1338_), .A3(new_n1335_), .ZN(new_n1341_));
  OAI21_X1   g0955(.A1(new_n1340_), .A2(new_n1341_), .B(new_n1334_), .ZN(new_n1342_));
  INV_X1     g0956(.I(new_n1341_), .ZN(new_n1343_));
  NAND3_X1   g0957(.A1(new_n1343_), .A2(\a[79] ), .A3(new_n1339_), .ZN(new_n1344_));
  NAND2_X1   g0958(.A1(new_n1342_), .A2(new_n1344_), .ZN(\f[79] ));
  NOR2_X1    g0959(.A1(\a[79] ), .A2(\b[79] ), .ZN(new_n1346_));
  AND2_X2    g0960(.A1(\a[79] ), .A2(\b[79] ), .Z(new_n1347_));
  NOR3_X1    g0961(.A1(new_n1337_), .A2(new_n1347_), .A3(new_n1338_), .ZN(new_n1348_));
  NOR2_X1    g0962(.A1(new_n1348_), .A2(new_n1346_), .ZN(new_n1349_));
  XOR2_X1    g0963(.A1(\a[80] ), .A2(\b[80] ), .Z(new_n1350_));
  NAND2_X1   g0964(.A1(new_n1349_), .A2(new_n1350_), .ZN(new_n1351_));
  INV_X1     g0965(.I(\a[80] ), .ZN(new_n1352_));
  INV_X1     g0966(.I(\b[80] ), .ZN(new_n1353_));
  NOR2_X1    g0967(.A1(new_n1352_), .A2(new_n1353_), .ZN(new_n1354_));
  NOR2_X1    g0968(.A1(\a[80] ), .A2(\b[80] ), .ZN(new_n1355_));
  NOR2_X1    g0969(.A1(new_n1354_), .A2(new_n1355_), .ZN(new_n1356_));
  OAI21_X1   g0970(.A1(new_n1349_), .A2(new_n1356_), .B(new_n1351_), .ZN(\f[80] ));
  NOR3_X1    g0971(.A1(new_n1348_), .A2(new_n1346_), .A3(new_n1354_), .ZN(new_n1358_));
  XOR2_X1    g0972(.A1(\a[81] ), .A2(\b[81] ), .Z(new_n1359_));
  OAI21_X1   g0973(.A1(new_n1358_), .A2(new_n1355_), .B(new_n1359_), .ZN(new_n1360_));
  INV_X1     g0974(.I(new_n1355_), .ZN(new_n1361_));
  INV_X1     g0975(.I(new_n1346_), .ZN(new_n1362_));
  OR4_X2     g0976(.A1(\a[77] ), .A2(\a[78] ), .A3(\b[77] ), .A4(\b[78] ), .Z(new_n1363_));
  NAND2_X1   g0977(.A1(\a[79] ), .A2(\b[79] ), .ZN(new_n1364_));
  NAND3_X1   g0978(.A1(new_n1363_), .A2(new_n1336_), .A3(new_n1364_), .ZN(new_n1365_));
  INV_X1     g0979(.I(new_n1354_), .ZN(new_n1366_));
  NAND3_X1   g0980(.A1(new_n1365_), .A2(new_n1362_), .A3(new_n1366_), .ZN(new_n1367_));
  XNOR2_X1   g0981(.A1(\a[81] ), .A2(\b[81] ), .ZN(new_n1368_));
  NAND3_X1   g0982(.A1(new_n1367_), .A2(new_n1361_), .A3(new_n1368_), .ZN(new_n1369_));
  NAND2_X1   g0983(.A1(new_n1369_), .A2(new_n1360_), .ZN(\f[81] ));
  INV_X1     g0984(.I(\a[82] ), .ZN(new_n1371_));
  INV_X1     g0985(.I(\b[82] ), .ZN(new_n1372_));
  NAND2_X1   g0986(.A1(\a[81] ), .A2(\b[81] ), .ZN(new_n1373_));
  INV_X1     g0987(.I(new_n1373_), .ZN(new_n1374_));
  NOR4_X1    g0988(.A1(\a[80] ), .A2(\a[81] ), .A3(\b[80] ), .A4(\b[81] ), .ZN(new_n1375_));
  OAI21_X1   g0989(.A1(new_n1374_), .A2(new_n1375_), .B(new_n1372_), .ZN(new_n1376_));
  INV_X1     g0990(.I(new_n1376_), .ZN(new_n1377_));
  NOR3_X1    g0991(.A1(new_n1374_), .A2(new_n1375_), .A3(new_n1372_), .ZN(new_n1378_));
  OAI21_X1   g0992(.A1(new_n1377_), .A2(new_n1378_), .B(new_n1371_), .ZN(new_n1379_));
  INV_X1     g0993(.I(new_n1378_), .ZN(new_n1380_));
  NAND3_X1   g0994(.A1(new_n1380_), .A2(\a[82] ), .A3(new_n1376_), .ZN(new_n1381_));
  NAND2_X1   g0995(.A1(new_n1379_), .A2(new_n1381_), .ZN(\f[82] ));
  NOR2_X1    g0996(.A1(\a[82] ), .A2(\b[82] ), .ZN(new_n1383_));
  AND2_X2    g0997(.A1(\a[82] ), .A2(\b[82] ), .Z(new_n1384_));
  NOR3_X1    g0998(.A1(new_n1374_), .A2(new_n1384_), .A3(new_n1375_), .ZN(new_n1385_));
  NOR2_X1    g0999(.A1(new_n1385_), .A2(new_n1383_), .ZN(new_n1386_));
  XOR2_X1    g1000(.A1(\a[83] ), .A2(\b[83] ), .Z(new_n1387_));
  NAND2_X1   g1001(.A1(new_n1386_), .A2(new_n1387_), .ZN(new_n1388_));
  INV_X1     g1002(.I(\a[83] ), .ZN(new_n1389_));
  INV_X1     g1003(.I(\b[83] ), .ZN(new_n1390_));
  NOR2_X1    g1004(.A1(new_n1389_), .A2(new_n1390_), .ZN(new_n1391_));
  NOR2_X1    g1005(.A1(\a[83] ), .A2(\b[83] ), .ZN(new_n1392_));
  NOR2_X1    g1006(.A1(new_n1391_), .A2(new_n1392_), .ZN(new_n1393_));
  OAI21_X1   g1007(.A1(new_n1386_), .A2(new_n1393_), .B(new_n1388_), .ZN(\f[83] ));
  NOR3_X1    g1008(.A1(new_n1385_), .A2(new_n1383_), .A3(new_n1391_), .ZN(new_n1395_));
  XOR2_X1    g1009(.A1(\a[84] ), .A2(\b[84] ), .Z(new_n1396_));
  OAI21_X1   g1010(.A1(new_n1395_), .A2(new_n1392_), .B(new_n1396_), .ZN(new_n1397_));
  INV_X1     g1011(.I(new_n1392_), .ZN(new_n1398_));
  INV_X1     g1012(.I(new_n1383_), .ZN(new_n1399_));
  OR4_X2     g1013(.A1(\a[80] ), .A2(\a[81] ), .A3(\b[80] ), .A4(\b[81] ), .Z(new_n1400_));
  NAND2_X1   g1014(.A1(\a[82] ), .A2(\b[82] ), .ZN(new_n1401_));
  NAND3_X1   g1015(.A1(new_n1400_), .A2(new_n1373_), .A3(new_n1401_), .ZN(new_n1402_));
  INV_X1     g1016(.I(new_n1391_), .ZN(new_n1403_));
  NAND3_X1   g1017(.A1(new_n1402_), .A2(new_n1399_), .A3(new_n1403_), .ZN(new_n1404_));
  XNOR2_X1   g1018(.A1(\a[84] ), .A2(\b[84] ), .ZN(new_n1405_));
  NAND3_X1   g1019(.A1(new_n1404_), .A2(new_n1398_), .A3(new_n1405_), .ZN(new_n1406_));
  NAND2_X1   g1020(.A1(new_n1406_), .A2(new_n1397_), .ZN(\f[84] ));
  INV_X1     g1021(.I(\a[85] ), .ZN(new_n1408_));
  INV_X1     g1022(.I(\b[85] ), .ZN(new_n1409_));
  NAND2_X1   g1023(.A1(\a[84] ), .A2(\b[84] ), .ZN(new_n1410_));
  INV_X1     g1024(.I(new_n1410_), .ZN(new_n1411_));
  NOR4_X1    g1025(.A1(\a[83] ), .A2(\a[84] ), .A3(\b[83] ), .A4(\b[84] ), .ZN(new_n1412_));
  OAI21_X1   g1026(.A1(new_n1411_), .A2(new_n1412_), .B(new_n1409_), .ZN(new_n1413_));
  INV_X1     g1027(.I(new_n1413_), .ZN(new_n1414_));
  NOR3_X1    g1028(.A1(new_n1411_), .A2(new_n1412_), .A3(new_n1409_), .ZN(new_n1415_));
  OAI21_X1   g1029(.A1(new_n1414_), .A2(new_n1415_), .B(new_n1408_), .ZN(new_n1416_));
  INV_X1     g1030(.I(new_n1415_), .ZN(new_n1417_));
  NAND3_X1   g1031(.A1(new_n1417_), .A2(\a[85] ), .A3(new_n1413_), .ZN(new_n1418_));
  NAND2_X1   g1032(.A1(new_n1416_), .A2(new_n1418_), .ZN(\f[85] ));
  NOR2_X1    g1033(.A1(\a[85] ), .A2(\b[85] ), .ZN(new_n1420_));
  AND2_X2    g1034(.A1(\a[85] ), .A2(\b[85] ), .Z(new_n1421_));
  NOR3_X1    g1035(.A1(new_n1411_), .A2(new_n1421_), .A3(new_n1412_), .ZN(new_n1422_));
  NOR2_X1    g1036(.A1(new_n1422_), .A2(new_n1420_), .ZN(new_n1423_));
  XOR2_X1    g1037(.A1(\a[86] ), .A2(\b[86] ), .Z(new_n1424_));
  NAND2_X1   g1038(.A1(new_n1423_), .A2(new_n1424_), .ZN(new_n1425_));
  INV_X1     g1039(.I(\a[86] ), .ZN(new_n1426_));
  INV_X1     g1040(.I(\b[86] ), .ZN(new_n1427_));
  NOR2_X1    g1041(.A1(new_n1426_), .A2(new_n1427_), .ZN(new_n1428_));
  NOR2_X1    g1042(.A1(\a[86] ), .A2(\b[86] ), .ZN(new_n1429_));
  NOR2_X1    g1043(.A1(new_n1428_), .A2(new_n1429_), .ZN(new_n1430_));
  OAI21_X1   g1044(.A1(new_n1423_), .A2(new_n1430_), .B(new_n1425_), .ZN(\f[86] ));
  NOR3_X1    g1045(.A1(new_n1422_), .A2(new_n1420_), .A3(new_n1428_), .ZN(new_n1432_));
  XOR2_X1    g1046(.A1(\a[87] ), .A2(\b[87] ), .Z(new_n1433_));
  OAI21_X1   g1047(.A1(new_n1432_), .A2(new_n1429_), .B(new_n1433_), .ZN(new_n1434_));
  INV_X1     g1048(.I(new_n1429_), .ZN(new_n1435_));
  INV_X1     g1049(.I(new_n1420_), .ZN(new_n1436_));
  OR4_X2     g1050(.A1(\a[83] ), .A2(\a[84] ), .A3(\b[83] ), .A4(\b[84] ), .Z(new_n1437_));
  NAND2_X1   g1051(.A1(\a[85] ), .A2(\b[85] ), .ZN(new_n1438_));
  NAND3_X1   g1052(.A1(new_n1437_), .A2(new_n1410_), .A3(new_n1438_), .ZN(new_n1439_));
  INV_X1     g1053(.I(new_n1428_), .ZN(new_n1440_));
  NAND3_X1   g1054(.A1(new_n1439_), .A2(new_n1436_), .A3(new_n1440_), .ZN(new_n1441_));
  XNOR2_X1   g1055(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n1442_));
  NAND3_X1   g1056(.A1(new_n1441_), .A2(new_n1435_), .A3(new_n1442_), .ZN(new_n1443_));
  NAND2_X1   g1057(.A1(new_n1443_), .A2(new_n1434_), .ZN(\f[87] ));
  INV_X1     g1058(.I(\a[88] ), .ZN(new_n1445_));
  INV_X1     g1059(.I(\b[88] ), .ZN(new_n1446_));
  NAND2_X1   g1060(.A1(\a[87] ), .A2(\b[87] ), .ZN(new_n1447_));
  INV_X1     g1061(.I(new_n1447_), .ZN(new_n1448_));
  NOR4_X1    g1062(.A1(\a[86] ), .A2(\a[87] ), .A3(\b[86] ), .A4(\b[87] ), .ZN(new_n1449_));
  OAI21_X1   g1063(.A1(new_n1448_), .A2(new_n1449_), .B(new_n1446_), .ZN(new_n1450_));
  INV_X1     g1064(.I(new_n1450_), .ZN(new_n1451_));
  NOR3_X1    g1065(.A1(new_n1448_), .A2(new_n1449_), .A3(new_n1446_), .ZN(new_n1452_));
  OAI21_X1   g1066(.A1(new_n1451_), .A2(new_n1452_), .B(new_n1445_), .ZN(new_n1453_));
  INV_X1     g1067(.I(new_n1452_), .ZN(new_n1454_));
  NAND3_X1   g1068(.A1(new_n1454_), .A2(\a[88] ), .A3(new_n1450_), .ZN(new_n1455_));
  NAND2_X1   g1069(.A1(new_n1453_), .A2(new_n1455_), .ZN(\f[88] ));
  NOR2_X1    g1070(.A1(\a[88] ), .A2(\b[88] ), .ZN(new_n1457_));
  AND2_X2    g1071(.A1(\a[88] ), .A2(\b[88] ), .Z(new_n1458_));
  NOR3_X1    g1072(.A1(new_n1448_), .A2(new_n1458_), .A3(new_n1449_), .ZN(new_n1459_));
  NOR2_X1    g1073(.A1(new_n1459_), .A2(new_n1457_), .ZN(new_n1460_));
  XOR2_X1    g1074(.A1(\a[89] ), .A2(\b[89] ), .Z(new_n1461_));
  NAND2_X1   g1075(.A1(new_n1460_), .A2(new_n1461_), .ZN(new_n1462_));
  INV_X1     g1076(.I(\a[89] ), .ZN(new_n1463_));
  INV_X1     g1077(.I(\b[89] ), .ZN(new_n1464_));
  NOR2_X1    g1078(.A1(new_n1463_), .A2(new_n1464_), .ZN(new_n1465_));
  NOR2_X1    g1079(.A1(\a[89] ), .A2(\b[89] ), .ZN(new_n1466_));
  NOR2_X1    g1080(.A1(new_n1465_), .A2(new_n1466_), .ZN(new_n1467_));
  OAI21_X1   g1081(.A1(new_n1460_), .A2(new_n1467_), .B(new_n1462_), .ZN(\f[89] ));
  NOR3_X1    g1082(.A1(new_n1459_), .A2(new_n1457_), .A3(new_n1465_), .ZN(new_n1469_));
  XOR2_X1    g1083(.A1(\a[90] ), .A2(\b[90] ), .Z(new_n1470_));
  OAI21_X1   g1084(.A1(new_n1469_), .A2(new_n1466_), .B(new_n1470_), .ZN(new_n1471_));
  INV_X1     g1085(.I(new_n1466_), .ZN(new_n1472_));
  INV_X1     g1086(.I(new_n1457_), .ZN(new_n1473_));
  OR4_X2     g1087(.A1(\a[86] ), .A2(\a[87] ), .A3(\b[86] ), .A4(\b[87] ), .Z(new_n1474_));
  NAND2_X1   g1088(.A1(\a[88] ), .A2(\b[88] ), .ZN(new_n1475_));
  NAND3_X1   g1089(.A1(new_n1474_), .A2(new_n1447_), .A3(new_n1475_), .ZN(new_n1476_));
  INV_X1     g1090(.I(new_n1465_), .ZN(new_n1477_));
  NAND3_X1   g1091(.A1(new_n1476_), .A2(new_n1473_), .A3(new_n1477_), .ZN(new_n1478_));
  XNOR2_X1   g1092(.A1(\a[90] ), .A2(\b[90] ), .ZN(new_n1479_));
  NAND3_X1   g1093(.A1(new_n1478_), .A2(new_n1472_), .A3(new_n1479_), .ZN(new_n1480_));
  NAND2_X1   g1094(.A1(new_n1480_), .A2(new_n1471_), .ZN(\f[90] ));
  INV_X1     g1095(.I(\a[91] ), .ZN(new_n1482_));
  INV_X1     g1096(.I(\b[91] ), .ZN(new_n1483_));
  NAND2_X1   g1097(.A1(\a[90] ), .A2(\b[90] ), .ZN(new_n1484_));
  INV_X1     g1098(.I(new_n1484_), .ZN(new_n1485_));
  NOR4_X1    g1099(.A1(\a[89] ), .A2(\a[90] ), .A3(\b[89] ), .A4(\b[90] ), .ZN(new_n1486_));
  OAI21_X1   g1100(.A1(new_n1485_), .A2(new_n1486_), .B(new_n1483_), .ZN(new_n1487_));
  INV_X1     g1101(.I(new_n1487_), .ZN(new_n1488_));
  NOR3_X1    g1102(.A1(new_n1485_), .A2(new_n1486_), .A3(new_n1483_), .ZN(new_n1489_));
  OAI21_X1   g1103(.A1(new_n1488_), .A2(new_n1489_), .B(new_n1482_), .ZN(new_n1490_));
  INV_X1     g1104(.I(new_n1489_), .ZN(new_n1491_));
  NAND3_X1   g1105(.A1(new_n1491_), .A2(\a[91] ), .A3(new_n1487_), .ZN(new_n1492_));
  NAND2_X1   g1106(.A1(new_n1490_), .A2(new_n1492_), .ZN(\f[91] ));
  NOR2_X1    g1107(.A1(\a[91] ), .A2(\b[91] ), .ZN(new_n1494_));
  AND2_X2    g1108(.A1(\a[91] ), .A2(\b[91] ), .Z(new_n1495_));
  NOR3_X1    g1109(.A1(new_n1485_), .A2(new_n1495_), .A3(new_n1486_), .ZN(new_n1496_));
  NOR2_X1    g1110(.A1(new_n1496_), .A2(new_n1494_), .ZN(new_n1497_));
  XOR2_X1    g1111(.A1(\a[92] ), .A2(\b[92] ), .Z(new_n1498_));
  NAND2_X1   g1112(.A1(new_n1497_), .A2(new_n1498_), .ZN(new_n1499_));
  INV_X1     g1113(.I(\a[92] ), .ZN(new_n1500_));
  INV_X1     g1114(.I(\b[92] ), .ZN(new_n1501_));
  NOR2_X1    g1115(.A1(new_n1500_), .A2(new_n1501_), .ZN(new_n1502_));
  NOR2_X1    g1116(.A1(\a[92] ), .A2(\b[92] ), .ZN(new_n1503_));
  NOR2_X1    g1117(.A1(new_n1502_), .A2(new_n1503_), .ZN(new_n1504_));
  OAI21_X1   g1118(.A1(new_n1497_), .A2(new_n1504_), .B(new_n1499_), .ZN(\f[92] ));
  NOR3_X1    g1119(.A1(new_n1496_), .A2(new_n1494_), .A3(new_n1502_), .ZN(new_n1506_));
  XOR2_X1    g1120(.A1(\a[93] ), .A2(\b[93] ), .Z(new_n1507_));
  OAI21_X1   g1121(.A1(new_n1506_), .A2(new_n1503_), .B(new_n1507_), .ZN(new_n1508_));
  INV_X1     g1122(.I(new_n1503_), .ZN(new_n1509_));
  INV_X1     g1123(.I(new_n1494_), .ZN(new_n1510_));
  OR4_X2     g1124(.A1(\a[89] ), .A2(\a[90] ), .A3(\b[89] ), .A4(\b[90] ), .Z(new_n1511_));
  NAND2_X1   g1125(.A1(\a[91] ), .A2(\b[91] ), .ZN(new_n1512_));
  NAND3_X1   g1126(.A1(new_n1511_), .A2(new_n1484_), .A3(new_n1512_), .ZN(new_n1513_));
  INV_X1     g1127(.I(new_n1502_), .ZN(new_n1514_));
  NAND3_X1   g1128(.A1(new_n1513_), .A2(new_n1510_), .A3(new_n1514_), .ZN(new_n1515_));
  XNOR2_X1   g1129(.A1(\a[93] ), .A2(\b[93] ), .ZN(new_n1516_));
  NAND3_X1   g1130(.A1(new_n1515_), .A2(new_n1509_), .A3(new_n1516_), .ZN(new_n1517_));
  NAND2_X1   g1131(.A1(new_n1517_), .A2(new_n1508_), .ZN(\f[93] ));
  INV_X1     g1132(.I(\a[94] ), .ZN(new_n1519_));
  INV_X1     g1133(.I(\b[94] ), .ZN(new_n1520_));
  NAND2_X1   g1134(.A1(\a[93] ), .A2(\b[93] ), .ZN(new_n1521_));
  INV_X1     g1135(.I(new_n1521_), .ZN(new_n1522_));
  NOR4_X1    g1136(.A1(\a[92] ), .A2(\a[93] ), .A3(\b[92] ), .A4(\b[93] ), .ZN(new_n1523_));
  OAI21_X1   g1137(.A1(new_n1522_), .A2(new_n1523_), .B(new_n1520_), .ZN(new_n1524_));
  INV_X1     g1138(.I(new_n1524_), .ZN(new_n1525_));
  NOR3_X1    g1139(.A1(new_n1522_), .A2(new_n1523_), .A3(new_n1520_), .ZN(new_n1526_));
  OAI21_X1   g1140(.A1(new_n1525_), .A2(new_n1526_), .B(new_n1519_), .ZN(new_n1527_));
  INV_X1     g1141(.I(new_n1526_), .ZN(new_n1528_));
  NAND3_X1   g1142(.A1(new_n1528_), .A2(\a[94] ), .A3(new_n1524_), .ZN(new_n1529_));
  NAND2_X1   g1143(.A1(new_n1527_), .A2(new_n1529_), .ZN(\f[94] ));
  NOR2_X1    g1144(.A1(\a[94] ), .A2(\b[94] ), .ZN(new_n1531_));
  AND2_X2    g1145(.A1(\a[94] ), .A2(\b[94] ), .Z(new_n1532_));
  NOR3_X1    g1146(.A1(new_n1522_), .A2(new_n1532_), .A3(new_n1523_), .ZN(new_n1533_));
  NOR2_X1    g1147(.A1(new_n1533_), .A2(new_n1531_), .ZN(new_n1534_));
  XOR2_X1    g1148(.A1(\a[95] ), .A2(\b[95] ), .Z(new_n1535_));
  NAND2_X1   g1149(.A1(new_n1534_), .A2(new_n1535_), .ZN(new_n1536_));
  INV_X1     g1150(.I(\a[95] ), .ZN(new_n1537_));
  INV_X1     g1151(.I(\b[95] ), .ZN(new_n1538_));
  NOR2_X1    g1152(.A1(new_n1537_), .A2(new_n1538_), .ZN(new_n1539_));
  NOR2_X1    g1153(.A1(\a[95] ), .A2(\b[95] ), .ZN(new_n1540_));
  NOR2_X1    g1154(.A1(new_n1539_), .A2(new_n1540_), .ZN(new_n1541_));
  OAI21_X1   g1155(.A1(new_n1534_), .A2(new_n1541_), .B(new_n1536_), .ZN(\f[95] ));
  NOR3_X1    g1156(.A1(new_n1533_), .A2(new_n1531_), .A3(new_n1539_), .ZN(new_n1543_));
  XOR2_X1    g1157(.A1(\a[96] ), .A2(\b[96] ), .Z(new_n1544_));
  OAI21_X1   g1158(.A1(new_n1543_), .A2(new_n1540_), .B(new_n1544_), .ZN(new_n1545_));
  INV_X1     g1159(.I(new_n1540_), .ZN(new_n1546_));
  INV_X1     g1160(.I(new_n1531_), .ZN(new_n1547_));
  OR4_X2     g1161(.A1(\a[92] ), .A2(\a[93] ), .A3(\b[92] ), .A4(\b[93] ), .Z(new_n1548_));
  NAND2_X1   g1162(.A1(\a[94] ), .A2(\b[94] ), .ZN(new_n1549_));
  NAND3_X1   g1163(.A1(new_n1548_), .A2(new_n1521_), .A3(new_n1549_), .ZN(new_n1550_));
  INV_X1     g1164(.I(new_n1539_), .ZN(new_n1551_));
  NAND3_X1   g1165(.A1(new_n1550_), .A2(new_n1547_), .A3(new_n1551_), .ZN(new_n1552_));
  XNOR2_X1   g1166(.A1(\a[96] ), .A2(\b[96] ), .ZN(new_n1553_));
  NAND3_X1   g1167(.A1(new_n1552_), .A2(new_n1546_), .A3(new_n1553_), .ZN(new_n1554_));
  NAND2_X1   g1168(.A1(new_n1554_), .A2(new_n1545_), .ZN(\f[96] ));
  INV_X1     g1169(.I(\a[97] ), .ZN(new_n1556_));
  INV_X1     g1170(.I(\b[97] ), .ZN(new_n1557_));
  NAND2_X1   g1171(.A1(\a[96] ), .A2(\b[96] ), .ZN(new_n1558_));
  INV_X1     g1172(.I(new_n1558_), .ZN(new_n1559_));
  NOR4_X1    g1173(.A1(\a[95] ), .A2(\a[96] ), .A3(\b[95] ), .A4(\b[96] ), .ZN(new_n1560_));
  OAI21_X1   g1174(.A1(new_n1559_), .A2(new_n1560_), .B(new_n1557_), .ZN(new_n1561_));
  INV_X1     g1175(.I(new_n1561_), .ZN(new_n1562_));
  NOR3_X1    g1176(.A1(new_n1559_), .A2(new_n1560_), .A3(new_n1557_), .ZN(new_n1563_));
  OAI21_X1   g1177(.A1(new_n1562_), .A2(new_n1563_), .B(new_n1556_), .ZN(new_n1564_));
  INV_X1     g1178(.I(new_n1563_), .ZN(new_n1565_));
  NAND3_X1   g1179(.A1(new_n1565_), .A2(\a[97] ), .A3(new_n1561_), .ZN(new_n1566_));
  NAND2_X1   g1180(.A1(new_n1564_), .A2(new_n1566_), .ZN(\f[97] ));
  NOR2_X1    g1181(.A1(\a[97] ), .A2(\b[97] ), .ZN(new_n1568_));
  AND2_X2    g1182(.A1(\a[97] ), .A2(\b[97] ), .Z(new_n1569_));
  NOR3_X1    g1183(.A1(new_n1559_), .A2(new_n1569_), .A3(new_n1560_), .ZN(new_n1570_));
  NOR2_X1    g1184(.A1(new_n1570_), .A2(new_n1568_), .ZN(new_n1571_));
  XOR2_X1    g1185(.A1(\a[98] ), .A2(\b[98] ), .Z(new_n1572_));
  NAND2_X1   g1186(.A1(new_n1571_), .A2(new_n1572_), .ZN(new_n1573_));
  INV_X1     g1187(.I(\a[98] ), .ZN(new_n1574_));
  INV_X1     g1188(.I(\b[98] ), .ZN(new_n1575_));
  NOR2_X1    g1189(.A1(new_n1574_), .A2(new_n1575_), .ZN(new_n1576_));
  NOR2_X1    g1190(.A1(\a[98] ), .A2(\b[98] ), .ZN(new_n1577_));
  NOR2_X1    g1191(.A1(new_n1576_), .A2(new_n1577_), .ZN(new_n1578_));
  OAI21_X1   g1192(.A1(new_n1571_), .A2(new_n1578_), .B(new_n1573_), .ZN(\f[98] ));
  NOR3_X1    g1193(.A1(new_n1570_), .A2(new_n1568_), .A3(new_n1576_), .ZN(new_n1580_));
  XOR2_X1    g1194(.A1(\a[99] ), .A2(\b[99] ), .Z(new_n1581_));
  OAI21_X1   g1195(.A1(new_n1580_), .A2(new_n1577_), .B(new_n1581_), .ZN(new_n1582_));
  INV_X1     g1196(.I(new_n1577_), .ZN(new_n1583_));
  INV_X1     g1197(.I(new_n1568_), .ZN(new_n1584_));
  OR4_X2     g1198(.A1(\a[95] ), .A2(\a[96] ), .A3(\b[95] ), .A4(\b[96] ), .Z(new_n1585_));
  NAND2_X1   g1199(.A1(\a[97] ), .A2(\b[97] ), .ZN(new_n1586_));
  NAND3_X1   g1200(.A1(new_n1585_), .A2(new_n1558_), .A3(new_n1586_), .ZN(new_n1587_));
  INV_X1     g1201(.I(new_n1576_), .ZN(new_n1588_));
  NAND3_X1   g1202(.A1(new_n1587_), .A2(new_n1584_), .A3(new_n1588_), .ZN(new_n1589_));
  XNOR2_X1   g1203(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n1590_));
  NAND3_X1   g1204(.A1(new_n1589_), .A2(new_n1583_), .A3(new_n1590_), .ZN(new_n1591_));
  NAND2_X1   g1205(.A1(new_n1591_), .A2(new_n1582_), .ZN(\f[99] ));
  INV_X1     g1206(.I(\a[100] ), .ZN(new_n1593_));
  INV_X1     g1207(.I(\b[100] ), .ZN(new_n1594_));
  NAND2_X1   g1208(.A1(\a[99] ), .A2(\b[99] ), .ZN(new_n1595_));
  INV_X1     g1209(.I(new_n1595_), .ZN(new_n1596_));
  NOR4_X1    g1210(.A1(\a[98] ), .A2(\a[99] ), .A3(\b[98] ), .A4(\b[99] ), .ZN(new_n1597_));
  OAI21_X1   g1211(.A1(new_n1596_), .A2(new_n1597_), .B(new_n1594_), .ZN(new_n1598_));
  INV_X1     g1212(.I(new_n1598_), .ZN(new_n1599_));
  NOR3_X1    g1213(.A1(new_n1596_), .A2(new_n1597_), .A3(new_n1594_), .ZN(new_n1600_));
  OAI21_X1   g1214(.A1(new_n1599_), .A2(new_n1600_), .B(new_n1593_), .ZN(new_n1601_));
  INV_X1     g1215(.I(new_n1600_), .ZN(new_n1602_));
  NAND3_X1   g1216(.A1(new_n1602_), .A2(\a[100] ), .A3(new_n1598_), .ZN(new_n1603_));
  NAND2_X1   g1217(.A1(new_n1601_), .A2(new_n1603_), .ZN(\f[100] ));
  NOR2_X1    g1218(.A1(\a[100] ), .A2(\b[100] ), .ZN(new_n1605_));
  AND2_X2    g1219(.A1(\a[100] ), .A2(\b[100] ), .Z(new_n1606_));
  NOR3_X1    g1220(.A1(new_n1596_), .A2(new_n1606_), .A3(new_n1597_), .ZN(new_n1607_));
  NOR2_X1    g1221(.A1(new_n1607_), .A2(new_n1605_), .ZN(new_n1608_));
  XOR2_X1    g1222(.A1(\a[101] ), .A2(\b[101] ), .Z(new_n1609_));
  NAND2_X1   g1223(.A1(new_n1608_), .A2(new_n1609_), .ZN(new_n1610_));
  INV_X1     g1224(.I(\a[101] ), .ZN(new_n1611_));
  INV_X1     g1225(.I(\b[101] ), .ZN(new_n1612_));
  NOR2_X1    g1226(.A1(new_n1611_), .A2(new_n1612_), .ZN(new_n1613_));
  NOR2_X1    g1227(.A1(\a[101] ), .A2(\b[101] ), .ZN(new_n1614_));
  NOR2_X1    g1228(.A1(new_n1613_), .A2(new_n1614_), .ZN(new_n1615_));
  OAI21_X1   g1229(.A1(new_n1608_), .A2(new_n1615_), .B(new_n1610_), .ZN(\f[101] ));
  NOR3_X1    g1230(.A1(new_n1607_), .A2(new_n1605_), .A3(new_n1613_), .ZN(new_n1617_));
  XOR2_X1    g1231(.A1(\a[102] ), .A2(\b[102] ), .Z(new_n1618_));
  OAI21_X1   g1232(.A1(new_n1617_), .A2(new_n1614_), .B(new_n1618_), .ZN(new_n1619_));
  INV_X1     g1233(.I(new_n1614_), .ZN(new_n1620_));
  INV_X1     g1234(.I(new_n1605_), .ZN(new_n1621_));
  OR4_X2     g1235(.A1(\a[98] ), .A2(\a[99] ), .A3(\b[98] ), .A4(\b[99] ), .Z(new_n1622_));
  NAND2_X1   g1236(.A1(\a[100] ), .A2(\b[100] ), .ZN(new_n1623_));
  NAND3_X1   g1237(.A1(new_n1622_), .A2(new_n1595_), .A3(new_n1623_), .ZN(new_n1624_));
  INV_X1     g1238(.I(new_n1613_), .ZN(new_n1625_));
  NAND3_X1   g1239(.A1(new_n1624_), .A2(new_n1621_), .A3(new_n1625_), .ZN(new_n1626_));
  XNOR2_X1   g1240(.A1(\a[102] ), .A2(\b[102] ), .ZN(new_n1627_));
  NAND3_X1   g1241(.A1(new_n1626_), .A2(new_n1620_), .A3(new_n1627_), .ZN(new_n1628_));
  NAND2_X1   g1242(.A1(new_n1628_), .A2(new_n1619_), .ZN(\f[102] ));
  INV_X1     g1243(.I(\a[103] ), .ZN(new_n1630_));
  INV_X1     g1244(.I(\b[103] ), .ZN(new_n1631_));
  NAND2_X1   g1245(.A1(\a[102] ), .A2(\b[102] ), .ZN(new_n1632_));
  INV_X1     g1246(.I(new_n1632_), .ZN(new_n1633_));
  NOR4_X1    g1247(.A1(\a[101] ), .A2(\a[102] ), .A3(\b[101] ), .A4(\b[102] ), .ZN(new_n1634_));
  OAI21_X1   g1248(.A1(new_n1633_), .A2(new_n1634_), .B(new_n1631_), .ZN(new_n1635_));
  INV_X1     g1249(.I(new_n1635_), .ZN(new_n1636_));
  NOR3_X1    g1250(.A1(new_n1633_), .A2(new_n1634_), .A3(new_n1631_), .ZN(new_n1637_));
  OAI21_X1   g1251(.A1(new_n1636_), .A2(new_n1637_), .B(new_n1630_), .ZN(new_n1638_));
  INV_X1     g1252(.I(new_n1637_), .ZN(new_n1639_));
  NAND3_X1   g1253(.A1(new_n1639_), .A2(\a[103] ), .A3(new_n1635_), .ZN(new_n1640_));
  NAND2_X1   g1254(.A1(new_n1638_), .A2(new_n1640_), .ZN(\f[103] ));
  NOR2_X1    g1255(.A1(\a[103] ), .A2(\b[103] ), .ZN(new_n1642_));
  AND2_X2    g1256(.A1(\a[103] ), .A2(\b[103] ), .Z(new_n1643_));
  NOR3_X1    g1257(.A1(new_n1633_), .A2(new_n1643_), .A3(new_n1634_), .ZN(new_n1644_));
  NOR2_X1    g1258(.A1(new_n1644_), .A2(new_n1642_), .ZN(new_n1645_));
  XOR2_X1    g1259(.A1(\a[104] ), .A2(\b[104] ), .Z(new_n1646_));
  NAND2_X1   g1260(.A1(new_n1645_), .A2(new_n1646_), .ZN(new_n1647_));
  INV_X1     g1261(.I(\a[104] ), .ZN(new_n1648_));
  INV_X1     g1262(.I(\b[104] ), .ZN(new_n1649_));
  NOR2_X1    g1263(.A1(new_n1648_), .A2(new_n1649_), .ZN(new_n1650_));
  NOR2_X1    g1264(.A1(\a[104] ), .A2(\b[104] ), .ZN(new_n1651_));
  NOR2_X1    g1265(.A1(new_n1650_), .A2(new_n1651_), .ZN(new_n1652_));
  OAI21_X1   g1266(.A1(new_n1645_), .A2(new_n1652_), .B(new_n1647_), .ZN(\f[104] ));
  NOR3_X1    g1267(.A1(new_n1644_), .A2(new_n1642_), .A3(new_n1650_), .ZN(new_n1654_));
  XOR2_X1    g1268(.A1(\a[105] ), .A2(\b[105] ), .Z(new_n1655_));
  OAI21_X1   g1269(.A1(new_n1654_), .A2(new_n1651_), .B(new_n1655_), .ZN(new_n1656_));
  INV_X1     g1270(.I(new_n1651_), .ZN(new_n1657_));
  INV_X1     g1271(.I(new_n1642_), .ZN(new_n1658_));
  OR4_X2     g1272(.A1(\a[101] ), .A2(\a[102] ), .A3(\b[101] ), .A4(\b[102] ), .Z(new_n1659_));
  NAND2_X1   g1273(.A1(\a[103] ), .A2(\b[103] ), .ZN(new_n1660_));
  NAND3_X1   g1274(.A1(new_n1659_), .A2(new_n1632_), .A3(new_n1660_), .ZN(new_n1661_));
  INV_X1     g1275(.I(new_n1650_), .ZN(new_n1662_));
  NAND3_X1   g1276(.A1(new_n1661_), .A2(new_n1658_), .A3(new_n1662_), .ZN(new_n1663_));
  XNOR2_X1   g1277(.A1(\a[105] ), .A2(\b[105] ), .ZN(new_n1664_));
  NAND3_X1   g1278(.A1(new_n1663_), .A2(new_n1657_), .A3(new_n1664_), .ZN(new_n1665_));
  NAND2_X1   g1279(.A1(new_n1665_), .A2(new_n1656_), .ZN(\f[105] ));
  INV_X1     g1280(.I(\a[106] ), .ZN(new_n1667_));
  INV_X1     g1281(.I(\b[106] ), .ZN(new_n1668_));
  NAND2_X1   g1282(.A1(\a[105] ), .A2(\b[105] ), .ZN(new_n1669_));
  INV_X1     g1283(.I(new_n1669_), .ZN(new_n1670_));
  NOR4_X1    g1284(.A1(\a[104] ), .A2(\a[105] ), .A3(\b[104] ), .A4(\b[105] ), .ZN(new_n1671_));
  OAI21_X1   g1285(.A1(new_n1670_), .A2(new_n1671_), .B(new_n1668_), .ZN(new_n1672_));
  INV_X1     g1286(.I(new_n1672_), .ZN(new_n1673_));
  NOR3_X1    g1287(.A1(new_n1670_), .A2(new_n1671_), .A3(new_n1668_), .ZN(new_n1674_));
  OAI21_X1   g1288(.A1(new_n1673_), .A2(new_n1674_), .B(new_n1667_), .ZN(new_n1675_));
  INV_X1     g1289(.I(new_n1674_), .ZN(new_n1676_));
  NAND3_X1   g1290(.A1(new_n1676_), .A2(\a[106] ), .A3(new_n1672_), .ZN(new_n1677_));
  NAND2_X1   g1291(.A1(new_n1675_), .A2(new_n1677_), .ZN(\f[106] ));
  NOR2_X1    g1292(.A1(\a[106] ), .A2(\b[106] ), .ZN(new_n1679_));
  AND2_X2    g1293(.A1(\a[106] ), .A2(\b[106] ), .Z(new_n1680_));
  NOR3_X1    g1294(.A1(new_n1670_), .A2(new_n1680_), .A3(new_n1671_), .ZN(new_n1681_));
  NOR2_X1    g1295(.A1(new_n1681_), .A2(new_n1679_), .ZN(new_n1682_));
  XOR2_X1    g1296(.A1(\a[107] ), .A2(\b[107] ), .Z(new_n1683_));
  NAND2_X1   g1297(.A1(new_n1682_), .A2(new_n1683_), .ZN(new_n1684_));
  INV_X1     g1298(.I(\a[107] ), .ZN(new_n1685_));
  INV_X1     g1299(.I(\b[107] ), .ZN(new_n1686_));
  NOR2_X1    g1300(.A1(new_n1685_), .A2(new_n1686_), .ZN(new_n1687_));
  NOR2_X1    g1301(.A1(\a[107] ), .A2(\b[107] ), .ZN(new_n1688_));
  NOR2_X1    g1302(.A1(new_n1687_), .A2(new_n1688_), .ZN(new_n1689_));
  OAI21_X1   g1303(.A1(new_n1682_), .A2(new_n1689_), .B(new_n1684_), .ZN(\f[107] ));
  NOR3_X1    g1304(.A1(new_n1681_), .A2(new_n1679_), .A3(new_n1687_), .ZN(new_n1691_));
  XOR2_X1    g1305(.A1(\a[108] ), .A2(\b[108] ), .Z(new_n1692_));
  OAI21_X1   g1306(.A1(new_n1691_), .A2(new_n1688_), .B(new_n1692_), .ZN(new_n1693_));
  INV_X1     g1307(.I(new_n1688_), .ZN(new_n1694_));
  INV_X1     g1308(.I(new_n1679_), .ZN(new_n1695_));
  OR4_X2     g1309(.A1(\a[104] ), .A2(\a[105] ), .A3(\b[104] ), .A4(\b[105] ), .Z(new_n1696_));
  NAND2_X1   g1310(.A1(\a[106] ), .A2(\b[106] ), .ZN(new_n1697_));
  NAND3_X1   g1311(.A1(new_n1696_), .A2(new_n1669_), .A3(new_n1697_), .ZN(new_n1698_));
  INV_X1     g1312(.I(new_n1687_), .ZN(new_n1699_));
  NAND3_X1   g1313(.A1(new_n1698_), .A2(new_n1695_), .A3(new_n1699_), .ZN(new_n1700_));
  XNOR2_X1   g1314(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1701_));
  NAND3_X1   g1315(.A1(new_n1700_), .A2(new_n1694_), .A3(new_n1701_), .ZN(new_n1702_));
  NAND2_X1   g1316(.A1(new_n1702_), .A2(new_n1693_), .ZN(\f[108] ));
  INV_X1     g1317(.I(\a[109] ), .ZN(new_n1704_));
  INV_X1     g1318(.I(\b[109] ), .ZN(new_n1705_));
  NAND2_X1   g1319(.A1(\a[108] ), .A2(\b[108] ), .ZN(new_n1706_));
  INV_X1     g1320(.I(new_n1706_), .ZN(new_n1707_));
  NOR4_X1    g1321(.A1(\a[107] ), .A2(\a[108] ), .A3(\b[107] ), .A4(\b[108] ), .ZN(new_n1708_));
  OAI21_X1   g1322(.A1(new_n1707_), .A2(new_n1708_), .B(new_n1705_), .ZN(new_n1709_));
  INV_X1     g1323(.I(new_n1709_), .ZN(new_n1710_));
  NOR3_X1    g1324(.A1(new_n1707_), .A2(new_n1708_), .A3(new_n1705_), .ZN(new_n1711_));
  OAI21_X1   g1325(.A1(new_n1710_), .A2(new_n1711_), .B(new_n1704_), .ZN(new_n1712_));
  INV_X1     g1326(.I(new_n1711_), .ZN(new_n1713_));
  NAND3_X1   g1327(.A1(new_n1713_), .A2(\a[109] ), .A3(new_n1709_), .ZN(new_n1714_));
  NAND2_X1   g1328(.A1(new_n1712_), .A2(new_n1714_), .ZN(\f[109] ));
  NOR2_X1    g1329(.A1(\a[109] ), .A2(\b[109] ), .ZN(new_n1716_));
  AND2_X2    g1330(.A1(\a[109] ), .A2(\b[109] ), .Z(new_n1717_));
  NOR3_X1    g1331(.A1(new_n1707_), .A2(new_n1717_), .A3(new_n1708_), .ZN(new_n1718_));
  NOR2_X1    g1332(.A1(new_n1718_), .A2(new_n1716_), .ZN(new_n1719_));
  XOR2_X1    g1333(.A1(\a[110] ), .A2(\b[110] ), .Z(new_n1720_));
  NAND2_X1   g1334(.A1(new_n1719_), .A2(new_n1720_), .ZN(new_n1721_));
  INV_X1     g1335(.I(\a[110] ), .ZN(new_n1722_));
  INV_X1     g1336(.I(\b[110] ), .ZN(new_n1723_));
  NOR2_X1    g1337(.A1(new_n1722_), .A2(new_n1723_), .ZN(new_n1724_));
  NOR2_X1    g1338(.A1(\a[110] ), .A2(\b[110] ), .ZN(new_n1725_));
  NOR2_X1    g1339(.A1(new_n1724_), .A2(new_n1725_), .ZN(new_n1726_));
  OAI21_X1   g1340(.A1(new_n1719_), .A2(new_n1726_), .B(new_n1721_), .ZN(\f[110] ));
  NOR3_X1    g1341(.A1(new_n1718_), .A2(new_n1716_), .A3(new_n1724_), .ZN(new_n1728_));
  XOR2_X1    g1342(.A1(\a[111] ), .A2(\b[111] ), .Z(new_n1729_));
  OAI21_X1   g1343(.A1(new_n1728_), .A2(new_n1725_), .B(new_n1729_), .ZN(new_n1730_));
  INV_X1     g1344(.I(new_n1725_), .ZN(new_n1731_));
  INV_X1     g1345(.I(new_n1716_), .ZN(new_n1732_));
  OR4_X2     g1346(.A1(\a[107] ), .A2(\a[108] ), .A3(\b[107] ), .A4(\b[108] ), .Z(new_n1733_));
  NAND2_X1   g1347(.A1(\a[109] ), .A2(\b[109] ), .ZN(new_n1734_));
  NAND3_X1   g1348(.A1(new_n1733_), .A2(new_n1706_), .A3(new_n1734_), .ZN(new_n1735_));
  INV_X1     g1349(.I(new_n1724_), .ZN(new_n1736_));
  NAND3_X1   g1350(.A1(new_n1735_), .A2(new_n1732_), .A3(new_n1736_), .ZN(new_n1737_));
  XNOR2_X1   g1351(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1738_));
  NAND3_X1   g1352(.A1(new_n1737_), .A2(new_n1731_), .A3(new_n1738_), .ZN(new_n1739_));
  NAND2_X1   g1353(.A1(new_n1739_), .A2(new_n1730_), .ZN(\f[111] ));
  INV_X1     g1354(.I(\a[112] ), .ZN(new_n1741_));
  INV_X1     g1355(.I(\b[112] ), .ZN(new_n1742_));
  NAND2_X1   g1356(.A1(\a[111] ), .A2(\b[111] ), .ZN(new_n1743_));
  INV_X1     g1357(.I(new_n1743_), .ZN(new_n1744_));
  NOR4_X1    g1358(.A1(\a[110] ), .A2(\a[111] ), .A3(\b[110] ), .A4(\b[111] ), .ZN(new_n1745_));
  OAI21_X1   g1359(.A1(new_n1744_), .A2(new_n1745_), .B(new_n1742_), .ZN(new_n1746_));
  INV_X1     g1360(.I(new_n1746_), .ZN(new_n1747_));
  NOR3_X1    g1361(.A1(new_n1744_), .A2(new_n1745_), .A3(new_n1742_), .ZN(new_n1748_));
  OAI21_X1   g1362(.A1(new_n1747_), .A2(new_n1748_), .B(new_n1741_), .ZN(new_n1749_));
  INV_X1     g1363(.I(new_n1748_), .ZN(new_n1750_));
  NAND3_X1   g1364(.A1(new_n1750_), .A2(\a[112] ), .A3(new_n1746_), .ZN(new_n1751_));
  NAND2_X1   g1365(.A1(new_n1749_), .A2(new_n1751_), .ZN(\f[112] ));
  NOR2_X1    g1366(.A1(\a[112] ), .A2(\b[112] ), .ZN(new_n1753_));
  AND2_X2    g1367(.A1(\a[112] ), .A2(\b[112] ), .Z(new_n1754_));
  NOR3_X1    g1368(.A1(new_n1744_), .A2(new_n1754_), .A3(new_n1745_), .ZN(new_n1755_));
  NOR2_X1    g1369(.A1(new_n1755_), .A2(new_n1753_), .ZN(new_n1756_));
  XOR2_X1    g1370(.A1(\a[113] ), .A2(\b[113] ), .Z(new_n1757_));
  NAND2_X1   g1371(.A1(new_n1756_), .A2(new_n1757_), .ZN(new_n1758_));
  INV_X1     g1372(.I(\a[113] ), .ZN(new_n1759_));
  INV_X1     g1373(.I(\b[113] ), .ZN(new_n1760_));
  NOR2_X1    g1374(.A1(new_n1759_), .A2(new_n1760_), .ZN(new_n1761_));
  NOR2_X1    g1375(.A1(\a[113] ), .A2(\b[113] ), .ZN(new_n1762_));
  NOR2_X1    g1376(.A1(new_n1761_), .A2(new_n1762_), .ZN(new_n1763_));
  OAI21_X1   g1377(.A1(new_n1756_), .A2(new_n1763_), .B(new_n1758_), .ZN(\f[113] ));
  NOR3_X1    g1378(.A1(new_n1755_), .A2(new_n1753_), .A3(new_n1761_), .ZN(new_n1765_));
  XOR2_X1    g1379(.A1(\a[114] ), .A2(\b[114] ), .Z(new_n1766_));
  OAI21_X1   g1380(.A1(new_n1765_), .A2(new_n1762_), .B(new_n1766_), .ZN(new_n1767_));
  INV_X1     g1381(.I(new_n1762_), .ZN(new_n1768_));
  INV_X1     g1382(.I(new_n1753_), .ZN(new_n1769_));
  OR4_X2     g1383(.A1(\a[110] ), .A2(\a[111] ), .A3(\b[110] ), .A4(\b[111] ), .Z(new_n1770_));
  NAND2_X1   g1384(.A1(\a[112] ), .A2(\b[112] ), .ZN(new_n1771_));
  NAND3_X1   g1385(.A1(new_n1770_), .A2(new_n1743_), .A3(new_n1771_), .ZN(new_n1772_));
  INV_X1     g1386(.I(new_n1761_), .ZN(new_n1773_));
  NAND3_X1   g1387(.A1(new_n1772_), .A2(new_n1769_), .A3(new_n1773_), .ZN(new_n1774_));
  XNOR2_X1   g1388(.A1(\a[114] ), .A2(\b[114] ), .ZN(new_n1775_));
  NAND3_X1   g1389(.A1(new_n1774_), .A2(new_n1768_), .A3(new_n1775_), .ZN(new_n1776_));
  NAND2_X1   g1390(.A1(new_n1776_), .A2(new_n1767_), .ZN(\f[114] ));
  INV_X1     g1391(.I(\a[115] ), .ZN(new_n1778_));
  INV_X1     g1392(.I(\b[115] ), .ZN(new_n1779_));
  NAND2_X1   g1393(.A1(\a[114] ), .A2(\b[114] ), .ZN(new_n1780_));
  INV_X1     g1394(.I(new_n1780_), .ZN(new_n1781_));
  NOR4_X1    g1395(.A1(\a[113] ), .A2(\a[114] ), .A3(\b[113] ), .A4(\b[114] ), .ZN(new_n1782_));
  OAI21_X1   g1396(.A1(new_n1781_), .A2(new_n1782_), .B(new_n1779_), .ZN(new_n1783_));
  INV_X1     g1397(.I(new_n1783_), .ZN(new_n1784_));
  NOR3_X1    g1398(.A1(new_n1781_), .A2(new_n1782_), .A3(new_n1779_), .ZN(new_n1785_));
  OAI21_X1   g1399(.A1(new_n1784_), .A2(new_n1785_), .B(new_n1778_), .ZN(new_n1786_));
  INV_X1     g1400(.I(new_n1785_), .ZN(new_n1787_));
  NAND3_X1   g1401(.A1(new_n1787_), .A2(\a[115] ), .A3(new_n1783_), .ZN(new_n1788_));
  NAND2_X1   g1402(.A1(new_n1786_), .A2(new_n1788_), .ZN(\f[115] ));
  NOR2_X1    g1403(.A1(\a[115] ), .A2(\b[115] ), .ZN(new_n1790_));
  AND2_X2    g1404(.A1(\a[115] ), .A2(\b[115] ), .Z(new_n1791_));
  NOR3_X1    g1405(.A1(new_n1781_), .A2(new_n1791_), .A3(new_n1782_), .ZN(new_n1792_));
  NOR2_X1    g1406(.A1(new_n1792_), .A2(new_n1790_), .ZN(new_n1793_));
  XOR2_X1    g1407(.A1(\a[116] ), .A2(\b[116] ), .Z(new_n1794_));
  NAND2_X1   g1408(.A1(new_n1793_), .A2(new_n1794_), .ZN(new_n1795_));
  INV_X1     g1409(.I(\a[116] ), .ZN(new_n1796_));
  INV_X1     g1410(.I(\b[116] ), .ZN(new_n1797_));
  NOR2_X1    g1411(.A1(new_n1796_), .A2(new_n1797_), .ZN(new_n1798_));
  NOR2_X1    g1412(.A1(\a[116] ), .A2(\b[116] ), .ZN(new_n1799_));
  NOR2_X1    g1413(.A1(new_n1798_), .A2(new_n1799_), .ZN(new_n1800_));
  OAI21_X1   g1414(.A1(new_n1793_), .A2(new_n1800_), .B(new_n1795_), .ZN(\f[116] ));
  NOR3_X1    g1415(.A1(new_n1792_), .A2(new_n1790_), .A3(new_n1798_), .ZN(new_n1802_));
  XOR2_X1    g1416(.A1(\a[117] ), .A2(\b[117] ), .Z(new_n1803_));
  OAI21_X1   g1417(.A1(new_n1802_), .A2(new_n1799_), .B(new_n1803_), .ZN(new_n1804_));
  INV_X1     g1418(.I(new_n1799_), .ZN(new_n1805_));
  INV_X1     g1419(.I(new_n1790_), .ZN(new_n1806_));
  OR4_X2     g1420(.A1(\a[113] ), .A2(\a[114] ), .A3(\b[113] ), .A4(\b[114] ), .Z(new_n1807_));
  NAND2_X1   g1421(.A1(\a[115] ), .A2(\b[115] ), .ZN(new_n1808_));
  NAND3_X1   g1422(.A1(new_n1807_), .A2(new_n1780_), .A3(new_n1808_), .ZN(new_n1809_));
  INV_X1     g1423(.I(new_n1798_), .ZN(new_n1810_));
  NAND3_X1   g1424(.A1(new_n1809_), .A2(new_n1806_), .A3(new_n1810_), .ZN(new_n1811_));
  XNOR2_X1   g1425(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1812_));
  NAND3_X1   g1426(.A1(new_n1811_), .A2(new_n1805_), .A3(new_n1812_), .ZN(new_n1813_));
  NAND2_X1   g1427(.A1(new_n1813_), .A2(new_n1804_), .ZN(\f[117] ));
  INV_X1     g1428(.I(\a[118] ), .ZN(new_n1815_));
  INV_X1     g1429(.I(\b[118] ), .ZN(new_n1816_));
  NAND2_X1   g1430(.A1(\a[117] ), .A2(\b[117] ), .ZN(new_n1817_));
  INV_X1     g1431(.I(new_n1817_), .ZN(new_n1818_));
  NOR4_X1    g1432(.A1(\a[116] ), .A2(\a[117] ), .A3(\b[116] ), .A4(\b[117] ), .ZN(new_n1819_));
  OAI21_X1   g1433(.A1(new_n1818_), .A2(new_n1819_), .B(new_n1816_), .ZN(new_n1820_));
  INV_X1     g1434(.I(new_n1820_), .ZN(new_n1821_));
  NOR3_X1    g1435(.A1(new_n1818_), .A2(new_n1819_), .A3(new_n1816_), .ZN(new_n1822_));
  OAI21_X1   g1436(.A1(new_n1821_), .A2(new_n1822_), .B(new_n1815_), .ZN(new_n1823_));
  INV_X1     g1437(.I(new_n1822_), .ZN(new_n1824_));
  NAND3_X1   g1438(.A1(new_n1824_), .A2(\a[118] ), .A3(new_n1820_), .ZN(new_n1825_));
  NAND2_X1   g1439(.A1(new_n1823_), .A2(new_n1825_), .ZN(\f[118] ));
  NOR2_X1    g1440(.A1(\a[118] ), .A2(\b[118] ), .ZN(new_n1827_));
  AND2_X2    g1441(.A1(\a[118] ), .A2(\b[118] ), .Z(new_n1828_));
  NOR3_X1    g1442(.A1(new_n1818_), .A2(new_n1828_), .A3(new_n1819_), .ZN(new_n1829_));
  NOR2_X1    g1443(.A1(new_n1829_), .A2(new_n1827_), .ZN(new_n1830_));
  XOR2_X1    g1444(.A1(\a[119] ), .A2(\b[119] ), .Z(new_n1831_));
  NAND2_X1   g1445(.A1(new_n1830_), .A2(new_n1831_), .ZN(new_n1832_));
  INV_X1     g1446(.I(\a[119] ), .ZN(new_n1833_));
  INV_X1     g1447(.I(\b[119] ), .ZN(new_n1834_));
  NOR2_X1    g1448(.A1(new_n1833_), .A2(new_n1834_), .ZN(new_n1835_));
  NOR2_X1    g1449(.A1(\a[119] ), .A2(\b[119] ), .ZN(new_n1836_));
  NOR2_X1    g1450(.A1(new_n1835_), .A2(new_n1836_), .ZN(new_n1837_));
  OAI21_X1   g1451(.A1(new_n1830_), .A2(new_n1837_), .B(new_n1832_), .ZN(\f[119] ));
  NOR3_X1    g1452(.A1(new_n1829_), .A2(new_n1827_), .A3(new_n1835_), .ZN(new_n1839_));
  XOR2_X1    g1453(.A1(\a[120] ), .A2(\b[120] ), .Z(new_n1840_));
  OAI21_X1   g1454(.A1(new_n1839_), .A2(new_n1836_), .B(new_n1840_), .ZN(new_n1841_));
  INV_X1     g1455(.I(new_n1836_), .ZN(new_n1842_));
  INV_X1     g1456(.I(new_n1827_), .ZN(new_n1843_));
  OR4_X2     g1457(.A1(\a[116] ), .A2(\a[117] ), .A3(\b[116] ), .A4(\b[117] ), .Z(new_n1844_));
  NAND2_X1   g1458(.A1(\a[118] ), .A2(\b[118] ), .ZN(new_n1845_));
  NAND3_X1   g1459(.A1(new_n1844_), .A2(new_n1817_), .A3(new_n1845_), .ZN(new_n1846_));
  INV_X1     g1460(.I(new_n1835_), .ZN(new_n1847_));
  NAND3_X1   g1461(.A1(new_n1846_), .A2(new_n1843_), .A3(new_n1847_), .ZN(new_n1848_));
  XNOR2_X1   g1462(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1849_));
  NAND3_X1   g1463(.A1(new_n1848_), .A2(new_n1842_), .A3(new_n1849_), .ZN(new_n1850_));
  NAND2_X1   g1464(.A1(new_n1850_), .A2(new_n1841_), .ZN(\f[120] ));
  INV_X1     g1465(.I(\a[121] ), .ZN(new_n1852_));
  INV_X1     g1466(.I(\b[121] ), .ZN(new_n1853_));
  NAND2_X1   g1467(.A1(\a[120] ), .A2(\b[120] ), .ZN(new_n1854_));
  INV_X1     g1468(.I(new_n1854_), .ZN(new_n1855_));
  NOR4_X1    g1469(.A1(\a[119] ), .A2(\a[120] ), .A3(\b[119] ), .A4(\b[120] ), .ZN(new_n1856_));
  OAI21_X1   g1470(.A1(new_n1855_), .A2(new_n1856_), .B(new_n1853_), .ZN(new_n1857_));
  INV_X1     g1471(.I(new_n1857_), .ZN(new_n1858_));
  NOR3_X1    g1472(.A1(new_n1855_), .A2(new_n1856_), .A3(new_n1853_), .ZN(new_n1859_));
  OAI21_X1   g1473(.A1(new_n1858_), .A2(new_n1859_), .B(new_n1852_), .ZN(new_n1860_));
  INV_X1     g1474(.I(new_n1859_), .ZN(new_n1861_));
  NAND3_X1   g1475(.A1(new_n1861_), .A2(\a[121] ), .A3(new_n1857_), .ZN(new_n1862_));
  NAND2_X1   g1476(.A1(new_n1860_), .A2(new_n1862_), .ZN(\f[121] ));
  NOR2_X1    g1477(.A1(\a[121] ), .A2(\b[121] ), .ZN(new_n1864_));
  AND2_X2    g1478(.A1(\a[121] ), .A2(\b[121] ), .Z(new_n1865_));
  NOR3_X1    g1479(.A1(new_n1855_), .A2(new_n1865_), .A3(new_n1856_), .ZN(new_n1866_));
  NOR2_X1    g1480(.A1(new_n1866_), .A2(new_n1864_), .ZN(new_n1867_));
  XOR2_X1    g1481(.A1(\a[122] ), .A2(\b[122] ), .Z(new_n1868_));
  NAND2_X1   g1482(.A1(new_n1867_), .A2(new_n1868_), .ZN(new_n1869_));
  INV_X1     g1483(.I(\a[122] ), .ZN(new_n1870_));
  INV_X1     g1484(.I(\b[122] ), .ZN(new_n1871_));
  NOR2_X1    g1485(.A1(new_n1870_), .A2(new_n1871_), .ZN(new_n1872_));
  NOR2_X1    g1486(.A1(\a[122] ), .A2(\b[122] ), .ZN(new_n1873_));
  NOR2_X1    g1487(.A1(new_n1872_), .A2(new_n1873_), .ZN(new_n1874_));
  OAI21_X1   g1488(.A1(new_n1867_), .A2(new_n1874_), .B(new_n1869_), .ZN(\f[122] ));
  NOR3_X1    g1489(.A1(new_n1866_), .A2(new_n1864_), .A3(new_n1872_), .ZN(new_n1876_));
  XOR2_X1    g1490(.A1(\a[123] ), .A2(\b[123] ), .Z(new_n1877_));
  OAI21_X1   g1491(.A1(new_n1876_), .A2(new_n1873_), .B(new_n1877_), .ZN(new_n1878_));
  INV_X1     g1492(.I(new_n1873_), .ZN(new_n1879_));
  INV_X1     g1493(.I(new_n1864_), .ZN(new_n1880_));
  OR4_X2     g1494(.A1(\a[119] ), .A2(\a[120] ), .A3(\b[119] ), .A4(\b[120] ), .Z(new_n1881_));
  NAND2_X1   g1495(.A1(\a[121] ), .A2(\b[121] ), .ZN(new_n1882_));
  NAND3_X1   g1496(.A1(new_n1881_), .A2(new_n1854_), .A3(new_n1882_), .ZN(new_n1883_));
  INV_X1     g1497(.I(new_n1872_), .ZN(new_n1884_));
  NAND3_X1   g1498(.A1(new_n1883_), .A2(new_n1880_), .A3(new_n1884_), .ZN(new_n1885_));
  XNOR2_X1   g1499(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1886_));
  NAND3_X1   g1500(.A1(new_n1885_), .A2(new_n1879_), .A3(new_n1886_), .ZN(new_n1887_));
  NAND2_X1   g1501(.A1(new_n1887_), .A2(new_n1878_), .ZN(\f[123] ));
  INV_X1     g1502(.I(\a[124] ), .ZN(new_n1889_));
  INV_X1     g1503(.I(\b[124] ), .ZN(new_n1890_));
  NAND2_X1   g1504(.A1(\a[123] ), .A2(\b[123] ), .ZN(new_n1891_));
  INV_X1     g1505(.I(new_n1891_), .ZN(new_n1892_));
  NOR4_X1    g1506(.A1(\a[122] ), .A2(\a[123] ), .A3(\b[122] ), .A4(\b[123] ), .ZN(new_n1893_));
  OAI21_X1   g1507(.A1(new_n1892_), .A2(new_n1893_), .B(new_n1890_), .ZN(new_n1894_));
  INV_X1     g1508(.I(new_n1894_), .ZN(new_n1895_));
  NOR3_X1    g1509(.A1(new_n1892_), .A2(new_n1893_), .A3(new_n1890_), .ZN(new_n1896_));
  OAI21_X1   g1510(.A1(new_n1895_), .A2(new_n1896_), .B(new_n1889_), .ZN(new_n1897_));
  INV_X1     g1511(.I(new_n1896_), .ZN(new_n1898_));
  NAND3_X1   g1512(.A1(new_n1898_), .A2(\a[124] ), .A3(new_n1894_), .ZN(new_n1899_));
  NAND2_X1   g1513(.A1(new_n1897_), .A2(new_n1899_), .ZN(\f[124] ));
  NOR2_X1    g1514(.A1(\a[124] ), .A2(\b[124] ), .ZN(new_n1901_));
  AND2_X2    g1515(.A1(\a[124] ), .A2(\b[124] ), .Z(new_n1902_));
  NOR3_X1    g1516(.A1(new_n1892_), .A2(new_n1902_), .A3(new_n1893_), .ZN(new_n1903_));
  NOR2_X1    g1517(.A1(new_n1903_), .A2(new_n1901_), .ZN(new_n1904_));
  XOR2_X1    g1518(.A1(\a[125] ), .A2(\b[125] ), .Z(new_n1905_));
  NAND2_X1   g1519(.A1(new_n1904_), .A2(new_n1905_), .ZN(new_n1906_));
  INV_X1     g1520(.I(\a[125] ), .ZN(new_n1907_));
  INV_X1     g1521(.I(\b[125] ), .ZN(new_n1908_));
  NOR2_X1    g1522(.A1(new_n1907_), .A2(new_n1908_), .ZN(new_n1909_));
  NOR2_X1    g1523(.A1(\a[125] ), .A2(\b[125] ), .ZN(new_n1910_));
  NOR2_X1    g1524(.A1(new_n1909_), .A2(new_n1910_), .ZN(new_n1911_));
  OAI21_X1   g1525(.A1(new_n1904_), .A2(new_n1911_), .B(new_n1906_), .ZN(\f[125] ));
  NOR3_X1    g1526(.A1(new_n1903_), .A2(new_n1901_), .A3(new_n1909_), .ZN(new_n1913_));
  XOR2_X1    g1527(.A1(\a[126] ), .A2(\b[126] ), .Z(new_n1914_));
  OAI21_X1   g1528(.A1(new_n1913_), .A2(new_n1910_), .B(new_n1914_), .ZN(new_n1915_));
  INV_X1     g1529(.I(new_n1910_), .ZN(new_n1916_));
  INV_X1     g1530(.I(new_n1901_), .ZN(new_n1917_));
  OR4_X2     g1531(.A1(\a[122] ), .A2(\a[123] ), .A3(\b[122] ), .A4(\b[123] ), .Z(new_n1918_));
  NAND2_X1   g1532(.A1(\a[124] ), .A2(\b[124] ), .ZN(new_n1919_));
  NAND3_X1   g1533(.A1(new_n1918_), .A2(new_n1891_), .A3(new_n1919_), .ZN(new_n1920_));
  INV_X1     g1534(.I(new_n1909_), .ZN(new_n1921_));
  NAND3_X1   g1535(.A1(new_n1920_), .A2(new_n1917_), .A3(new_n1921_), .ZN(new_n1922_));
  XNOR2_X1   g1536(.A1(\a[126] ), .A2(\b[126] ), .ZN(new_n1923_));
  NAND3_X1   g1537(.A1(new_n1922_), .A2(new_n1916_), .A3(new_n1923_), .ZN(new_n1924_));
  NAND2_X1   g1538(.A1(new_n1924_), .A2(new_n1915_), .ZN(\f[126] ));
  INV_X1     g1539(.I(\a[127] ), .ZN(new_n1926_));
  INV_X1     g1540(.I(\b[127] ), .ZN(new_n1927_));
  AND2_X2    g1541(.A1(\a[126] ), .A2(\b[126] ), .Z(new_n1928_));
  NOR4_X1    g1542(.A1(\a[125] ), .A2(\a[126] ), .A3(\b[125] ), .A4(\b[126] ), .ZN(new_n1929_));
  OAI21_X1   g1543(.A1(new_n1928_), .A2(new_n1929_), .B(new_n1927_), .ZN(new_n1930_));
  INV_X1     g1544(.I(new_n1930_), .ZN(new_n1931_));
  NOR3_X1    g1545(.A1(new_n1928_), .A2(new_n1929_), .A3(new_n1927_), .ZN(new_n1932_));
  OAI21_X1   g1546(.A1(new_n1931_), .A2(new_n1932_), .B(new_n1926_), .ZN(new_n1933_));
  INV_X1     g1547(.I(new_n1932_), .ZN(new_n1934_));
  NAND3_X1   g1548(.A1(new_n1934_), .A2(\a[127] ), .A3(new_n1930_), .ZN(new_n1935_));
  NAND2_X1   g1549(.A1(new_n1933_), .A2(new_n1935_), .ZN(\f[127] ));
  NOR2_X1    g1550(.A1(new_n1928_), .A2(new_n1929_), .ZN(new_n1937_));
  NOR2_X1    g1551(.A1(\a[127] ), .A2(\b[127] ), .ZN(new_n1938_));
  NAND2_X1   g1552(.A1(\a[127] ), .A2(\b[127] ), .ZN(new_n1939_));
  AOI21_X1   g1553(.A1(new_n1937_), .A2(new_n1939_), .B(new_n1938_), .ZN(cOut));
endmodule


