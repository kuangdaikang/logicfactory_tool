// Benchmark "priority" written by ABC on Mon Sep 11 23:34:22 2023

module priority ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_,
    new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1317_, new_n1318_, new_n1319_;
  INV_X1     g0000(.I(\A[127] ), .ZN(new_n137_));
  AOI21_X1   g0001(.A1(new_n137_), .A2(\A[126] ), .B(\A[124] ), .ZN(new_n138_));
  INV_X1     g0002(.I(\A[125] ), .ZN(new_n139_));
  OAI21_X1   g0003(.A1(new_n139_), .A2(\A[126] ), .B(new_n137_), .ZN(new_n140_));
  AOI21_X1   g0004(.A1(new_n140_), .A2(\A[124] ), .B(new_n138_), .ZN(new_n141_));
  NOR2_X1    g0005(.A1(new_n141_), .A2(\A[122] ), .ZN(new_n142_));
  INV_X1     g0006(.I(\A[123] ), .ZN(new_n143_));
  NAND2_X1   g0007(.A1(new_n140_), .A2(new_n143_), .ZN(new_n144_));
  OAI21_X1   g0008(.A1(new_n141_), .A2(new_n143_), .B(new_n144_), .ZN(new_n145_));
  AOI21_X1   g0009(.A1(new_n145_), .A2(\A[122] ), .B(new_n142_), .ZN(new_n146_));
  NOR2_X1    g0010(.A1(new_n146_), .A2(\A[120] ), .ZN(new_n147_));
  INV_X1     g0011(.I(\A[121] ), .ZN(new_n148_));
  NAND2_X1   g0012(.A1(new_n145_), .A2(new_n148_), .ZN(new_n149_));
  OAI21_X1   g0013(.A1(new_n146_), .A2(new_n148_), .B(new_n149_), .ZN(new_n150_));
  AOI21_X1   g0014(.A1(new_n150_), .A2(\A[120] ), .B(new_n147_), .ZN(new_n151_));
  NOR2_X1    g0015(.A1(new_n151_), .A2(\A[118] ), .ZN(new_n152_));
  INV_X1     g0016(.I(\A[119] ), .ZN(new_n153_));
  NAND2_X1   g0017(.A1(new_n150_), .A2(new_n153_), .ZN(new_n154_));
  OAI21_X1   g0018(.A1(new_n151_), .A2(new_n153_), .B(new_n154_), .ZN(new_n155_));
  AOI21_X1   g0019(.A1(new_n155_), .A2(\A[118] ), .B(new_n152_), .ZN(new_n156_));
  NOR2_X1    g0020(.A1(new_n156_), .A2(\A[116] ), .ZN(new_n157_));
  INV_X1     g0021(.I(new_n157_), .ZN(new_n158_));
  INV_X1     g0022(.I(\A[117] ), .ZN(new_n159_));
  NAND2_X1   g0023(.A1(new_n155_), .A2(new_n159_), .ZN(new_n160_));
  OAI21_X1   g0024(.A1(new_n156_), .A2(new_n159_), .B(new_n160_), .ZN(new_n161_));
  NAND2_X1   g0025(.A1(new_n161_), .A2(\A[116] ), .ZN(new_n162_));
  AOI21_X1   g0026(.A1(new_n162_), .A2(new_n158_), .B(\A[114] ), .ZN(new_n163_));
  INV_X1     g0027(.I(new_n163_), .ZN(new_n164_));
  INV_X1     g0028(.I(\A[115] ), .ZN(new_n165_));
  AOI21_X1   g0029(.A1(new_n161_), .A2(\A[116] ), .B(new_n157_), .ZN(new_n166_));
  NAND2_X1   g0030(.A1(new_n161_), .A2(new_n165_), .ZN(new_n167_));
  OAI21_X1   g0031(.A1(new_n166_), .A2(new_n165_), .B(new_n167_), .ZN(new_n168_));
  NAND2_X1   g0032(.A1(new_n168_), .A2(\A[114] ), .ZN(new_n169_));
  AOI21_X1   g0033(.A1(new_n169_), .A2(new_n164_), .B(\A[112] ), .ZN(new_n170_));
  INV_X1     g0034(.I(new_n170_), .ZN(new_n171_));
  INV_X1     g0035(.I(\A[113] ), .ZN(new_n172_));
  NAND2_X1   g0036(.A1(new_n168_), .A2(new_n172_), .ZN(new_n173_));
  INV_X1     g0037(.I(new_n173_), .ZN(new_n174_));
  AOI21_X1   g0038(.A1(new_n169_), .A2(new_n164_), .B(new_n172_), .ZN(new_n175_));
  OAI21_X1   g0039(.A1(new_n175_), .A2(new_n174_), .B(\A[112] ), .ZN(new_n176_));
  AOI21_X1   g0040(.A1(new_n176_), .A2(new_n171_), .B(\A[110] ), .ZN(new_n177_));
  INV_X1     g0041(.I(new_n177_), .ZN(new_n178_));
  INV_X1     g0042(.I(\A[111] ), .ZN(new_n179_));
  OAI21_X1   g0043(.A1(new_n175_), .A2(new_n174_), .B(new_n179_), .ZN(new_n180_));
  INV_X1     g0044(.I(new_n180_), .ZN(new_n181_));
  AOI21_X1   g0045(.A1(new_n176_), .A2(new_n171_), .B(new_n179_), .ZN(new_n182_));
  OAI21_X1   g0046(.A1(new_n182_), .A2(new_n181_), .B(\A[110] ), .ZN(new_n183_));
  AOI21_X1   g0047(.A1(new_n183_), .A2(new_n178_), .B(\A[108] ), .ZN(new_n184_));
  INV_X1     g0048(.I(new_n184_), .ZN(new_n185_));
  INV_X1     g0049(.I(\A[109] ), .ZN(new_n186_));
  OAI21_X1   g0050(.A1(new_n182_), .A2(new_n181_), .B(new_n186_), .ZN(new_n187_));
  INV_X1     g0051(.I(new_n187_), .ZN(new_n188_));
  AOI21_X1   g0052(.A1(new_n183_), .A2(new_n178_), .B(new_n186_), .ZN(new_n189_));
  OAI21_X1   g0053(.A1(new_n189_), .A2(new_n188_), .B(\A[108] ), .ZN(new_n190_));
  AOI21_X1   g0054(.A1(new_n190_), .A2(new_n185_), .B(\A[106] ), .ZN(new_n191_));
  INV_X1     g0055(.I(new_n191_), .ZN(new_n192_));
  INV_X1     g0056(.I(\A[107] ), .ZN(new_n193_));
  OAI21_X1   g0057(.A1(new_n189_), .A2(new_n188_), .B(new_n193_), .ZN(new_n194_));
  INV_X1     g0058(.I(new_n194_), .ZN(new_n195_));
  AOI21_X1   g0059(.A1(new_n190_), .A2(new_n185_), .B(new_n193_), .ZN(new_n196_));
  OAI21_X1   g0060(.A1(new_n196_), .A2(new_n195_), .B(\A[106] ), .ZN(new_n197_));
  AOI21_X1   g0061(.A1(new_n197_), .A2(new_n192_), .B(\A[104] ), .ZN(new_n198_));
  INV_X1     g0062(.I(new_n198_), .ZN(new_n199_));
  INV_X1     g0063(.I(\A[105] ), .ZN(new_n200_));
  OAI21_X1   g0064(.A1(new_n196_), .A2(new_n195_), .B(new_n200_), .ZN(new_n201_));
  INV_X1     g0065(.I(new_n201_), .ZN(new_n202_));
  AOI21_X1   g0066(.A1(new_n197_), .A2(new_n192_), .B(new_n200_), .ZN(new_n203_));
  OAI21_X1   g0067(.A1(new_n203_), .A2(new_n202_), .B(\A[104] ), .ZN(new_n204_));
  AOI21_X1   g0068(.A1(new_n204_), .A2(new_n199_), .B(\A[102] ), .ZN(new_n205_));
  INV_X1     g0069(.I(new_n205_), .ZN(new_n206_));
  INV_X1     g0070(.I(\A[103] ), .ZN(new_n207_));
  OAI21_X1   g0071(.A1(new_n203_), .A2(new_n202_), .B(new_n207_), .ZN(new_n208_));
  INV_X1     g0072(.I(new_n208_), .ZN(new_n209_));
  AOI21_X1   g0073(.A1(new_n204_), .A2(new_n199_), .B(new_n207_), .ZN(new_n210_));
  OAI21_X1   g0074(.A1(new_n210_), .A2(new_n209_), .B(\A[102] ), .ZN(new_n211_));
  AOI21_X1   g0075(.A1(new_n211_), .A2(new_n206_), .B(\A[100] ), .ZN(new_n212_));
  INV_X1     g0076(.I(new_n212_), .ZN(new_n213_));
  INV_X1     g0077(.I(\A[101] ), .ZN(new_n214_));
  OAI21_X1   g0078(.A1(new_n210_), .A2(new_n209_), .B(new_n214_), .ZN(new_n215_));
  INV_X1     g0079(.I(new_n215_), .ZN(new_n216_));
  AOI21_X1   g0080(.A1(new_n211_), .A2(new_n206_), .B(new_n214_), .ZN(new_n217_));
  OAI21_X1   g0081(.A1(new_n217_), .A2(new_n216_), .B(\A[100] ), .ZN(new_n218_));
  AOI21_X1   g0082(.A1(new_n218_), .A2(new_n213_), .B(\A[98] ), .ZN(new_n219_));
  INV_X1     g0083(.I(new_n219_), .ZN(new_n220_));
  INV_X1     g0084(.I(\A[99] ), .ZN(new_n221_));
  OAI21_X1   g0085(.A1(new_n217_), .A2(new_n216_), .B(new_n221_), .ZN(new_n222_));
  INV_X1     g0086(.I(new_n222_), .ZN(new_n223_));
  AOI21_X1   g0087(.A1(new_n218_), .A2(new_n213_), .B(new_n221_), .ZN(new_n224_));
  OAI21_X1   g0088(.A1(new_n224_), .A2(new_n223_), .B(\A[98] ), .ZN(new_n225_));
  AOI21_X1   g0089(.A1(new_n225_), .A2(new_n220_), .B(\A[96] ), .ZN(new_n226_));
  INV_X1     g0090(.I(new_n226_), .ZN(new_n227_));
  INV_X1     g0091(.I(\A[97] ), .ZN(new_n228_));
  OAI21_X1   g0092(.A1(new_n224_), .A2(new_n223_), .B(new_n228_), .ZN(new_n229_));
  INV_X1     g0093(.I(new_n229_), .ZN(new_n230_));
  AOI21_X1   g0094(.A1(new_n225_), .A2(new_n220_), .B(new_n228_), .ZN(new_n231_));
  OAI21_X1   g0095(.A1(new_n231_), .A2(new_n230_), .B(\A[96] ), .ZN(new_n232_));
  AOI21_X1   g0096(.A1(new_n232_), .A2(new_n227_), .B(\A[94] ), .ZN(new_n233_));
  INV_X1     g0097(.I(new_n233_), .ZN(new_n234_));
  INV_X1     g0098(.I(\A[95] ), .ZN(new_n235_));
  OAI21_X1   g0099(.A1(new_n231_), .A2(new_n230_), .B(new_n235_), .ZN(new_n236_));
  INV_X1     g0100(.I(new_n236_), .ZN(new_n237_));
  AOI21_X1   g0101(.A1(new_n232_), .A2(new_n227_), .B(new_n235_), .ZN(new_n238_));
  OAI21_X1   g0102(.A1(new_n238_), .A2(new_n237_), .B(\A[94] ), .ZN(new_n239_));
  AOI21_X1   g0103(.A1(new_n239_), .A2(new_n234_), .B(\A[92] ), .ZN(new_n240_));
  INV_X1     g0104(.I(new_n240_), .ZN(new_n241_));
  INV_X1     g0105(.I(\A[93] ), .ZN(new_n242_));
  OAI21_X1   g0106(.A1(new_n238_), .A2(new_n237_), .B(new_n242_), .ZN(new_n243_));
  INV_X1     g0107(.I(new_n243_), .ZN(new_n244_));
  AOI21_X1   g0108(.A1(new_n239_), .A2(new_n234_), .B(new_n242_), .ZN(new_n245_));
  OAI21_X1   g0109(.A1(new_n245_), .A2(new_n244_), .B(\A[92] ), .ZN(new_n246_));
  AOI21_X1   g0110(.A1(new_n246_), .A2(new_n241_), .B(\A[90] ), .ZN(new_n247_));
  INV_X1     g0111(.I(new_n247_), .ZN(new_n248_));
  INV_X1     g0112(.I(\A[91] ), .ZN(new_n249_));
  OAI21_X1   g0113(.A1(new_n245_), .A2(new_n244_), .B(new_n249_), .ZN(new_n250_));
  INV_X1     g0114(.I(new_n250_), .ZN(new_n251_));
  AOI21_X1   g0115(.A1(new_n246_), .A2(new_n241_), .B(new_n249_), .ZN(new_n252_));
  OAI21_X1   g0116(.A1(new_n252_), .A2(new_n251_), .B(\A[90] ), .ZN(new_n253_));
  AOI21_X1   g0117(.A1(new_n253_), .A2(new_n248_), .B(\A[88] ), .ZN(new_n254_));
  INV_X1     g0118(.I(new_n254_), .ZN(new_n255_));
  INV_X1     g0119(.I(\A[89] ), .ZN(new_n256_));
  OAI21_X1   g0120(.A1(new_n252_), .A2(new_n251_), .B(new_n256_), .ZN(new_n257_));
  INV_X1     g0121(.I(new_n257_), .ZN(new_n258_));
  AOI21_X1   g0122(.A1(new_n253_), .A2(new_n248_), .B(new_n256_), .ZN(new_n259_));
  OAI21_X1   g0123(.A1(new_n259_), .A2(new_n258_), .B(\A[88] ), .ZN(new_n260_));
  AOI21_X1   g0124(.A1(new_n260_), .A2(new_n255_), .B(\A[86] ), .ZN(new_n261_));
  INV_X1     g0125(.I(new_n261_), .ZN(new_n262_));
  INV_X1     g0126(.I(\A[87] ), .ZN(new_n263_));
  OAI21_X1   g0127(.A1(new_n259_), .A2(new_n258_), .B(new_n263_), .ZN(new_n264_));
  INV_X1     g0128(.I(new_n264_), .ZN(new_n265_));
  AOI21_X1   g0129(.A1(new_n260_), .A2(new_n255_), .B(new_n263_), .ZN(new_n266_));
  OAI21_X1   g0130(.A1(new_n266_), .A2(new_n265_), .B(\A[86] ), .ZN(new_n267_));
  AOI21_X1   g0131(.A1(new_n267_), .A2(new_n262_), .B(\A[84] ), .ZN(new_n268_));
  INV_X1     g0132(.I(new_n268_), .ZN(new_n269_));
  INV_X1     g0133(.I(\A[85] ), .ZN(new_n270_));
  OAI21_X1   g0134(.A1(new_n266_), .A2(new_n265_), .B(new_n270_), .ZN(new_n271_));
  INV_X1     g0135(.I(new_n271_), .ZN(new_n272_));
  AOI21_X1   g0136(.A1(new_n267_), .A2(new_n262_), .B(new_n270_), .ZN(new_n273_));
  OAI21_X1   g0137(.A1(new_n273_), .A2(new_n272_), .B(\A[84] ), .ZN(new_n274_));
  AOI21_X1   g0138(.A1(new_n274_), .A2(new_n269_), .B(\A[82] ), .ZN(new_n275_));
  INV_X1     g0139(.I(new_n275_), .ZN(new_n276_));
  INV_X1     g0140(.I(\A[83] ), .ZN(new_n277_));
  OAI21_X1   g0141(.A1(new_n273_), .A2(new_n272_), .B(new_n277_), .ZN(new_n278_));
  INV_X1     g0142(.I(new_n278_), .ZN(new_n279_));
  AOI21_X1   g0143(.A1(new_n274_), .A2(new_n269_), .B(new_n277_), .ZN(new_n280_));
  OAI21_X1   g0144(.A1(new_n280_), .A2(new_n279_), .B(\A[82] ), .ZN(new_n281_));
  AOI21_X1   g0145(.A1(new_n281_), .A2(new_n276_), .B(\A[80] ), .ZN(new_n282_));
  INV_X1     g0146(.I(new_n282_), .ZN(new_n283_));
  INV_X1     g0147(.I(\A[81] ), .ZN(new_n284_));
  OAI21_X1   g0148(.A1(new_n280_), .A2(new_n279_), .B(new_n284_), .ZN(new_n285_));
  INV_X1     g0149(.I(new_n285_), .ZN(new_n286_));
  AOI21_X1   g0150(.A1(new_n281_), .A2(new_n276_), .B(new_n284_), .ZN(new_n287_));
  OAI21_X1   g0151(.A1(new_n287_), .A2(new_n286_), .B(\A[80] ), .ZN(new_n288_));
  AOI21_X1   g0152(.A1(new_n288_), .A2(new_n283_), .B(\A[78] ), .ZN(new_n289_));
  INV_X1     g0153(.I(new_n289_), .ZN(new_n290_));
  INV_X1     g0154(.I(\A[79] ), .ZN(new_n291_));
  OAI21_X1   g0155(.A1(new_n287_), .A2(new_n286_), .B(new_n291_), .ZN(new_n292_));
  INV_X1     g0156(.I(new_n292_), .ZN(new_n293_));
  AOI21_X1   g0157(.A1(new_n288_), .A2(new_n283_), .B(new_n291_), .ZN(new_n294_));
  OAI21_X1   g0158(.A1(new_n294_), .A2(new_n293_), .B(\A[78] ), .ZN(new_n295_));
  AOI21_X1   g0159(.A1(new_n295_), .A2(new_n290_), .B(\A[76] ), .ZN(new_n296_));
  INV_X1     g0160(.I(new_n296_), .ZN(new_n297_));
  INV_X1     g0161(.I(\A[77] ), .ZN(new_n298_));
  OAI21_X1   g0162(.A1(new_n294_), .A2(new_n293_), .B(new_n298_), .ZN(new_n299_));
  INV_X1     g0163(.I(new_n299_), .ZN(new_n300_));
  AOI21_X1   g0164(.A1(new_n295_), .A2(new_n290_), .B(new_n298_), .ZN(new_n301_));
  OAI21_X1   g0165(.A1(new_n301_), .A2(new_n300_), .B(\A[76] ), .ZN(new_n302_));
  AOI21_X1   g0166(.A1(new_n302_), .A2(new_n297_), .B(\A[74] ), .ZN(new_n303_));
  INV_X1     g0167(.I(new_n303_), .ZN(new_n304_));
  INV_X1     g0168(.I(\A[75] ), .ZN(new_n305_));
  OAI21_X1   g0169(.A1(new_n301_), .A2(new_n300_), .B(new_n305_), .ZN(new_n306_));
  INV_X1     g0170(.I(new_n306_), .ZN(new_n307_));
  AOI21_X1   g0171(.A1(new_n302_), .A2(new_n297_), .B(new_n305_), .ZN(new_n308_));
  OAI21_X1   g0172(.A1(new_n308_), .A2(new_n307_), .B(\A[74] ), .ZN(new_n309_));
  AOI21_X1   g0173(.A1(new_n309_), .A2(new_n304_), .B(\A[72] ), .ZN(new_n310_));
  INV_X1     g0174(.I(new_n310_), .ZN(new_n311_));
  INV_X1     g0175(.I(\A[73] ), .ZN(new_n312_));
  OAI21_X1   g0176(.A1(new_n308_), .A2(new_n307_), .B(new_n312_), .ZN(new_n313_));
  INV_X1     g0177(.I(new_n313_), .ZN(new_n314_));
  AOI21_X1   g0178(.A1(new_n309_), .A2(new_n304_), .B(new_n312_), .ZN(new_n315_));
  OAI21_X1   g0179(.A1(new_n315_), .A2(new_n314_), .B(\A[72] ), .ZN(new_n316_));
  AOI21_X1   g0180(.A1(new_n316_), .A2(new_n311_), .B(\A[70] ), .ZN(new_n317_));
  INV_X1     g0181(.I(new_n317_), .ZN(new_n318_));
  INV_X1     g0182(.I(\A[71] ), .ZN(new_n319_));
  OAI21_X1   g0183(.A1(new_n315_), .A2(new_n314_), .B(new_n319_), .ZN(new_n320_));
  INV_X1     g0184(.I(new_n320_), .ZN(new_n321_));
  AOI21_X1   g0185(.A1(new_n316_), .A2(new_n311_), .B(new_n319_), .ZN(new_n322_));
  OAI21_X1   g0186(.A1(new_n322_), .A2(new_n321_), .B(\A[70] ), .ZN(new_n323_));
  AOI21_X1   g0187(.A1(new_n323_), .A2(new_n318_), .B(\A[68] ), .ZN(new_n324_));
  INV_X1     g0188(.I(new_n324_), .ZN(new_n325_));
  INV_X1     g0189(.I(\A[69] ), .ZN(new_n326_));
  OAI21_X1   g0190(.A1(new_n322_), .A2(new_n321_), .B(new_n326_), .ZN(new_n327_));
  INV_X1     g0191(.I(new_n327_), .ZN(new_n328_));
  AOI21_X1   g0192(.A1(new_n323_), .A2(new_n318_), .B(new_n326_), .ZN(new_n329_));
  OAI21_X1   g0193(.A1(new_n329_), .A2(new_n328_), .B(\A[68] ), .ZN(new_n330_));
  AOI21_X1   g0194(.A1(new_n330_), .A2(new_n325_), .B(\A[66] ), .ZN(new_n331_));
  INV_X1     g0195(.I(new_n331_), .ZN(new_n332_));
  INV_X1     g0196(.I(\A[67] ), .ZN(new_n333_));
  OAI21_X1   g0197(.A1(new_n329_), .A2(new_n328_), .B(new_n333_), .ZN(new_n334_));
  INV_X1     g0198(.I(new_n334_), .ZN(new_n335_));
  AOI21_X1   g0199(.A1(new_n330_), .A2(new_n325_), .B(new_n333_), .ZN(new_n336_));
  OAI21_X1   g0200(.A1(new_n336_), .A2(new_n335_), .B(\A[66] ), .ZN(new_n337_));
  AOI21_X1   g0201(.A1(new_n337_), .A2(new_n332_), .B(\A[64] ), .ZN(new_n338_));
  INV_X1     g0202(.I(new_n338_), .ZN(new_n339_));
  INV_X1     g0203(.I(\A[65] ), .ZN(new_n340_));
  OAI21_X1   g0204(.A1(new_n336_), .A2(new_n335_), .B(new_n340_), .ZN(new_n341_));
  INV_X1     g0205(.I(new_n341_), .ZN(new_n342_));
  AOI21_X1   g0206(.A1(new_n337_), .A2(new_n332_), .B(new_n340_), .ZN(new_n343_));
  OAI21_X1   g0207(.A1(new_n343_), .A2(new_n342_), .B(\A[64] ), .ZN(new_n344_));
  AOI21_X1   g0208(.A1(new_n344_), .A2(new_n339_), .B(\A[62] ), .ZN(new_n345_));
  INV_X1     g0209(.I(new_n345_), .ZN(new_n346_));
  INV_X1     g0210(.I(\A[63] ), .ZN(new_n347_));
  OAI21_X1   g0211(.A1(new_n343_), .A2(new_n342_), .B(new_n347_), .ZN(new_n348_));
  INV_X1     g0212(.I(new_n348_), .ZN(new_n349_));
  AOI21_X1   g0213(.A1(new_n344_), .A2(new_n339_), .B(new_n347_), .ZN(new_n350_));
  OAI21_X1   g0214(.A1(new_n350_), .A2(new_n349_), .B(\A[62] ), .ZN(new_n351_));
  AOI21_X1   g0215(.A1(new_n351_), .A2(new_n346_), .B(\A[60] ), .ZN(new_n352_));
  INV_X1     g0216(.I(new_n352_), .ZN(new_n353_));
  INV_X1     g0217(.I(\A[61] ), .ZN(new_n354_));
  OAI21_X1   g0218(.A1(new_n350_), .A2(new_n349_), .B(new_n354_), .ZN(new_n355_));
  INV_X1     g0219(.I(new_n355_), .ZN(new_n356_));
  AOI21_X1   g0220(.A1(new_n351_), .A2(new_n346_), .B(new_n354_), .ZN(new_n357_));
  OAI21_X1   g0221(.A1(new_n357_), .A2(new_n356_), .B(\A[60] ), .ZN(new_n358_));
  AOI21_X1   g0222(.A1(new_n358_), .A2(new_n353_), .B(\A[58] ), .ZN(new_n359_));
  INV_X1     g0223(.I(new_n359_), .ZN(new_n360_));
  INV_X1     g0224(.I(\A[59] ), .ZN(new_n361_));
  OAI21_X1   g0225(.A1(new_n357_), .A2(new_n356_), .B(new_n361_), .ZN(new_n362_));
  INV_X1     g0226(.I(new_n362_), .ZN(new_n363_));
  AOI21_X1   g0227(.A1(new_n358_), .A2(new_n353_), .B(new_n361_), .ZN(new_n364_));
  OAI21_X1   g0228(.A1(new_n364_), .A2(new_n363_), .B(\A[58] ), .ZN(new_n365_));
  AOI21_X1   g0229(.A1(new_n365_), .A2(new_n360_), .B(\A[56] ), .ZN(new_n366_));
  INV_X1     g0230(.I(new_n366_), .ZN(new_n367_));
  INV_X1     g0231(.I(\A[57] ), .ZN(new_n368_));
  OAI21_X1   g0232(.A1(new_n364_), .A2(new_n363_), .B(new_n368_), .ZN(new_n369_));
  INV_X1     g0233(.I(new_n369_), .ZN(new_n370_));
  AOI21_X1   g0234(.A1(new_n365_), .A2(new_n360_), .B(new_n368_), .ZN(new_n371_));
  OAI21_X1   g0235(.A1(new_n371_), .A2(new_n370_), .B(\A[56] ), .ZN(new_n372_));
  AOI21_X1   g0236(.A1(new_n372_), .A2(new_n367_), .B(\A[54] ), .ZN(new_n373_));
  INV_X1     g0237(.I(new_n373_), .ZN(new_n374_));
  INV_X1     g0238(.I(\A[55] ), .ZN(new_n375_));
  OAI21_X1   g0239(.A1(new_n371_), .A2(new_n370_), .B(new_n375_), .ZN(new_n376_));
  INV_X1     g0240(.I(new_n376_), .ZN(new_n377_));
  AOI21_X1   g0241(.A1(new_n372_), .A2(new_n367_), .B(new_n375_), .ZN(new_n378_));
  OAI21_X1   g0242(.A1(new_n378_), .A2(new_n377_), .B(\A[54] ), .ZN(new_n379_));
  AOI21_X1   g0243(.A1(new_n379_), .A2(new_n374_), .B(\A[52] ), .ZN(new_n380_));
  INV_X1     g0244(.I(new_n380_), .ZN(new_n381_));
  INV_X1     g0245(.I(\A[53] ), .ZN(new_n382_));
  OAI21_X1   g0246(.A1(new_n378_), .A2(new_n377_), .B(new_n382_), .ZN(new_n383_));
  INV_X1     g0247(.I(new_n383_), .ZN(new_n384_));
  AOI21_X1   g0248(.A1(new_n379_), .A2(new_n374_), .B(new_n382_), .ZN(new_n385_));
  OAI21_X1   g0249(.A1(new_n385_), .A2(new_n384_), .B(\A[52] ), .ZN(new_n386_));
  AOI21_X1   g0250(.A1(new_n386_), .A2(new_n381_), .B(\A[50] ), .ZN(new_n387_));
  INV_X1     g0251(.I(new_n387_), .ZN(new_n388_));
  INV_X1     g0252(.I(\A[51] ), .ZN(new_n389_));
  OAI21_X1   g0253(.A1(new_n385_), .A2(new_n384_), .B(new_n389_), .ZN(new_n390_));
  INV_X1     g0254(.I(new_n390_), .ZN(new_n391_));
  AOI21_X1   g0255(.A1(new_n386_), .A2(new_n381_), .B(new_n389_), .ZN(new_n392_));
  OAI21_X1   g0256(.A1(new_n392_), .A2(new_n391_), .B(\A[50] ), .ZN(new_n393_));
  AOI21_X1   g0257(.A1(new_n393_), .A2(new_n388_), .B(\A[48] ), .ZN(new_n394_));
  INV_X1     g0258(.I(new_n394_), .ZN(new_n395_));
  INV_X1     g0259(.I(\A[49] ), .ZN(new_n396_));
  OAI21_X1   g0260(.A1(new_n392_), .A2(new_n391_), .B(new_n396_), .ZN(new_n397_));
  INV_X1     g0261(.I(new_n397_), .ZN(new_n398_));
  AOI21_X1   g0262(.A1(new_n393_), .A2(new_n388_), .B(new_n396_), .ZN(new_n399_));
  OAI21_X1   g0263(.A1(new_n399_), .A2(new_n398_), .B(\A[48] ), .ZN(new_n400_));
  AOI21_X1   g0264(.A1(new_n400_), .A2(new_n395_), .B(\A[46] ), .ZN(new_n401_));
  INV_X1     g0265(.I(new_n401_), .ZN(new_n402_));
  INV_X1     g0266(.I(\A[47] ), .ZN(new_n403_));
  OAI21_X1   g0267(.A1(new_n399_), .A2(new_n398_), .B(new_n403_), .ZN(new_n404_));
  INV_X1     g0268(.I(new_n404_), .ZN(new_n405_));
  AOI21_X1   g0269(.A1(new_n400_), .A2(new_n395_), .B(new_n403_), .ZN(new_n406_));
  OAI21_X1   g0270(.A1(new_n406_), .A2(new_n405_), .B(\A[46] ), .ZN(new_n407_));
  AOI21_X1   g0271(.A1(new_n407_), .A2(new_n402_), .B(\A[44] ), .ZN(new_n408_));
  INV_X1     g0272(.I(new_n408_), .ZN(new_n409_));
  INV_X1     g0273(.I(\A[45] ), .ZN(new_n410_));
  OAI21_X1   g0274(.A1(new_n406_), .A2(new_n405_), .B(new_n410_), .ZN(new_n411_));
  INV_X1     g0275(.I(new_n411_), .ZN(new_n412_));
  AOI21_X1   g0276(.A1(new_n407_), .A2(new_n402_), .B(new_n410_), .ZN(new_n413_));
  OAI21_X1   g0277(.A1(new_n413_), .A2(new_n412_), .B(\A[44] ), .ZN(new_n414_));
  AOI21_X1   g0278(.A1(new_n414_), .A2(new_n409_), .B(\A[42] ), .ZN(new_n415_));
  INV_X1     g0279(.I(new_n415_), .ZN(new_n416_));
  INV_X1     g0280(.I(\A[43] ), .ZN(new_n417_));
  OAI21_X1   g0281(.A1(new_n413_), .A2(new_n412_), .B(new_n417_), .ZN(new_n418_));
  INV_X1     g0282(.I(new_n418_), .ZN(new_n419_));
  AOI21_X1   g0283(.A1(new_n414_), .A2(new_n409_), .B(new_n417_), .ZN(new_n420_));
  OAI21_X1   g0284(.A1(new_n420_), .A2(new_n419_), .B(\A[42] ), .ZN(new_n421_));
  AOI21_X1   g0285(.A1(new_n421_), .A2(new_n416_), .B(\A[40] ), .ZN(new_n422_));
  INV_X1     g0286(.I(new_n422_), .ZN(new_n423_));
  INV_X1     g0287(.I(\A[41] ), .ZN(new_n424_));
  OAI21_X1   g0288(.A1(new_n420_), .A2(new_n419_), .B(new_n424_), .ZN(new_n425_));
  INV_X1     g0289(.I(new_n425_), .ZN(new_n426_));
  AOI21_X1   g0290(.A1(new_n421_), .A2(new_n416_), .B(new_n424_), .ZN(new_n427_));
  OAI21_X1   g0291(.A1(new_n427_), .A2(new_n426_), .B(\A[40] ), .ZN(new_n428_));
  AOI21_X1   g0292(.A1(new_n428_), .A2(new_n423_), .B(\A[38] ), .ZN(new_n429_));
  INV_X1     g0293(.I(new_n429_), .ZN(new_n430_));
  INV_X1     g0294(.I(\A[39] ), .ZN(new_n431_));
  OAI21_X1   g0295(.A1(new_n427_), .A2(new_n426_), .B(new_n431_), .ZN(new_n432_));
  INV_X1     g0296(.I(new_n432_), .ZN(new_n433_));
  AOI21_X1   g0297(.A1(new_n428_), .A2(new_n423_), .B(new_n431_), .ZN(new_n434_));
  OAI21_X1   g0298(.A1(new_n434_), .A2(new_n433_), .B(\A[38] ), .ZN(new_n435_));
  AOI21_X1   g0299(.A1(new_n435_), .A2(new_n430_), .B(\A[36] ), .ZN(new_n436_));
  INV_X1     g0300(.I(new_n436_), .ZN(new_n437_));
  INV_X1     g0301(.I(\A[37] ), .ZN(new_n438_));
  OAI21_X1   g0302(.A1(new_n434_), .A2(new_n433_), .B(new_n438_), .ZN(new_n439_));
  INV_X1     g0303(.I(new_n439_), .ZN(new_n440_));
  AOI21_X1   g0304(.A1(new_n435_), .A2(new_n430_), .B(new_n438_), .ZN(new_n441_));
  OAI21_X1   g0305(.A1(new_n441_), .A2(new_n440_), .B(\A[36] ), .ZN(new_n442_));
  AOI21_X1   g0306(.A1(new_n442_), .A2(new_n437_), .B(\A[34] ), .ZN(new_n443_));
  INV_X1     g0307(.I(new_n443_), .ZN(new_n444_));
  INV_X1     g0308(.I(\A[35] ), .ZN(new_n445_));
  OAI21_X1   g0309(.A1(new_n441_), .A2(new_n440_), .B(new_n445_), .ZN(new_n446_));
  INV_X1     g0310(.I(new_n446_), .ZN(new_n447_));
  AOI21_X1   g0311(.A1(new_n442_), .A2(new_n437_), .B(new_n445_), .ZN(new_n448_));
  OAI21_X1   g0312(.A1(new_n448_), .A2(new_n447_), .B(\A[34] ), .ZN(new_n449_));
  AOI21_X1   g0313(.A1(new_n449_), .A2(new_n444_), .B(\A[32] ), .ZN(new_n450_));
  INV_X1     g0314(.I(new_n450_), .ZN(new_n451_));
  INV_X1     g0315(.I(\A[33] ), .ZN(new_n452_));
  OAI21_X1   g0316(.A1(new_n448_), .A2(new_n447_), .B(new_n452_), .ZN(new_n453_));
  INV_X1     g0317(.I(new_n453_), .ZN(new_n454_));
  AOI21_X1   g0318(.A1(new_n449_), .A2(new_n444_), .B(new_n452_), .ZN(new_n455_));
  OAI21_X1   g0319(.A1(new_n455_), .A2(new_n454_), .B(\A[32] ), .ZN(new_n456_));
  AOI21_X1   g0320(.A1(new_n456_), .A2(new_n451_), .B(\A[30] ), .ZN(new_n457_));
  INV_X1     g0321(.I(new_n457_), .ZN(new_n458_));
  INV_X1     g0322(.I(\A[31] ), .ZN(new_n459_));
  OAI21_X1   g0323(.A1(new_n455_), .A2(new_n454_), .B(new_n459_), .ZN(new_n460_));
  INV_X1     g0324(.I(new_n460_), .ZN(new_n461_));
  AOI21_X1   g0325(.A1(new_n456_), .A2(new_n451_), .B(new_n459_), .ZN(new_n462_));
  OAI21_X1   g0326(.A1(new_n462_), .A2(new_n461_), .B(\A[30] ), .ZN(new_n463_));
  AOI21_X1   g0327(.A1(new_n463_), .A2(new_n458_), .B(\A[28] ), .ZN(new_n464_));
  INV_X1     g0328(.I(new_n464_), .ZN(new_n465_));
  INV_X1     g0329(.I(\A[29] ), .ZN(new_n466_));
  OAI21_X1   g0330(.A1(new_n462_), .A2(new_n461_), .B(new_n466_), .ZN(new_n467_));
  INV_X1     g0331(.I(new_n467_), .ZN(new_n468_));
  AOI21_X1   g0332(.A1(new_n463_), .A2(new_n458_), .B(new_n466_), .ZN(new_n469_));
  OAI21_X1   g0333(.A1(new_n469_), .A2(new_n468_), .B(\A[28] ), .ZN(new_n470_));
  AOI21_X1   g0334(.A1(new_n470_), .A2(new_n465_), .B(\A[26] ), .ZN(new_n471_));
  INV_X1     g0335(.I(new_n471_), .ZN(new_n472_));
  INV_X1     g0336(.I(\A[27] ), .ZN(new_n473_));
  OAI21_X1   g0337(.A1(new_n469_), .A2(new_n468_), .B(new_n473_), .ZN(new_n474_));
  INV_X1     g0338(.I(new_n474_), .ZN(new_n475_));
  AOI21_X1   g0339(.A1(new_n470_), .A2(new_n465_), .B(new_n473_), .ZN(new_n476_));
  OAI21_X1   g0340(.A1(new_n476_), .A2(new_n475_), .B(\A[26] ), .ZN(new_n477_));
  AOI21_X1   g0341(.A1(new_n477_), .A2(new_n472_), .B(\A[24] ), .ZN(new_n478_));
  INV_X1     g0342(.I(new_n478_), .ZN(new_n479_));
  INV_X1     g0343(.I(\A[25] ), .ZN(new_n480_));
  OAI21_X1   g0344(.A1(new_n476_), .A2(new_n475_), .B(new_n480_), .ZN(new_n481_));
  INV_X1     g0345(.I(new_n481_), .ZN(new_n482_));
  AOI21_X1   g0346(.A1(new_n477_), .A2(new_n472_), .B(new_n480_), .ZN(new_n483_));
  OAI21_X1   g0347(.A1(new_n483_), .A2(new_n482_), .B(\A[24] ), .ZN(new_n484_));
  AOI21_X1   g0348(.A1(new_n484_), .A2(new_n479_), .B(\A[22] ), .ZN(new_n485_));
  INV_X1     g0349(.I(new_n485_), .ZN(new_n486_));
  INV_X1     g0350(.I(\A[23] ), .ZN(new_n487_));
  OAI21_X1   g0351(.A1(new_n483_), .A2(new_n482_), .B(new_n487_), .ZN(new_n488_));
  INV_X1     g0352(.I(new_n488_), .ZN(new_n489_));
  AOI21_X1   g0353(.A1(new_n484_), .A2(new_n479_), .B(new_n487_), .ZN(new_n490_));
  OAI21_X1   g0354(.A1(new_n490_), .A2(new_n489_), .B(\A[22] ), .ZN(new_n491_));
  AOI21_X1   g0355(.A1(new_n491_), .A2(new_n486_), .B(\A[20] ), .ZN(new_n492_));
  INV_X1     g0356(.I(new_n492_), .ZN(new_n493_));
  INV_X1     g0357(.I(\A[21] ), .ZN(new_n494_));
  OAI21_X1   g0358(.A1(new_n490_), .A2(new_n489_), .B(new_n494_), .ZN(new_n495_));
  INV_X1     g0359(.I(new_n495_), .ZN(new_n496_));
  AOI21_X1   g0360(.A1(new_n491_), .A2(new_n486_), .B(new_n494_), .ZN(new_n497_));
  OAI21_X1   g0361(.A1(new_n497_), .A2(new_n496_), .B(\A[20] ), .ZN(new_n498_));
  AOI21_X1   g0362(.A1(new_n498_), .A2(new_n493_), .B(\A[18] ), .ZN(new_n499_));
  INV_X1     g0363(.I(new_n499_), .ZN(new_n500_));
  INV_X1     g0364(.I(\A[19] ), .ZN(new_n501_));
  OAI21_X1   g0365(.A1(new_n497_), .A2(new_n496_), .B(new_n501_), .ZN(new_n502_));
  INV_X1     g0366(.I(new_n502_), .ZN(new_n503_));
  AOI21_X1   g0367(.A1(new_n498_), .A2(new_n493_), .B(new_n501_), .ZN(new_n504_));
  OAI21_X1   g0368(.A1(new_n504_), .A2(new_n503_), .B(\A[18] ), .ZN(new_n505_));
  AOI21_X1   g0369(.A1(new_n505_), .A2(new_n500_), .B(\A[16] ), .ZN(new_n506_));
  INV_X1     g0370(.I(new_n506_), .ZN(new_n507_));
  INV_X1     g0371(.I(\A[17] ), .ZN(new_n508_));
  OAI21_X1   g0372(.A1(new_n504_), .A2(new_n503_), .B(new_n508_), .ZN(new_n509_));
  INV_X1     g0373(.I(new_n509_), .ZN(new_n510_));
  AOI21_X1   g0374(.A1(new_n505_), .A2(new_n500_), .B(new_n508_), .ZN(new_n511_));
  OAI21_X1   g0375(.A1(new_n511_), .A2(new_n510_), .B(\A[16] ), .ZN(new_n512_));
  AOI21_X1   g0376(.A1(new_n512_), .A2(new_n507_), .B(\A[14] ), .ZN(new_n513_));
  INV_X1     g0377(.I(new_n513_), .ZN(new_n514_));
  INV_X1     g0378(.I(\A[15] ), .ZN(new_n515_));
  OAI21_X1   g0379(.A1(new_n511_), .A2(new_n510_), .B(new_n515_), .ZN(new_n516_));
  INV_X1     g0380(.I(new_n516_), .ZN(new_n517_));
  AOI21_X1   g0381(.A1(new_n512_), .A2(new_n507_), .B(new_n515_), .ZN(new_n518_));
  OAI21_X1   g0382(.A1(new_n518_), .A2(new_n517_), .B(\A[14] ), .ZN(new_n519_));
  AOI21_X1   g0383(.A1(new_n519_), .A2(new_n514_), .B(\A[12] ), .ZN(new_n520_));
  INV_X1     g0384(.I(new_n520_), .ZN(new_n521_));
  INV_X1     g0385(.I(\A[13] ), .ZN(new_n522_));
  OAI21_X1   g0386(.A1(new_n518_), .A2(new_n517_), .B(new_n522_), .ZN(new_n523_));
  INV_X1     g0387(.I(new_n523_), .ZN(new_n524_));
  AOI21_X1   g0388(.A1(new_n519_), .A2(new_n514_), .B(new_n522_), .ZN(new_n525_));
  OAI21_X1   g0389(.A1(new_n525_), .A2(new_n524_), .B(\A[12] ), .ZN(new_n526_));
  AOI21_X1   g0390(.A1(new_n526_), .A2(new_n521_), .B(\A[10] ), .ZN(new_n527_));
  INV_X1     g0391(.I(new_n527_), .ZN(new_n528_));
  INV_X1     g0392(.I(\A[11] ), .ZN(new_n529_));
  OAI21_X1   g0393(.A1(new_n525_), .A2(new_n524_), .B(new_n529_), .ZN(new_n530_));
  INV_X1     g0394(.I(new_n530_), .ZN(new_n531_));
  AOI21_X1   g0395(.A1(new_n526_), .A2(new_n521_), .B(new_n529_), .ZN(new_n532_));
  OAI21_X1   g0396(.A1(new_n532_), .A2(new_n531_), .B(\A[10] ), .ZN(new_n533_));
  AOI21_X1   g0397(.A1(new_n533_), .A2(new_n528_), .B(\A[8] ), .ZN(new_n534_));
  INV_X1     g0398(.I(new_n534_), .ZN(new_n535_));
  INV_X1     g0399(.I(\A[9] ), .ZN(new_n536_));
  OAI21_X1   g0400(.A1(new_n532_), .A2(new_n531_), .B(new_n536_), .ZN(new_n537_));
  INV_X1     g0401(.I(new_n537_), .ZN(new_n538_));
  AOI21_X1   g0402(.A1(new_n533_), .A2(new_n528_), .B(new_n536_), .ZN(new_n539_));
  OAI21_X1   g0403(.A1(new_n539_), .A2(new_n538_), .B(\A[8] ), .ZN(new_n540_));
  AOI21_X1   g0404(.A1(new_n540_), .A2(new_n535_), .B(\A[6] ), .ZN(new_n541_));
  INV_X1     g0405(.I(new_n541_), .ZN(new_n542_));
  INV_X1     g0406(.I(\A[7] ), .ZN(new_n543_));
  OAI21_X1   g0407(.A1(new_n539_), .A2(new_n538_), .B(new_n543_), .ZN(new_n544_));
  INV_X1     g0408(.I(new_n544_), .ZN(new_n545_));
  AOI21_X1   g0409(.A1(new_n540_), .A2(new_n535_), .B(new_n543_), .ZN(new_n546_));
  OAI21_X1   g0410(.A1(new_n546_), .A2(new_n545_), .B(\A[6] ), .ZN(new_n547_));
  AOI21_X1   g0411(.A1(new_n547_), .A2(new_n542_), .B(\A[4] ), .ZN(new_n548_));
  INV_X1     g0412(.I(\A[5] ), .ZN(new_n549_));
  AOI21_X1   g0413(.A1(new_n168_), .A2(\A[114] ), .B(new_n163_), .ZN(new_n550_));
  OAI21_X1   g0414(.A1(new_n550_), .A2(new_n172_), .B(new_n173_), .ZN(new_n551_));
  AOI21_X1   g0415(.A1(new_n551_), .A2(\A[112] ), .B(new_n170_), .ZN(new_n552_));
  OAI21_X1   g0416(.A1(new_n552_), .A2(new_n179_), .B(new_n180_), .ZN(new_n553_));
  AOI21_X1   g0417(.A1(new_n553_), .A2(\A[110] ), .B(new_n177_), .ZN(new_n554_));
  OAI21_X1   g0418(.A1(new_n554_), .A2(new_n186_), .B(new_n187_), .ZN(new_n555_));
  AOI21_X1   g0419(.A1(new_n555_), .A2(\A[108] ), .B(new_n184_), .ZN(new_n556_));
  OAI21_X1   g0420(.A1(new_n556_), .A2(new_n193_), .B(new_n194_), .ZN(new_n557_));
  AOI21_X1   g0421(.A1(new_n557_), .A2(\A[106] ), .B(new_n191_), .ZN(new_n558_));
  OAI21_X1   g0422(.A1(new_n558_), .A2(new_n200_), .B(new_n201_), .ZN(new_n559_));
  AOI21_X1   g0423(.A1(new_n559_), .A2(\A[104] ), .B(new_n198_), .ZN(new_n560_));
  OAI21_X1   g0424(.A1(new_n560_), .A2(new_n207_), .B(new_n208_), .ZN(new_n561_));
  AOI21_X1   g0425(.A1(new_n561_), .A2(\A[102] ), .B(new_n205_), .ZN(new_n562_));
  OAI21_X1   g0426(.A1(new_n562_), .A2(new_n214_), .B(new_n215_), .ZN(new_n563_));
  AOI21_X1   g0427(.A1(new_n563_), .A2(\A[100] ), .B(new_n212_), .ZN(new_n564_));
  OAI21_X1   g0428(.A1(new_n564_), .A2(new_n221_), .B(new_n222_), .ZN(new_n565_));
  AOI21_X1   g0429(.A1(new_n565_), .A2(\A[98] ), .B(new_n219_), .ZN(new_n566_));
  OAI21_X1   g0430(.A1(new_n566_), .A2(new_n228_), .B(new_n229_), .ZN(new_n567_));
  AOI21_X1   g0431(.A1(new_n567_), .A2(\A[96] ), .B(new_n226_), .ZN(new_n568_));
  OAI21_X1   g0432(.A1(new_n568_), .A2(new_n235_), .B(new_n236_), .ZN(new_n569_));
  AOI21_X1   g0433(.A1(new_n569_), .A2(\A[94] ), .B(new_n233_), .ZN(new_n570_));
  OAI21_X1   g0434(.A1(new_n570_), .A2(new_n242_), .B(new_n243_), .ZN(new_n571_));
  AOI21_X1   g0435(.A1(new_n571_), .A2(\A[92] ), .B(new_n240_), .ZN(new_n572_));
  OAI21_X1   g0436(.A1(new_n572_), .A2(new_n249_), .B(new_n250_), .ZN(new_n573_));
  AOI21_X1   g0437(.A1(new_n573_), .A2(\A[90] ), .B(new_n247_), .ZN(new_n574_));
  OAI21_X1   g0438(.A1(new_n574_), .A2(new_n256_), .B(new_n257_), .ZN(new_n575_));
  AOI21_X1   g0439(.A1(new_n575_), .A2(\A[88] ), .B(new_n254_), .ZN(new_n576_));
  OAI21_X1   g0440(.A1(new_n576_), .A2(new_n263_), .B(new_n264_), .ZN(new_n577_));
  AOI21_X1   g0441(.A1(new_n577_), .A2(\A[86] ), .B(new_n261_), .ZN(new_n578_));
  OAI21_X1   g0442(.A1(new_n578_), .A2(new_n270_), .B(new_n271_), .ZN(new_n579_));
  AOI21_X1   g0443(.A1(new_n579_), .A2(\A[84] ), .B(new_n268_), .ZN(new_n580_));
  OAI21_X1   g0444(.A1(new_n580_), .A2(new_n277_), .B(new_n278_), .ZN(new_n581_));
  AOI21_X1   g0445(.A1(new_n581_), .A2(\A[82] ), .B(new_n275_), .ZN(new_n582_));
  OAI21_X1   g0446(.A1(new_n582_), .A2(new_n284_), .B(new_n285_), .ZN(new_n583_));
  AOI21_X1   g0447(.A1(new_n583_), .A2(\A[80] ), .B(new_n282_), .ZN(new_n584_));
  OAI21_X1   g0448(.A1(new_n584_), .A2(new_n291_), .B(new_n292_), .ZN(new_n585_));
  AOI21_X1   g0449(.A1(new_n585_), .A2(\A[78] ), .B(new_n289_), .ZN(new_n586_));
  OAI21_X1   g0450(.A1(new_n586_), .A2(new_n298_), .B(new_n299_), .ZN(new_n587_));
  AOI21_X1   g0451(.A1(new_n587_), .A2(\A[76] ), .B(new_n296_), .ZN(new_n588_));
  OAI21_X1   g0452(.A1(new_n588_), .A2(new_n305_), .B(new_n306_), .ZN(new_n589_));
  AOI21_X1   g0453(.A1(new_n589_), .A2(\A[74] ), .B(new_n303_), .ZN(new_n590_));
  OAI21_X1   g0454(.A1(new_n590_), .A2(new_n312_), .B(new_n313_), .ZN(new_n591_));
  AOI21_X1   g0455(.A1(new_n591_), .A2(\A[72] ), .B(new_n310_), .ZN(new_n592_));
  OAI21_X1   g0456(.A1(new_n592_), .A2(new_n319_), .B(new_n320_), .ZN(new_n593_));
  AOI21_X1   g0457(.A1(new_n593_), .A2(\A[70] ), .B(new_n317_), .ZN(new_n594_));
  OAI21_X1   g0458(.A1(new_n594_), .A2(new_n326_), .B(new_n327_), .ZN(new_n595_));
  AOI21_X1   g0459(.A1(new_n595_), .A2(\A[68] ), .B(new_n324_), .ZN(new_n596_));
  OAI21_X1   g0460(.A1(new_n596_), .A2(new_n333_), .B(new_n334_), .ZN(new_n597_));
  AOI21_X1   g0461(.A1(new_n597_), .A2(\A[66] ), .B(new_n331_), .ZN(new_n598_));
  OAI21_X1   g0462(.A1(new_n598_), .A2(new_n340_), .B(new_n341_), .ZN(new_n599_));
  AOI21_X1   g0463(.A1(new_n599_), .A2(\A[64] ), .B(new_n338_), .ZN(new_n600_));
  OAI21_X1   g0464(.A1(new_n600_), .A2(new_n347_), .B(new_n348_), .ZN(new_n601_));
  AOI21_X1   g0465(.A1(new_n601_), .A2(\A[62] ), .B(new_n345_), .ZN(new_n602_));
  OAI21_X1   g0466(.A1(new_n602_), .A2(new_n354_), .B(new_n355_), .ZN(new_n603_));
  AOI21_X1   g0467(.A1(new_n603_), .A2(\A[60] ), .B(new_n352_), .ZN(new_n604_));
  OAI21_X1   g0468(.A1(new_n604_), .A2(new_n361_), .B(new_n362_), .ZN(new_n605_));
  AOI21_X1   g0469(.A1(new_n605_), .A2(\A[58] ), .B(new_n359_), .ZN(new_n606_));
  OAI21_X1   g0470(.A1(new_n606_), .A2(new_n368_), .B(new_n369_), .ZN(new_n607_));
  AOI21_X1   g0471(.A1(new_n607_), .A2(\A[56] ), .B(new_n366_), .ZN(new_n608_));
  OAI21_X1   g0472(.A1(new_n608_), .A2(new_n375_), .B(new_n376_), .ZN(new_n609_));
  AOI21_X1   g0473(.A1(new_n609_), .A2(\A[54] ), .B(new_n373_), .ZN(new_n610_));
  OAI21_X1   g0474(.A1(new_n610_), .A2(new_n382_), .B(new_n383_), .ZN(new_n611_));
  AOI21_X1   g0475(.A1(new_n611_), .A2(\A[52] ), .B(new_n380_), .ZN(new_n612_));
  OAI21_X1   g0476(.A1(new_n612_), .A2(new_n389_), .B(new_n390_), .ZN(new_n613_));
  AOI21_X1   g0477(.A1(new_n613_), .A2(\A[50] ), .B(new_n387_), .ZN(new_n614_));
  OAI21_X1   g0478(.A1(new_n614_), .A2(new_n396_), .B(new_n397_), .ZN(new_n615_));
  AOI21_X1   g0479(.A1(new_n615_), .A2(\A[48] ), .B(new_n394_), .ZN(new_n616_));
  OAI21_X1   g0480(.A1(new_n616_), .A2(new_n403_), .B(new_n404_), .ZN(new_n617_));
  AOI21_X1   g0481(.A1(new_n617_), .A2(\A[46] ), .B(new_n401_), .ZN(new_n618_));
  OAI21_X1   g0482(.A1(new_n618_), .A2(new_n410_), .B(new_n411_), .ZN(new_n619_));
  AOI21_X1   g0483(.A1(new_n619_), .A2(\A[44] ), .B(new_n408_), .ZN(new_n620_));
  OAI21_X1   g0484(.A1(new_n620_), .A2(new_n417_), .B(new_n418_), .ZN(new_n621_));
  AOI21_X1   g0485(.A1(new_n621_), .A2(\A[42] ), .B(new_n415_), .ZN(new_n622_));
  OAI21_X1   g0486(.A1(new_n622_), .A2(new_n424_), .B(new_n425_), .ZN(new_n623_));
  AOI21_X1   g0487(.A1(new_n623_), .A2(\A[40] ), .B(new_n422_), .ZN(new_n624_));
  OAI21_X1   g0488(.A1(new_n624_), .A2(new_n431_), .B(new_n432_), .ZN(new_n625_));
  AOI21_X1   g0489(.A1(new_n625_), .A2(\A[38] ), .B(new_n429_), .ZN(new_n626_));
  OAI21_X1   g0490(.A1(new_n626_), .A2(new_n438_), .B(new_n439_), .ZN(new_n627_));
  AOI21_X1   g0491(.A1(new_n627_), .A2(\A[36] ), .B(new_n436_), .ZN(new_n628_));
  OAI21_X1   g0492(.A1(new_n628_), .A2(new_n445_), .B(new_n446_), .ZN(new_n629_));
  AOI21_X1   g0493(.A1(new_n629_), .A2(\A[34] ), .B(new_n443_), .ZN(new_n630_));
  OAI21_X1   g0494(.A1(new_n630_), .A2(new_n452_), .B(new_n453_), .ZN(new_n631_));
  AOI21_X1   g0495(.A1(new_n631_), .A2(\A[32] ), .B(new_n450_), .ZN(new_n632_));
  OAI21_X1   g0496(.A1(new_n632_), .A2(new_n459_), .B(new_n460_), .ZN(new_n633_));
  AOI21_X1   g0497(.A1(new_n633_), .A2(\A[30] ), .B(new_n457_), .ZN(new_n634_));
  OAI21_X1   g0498(.A1(new_n634_), .A2(new_n466_), .B(new_n467_), .ZN(new_n635_));
  AOI21_X1   g0499(.A1(new_n635_), .A2(\A[28] ), .B(new_n464_), .ZN(new_n636_));
  OAI21_X1   g0500(.A1(new_n636_), .A2(new_n473_), .B(new_n474_), .ZN(new_n637_));
  AOI21_X1   g0501(.A1(new_n637_), .A2(\A[26] ), .B(new_n471_), .ZN(new_n638_));
  OAI21_X1   g0502(.A1(new_n638_), .A2(new_n480_), .B(new_n481_), .ZN(new_n639_));
  AOI21_X1   g0503(.A1(new_n639_), .A2(\A[24] ), .B(new_n478_), .ZN(new_n640_));
  OAI21_X1   g0504(.A1(new_n640_), .A2(new_n487_), .B(new_n488_), .ZN(new_n641_));
  AOI21_X1   g0505(.A1(new_n641_), .A2(\A[22] ), .B(new_n485_), .ZN(new_n642_));
  OAI21_X1   g0506(.A1(new_n642_), .A2(new_n494_), .B(new_n495_), .ZN(new_n643_));
  AOI21_X1   g0507(.A1(new_n643_), .A2(\A[20] ), .B(new_n492_), .ZN(new_n644_));
  OAI21_X1   g0508(.A1(new_n644_), .A2(new_n501_), .B(new_n502_), .ZN(new_n645_));
  AOI21_X1   g0509(.A1(new_n645_), .A2(\A[18] ), .B(new_n499_), .ZN(new_n646_));
  OAI21_X1   g0510(.A1(new_n646_), .A2(new_n508_), .B(new_n509_), .ZN(new_n647_));
  AOI21_X1   g0511(.A1(new_n647_), .A2(\A[16] ), .B(new_n506_), .ZN(new_n648_));
  OAI21_X1   g0512(.A1(new_n648_), .A2(new_n515_), .B(new_n516_), .ZN(new_n649_));
  AOI21_X1   g0513(.A1(new_n649_), .A2(\A[14] ), .B(new_n513_), .ZN(new_n650_));
  OAI21_X1   g0514(.A1(new_n650_), .A2(new_n522_), .B(new_n523_), .ZN(new_n651_));
  AOI21_X1   g0515(.A1(new_n651_), .A2(\A[12] ), .B(new_n520_), .ZN(new_n652_));
  OAI21_X1   g0516(.A1(new_n652_), .A2(new_n529_), .B(new_n530_), .ZN(new_n653_));
  AOI21_X1   g0517(.A1(new_n653_), .A2(\A[10] ), .B(new_n527_), .ZN(new_n654_));
  OAI21_X1   g0518(.A1(new_n654_), .A2(new_n536_), .B(new_n537_), .ZN(new_n655_));
  AOI21_X1   g0519(.A1(new_n655_), .A2(\A[8] ), .B(new_n534_), .ZN(new_n656_));
  OAI21_X1   g0520(.A1(new_n656_), .A2(new_n543_), .B(new_n544_), .ZN(new_n657_));
  AOI21_X1   g0521(.A1(new_n657_), .A2(\A[6] ), .B(new_n541_), .ZN(new_n658_));
  OAI21_X1   g0522(.A1(new_n546_), .A2(new_n545_), .B(new_n549_), .ZN(new_n659_));
  OAI21_X1   g0523(.A1(new_n658_), .A2(new_n549_), .B(new_n659_), .ZN(new_n660_));
  AOI21_X1   g0524(.A1(new_n660_), .A2(\A[4] ), .B(new_n548_), .ZN(new_n661_));
  INV_X1     g0525(.I(\A[1] ), .ZN(new_n662_));
  NOR2_X1    g0526(.A1(new_n662_), .A2(\A[2] ), .ZN(new_n663_));
  INV_X1     g0527(.I(\A[4] ), .ZN(new_n664_));
  INV_X1     g0528(.I(\A[6] ), .ZN(new_n665_));
  INV_X1     g0529(.I(\A[8] ), .ZN(new_n666_));
  INV_X1     g0530(.I(\A[10] ), .ZN(new_n667_));
  INV_X1     g0531(.I(\A[12] ), .ZN(new_n668_));
  INV_X1     g0532(.I(\A[14] ), .ZN(new_n669_));
  INV_X1     g0533(.I(\A[16] ), .ZN(new_n670_));
  INV_X1     g0534(.I(\A[18] ), .ZN(new_n671_));
  INV_X1     g0535(.I(\A[20] ), .ZN(new_n672_));
  INV_X1     g0536(.I(\A[22] ), .ZN(new_n673_));
  INV_X1     g0537(.I(\A[24] ), .ZN(new_n674_));
  INV_X1     g0538(.I(\A[26] ), .ZN(new_n675_));
  INV_X1     g0539(.I(\A[28] ), .ZN(new_n676_));
  INV_X1     g0540(.I(\A[30] ), .ZN(new_n677_));
  INV_X1     g0541(.I(\A[32] ), .ZN(new_n678_));
  INV_X1     g0542(.I(\A[34] ), .ZN(new_n679_));
  INV_X1     g0543(.I(\A[36] ), .ZN(new_n680_));
  INV_X1     g0544(.I(\A[38] ), .ZN(new_n681_));
  INV_X1     g0545(.I(\A[40] ), .ZN(new_n682_));
  INV_X1     g0546(.I(\A[42] ), .ZN(new_n683_));
  INV_X1     g0547(.I(\A[44] ), .ZN(new_n684_));
  INV_X1     g0548(.I(\A[46] ), .ZN(new_n685_));
  INV_X1     g0549(.I(\A[48] ), .ZN(new_n686_));
  INV_X1     g0550(.I(\A[50] ), .ZN(new_n687_));
  INV_X1     g0551(.I(\A[52] ), .ZN(new_n688_));
  INV_X1     g0552(.I(\A[54] ), .ZN(new_n689_));
  INV_X1     g0553(.I(\A[56] ), .ZN(new_n690_));
  INV_X1     g0554(.I(\A[58] ), .ZN(new_n691_));
  INV_X1     g0555(.I(\A[60] ), .ZN(new_n692_));
  INV_X1     g0556(.I(\A[62] ), .ZN(new_n693_));
  INV_X1     g0557(.I(\A[64] ), .ZN(new_n694_));
  INV_X1     g0558(.I(\A[66] ), .ZN(new_n695_));
  INV_X1     g0559(.I(\A[68] ), .ZN(new_n696_));
  INV_X1     g0560(.I(\A[70] ), .ZN(new_n697_));
  INV_X1     g0561(.I(\A[72] ), .ZN(new_n698_));
  INV_X1     g0562(.I(\A[74] ), .ZN(new_n699_));
  INV_X1     g0563(.I(\A[76] ), .ZN(new_n700_));
  INV_X1     g0564(.I(\A[78] ), .ZN(new_n701_));
  INV_X1     g0565(.I(\A[80] ), .ZN(new_n702_));
  INV_X1     g0566(.I(\A[82] ), .ZN(new_n703_));
  INV_X1     g0567(.I(\A[84] ), .ZN(new_n704_));
  INV_X1     g0568(.I(\A[86] ), .ZN(new_n705_));
  INV_X1     g0569(.I(\A[88] ), .ZN(new_n706_));
  INV_X1     g0570(.I(\A[90] ), .ZN(new_n707_));
  INV_X1     g0571(.I(\A[92] ), .ZN(new_n708_));
  INV_X1     g0572(.I(\A[94] ), .ZN(new_n709_));
  INV_X1     g0573(.I(\A[96] ), .ZN(new_n710_));
  INV_X1     g0574(.I(\A[98] ), .ZN(new_n711_));
  INV_X1     g0575(.I(\A[100] ), .ZN(new_n712_));
  INV_X1     g0576(.I(\A[102] ), .ZN(new_n713_));
  INV_X1     g0577(.I(\A[104] ), .ZN(new_n714_));
  INV_X1     g0578(.I(\A[106] ), .ZN(new_n715_));
  INV_X1     g0579(.I(\A[108] ), .ZN(new_n716_));
  INV_X1     g0580(.I(\A[110] ), .ZN(new_n717_));
  INV_X1     g0581(.I(\A[112] ), .ZN(new_n718_));
  INV_X1     g0582(.I(\A[114] ), .ZN(new_n719_));
  INV_X1     g0583(.I(\A[116] ), .ZN(new_n720_));
  INV_X1     g0584(.I(\A[118] ), .ZN(new_n721_));
  INV_X1     g0585(.I(\A[120] ), .ZN(new_n722_));
  INV_X1     g0586(.I(\A[122] ), .ZN(new_n723_));
  INV_X1     g0587(.I(\A[124] ), .ZN(new_n724_));
  INV_X1     g0588(.I(\A[126] ), .ZN(new_n725_));
  AOI21_X1   g0589(.A1(new_n725_), .A2(\A[125] ), .B(\A[127] ), .ZN(new_n726_));
  NOR2_X1    g0590(.A1(new_n726_), .A2(new_n724_), .ZN(new_n727_));
  OAI21_X1   g0591(.A1(new_n727_), .A2(new_n138_), .B(\A[123] ), .ZN(new_n728_));
  AOI21_X1   g0592(.A1(new_n728_), .A2(new_n144_), .B(new_n723_), .ZN(new_n729_));
  OAI21_X1   g0593(.A1(new_n729_), .A2(new_n142_), .B(\A[121] ), .ZN(new_n730_));
  AOI21_X1   g0594(.A1(new_n730_), .A2(new_n149_), .B(new_n722_), .ZN(new_n731_));
  OAI21_X1   g0595(.A1(new_n731_), .A2(new_n147_), .B(\A[119] ), .ZN(new_n732_));
  AOI21_X1   g0596(.A1(new_n732_), .A2(new_n154_), .B(new_n721_), .ZN(new_n733_));
  OAI21_X1   g0597(.A1(new_n733_), .A2(new_n152_), .B(\A[117] ), .ZN(new_n734_));
  AOI21_X1   g0598(.A1(new_n734_), .A2(new_n160_), .B(new_n720_), .ZN(new_n735_));
  OAI21_X1   g0599(.A1(new_n735_), .A2(new_n157_), .B(\A[115] ), .ZN(new_n736_));
  AOI21_X1   g0600(.A1(new_n736_), .A2(new_n167_), .B(new_n719_), .ZN(new_n737_));
  OAI21_X1   g0601(.A1(new_n737_), .A2(new_n163_), .B(\A[113] ), .ZN(new_n738_));
  AOI21_X1   g0602(.A1(new_n738_), .A2(new_n173_), .B(new_n718_), .ZN(new_n739_));
  OAI21_X1   g0603(.A1(new_n739_), .A2(new_n170_), .B(\A[111] ), .ZN(new_n740_));
  AOI21_X1   g0604(.A1(new_n740_), .A2(new_n180_), .B(new_n717_), .ZN(new_n741_));
  OAI21_X1   g0605(.A1(new_n741_), .A2(new_n177_), .B(\A[109] ), .ZN(new_n742_));
  AOI21_X1   g0606(.A1(new_n742_), .A2(new_n187_), .B(new_n716_), .ZN(new_n743_));
  OAI21_X1   g0607(.A1(new_n743_), .A2(new_n184_), .B(\A[107] ), .ZN(new_n744_));
  AOI21_X1   g0608(.A1(new_n744_), .A2(new_n194_), .B(new_n715_), .ZN(new_n745_));
  OAI21_X1   g0609(.A1(new_n745_), .A2(new_n191_), .B(\A[105] ), .ZN(new_n746_));
  AOI21_X1   g0610(.A1(new_n746_), .A2(new_n201_), .B(new_n714_), .ZN(new_n747_));
  OAI21_X1   g0611(.A1(new_n747_), .A2(new_n198_), .B(\A[103] ), .ZN(new_n748_));
  AOI21_X1   g0612(.A1(new_n748_), .A2(new_n208_), .B(new_n713_), .ZN(new_n749_));
  OAI21_X1   g0613(.A1(new_n749_), .A2(new_n205_), .B(\A[101] ), .ZN(new_n750_));
  AOI21_X1   g0614(.A1(new_n750_), .A2(new_n215_), .B(new_n712_), .ZN(new_n751_));
  OAI21_X1   g0615(.A1(new_n751_), .A2(new_n212_), .B(\A[99] ), .ZN(new_n752_));
  AOI21_X1   g0616(.A1(new_n752_), .A2(new_n222_), .B(new_n711_), .ZN(new_n753_));
  OAI21_X1   g0617(.A1(new_n753_), .A2(new_n219_), .B(\A[97] ), .ZN(new_n754_));
  AOI21_X1   g0618(.A1(new_n754_), .A2(new_n229_), .B(new_n710_), .ZN(new_n755_));
  OAI21_X1   g0619(.A1(new_n755_), .A2(new_n226_), .B(\A[95] ), .ZN(new_n756_));
  AOI21_X1   g0620(.A1(new_n756_), .A2(new_n236_), .B(new_n709_), .ZN(new_n757_));
  OAI21_X1   g0621(.A1(new_n757_), .A2(new_n233_), .B(\A[93] ), .ZN(new_n758_));
  AOI21_X1   g0622(.A1(new_n758_), .A2(new_n243_), .B(new_n708_), .ZN(new_n759_));
  OAI21_X1   g0623(.A1(new_n759_), .A2(new_n240_), .B(\A[91] ), .ZN(new_n760_));
  AOI21_X1   g0624(.A1(new_n760_), .A2(new_n250_), .B(new_n707_), .ZN(new_n761_));
  OAI21_X1   g0625(.A1(new_n761_), .A2(new_n247_), .B(\A[89] ), .ZN(new_n762_));
  AOI21_X1   g0626(.A1(new_n762_), .A2(new_n257_), .B(new_n706_), .ZN(new_n763_));
  OAI21_X1   g0627(.A1(new_n763_), .A2(new_n254_), .B(\A[87] ), .ZN(new_n764_));
  AOI21_X1   g0628(.A1(new_n764_), .A2(new_n264_), .B(new_n705_), .ZN(new_n765_));
  OAI21_X1   g0629(.A1(new_n765_), .A2(new_n261_), .B(\A[85] ), .ZN(new_n766_));
  AOI21_X1   g0630(.A1(new_n766_), .A2(new_n271_), .B(new_n704_), .ZN(new_n767_));
  OAI21_X1   g0631(.A1(new_n767_), .A2(new_n268_), .B(\A[83] ), .ZN(new_n768_));
  AOI21_X1   g0632(.A1(new_n768_), .A2(new_n278_), .B(new_n703_), .ZN(new_n769_));
  OAI21_X1   g0633(.A1(new_n769_), .A2(new_n275_), .B(\A[81] ), .ZN(new_n770_));
  AOI21_X1   g0634(.A1(new_n770_), .A2(new_n285_), .B(new_n702_), .ZN(new_n771_));
  OAI21_X1   g0635(.A1(new_n771_), .A2(new_n282_), .B(\A[79] ), .ZN(new_n772_));
  AOI21_X1   g0636(.A1(new_n772_), .A2(new_n292_), .B(new_n701_), .ZN(new_n773_));
  OAI21_X1   g0637(.A1(new_n773_), .A2(new_n289_), .B(\A[77] ), .ZN(new_n774_));
  AOI21_X1   g0638(.A1(new_n774_), .A2(new_n299_), .B(new_n700_), .ZN(new_n775_));
  OAI21_X1   g0639(.A1(new_n775_), .A2(new_n296_), .B(\A[75] ), .ZN(new_n776_));
  AOI21_X1   g0640(.A1(new_n776_), .A2(new_n306_), .B(new_n699_), .ZN(new_n777_));
  OAI21_X1   g0641(.A1(new_n777_), .A2(new_n303_), .B(\A[73] ), .ZN(new_n778_));
  AOI21_X1   g0642(.A1(new_n778_), .A2(new_n313_), .B(new_n698_), .ZN(new_n779_));
  OAI21_X1   g0643(.A1(new_n779_), .A2(new_n310_), .B(\A[71] ), .ZN(new_n780_));
  AOI21_X1   g0644(.A1(new_n780_), .A2(new_n320_), .B(new_n697_), .ZN(new_n781_));
  OAI21_X1   g0645(.A1(new_n781_), .A2(new_n317_), .B(\A[69] ), .ZN(new_n782_));
  AOI21_X1   g0646(.A1(new_n782_), .A2(new_n327_), .B(new_n696_), .ZN(new_n783_));
  OAI21_X1   g0647(.A1(new_n783_), .A2(new_n324_), .B(\A[67] ), .ZN(new_n784_));
  AOI21_X1   g0648(.A1(new_n784_), .A2(new_n334_), .B(new_n695_), .ZN(new_n785_));
  OAI21_X1   g0649(.A1(new_n785_), .A2(new_n331_), .B(\A[65] ), .ZN(new_n786_));
  AOI21_X1   g0650(.A1(new_n786_), .A2(new_n341_), .B(new_n694_), .ZN(new_n787_));
  OAI21_X1   g0651(.A1(new_n787_), .A2(new_n338_), .B(\A[63] ), .ZN(new_n788_));
  AOI21_X1   g0652(.A1(new_n788_), .A2(new_n348_), .B(new_n693_), .ZN(new_n789_));
  OAI21_X1   g0653(.A1(new_n789_), .A2(new_n345_), .B(\A[61] ), .ZN(new_n790_));
  AOI21_X1   g0654(.A1(new_n790_), .A2(new_n355_), .B(new_n692_), .ZN(new_n791_));
  OAI21_X1   g0655(.A1(new_n791_), .A2(new_n352_), .B(\A[59] ), .ZN(new_n792_));
  AOI21_X1   g0656(.A1(new_n792_), .A2(new_n362_), .B(new_n691_), .ZN(new_n793_));
  OAI21_X1   g0657(.A1(new_n793_), .A2(new_n359_), .B(\A[57] ), .ZN(new_n794_));
  AOI21_X1   g0658(.A1(new_n794_), .A2(new_n369_), .B(new_n690_), .ZN(new_n795_));
  OAI21_X1   g0659(.A1(new_n795_), .A2(new_n366_), .B(\A[55] ), .ZN(new_n796_));
  AOI21_X1   g0660(.A1(new_n796_), .A2(new_n376_), .B(new_n689_), .ZN(new_n797_));
  OAI21_X1   g0661(.A1(new_n797_), .A2(new_n373_), .B(\A[53] ), .ZN(new_n798_));
  AOI21_X1   g0662(.A1(new_n798_), .A2(new_n383_), .B(new_n688_), .ZN(new_n799_));
  OAI21_X1   g0663(.A1(new_n799_), .A2(new_n380_), .B(\A[51] ), .ZN(new_n800_));
  AOI21_X1   g0664(.A1(new_n800_), .A2(new_n390_), .B(new_n687_), .ZN(new_n801_));
  OAI21_X1   g0665(.A1(new_n801_), .A2(new_n387_), .B(\A[49] ), .ZN(new_n802_));
  AOI21_X1   g0666(.A1(new_n802_), .A2(new_n397_), .B(new_n686_), .ZN(new_n803_));
  OAI21_X1   g0667(.A1(new_n803_), .A2(new_n394_), .B(\A[47] ), .ZN(new_n804_));
  AOI21_X1   g0668(.A1(new_n804_), .A2(new_n404_), .B(new_n685_), .ZN(new_n805_));
  OAI21_X1   g0669(.A1(new_n805_), .A2(new_n401_), .B(\A[45] ), .ZN(new_n806_));
  AOI21_X1   g0670(.A1(new_n806_), .A2(new_n411_), .B(new_n684_), .ZN(new_n807_));
  OAI21_X1   g0671(.A1(new_n807_), .A2(new_n408_), .B(\A[43] ), .ZN(new_n808_));
  AOI21_X1   g0672(.A1(new_n808_), .A2(new_n418_), .B(new_n683_), .ZN(new_n809_));
  OAI21_X1   g0673(.A1(new_n809_), .A2(new_n415_), .B(\A[41] ), .ZN(new_n810_));
  AOI21_X1   g0674(.A1(new_n810_), .A2(new_n425_), .B(new_n682_), .ZN(new_n811_));
  OAI21_X1   g0675(.A1(new_n811_), .A2(new_n422_), .B(\A[39] ), .ZN(new_n812_));
  AOI21_X1   g0676(.A1(new_n812_), .A2(new_n432_), .B(new_n681_), .ZN(new_n813_));
  OAI21_X1   g0677(.A1(new_n813_), .A2(new_n429_), .B(\A[37] ), .ZN(new_n814_));
  AOI21_X1   g0678(.A1(new_n814_), .A2(new_n439_), .B(new_n680_), .ZN(new_n815_));
  OAI21_X1   g0679(.A1(new_n815_), .A2(new_n436_), .B(\A[35] ), .ZN(new_n816_));
  AOI21_X1   g0680(.A1(new_n816_), .A2(new_n446_), .B(new_n679_), .ZN(new_n817_));
  OAI21_X1   g0681(.A1(new_n817_), .A2(new_n443_), .B(\A[33] ), .ZN(new_n818_));
  AOI21_X1   g0682(.A1(new_n818_), .A2(new_n453_), .B(new_n678_), .ZN(new_n819_));
  OAI21_X1   g0683(.A1(new_n819_), .A2(new_n450_), .B(\A[31] ), .ZN(new_n820_));
  AOI21_X1   g0684(.A1(new_n820_), .A2(new_n460_), .B(new_n677_), .ZN(new_n821_));
  OAI21_X1   g0685(.A1(new_n821_), .A2(new_n457_), .B(\A[29] ), .ZN(new_n822_));
  AOI21_X1   g0686(.A1(new_n822_), .A2(new_n467_), .B(new_n676_), .ZN(new_n823_));
  OAI21_X1   g0687(.A1(new_n823_), .A2(new_n464_), .B(\A[27] ), .ZN(new_n824_));
  AOI21_X1   g0688(.A1(new_n824_), .A2(new_n474_), .B(new_n675_), .ZN(new_n825_));
  OAI21_X1   g0689(.A1(new_n825_), .A2(new_n471_), .B(\A[25] ), .ZN(new_n826_));
  AOI21_X1   g0690(.A1(new_n826_), .A2(new_n481_), .B(new_n674_), .ZN(new_n827_));
  OAI21_X1   g0691(.A1(new_n827_), .A2(new_n478_), .B(\A[23] ), .ZN(new_n828_));
  AOI21_X1   g0692(.A1(new_n828_), .A2(new_n488_), .B(new_n673_), .ZN(new_n829_));
  OAI21_X1   g0693(.A1(new_n829_), .A2(new_n485_), .B(\A[21] ), .ZN(new_n830_));
  AOI21_X1   g0694(.A1(new_n830_), .A2(new_n495_), .B(new_n672_), .ZN(new_n831_));
  OAI21_X1   g0695(.A1(new_n831_), .A2(new_n492_), .B(\A[19] ), .ZN(new_n832_));
  AOI21_X1   g0696(.A1(new_n832_), .A2(new_n502_), .B(new_n671_), .ZN(new_n833_));
  OAI21_X1   g0697(.A1(new_n833_), .A2(new_n499_), .B(\A[17] ), .ZN(new_n834_));
  AOI21_X1   g0698(.A1(new_n834_), .A2(new_n509_), .B(new_n670_), .ZN(new_n835_));
  OAI21_X1   g0699(.A1(new_n835_), .A2(new_n506_), .B(\A[15] ), .ZN(new_n836_));
  AOI21_X1   g0700(.A1(new_n836_), .A2(new_n516_), .B(new_n669_), .ZN(new_n837_));
  OAI21_X1   g0701(.A1(new_n837_), .A2(new_n513_), .B(\A[13] ), .ZN(new_n838_));
  AOI21_X1   g0702(.A1(new_n838_), .A2(new_n523_), .B(new_n668_), .ZN(new_n839_));
  OAI21_X1   g0703(.A1(new_n839_), .A2(new_n520_), .B(\A[11] ), .ZN(new_n840_));
  AOI21_X1   g0704(.A1(new_n840_), .A2(new_n530_), .B(new_n667_), .ZN(new_n841_));
  OAI21_X1   g0705(.A1(new_n841_), .A2(new_n527_), .B(\A[9] ), .ZN(new_n842_));
  AOI21_X1   g0706(.A1(new_n842_), .A2(new_n537_), .B(new_n666_), .ZN(new_n843_));
  OAI21_X1   g0707(.A1(new_n843_), .A2(new_n534_), .B(\A[7] ), .ZN(new_n844_));
  AOI21_X1   g0708(.A1(new_n844_), .A2(new_n544_), .B(new_n665_), .ZN(new_n845_));
  OAI21_X1   g0709(.A1(new_n845_), .A2(new_n541_), .B(\A[5] ), .ZN(new_n846_));
  AOI21_X1   g0710(.A1(new_n846_), .A2(new_n659_), .B(new_n664_), .ZN(new_n847_));
  OAI21_X1   g0711(.A1(new_n847_), .A2(new_n548_), .B(\A[3] ), .ZN(new_n848_));
  INV_X1     g0712(.I(\A[3] ), .ZN(new_n849_));
  AOI21_X1   g0713(.A1(new_n660_), .A2(new_n849_), .B(new_n663_), .ZN(new_n850_));
  AOI22_X1   g0714(.A1(new_n848_), .A2(new_n850_), .B1(new_n661_), .B2(new_n663_), .ZN(\P[0] ));
  NOR2_X1    g0715(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n852_));
  INV_X1     g0716(.I(new_n852_), .ZN(new_n853_));
  NOR2_X1    g0717(.A1(\A[18] ), .A2(\A[19] ), .ZN(new_n854_));
  INV_X1     g0718(.I(new_n854_), .ZN(new_n855_));
  NOR2_X1    g0719(.A1(\A[22] ), .A2(\A[23] ), .ZN(new_n856_));
  INV_X1     g0720(.I(new_n856_), .ZN(new_n857_));
  NOR2_X1    g0721(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n858_));
  INV_X1     g0722(.I(new_n858_), .ZN(new_n859_));
  NOR2_X1    g0723(.A1(\A[30] ), .A2(\A[31] ), .ZN(new_n860_));
  INV_X1     g0724(.I(new_n860_), .ZN(new_n861_));
  NOR2_X1    g0725(.A1(\A[34] ), .A2(\A[35] ), .ZN(new_n862_));
  INV_X1     g0726(.I(new_n862_), .ZN(new_n863_));
  NOR2_X1    g0727(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n864_));
  INV_X1     g0728(.I(new_n864_), .ZN(new_n865_));
  NOR2_X1    g0729(.A1(\A[42] ), .A2(\A[43] ), .ZN(new_n866_));
  INV_X1     g0730(.I(new_n866_), .ZN(new_n867_));
  NOR2_X1    g0731(.A1(\A[46] ), .A2(\A[47] ), .ZN(new_n868_));
  INV_X1     g0732(.I(new_n868_), .ZN(new_n869_));
  NOR2_X1    g0733(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n870_));
  INV_X1     g0734(.I(new_n870_), .ZN(new_n871_));
  NOR2_X1    g0735(.A1(\A[54] ), .A2(\A[55] ), .ZN(new_n872_));
  INV_X1     g0736(.I(new_n872_), .ZN(new_n873_));
  NOR2_X1    g0737(.A1(\A[58] ), .A2(\A[59] ), .ZN(new_n874_));
  INV_X1     g0738(.I(new_n874_), .ZN(new_n875_));
  NOR2_X1    g0739(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n876_));
  INV_X1     g0740(.I(new_n876_), .ZN(new_n877_));
  NOR2_X1    g0741(.A1(\A[66] ), .A2(\A[67] ), .ZN(new_n878_));
  INV_X1     g0742(.I(new_n878_), .ZN(new_n879_));
  NOR2_X1    g0743(.A1(\A[70] ), .A2(\A[71] ), .ZN(new_n880_));
  INV_X1     g0744(.I(new_n880_), .ZN(new_n881_));
  NOR2_X1    g0745(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n882_));
  INV_X1     g0746(.I(new_n882_), .ZN(new_n883_));
  NOR2_X1    g0747(.A1(\A[78] ), .A2(\A[79] ), .ZN(new_n884_));
  INV_X1     g0748(.I(new_n884_), .ZN(new_n885_));
  NOR2_X1    g0749(.A1(\A[82] ), .A2(\A[83] ), .ZN(new_n886_));
  INV_X1     g0750(.I(new_n886_), .ZN(new_n887_));
  NOR2_X1    g0751(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n888_));
  INV_X1     g0752(.I(new_n888_), .ZN(new_n889_));
  NOR2_X1    g0753(.A1(\A[90] ), .A2(\A[91] ), .ZN(new_n890_));
  INV_X1     g0754(.I(new_n890_), .ZN(new_n891_));
  NOR2_X1    g0755(.A1(\A[126] ), .A2(\A[127] ), .ZN(new_n892_));
  NAND2_X1   g0756(.A1(new_n723_), .A2(new_n143_), .ZN(new_n893_));
  NOR2_X1    g0757(.A1(\A[124] ), .A2(\A[125] ), .ZN(new_n894_));
  NAND2_X1   g0758(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1   g0759(.A1(new_n895_), .A2(new_n892_), .ZN(new_n896_));
  NAND2_X1   g0760(.A1(new_n896_), .A2(\A[120] ), .ZN(new_n897_));
  OAI21_X1   g0761(.A1(new_n893_), .A2(new_n148_), .B(new_n894_), .ZN(new_n898_));
  NAND2_X1   g0762(.A1(new_n898_), .A2(new_n892_), .ZN(new_n899_));
  NAND2_X1   g0763(.A1(new_n899_), .A2(new_n722_), .ZN(new_n900_));
  NAND2_X1   g0764(.A1(new_n900_), .A2(new_n897_), .ZN(new_n901_));
  NOR2_X1    g0765(.A1(\A[118] ), .A2(\A[119] ), .ZN(new_n902_));
  NOR2_X1    g0766(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1     g0767(.I(new_n902_), .ZN(new_n904_));
  NOR2_X1    g0768(.A1(new_n896_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1    g0769(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1    g0770(.A1(\A[114] ), .A2(\A[115] ), .ZN(new_n907_));
  INV_X1     g0771(.I(new_n907_), .ZN(new_n908_));
  NOR2_X1    g0772(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1    g0773(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n910_));
  NAND2_X1   g0774(.A1(new_n901_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1     g0775(.I(new_n910_), .ZN(new_n912_));
  NAND2_X1   g0776(.A1(new_n906_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1   g0777(.A1(new_n913_), .A2(new_n911_), .ZN(new_n914_));
  NOR2_X1    g0778(.A1(new_n914_), .A2(new_n907_), .ZN(new_n915_));
  NOR2_X1    g0779(.A1(new_n915_), .A2(new_n909_), .ZN(new_n916_));
  NOR2_X1    g0780(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n917_));
  INV_X1     g0781(.I(new_n917_), .ZN(new_n918_));
  NOR2_X1    g0782(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1    g0783(.A1(\A[112] ), .A2(\A[113] ), .ZN(new_n920_));
  NAND2_X1   g0784(.A1(new_n914_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1     g0785(.I(new_n920_), .ZN(new_n922_));
  NAND2_X1   g0786(.A1(new_n916_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1   g0787(.A1(new_n923_), .A2(new_n921_), .ZN(new_n924_));
  NOR2_X1    g0788(.A1(new_n924_), .A2(new_n917_), .ZN(new_n925_));
  NOR2_X1    g0789(.A1(new_n925_), .A2(new_n919_), .ZN(new_n926_));
  NOR2_X1    g0790(.A1(\A[106] ), .A2(\A[107] ), .ZN(new_n927_));
  INV_X1     g0791(.I(new_n927_), .ZN(new_n928_));
  NOR2_X1    g0792(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1    g0793(.A1(\A[108] ), .A2(\A[109] ), .ZN(new_n930_));
  NAND2_X1   g0794(.A1(new_n924_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1     g0795(.I(new_n930_), .ZN(new_n932_));
  NAND2_X1   g0796(.A1(new_n926_), .A2(new_n932_), .ZN(new_n933_));
  NAND2_X1   g0797(.A1(new_n933_), .A2(new_n931_), .ZN(new_n934_));
  NOR2_X1    g0798(.A1(new_n934_), .A2(new_n927_), .ZN(new_n935_));
  NOR2_X1    g0799(.A1(new_n935_), .A2(new_n929_), .ZN(new_n936_));
  NOR2_X1    g0800(.A1(\A[102] ), .A2(\A[103] ), .ZN(new_n937_));
  INV_X1     g0801(.I(new_n937_), .ZN(new_n938_));
  NOR2_X1    g0802(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1    g0803(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n940_));
  NAND2_X1   g0804(.A1(new_n934_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1     g0805(.I(new_n940_), .ZN(new_n942_));
  NAND2_X1   g0806(.A1(new_n936_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1   g0807(.A1(new_n943_), .A2(new_n941_), .ZN(new_n944_));
  NOR2_X1    g0808(.A1(new_n944_), .A2(new_n937_), .ZN(new_n945_));
  NOR2_X1    g0809(.A1(new_n945_), .A2(new_n939_), .ZN(new_n946_));
  NOR2_X1    g0810(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n947_));
  INV_X1     g0811(.I(new_n947_), .ZN(new_n948_));
  NOR2_X1    g0812(.A1(new_n946_), .A2(new_n948_), .ZN(new_n949_));
  NOR2_X1    g0813(.A1(\A[100] ), .A2(\A[101] ), .ZN(new_n950_));
  NAND2_X1   g0814(.A1(new_n944_), .A2(new_n950_), .ZN(new_n951_));
  INV_X1     g0815(.I(new_n950_), .ZN(new_n952_));
  NAND2_X1   g0816(.A1(new_n946_), .A2(new_n952_), .ZN(new_n953_));
  NAND2_X1   g0817(.A1(new_n953_), .A2(new_n951_), .ZN(new_n954_));
  NOR2_X1    g0818(.A1(new_n954_), .A2(new_n947_), .ZN(new_n955_));
  NOR2_X1    g0819(.A1(new_n955_), .A2(new_n949_), .ZN(new_n956_));
  NOR3_X1    g0820(.A1(new_n956_), .A2(\A[94] ), .A3(\A[95] ), .ZN(new_n957_));
  NOR2_X1    g0821(.A1(\A[94] ), .A2(\A[95] ), .ZN(new_n958_));
  NOR2_X1    g0822(.A1(\A[96] ), .A2(\A[97] ), .ZN(new_n959_));
  NAND2_X1   g0823(.A1(new_n954_), .A2(new_n959_), .ZN(new_n960_));
  INV_X1     g0824(.I(new_n959_), .ZN(new_n961_));
  NAND2_X1   g0825(.A1(new_n956_), .A2(new_n961_), .ZN(new_n962_));
  NAND2_X1   g0826(.A1(new_n962_), .A2(new_n960_), .ZN(new_n963_));
  NOR2_X1    g0827(.A1(new_n963_), .A2(new_n958_), .ZN(new_n964_));
  NOR2_X1    g0828(.A1(new_n964_), .A2(new_n957_), .ZN(new_n965_));
  NOR2_X1    g0829(.A1(new_n965_), .A2(new_n891_), .ZN(new_n966_));
  NOR2_X1    g0830(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n967_));
  NOR3_X1    g0831(.A1(new_n964_), .A2(new_n957_), .A3(new_n967_), .ZN(new_n968_));
  AOI21_X1   g0832(.A1(new_n963_), .A2(new_n967_), .B(new_n968_), .ZN(new_n969_));
  AOI21_X1   g0833(.A1(new_n969_), .A2(new_n891_), .B(new_n966_), .ZN(new_n970_));
  NOR2_X1    g0834(.A1(new_n970_), .A2(new_n889_), .ZN(new_n971_));
  NOR2_X1    g0835(.A1(\A[88] ), .A2(\A[89] ), .ZN(new_n972_));
  INV_X1     g0836(.I(new_n972_), .ZN(new_n973_));
  NOR2_X1    g0837(.A1(new_n969_), .A2(new_n973_), .ZN(new_n974_));
  AOI21_X1   g0838(.A1(new_n970_), .A2(new_n973_), .B(new_n974_), .ZN(new_n975_));
  AOI21_X1   g0839(.A1(new_n975_), .A2(new_n889_), .B(new_n971_), .ZN(new_n976_));
  NOR2_X1    g0840(.A1(new_n976_), .A2(new_n887_), .ZN(new_n977_));
  NOR2_X1    g0841(.A1(\A[84] ), .A2(\A[85] ), .ZN(new_n978_));
  INV_X1     g0842(.I(new_n978_), .ZN(new_n979_));
  NOR2_X1    g0843(.A1(new_n975_), .A2(new_n979_), .ZN(new_n980_));
  AOI21_X1   g0844(.A1(new_n976_), .A2(new_n979_), .B(new_n980_), .ZN(new_n981_));
  AOI21_X1   g0845(.A1(new_n981_), .A2(new_n887_), .B(new_n977_), .ZN(new_n982_));
  NOR2_X1    g0846(.A1(new_n982_), .A2(new_n885_), .ZN(new_n983_));
  NOR2_X1    g0847(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n984_));
  INV_X1     g0848(.I(new_n984_), .ZN(new_n985_));
  NOR2_X1    g0849(.A1(new_n981_), .A2(new_n985_), .ZN(new_n986_));
  AOI21_X1   g0850(.A1(new_n982_), .A2(new_n985_), .B(new_n986_), .ZN(new_n987_));
  AOI21_X1   g0851(.A1(new_n987_), .A2(new_n885_), .B(new_n983_), .ZN(new_n988_));
  NOR2_X1    g0852(.A1(new_n988_), .A2(new_n883_), .ZN(new_n989_));
  NOR2_X1    g0853(.A1(\A[76] ), .A2(\A[77] ), .ZN(new_n990_));
  INV_X1     g0854(.I(new_n990_), .ZN(new_n991_));
  NOR2_X1    g0855(.A1(new_n987_), .A2(new_n991_), .ZN(new_n992_));
  AOI21_X1   g0856(.A1(new_n988_), .A2(new_n991_), .B(new_n992_), .ZN(new_n993_));
  AOI21_X1   g0857(.A1(new_n993_), .A2(new_n883_), .B(new_n989_), .ZN(new_n994_));
  NOR2_X1    g0858(.A1(new_n994_), .A2(new_n881_), .ZN(new_n995_));
  NOR2_X1    g0859(.A1(\A[72] ), .A2(\A[73] ), .ZN(new_n996_));
  INV_X1     g0860(.I(new_n996_), .ZN(new_n997_));
  NOR2_X1    g0861(.A1(new_n993_), .A2(new_n997_), .ZN(new_n998_));
  AOI21_X1   g0862(.A1(new_n994_), .A2(new_n997_), .B(new_n998_), .ZN(new_n999_));
  AOI21_X1   g0863(.A1(new_n999_), .A2(new_n881_), .B(new_n995_), .ZN(new_n1000_));
  NOR2_X1    g0864(.A1(new_n1000_), .A2(new_n879_), .ZN(new_n1001_));
  NOR2_X1    g0865(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n1002_));
  INV_X1     g0866(.I(new_n1002_), .ZN(new_n1003_));
  NOR2_X1    g0867(.A1(new_n999_), .A2(new_n1003_), .ZN(new_n1004_));
  AOI21_X1   g0868(.A1(new_n1000_), .A2(new_n1003_), .B(new_n1004_), .ZN(new_n1005_));
  AOI21_X1   g0869(.A1(new_n1005_), .A2(new_n879_), .B(new_n1001_), .ZN(new_n1006_));
  NOR2_X1    g0870(.A1(new_n1006_), .A2(new_n877_), .ZN(new_n1007_));
  NOR2_X1    g0871(.A1(\A[64] ), .A2(\A[65] ), .ZN(new_n1008_));
  INV_X1     g0872(.I(new_n1008_), .ZN(new_n1009_));
  NOR2_X1    g0873(.A1(new_n1005_), .A2(new_n1009_), .ZN(new_n1010_));
  AOI21_X1   g0874(.A1(new_n1006_), .A2(new_n1009_), .B(new_n1010_), .ZN(new_n1011_));
  AOI21_X1   g0875(.A1(new_n1011_), .A2(new_n877_), .B(new_n1007_), .ZN(new_n1012_));
  NOR2_X1    g0876(.A1(new_n1012_), .A2(new_n875_), .ZN(new_n1013_));
  NOR2_X1    g0877(.A1(\A[60] ), .A2(\A[61] ), .ZN(new_n1014_));
  INV_X1     g0878(.I(new_n1014_), .ZN(new_n1015_));
  NOR2_X1    g0879(.A1(new_n1011_), .A2(new_n1015_), .ZN(new_n1016_));
  AOI21_X1   g0880(.A1(new_n1012_), .A2(new_n1015_), .B(new_n1016_), .ZN(new_n1017_));
  AOI21_X1   g0881(.A1(new_n1017_), .A2(new_n875_), .B(new_n1013_), .ZN(new_n1018_));
  NOR2_X1    g0882(.A1(new_n1018_), .A2(new_n873_), .ZN(new_n1019_));
  NOR2_X1    g0883(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n1020_));
  INV_X1     g0884(.I(new_n1020_), .ZN(new_n1021_));
  NOR2_X1    g0885(.A1(new_n1017_), .A2(new_n1021_), .ZN(new_n1022_));
  AOI21_X1   g0886(.A1(new_n1018_), .A2(new_n1021_), .B(new_n1022_), .ZN(new_n1023_));
  AOI21_X1   g0887(.A1(new_n1023_), .A2(new_n873_), .B(new_n1019_), .ZN(new_n1024_));
  NOR2_X1    g0888(.A1(new_n1024_), .A2(new_n871_), .ZN(new_n1025_));
  NOR2_X1    g0889(.A1(\A[52] ), .A2(\A[53] ), .ZN(new_n1026_));
  INV_X1     g0890(.I(new_n1026_), .ZN(new_n1027_));
  NOR2_X1    g0891(.A1(new_n1023_), .A2(new_n1027_), .ZN(new_n1028_));
  AOI21_X1   g0892(.A1(new_n1024_), .A2(new_n1027_), .B(new_n1028_), .ZN(new_n1029_));
  AOI21_X1   g0893(.A1(new_n1029_), .A2(new_n871_), .B(new_n1025_), .ZN(new_n1030_));
  NOR2_X1    g0894(.A1(new_n1030_), .A2(new_n869_), .ZN(new_n1031_));
  NOR2_X1    g0895(.A1(\A[48] ), .A2(\A[49] ), .ZN(new_n1032_));
  INV_X1     g0896(.I(new_n1032_), .ZN(new_n1033_));
  NOR2_X1    g0897(.A1(new_n1029_), .A2(new_n1033_), .ZN(new_n1034_));
  AOI21_X1   g0898(.A1(new_n1030_), .A2(new_n1033_), .B(new_n1034_), .ZN(new_n1035_));
  AOI21_X1   g0899(.A1(new_n1035_), .A2(new_n869_), .B(new_n1031_), .ZN(new_n1036_));
  NOR2_X1    g0900(.A1(new_n1036_), .A2(new_n867_), .ZN(new_n1037_));
  NOR2_X1    g0901(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n1038_));
  INV_X1     g0902(.I(new_n1038_), .ZN(new_n1039_));
  NOR2_X1    g0903(.A1(new_n1035_), .A2(new_n1039_), .ZN(new_n1040_));
  AOI21_X1   g0904(.A1(new_n1036_), .A2(new_n1039_), .B(new_n1040_), .ZN(new_n1041_));
  AOI21_X1   g0905(.A1(new_n1041_), .A2(new_n867_), .B(new_n1037_), .ZN(new_n1042_));
  NOR2_X1    g0906(.A1(new_n1042_), .A2(new_n865_), .ZN(new_n1043_));
  NOR2_X1    g0907(.A1(\A[40] ), .A2(\A[41] ), .ZN(new_n1044_));
  INV_X1     g0908(.I(new_n1044_), .ZN(new_n1045_));
  NOR2_X1    g0909(.A1(new_n1041_), .A2(new_n1045_), .ZN(new_n1046_));
  AOI21_X1   g0910(.A1(new_n1042_), .A2(new_n1045_), .B(new_n1046_), .ZN(new_n1047_));
  AOI21_X1   g0911(.A1(new_n1047_), .A2(new_n865_), .B(new_n1043_), .ZN(new_n1048_));
  NOR2_X1    g0912(.A1(new_n1048_), .A2(new_n863_), .ZN(new_n1049_));
  NOR2_X1    g0913(.A1(\A[36] ), .A2(\A[37] ), .ZN(new_n1050_));
  INV_X1     g0914(.I(new_n1050_), .ZN(new_n1051_));
  NOR2_X1    g0915(.A1(new_n1047_), .A2(new_n1051_), .ZN(new_n1052_));
  AOI21_X1   g0916(.A1(new_n1048_), .A2(new_n1051_), .B(new_n1052_), .ZN(new_n1053_));
  AOI21_X1   g0917(.A1(new_n1053_), .A2(new_n863_), .B(new_n1049_), .ZN(new_n1054_));
  NOR2_X1    g0918(.A1(new_n1054_), .A2(new_n861_), .ZN(new_n1055_));
  NOR2_X1    g0919(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n1056_));
  INV_X1     g0920(.I(new_n1056_), .ZN(new_n1057_));
  NOR2_X1    g0921(.A1(new_n1053_), .A2(new_n1057_), .ZN(new_n1058_));
  AOI21_X1   g0922(.A1(new_n1054_), .A2(new_n1057_), .B(new_n1058_), .ZN(new_n1059_));
  AOI21_X1   g0923(.A1(new_n1059_), .A2(new_n861_), .B(new_n1055_), .ZN(new_n1060_));
  NOR2_X1    g0924(.A1(new_n1060_), .A2(new_n859_), .ZN(new_n1061_));
  NOR2_X1    g0925(.A1(\A[28] ), .A2(\A[29] ), .ZN(new_n1062_));
  INV_X1     g0926(.I(new_n1062_), .ZN(new_n1063_));
  NOR2_X1    g0927(.A1(new_n1059_), .A2(new_n1063_), .ZN(new_n1064_));
  AOI21_X1   g0928(.A1(new_n1060_), .A2(new_n1063_), .B(new_n1064_), .ZN(new_n1065_));
  AOI21_X1   g0929(.A1(new_n1065_), .A2(new_n859_), .B(new_n1061_), .ZN(new_n1066_));
  NOR2_X1    g0930(.A1(new_n1066_), .A2(new_n857_), .ZN(new_n1067_));
  NOR2_X1    g0931(.A1(\A[24] ), .A2(\A[25] ), .ZN(new_n1068_));
  INV_X1     g0932(.I(new_n1068_), .ZN(new_n1069_));
  NOR2_X1    g0933(.A1(new_n1065_), .A2(new_n1069_), .ZN(new_n1070_));
  AOI21_X1   g0934(.A1(new_n1066_), .A2(new_n1069_), .B(new_n1070_), .ZN(new_n1071_));
  AOI21_X1   g0935(.A1(new_n1071_), .A2(new_n857_), .B(new_n1067_), .ZN(new_n1072_));
  NOR2_X1    g0936(.A1(new_n1072_), .A2(new_n855_), .ZN(new_n1073_));
  NOR2_X1    g0937(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n1074_));
  INV_X1     g0938(.I(new_n1074_), .ZN(new_n1075_));
  NOR2_X1    g0939(.A1(new_n1071_), .A2(new_n1075_), .ZN(new_n1076_));
  AOI21_X1   g0940(.A1(new_n1072_), .A2(new_n1075_), .B(new_n1076_), .ZN(new_n1077_));
  AOI21_X1   g0941(.A1(new_n1077_), .A2(new_n855_), .B(new_n1073_), .ZN(new_n1078_));
  NOR2_X1    g0942(.A1(new_n1078_), .A2(new_n853_), .ZN(new_n1079_));
  NOR2_X1    g0943(.A1(\A[16] ), .A2(\A[17] ), .ZN(new_n1080_));
  INV_X1     g0944(.I(new_n1080_), .ZN(new_n1081_));
  NOR2_X1    g0945(.A1(new_n1077_), .A2(new_n1081_), .ZN(new_n1082_));
  AOI21_X1   g0946(.A1(new_n1078_), .A2(new_n1081_), .B(new_n1082_), .ZN(new_n1083_));
  AOI21_X1   g0947(.A1(new_n1083_), .A2(new_n853_), .B(new_n1079_), .ZN(new_n1084_));
  NOR2_X1    g0948(.A1(\A[10] ), .A2(\A[11] ), .ZN(new_n1085_));
  INV_X1     g0949(.I(new_n1085_), .ZN(new_n1086_));
  OR2_X2     g0950(.A1(new_n1084_), .A2(new_n1086_), .Z(new_n1087_));
  NOR2_X1    g0951(.A1(\A[12] ), .A2(\A[13] ), .ZN(new_n1088_));
  INV_X1     g0952(.I(new_n1088_), .ZN(new_n1089_));
  OR2_X2     g0953(.A1(new_n1083_), .A2(new_n1089_), .Z(new_n1090_));
  NAND2_X1   g0954(.A1(new_n1084_), .A2(new_n1089_), .ZN(new_n1091_));
  NAND3_X1   g0955(.A1(new_n1091_), .A2(new_n1086_), .A3(new_n1090_), .ZN(new_n1092_));
  NAND2_X1   g0956(.A1(new_n1092_), .A2(new_n1087_), .ZN(new_n1093_));
  NOR2_X1    g0957(.A1(\A[6] ), .A2(\A[7] ), .ZN(new_n1094_));
  NAND2_X1   g0958(.A1(new_n1093_), .A2(new_n1094_), .ZN(new_n1095_));
  INV_X1     g0959(.I(new_n1094_), .ZN(new_n1096_));
  NAND2_X1   g0960(.A1(new_n1091_), .A2(new_n1090_), .ZN(new_n1097_));
  NOR2_X1    g0961(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n1098_));
  NAND2_X1   g0962(.A1(new_n1097_), .A2(new_n1098_), .ZN(new_n1099_));
  INV_X1     g0963(.I(new_n1098_), .ZN(new_n1100_));
  NAND3_X1   g0964(.A1(new_n1092_), .A2(new_n1087_), .A3(new_n1100_), .ZN(new_n1101_));
  NAND3_X1   g0965(.A1(new_n1101_), .A2(new_n1096_), .A3(new_n1099_), .ZN(new_n1102_));
  NAND2_X1   g0966(.A1(new_n1102_), .A2(new_n1095_), .ZN(new_n1103_));
  NOR2_X1    g0967(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n1104_));
  INV_X1     g0968(.I(new_n1104_), .ZN(new_n1105_));
  NAND3_X1   g0969(.A1(new_n1102_), .A2(new_n1095_), .A3(new_n1105_), .ZN(new_n1106_));
  NOR2_X1    g0970(.A1(\A[2] ), .A2(\A[3] ), .ZN(new_n1107_));
  NAND2_X1   g0971(.A1(new_n1101_), .A2(new_n1099_), .ZN(new_n1108_));
  AOI21_X1   g0972(.A1(new_n1108_), .A2(new_n1104_), .B(new_n1107_), .ZN(new_n1109_));
  AOI22_X1   g0973(.A1(new_n1106_), .A2(new_n1109_), .B1(new_n1103_), .B2(new_n1107_), .ZN(\P[1] ));
  NOR2_X1    g0974(.A1(new_n857_), .A2(new_n1075_), .ZN(new_n1111_));
  NAND2_X1   g0975(.A1(new_n958_), .A2(new_n967_), .ZN(new_n1112_));
  NAND2_X1   g0976(.A1(new_n892_), .A2(new_n894_), .ZN(new_n1113_));
  INV_X1     g0977(.I(new_n1113_), .ZN(new_n1114_));
  NOR3_X1    g0978(.A1(new_n893_), .A2(\A[120] ), .A3(\A[121] ), .ZN(new_n1115_));
  INV_X1     g0979(.I(new_n1115_), .ZN(new_n1116_));
  NOR2_X1    g0980(.A1(new_n904_), .A2(new_n912_), .ZN(new_n1117_));
  OAI21_X1   g0981(.A1(new_n1116_), .A2(new_n1117_), .B(new_n1114_), .ZN(new_n1118_));
  NOR2_X1    g0982(.A1(new_n918_), .A2(new_n932_), .ZN(new_n1119_));
  NOR2_X1    g0983(.A1(new_n922_), .A2(\A[114] ), .ZN(new_n1120_));
  NOR2_X1    g0984(.A1(new_n1118_), .A2(new_n1120_), .ZN(new_n1121_));
  NAND2_X1   g0985(.A1(new_n1117_), .A2(\A[115] ), .ZN(new_n1122_));
  NAND2_X1   g0986(.A1(new_n1114_), .A2(new_n1120_), .ZN(new_n1123_));
  AOI21_X1   g0987(.A1(new_n1115_), .A2(new_n1122_), .B(new_n1123_), .ZN(new_n1124_));
  NOR3_X1    g0988(.A1(new_n1121_), .A2(new_n1119_), .A3(new_n1124_), .ZN(new_n1125_));
  AOI21_X1   g0989(.A1(new_n1118_), .A2(new_n1119_), .B(new_n1125_), .ZN(new_n1126_));
  NOR2_X1    g0990(.A1(new_n938_), .A2(new_n952_), .ZN(new_n1127_));
  INV_X1     g0991(.I(new_n1127_), .ZN(new_n1128_));
  NOR2_X1    g0992(.A1(new_n1126_), .A2(new_n1128_), .ZN(new_n1129_));
  NOR2_X1    g0993(.A1(new_n1121_), .A2(new_n1124_), .ZN(new_n1130_));
  NOR2_X1    g0994(.A1(new_n928_), .A2(new_n942_), .ZN(new_n1131_));
  INV_X1     g0995(.I(new_n1131_), .ZN(new_n1132_));
  NAND2_X1   g0996(.A1(new_n1126_), .A2(new_n1132_), .ZN(new_n1133_));
  OAI21_X1   g0997(.A1(new_n1130_), .A2(new_n1132_), .B(new_n1133_), .ZN(new_n1134_));
  NOR2_X1    g0998(.A1(new_n1134_), .A2(new_n1127_), .ZN(new_n1135_));
  NOR2_X1    g0999(.A1(new_n1135_), .A2(new_n1129_), .ZN(new_n1136_));
  NOR2_X1    g1000(.A1(new_n1136_), .A2(new_n1112_), .ZN(new_n1137_));
  NOR2_X1    g1001(.A1(new_n948_), .A2(new_n961_), .ZN(new_n1138_));
  NAND2_X1   g1002(.A1(new_n1134_), .A2(new_n1138_), .ZN(new_n1139_));
  INV_X1     g1003(.I(new_n1138_), .ZN(new_n1140_));
  NAND2_X1   g1004(.A1(new_n1136_), .A2(new_n1140_), .ZN(new_n1141_));
  NAND2_X1   g1005(.A1(new_n1141_), .A2(new_n1139_), .ZN(new_n1142_));
  INV_X1     g1006(.I(new_n1142_), .ZN(new_n1143_));
  AOI21_X1   g1007(.A1(new_n1143_), .A2(new_n1112_), .B(new_n1137_), .ZN(new_n1144_));
  NOR2_X1    g1008(.A1(new_n889_), .A2(new_n979_), .ZN(new_n1145_));
  INV_X1     g1009(.I(new_n1145_), .ZN(new_n1146_));
  NOR2_X1    g1010(.A1(new_n1144_), .A2(new_n1146_), .ZN(new_n1147_));
  NOR2_X1    g1011(.A1(new_n891_), .A2(new_n973_), .ZN(new_n1148_));
  INV_X1     g1012(.I(new_n1148_), .ZN(new_n1149_));
  NAND2_X1   g1013(.A1(new_n1144_), .A2(new_n1149_), .ZN(new_n1150_));
  OAI21_X1   g1014(.A1(new_n1143_), .A2(new_n1149_), .B(new_n1150_), .ZN(new_n1151_));
  NOR2_X1    g1015(.A1(new_n1151_), .A2(new_n1145_), .ZN(new_n1152_));
  NOR2_X1    g1016(.A1(new_n1152_), .A2(new_n1147_), .ZN(new_n1153_));
  NOR2_X1    g1017(.A1(new_n885_), .A2(new_n991_), .ZN(new_n1154_));
  INV_X1     g1018(.I(new_n1154_), .ZN(new_n1155_));
  NOR2_X1    g1019(.A1(new_n1153_), .A2(new_n1155_), .ZN(new_n1156_));
  NOR2_X1    g1020(.A1(new_n887_), .A2(new_n985_), .ZN(new_n1157_));
  NAND2_X1   g1021(.A1(new_n1151_), .A2(new_n1157_), .ZN(new_n1158_));
  INV_X1     g1022(.I(new_n1157_), .ZN(new_n1159_));
  NAND2_X1   g1023(.A1(new_n1153_), .A2(new_n1159_), .ZN(new_n1160_));
  NAND2_X1   g1024(.A1(new_n1160_), .A2(new_n1158_), .ZN(new_n1161_));
  NOR2_X1    g1025(.A1(new_n1161_), .A2(new_n1154_), .ZN(new_n1162_));
  NOR2_X1    g1026(.A1(new_n1162_), .A2(new_n1156_), .ZN(new_n1163_));
  NOR2_X1    g1027(.A1(new_n881_), .A2(new_n1003_), .ZN(new_n1164_));
  INV_X1     g1028(.I(new_n1164_), .ZN(new_n1165_));
  NOR2_X1    g1029(.A1(new_n1163_), .A2(new_n1165_), .ZN(new_n1166_));
  NOR2_X1    g1030(.A1(new_n883_), .A2(new_n997_), .ZN(new_n1167_));
  NAND2_X1   g1031(.A1(new_n1161_), .A2(new_n1167_), .ZN(new_n1168_));
  INV_X1     g1032(.I(new_n1167_), .ZN(new_n1169_));
  NAND2_X1   g1033(.A1(new_n1163_), .A2(new_n1169_), .ZN(new_n1170_));
  NAND2_X1   g1034(.A1(new_n1170_), .A2(new_n1168_), .ZN(new_n1171_));
  NOR2_X1    g1035(.A1(new_n1171_), .A2(new_n1164_), .ZN(new_n1172_));
  NOR2_X1    g1036(.A1(new_n1172_), .A2(new_n1166_), .ZN(new_n1173_));
  NOR2_X1    g1037(.A1(new_n877_), .A2(new_n1015_), .ZN(new_n1174_));
  NOR2_X1    g1038(.A1(new_n879_), .A2(new_n1009_), .ZN(new_n1175_));
  NAND2_X1   g1039(.A1(new_n1171_), .A2(new_n1175_), .ZN(new_n1176_));
  INV_X1     g1040(.I(new_n1175_), .ZN(new_n1177_));
  NAND2_X1   g1041(.A1(new_n1173_), .A2(new_n1177_), .ZN(new_n1178_));
  NAND2_X1   g1042(.A1(new_n1178_), .A2(new_n1176_), .ZN(new_n1179_));
  MUX2_X1    g1043(.I0(new_n1179_), .I1(new_n1173_), .S(new_n1174_), .Z(new_n1180_));
  INV_X1     g1044(.I(new_n1180_), .ZN(new_n1181_));
  NOR2_X1    g1045(.A1(new_n873_), .A2(new_n1027_), .ZN(new_n1182_));
  NAND2_X1   g1046(.A1(new_n1181_), .A2(new_n1182_), .ZN(new_n1183_));
  NOR2_X1    g1047(.A1(new_n875_), .A2(new_n1021_), .ZN(new_n1184_));
  NAND2_X1   g1048(.A1(new_n1179_), .A2(new_n1184_), .ZN(new_n1185_));
  OAI21_X1   g1049(.A1(new_n1181_), .A2(new_n1184_), .B(new_n1185_), .ZN(new_n1186_));
  OR2_X2     g1050(.A1(new_n1186_), .A2(new_n1182_), .Z(new_n1187_));
  NAND2_X1   g1051(.A1(new_n1187_), .A2(new_n1183_), .ZN(new_n1188_));
  NOR2_X1    g1052(.A1(new_n869_), .A2(new_n1039_), .ZN(new_n1189_));
  NAND2_X1   g1053(.A1(new_n1188_), .A2(new_n1189_), .ZN(new_n1190_));
  INV_X1     g1054(.I(new_n1189_), .ZN(new_n1191_));
  NOR2_X1    g1055(.A1(new_n871_), .A2(new_n1033_), .ZN(new_n1192_));
  NAND2_X1   g1056(.A1(new_n1186_), .A2(new_n1192_), .ZN(new_n1193_));
  OR2_X2     g1057(.A1(new_n1188_), .A2(new_n1192_), .Z(new_n1194_));
  NAND3_X1   g1058(.A1(new_n1194_), .A2(new_n1191_), .A3(new_n1193_), .ZN(new_n1195_));
  NAND2_X1   g1059(.A1(new_n1195_), .A2(new_n1190_), .ZN(new_n1196_));
  NOR2_X1    g1060(.A1(new_n865_), .A2(new_n1051_), .ZN(new_n1197_));
  NAND2_X1   g1061(.A1(new_n1196_), .A2(new_n1197_), .ZN(new_n1198_));
  INV_X1     g1062(.I(new_n1197_), .ZN(new_n1199_));
  NAND2_X1   g1063(.A1(new_n1194_), .A2(new_n1193_), .ZN(new_n1200_));
  NOR2_X1    g1064(.A1(new_n867_), .A2(new_n1045_), .ZN(new_n1201_));
  NAND2_X1   g1065(.A1(new_n1200_), .A2(new_n1201_), .ZN(new_n1202_));
  INV_X1     g1066(.I(new_n1201_), .ZN(new_n1203_));
  NAND3_X1   g1067(.A1(new_n1195_), .A2(new_n1190_), .A3(new_n1203_), .ZN(new_n1204_));
  NAND3_X1   g1068(.A1(new_n1204_), .A2(new_n1199_), .A3(new_n1202_), .ZN(new_n1205_));
  NAND2_X1   g1069(.A1(new_n1205_), .A2(new_n1198_), .ZN(new_n1206_));
  NOR2_X1    g1070(.A1(new_n861_), .A2(new_n1063_), .ZN(new_n1207_));
  NAND2_X1   g1071(.A1(new_n1206_), .A2(new_n1207_), .ZN(new_n1208_));
  INV_X1     g1072(.I(new_n1207_), .ZN(new_n1209_));
  NAND2_X1   g1073(.A1(new_n1204_), .A2(new_n1202_), .ZN(new_n1210_));
  NOR2_X1    g1074(.A1(new_n863_), .A2(new_n1057_), .ZN(new_n1211_));
  NAND2_X1   g1075(.A1(new_n1210_), .A2(new_n1211_), .ZN(new_n1212_));
  INV_X1     g1076(.I(new_n1211_), .ZN(new_n1213_));
  NAND3_X1   g1077(.A1(new_n1205_), .A2(new_n1198_), .A3(new_n1213_), .ZN(new_n1214_));
  NAND3_X1   g1078(.A1(new_n1214_), .A2(new_n1209_), .A3(new_n1212_), .ZN(new_n1215_));
  NAND2_X1   g1079(.A1(new_n1215_), .A2(new_n1208_), .ZN(new_n1216_));
  NAND2_X1   g1080(.A1(new_n1216_), .A2(new_n1111_), .ZN(new_n1217_));
  NAND2_X1   g1081(.A1(new_n1214_), .A2(new_n1212_), .ZN(new_n1218_));
  NOR2_X1    g1082(.A1(new_n859_), .A2(new_n1069_), .ZN(new_n1219_));
  NAND2_X1   g1083(.A1(new_n1218_), .A2(new_n1219_), .ZN(new_n1220_));
  INV_X1     g1084(.I(new_n1219_), .ZN(new_n1221_));
  NAND3_X1   g1085(.A1(new_n1215_), .A2(new_n1208_), .A3(new_n1221_), .ZN(new_n1222_));
  NAND2_X1   g1086(.A1(new_n1222_), .A2(new_n1220_), .ZN(new_n1223_));
  OAI21_X1   g1087(.A1(new_n1223_), .A2(new_n1111_), .B(new_n1217_), .ZN(new_n1224_));
  NOR2_X1    g1088(.A1(new_n853_), .A2(new_n1089_), .ZN(new_n1225_));
  NOR2_X1    g1089(.A1(new_n855_), .A2(new_n1081_), .ZN(new_n1226_));
  NAND2_X1   g1090(.A1(new_n1223_), .A2(new_n1226_), .ZN(new_n1227_));
  OAI21_X1   g1091(.A1(new_n1224_), .A2(new_n1226_), .B(new_n1227_), .ZN(new_n1228_));
  NOR2_X1    g1092(.A1(new_n1228_), .A2(new_n1225_), .ZN(new_n1229_));
  AOI21_X1   g1093(.A1(new_n1224_), .A2(new_n1225_), .B(new_n1229_), .ZN(new_n1230_));
  INV_X1     g1094(.I(new_n1230_), .ZN(new_n1231_));
  NOR2_X1    g1095(.A1(new_n1086_), .A2(new_n1100_), .ZN(new_n1232_));
  NOR2_X1    g1096(.A1(new_n1096_), .A2(new_n1105_), .ZN(new_n1233_));
  AOI21_X1   g1097(.A1(new_n1228_), .A2(new_n1232_), .B(new_n1233_), .ZN(new_n1234_));
  OAI21_X1   g1098(.A1(new_n1231_), .A2(new_n1232_), .B(new_n1234_), .ZN(new_n1235_));
  NAND2_X1   g1099(.A1(new_n1231_), .A2(new_n1233_), .ZN(new_n1236_));
  NAND2_X1   g1100(.A1(new_n1235_), .A2(new_n1236_), .ZN(\P[2] ));
  NOR2_X1    g1101(.A1(new_n1149_), .A2(new_n1112_), .ZN(new_n1238_));
  INV_X1     g1102(.I(new_n1238_), .ZN(new_n1239_));
  NOR2_X1    g1103(.A1(new_n1116_), .A2(new_n1113_), .ZN(new_n1240_));
  INV_X1     g1104(.I(new_n1240_), .ZN(new_n1241_));
  NOR4_X1    g1105(.A1(new_n904_), .A2(new_n908_), .A3(new_n912_), .A4(new_n922_), .ZN(new_n1242_));
  NAND2_X1   g1106(.A1(new_n1119_), .A2(new_n1131_), .ZN(new_n1243_));
  AOI21_X1   g1107(.A1(new_n1243_), .A2(new_n1242_), .B(new_n1241_), .ZN(new_n1244_));
  NOR2_X1    g1108(.A1(new_n1244_), .A2(new_n1239_), .ZN(new_n1245_));
  INV_X1     g1109(.I(new_n1244_), .ZN(new_n1246_));
  NOR3_X1    g1110(.A1(new_n1140_), .A2(\A[102] ), .A3(new_n952_), .ZN(new_n1247_));
  NOR2_X1    g1111(.A1(new_n1246_), .A2(new_n1247_), .ZN(new_n1248_));
  OAI21_X1   g1112(.A1(new_n1243_), .A2(new_n207_), .B(new_n1242_), .ZN(new_n1249_));
  AND3_X2    g1113(.A1(new_n1249_), .A2(new_n1240_), .A3(new_n1247_), .Z(new_n1250_));
  NOR2_X1    g1114(.A1(new_n1248_), .A2(new_n1250_), .ZN(new_n1251_));
  AOI21_X1   g1115(.A1(new_n1251_), .A2(new_n1239_), .B(new_n1245_), .ZN(new_n1252_));
  NOR2_X1    g1116(.A1(new_n1155_), .A2(new_n1169_), .ZN(new_n1253_));
  INV_X1     g1117(.I(new_n1253_), .ZN(new_n1254_));
  NOR2_X1    g1118(.A1(new_n1252_), .A2(new_n1254_), .ZN(new_n1255_));
  NOR2_X1    g1119(.A1(new_n1146_), .A2(new_n1159_), .ZN(new_n1256_));
  INV_X1     g1120(.I(new_n1256_), .ZN(new_n1257_));
  NAND2_X1   g1121(.A1(new_n1252_), .A2(new_n1257_), .ZN(new_n1258_));
  OAI21_X1   g1122(.A1(new_n1251_), .A2(new_n1257_), .B(new_n1258_), .ZN(new_n1259_));
  NOR2_X1    g1123(.A1(new_n1259_), .A2(new_n1253_), .ZN(new_n1260_));
  NOR2_X1    g1124(.A1(new_n1260_), .A2(new_n1255_), .ZN(new_n1261_));
  NAND2_X1   g1125(.A1(new_n1174_), .A2(new_n1184_), .ZN(new_n1262_));
  NOR2_X1    g1126(.A1(new_n1261_), .A2(new_n1262_), .ZN(new_n1263_));
  INV_X1     g1127(.I(new_n1262_), .ZN(new_n1264_));
  NOR2_X1    g1128(.A1(new_n1165_), .A2(new_n1177_), .ZN(new_n1265_));
  NAND2_X1   g1129(.A1(new_n1259_), .A2(new_n1265_), .ZN(new_n1266_));
  INV_X1     g1130(.I(new_n1265_), .ZN(new_n1267_));
  NAND2_X1   g1131(.A1(new_n1261_), .A2(new_n1267_), .ZN(new_n1268_));
  NAND2_X1   g1132(.A1(new_n1268_), .A2(new_n1266_), .ZN(new_n1269_));
  NOR2_X1    g1133(.A1(new_n1269_), .A2(new_n1264_), .ZN(new_n1270_));
  NOR2_X1    g1134(.A1(new_n1270_), .A2(new_n1263_), .ZN(new_n1271_));
  NOR2_X1    g1135(.A1(new_n1191_), .A2(new_n1203_), .ZN(new_n1272_));
  NAND2_X1   g1136(.A1(new_n1182_), .A2(new_n1192_), .ZN(new_n1273_));
  INV_X1     g1137(.I(new_n1273_), .ZN(new_n1274_));
  NAND2_X1   g1138(.A1(new_n1269_), .A2(new_n1274_), .ZN(new_n1275_));
  NAND2_X1   g1139(.A1(new_n1271_), .A2(new_n1273_), .ZN(new_n1276_));
  NAND2_X1   g1140(.A1(new_n1276_), .A2(new_n1275_), .ZN(new_n1277_));
  MUX2_X1    g1141(.I0(new_n1277_), .I1(new_n1271_), .S(new_n1272_), .Z(new_n1278_));
  INV_X1     g1142(.I(new_n1278_), .ZN(new_n1279_));
  NOR2_X1    g1143(.A1(new_n1209_), .A2(new_n1221_), .ZN(new_n1280_));
  NOR2_X1    g1144(.A1(new_n1199_), .A2(new_n1213_), .ZN(new_n1281_));
  NAND2_X1   g1145(.A1(new_n1277_), .A2(new_n1281_), .ZN(new_n1282_));
  OAI21_X1   g1146(.A1(new_n1279_), .A2(new_n1281_), .B(new_n1282_), .ZN(new_n1283_));
  NOR2_X1    g1147(.A1(new_n1283_), .A2(new_n1280_), .ZN(new_n1284_));
  AOI21_X1   g1148(.A1(new_n1279_), .A2(new_n1280_), .B(new_n1284_), .ZN(new_n1285_));
  NAND2_X1   g1149(.A1(new_n1225_), .A2(new_n1232_), .ZN(new_n1286_));
  INV_X1     g1150(.I(new_n1285_), .ZN(new_n1287_));
  NOR4_X1    g1151(.A1(new_n857_), .A2(new_n855_), .A3(new_n1075_), .A4(new_n1081_), .ZN(new_n1288_));
  INV_X1     g1152(.I(new_n1286_), .ZN(new_n1289_));
  AOI21_X1   g1153(.A1(new_n1283_), .A2(new_n1288_), .B(new_n1289_), .ZN(new_n1290_));
  OAI21_X1   g1154(.A1(new_n1287_), .A2(new_n1288_), .B(new_n1290_), .ZN(new_n1291_));
  OAI21_X1   g1155(.A1(new_n1285_), .A2(new_n1286_), .B(new_n1291_), .ZN(\P[3] ));
  NAND2_X1   g1156(.A1(new_n1264_), .A2(new_n1274_), .ZN(new_n1293_));
  NAND2_X1   g1157(.A1(new_n1240_), .A2(new_n1242_), .ZN(new_n1294_));
  NOR3_X1    g1158(.A1(new_n1243_), .A2(new_n1128_), .A3(new_n1140_), .ZN(new_n1295_));
  NOR2_X1    g1159(.A1(new_n1257_), .A2(new_n1239_), .ZN(new_n1296_));
  INV_X1     g1160(.I(new_n1296_), .ZN(new_n1297_));
  AOI21_X1   g1161(.A1(new_n1297_), .A2(new_n1295_), .B(new_n1294_), .ZN(new_n1298_));
  NOR2_X1    g1162(.A1(new_n1298_), .A2(new_n1293_), .ZN(new_n1299_));
  NAND4_X1   g1163(.A1(new_n1265_), .A2(new_n701_), .A3(new_n1167_), .A4(new_n990_), .ZN(new_n1300_));
  OAI21_X1   g1164(.A1(new_n1297_), .A2(new_n291_), .B(new_n1295_), .ZN(new_n1301_));
  NOR2_X1    g1165(.A1(new_n1300_), .A2(new_n1294_), .ZN(new_n1302_));
  AOI22_X1   g1166(.A1(new_n1298_), .A2(new_n1300_), .B1(new_n1301_), .B2(new_n1302_), .ZN(new_n1303_));
  AOI21_X1   g1167(.A1(new_n1303_), .A2(new_n1293_), .B(new_n1299_), .ZN(new_n1304_));
  NAND2_X1   g1168(.A1(new_n1272_), .A2(new_n1281_), .ZN(new_n1305_));
  AND2_X2    g1169(.A1(new_n1304_), .A2(new_n1305_), .Z(new_n1306_));
  NAND2_X1   g1170(.A1(new_n1280_), .A2(new_n1288_), .ZN(new_n1307_));
  OAI21_X1   g1171(.A1(new_n1303_), .A2(new_n1305_), .B(new_n1307_), .ZN(new_n1308_));
  OAI22_X1   g1172(.A1(new_n1306_), .A2(new_n1308_), .B1(new_n1304_), .B2(new_n1307_), .ZN(\P[4] ));
  INV_X1     g1173(.I(new_n1295_), .ZN(new_n1310_));
  NOR2_X1    g1174(.A1(new_n1310_), .A2(new_n1294_), .ZN(new_n1311_));
  NOR3_X1    g1175(.A1(new_n1297_), .A2(new_n1254_), .A3(new_n1267_), .ZN(new_n1312_));
  INV_X1     g1176(.I(new_n1312_), .ZN(new_n1313_));
  NOR2_X1    g1177(.A1(new_n1305_), .A2(new_n1293_), .ZN(new_n1314_));
  OAI21_X1   g1178(.A1(new_n1313_), .A2(new_n1314_), .B(new_n1311_), .ZN(\P[5] ));
  NAND2_X1   g1179(.A1(new_n1312_), .A2(new_n1311_), .ZN(\P[6] ));
  NOR2_X1    g1180(.A1(\A[0] ), .A2(\A[1] ), .ZN(new_n1317_));
  NAND4_X1   g1181(.A1(new_n1289_), .A2(new_n1107_), .A3(new_n1233_), .A4(new_n1317_), .ZN(new_n1318_));
  NOR2_X1    g1182(.A1(new_n1318_), .A2(new_n1307_), .ZN(new_n1319_));
  NAND4_X1   g1183(.A1(new_n1312_), .A2(new_n1311_), .A3(new_n1314_), .A4(new_n1319_), .ZN(F));
endmodule


