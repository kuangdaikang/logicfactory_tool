// Benchmark "source.pla" written by ABC on Fri Feb 25 15:13:08 2022

module exp  ( 
    v0, v1, v2, v3, v4, v5, v6, v7,
    \v8.0 , \v8.1 , \v8.2 , \v8.3 , \v8.4 , \v8.5 , \v8.6 , \v8.7 , \v8.8 ,
    \v8.9 , \v8.10 , \v8.11 , \v8.12 , \v8.13 , \v8.14 , \v8.15 , \v8.16 ,
    \v8.17   );
  input  v0, v1, v2, v3, v4, v5, v6, v7;
  output \v8.0 , \v8.1 , \v8.2 , \v8.3 , \v8.4 , \v8.5 , \v8.6 , \v8.7 ,
    \v8.8 , \v8.9 , \v8.10 , \v8.11 , \v8.12 , \v8.13 , \v8.14 , \v8.15 ,
    \v8.16 , \v8.17 ;
  wire new_n28_, new_n29_, new_n30_, new_n31_, new_n32_, new_n33_, new_n34_,
    new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_, new_n41_,
    new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n48_, new_n49_,
    new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_,
    new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_,
    new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_;
  assign new_n28_ = ~v5 & v6;
  assign new_n29_ = v5 & ~v6;
  assign new_n30_ = ~new_n28_ & ~new_n29_;
  assign new_n31_ = v1 & ~new_n30_;
  assign new_n32_ = ~v1 & new_n28_;
  assign new_n33_ = ~new_n31_ & ~new_n32_;
  assign new_n34_ = ~v6 & v7;
  assign new_n35_ = ~v5 & new_n34_;
  assign new_n36_ = new_n33_ & ~new_n35_;
  assign new_n37_ = ~v2 & v6;
  assign new_n38_ = v1 & new_n37_;
  assign new_n39_ = v2 & ~v6;
  assign new_n40_ = ~v1 & new_n39_;
  assign new_n41_ = ~new_n38_ & ~new_n40_;
  assign new_n42_ = ~v7 & ~new_n41_;
  assign new_n43_ = v5 & new_n42_;
  assign new_n44_ = new_n36_ & ~new_n43_;
  assign new_n45_ = ~v4 & ~new_n44_;
  assign new_n46_ = ~v3 & new_n45_;
  assign \v8.0  = ~v0 & new_n46_;
  assign new_n48_ = ~v1 & ~v5;
  assign new_n49_ = ~v1 & ~new_n48_;
  assign new_n50_ = v6 & ~new_n49_;
  assign new_n51_ = ~v1 & new_n29_;
  assign new_n52_ = ~new_n50_ & ~new_n51_;
  assign new_n53_ = ~v4 & ~new_n52_;
  assign new_n54_ = v5 & v6;
  assign new_n55_ = ~v5 & ~v6;
  assign new_n56_ = ~new_n54_ & ~new_n55_;
  assign new_n57_ = v4 & ~new_n56_;
  assign new_n58_ = ~v1 & new_n57_;
  assign new_n59_ = ~new_n53_ & ~new_n58_;
  assign new_n60_ = v0 & ~new_n59_;
  assign new_n61_ = ~v4 & ~new_n33_;
  assign new_n62_ = ~v0 & new_n61_;
  assign new_n63_ = ~new_n60_ & ~new_n62_;
  assign new_n64_ = ~v2 & new_n28_;
  assign new_n65_ = v2 & new_n29_;
  assign new_n66_ = ~new_n64_ & ~new_n65_;
  assign new_n67_ = v4 & ~new_n66_;
  assign new_n68_ = ~v1 & new_n67_;
  assign new_n69_ = v0 & new_n68_;
  assign new_n70_ = new_n63_ & ~new_n69_;
  assign new_n71_ = ~v3 & ~new_n70_;
  assign new_n72_ = ~v1 & ~v2;
  assign new_n73_ = v0 & new_n72_;
  assign new_n74_ = v3 & ~v4;
  assign new_n75_ = new_n55_ & new_n74_;
  assign new_n76_ = new_n73_ & new_n75_;
  assign new_n77_ = ~new_n71_ & ~new_n76_;
  assign new_n78_ = ~v1 & new_n37_;
  assign new_n79_ = v1 & new_n39_;
  assign new_n80_ = ~new_n78_ & ~new_n79_;
  assign new_n81_ = v0 & ~new_n80_;
  assign new_n82_ = ~v0 & ~new_n41_;
  assign new_n83_ = ~new_n81_ & ~new_n82_;
  assign new_n84_ = ~v4 & ~new_n83_;
  assign new_n85_ = v0 & ~v1;
  assign new_n86_ = v4 & ~v6;
  assign new_n87_ = ~v2 & new_n86_;
  assign new_n88_ = new_n85_ & new_n87_;
  assign new_n89_ = ~new_n84_ & ~new_n88_;
  assign new_n90_ = v5 & ~new_n89_;
  assign new_n91_ = ~v1 & v6;
  assign new_n92_ = v1 & ~v6;
  assign new_n93_ = ~new_n91_ & ~new_n92_;
  assign new_n94_ = ~v5 & ~new_n93_;
  assign new_n95_ = v4 & new_n94_;
  assign new_n96_ = v2 & new_n95_;
  assign new_n97_ = v0 & new_n96_;
  assign new_n98_ = ~new_n90_ & ~new_n97_;
  assign new_n99_ = ~v7 & ~new_n98_;
  assign new_n100_ = ~v1 & v2;
  assign new_n101_ = v0 & new_n100_;
  assign new_n102_ = ~v4 & v5;
  assign new_n103_ = v6 & v7;
  assign new_n104_ = new_n102_ & new_n103_;
  assign new_n105_ = new_n101_ & new_n104_;
  assign new_n106_ = ~new_n99_ & ~new_n105_;
  assign new_n107_ = ~v3 & ~new_n106_;
  assign new_n108_ = ~v2 & v3;
  assign new_n109_ = new_n85_ & new_n108_;
  assign new_n110_ = ~v4 & ~v5;
  assign new_n111_ = v6 & ~v7;
  assign new_n112_ = new_n110_ & new_n111_;
  assign new_n113_ = new_n109_ & new_n112_;
  assign new_n114_ = ~new_n107_ & ~new_n113_;
  assign \v8.1  = ~new_n77_ | ~new_n114_;
  assign new_n116_ = v2 & v4;
  assign new_n117_ = ~v1 & new_n116_;
  assign new_n118_ = v1 & ~v2;
  assign new_n119_ = ~v4 & v6;
  assign new_n120_ = new_n118_ & new_n119_;
  assign new_n121_ = ~new_n117_ & ~new_n120_;
  assign new_n122_ = ~v4 & new_n34_;
  assign new_n123_ = new_n118_ & new_n122_;
  assign new_n124_ = new_n121_ & ~new_n123_;
  assign new_n125_ = v5 & ~new_n124_;
  assign new_n126_ = ~v5 & new_n103_;
  assign new_n127_ = new_n117_ & new_n126_;
  assign new_n128_ = ~new_n125_ & ~new_n127_;
  assign new_n129_ = ~v3 & ~new_n128_;
  assign \v8.2  = v0 & new_n129_;
  assign new_n131_ = v4 & v6;
  assign new_n132_ = ~v4 & ~v6;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_ = v2 & ~new_n133_;
  assign new_n135_ = ~v2 & new_n132_;
  assign new_n136_ = ~new_n134_ & ~new_n135_;
  assign new_n137_ = ~v5 & ~new_n136_;
  assign new_n138_ = ~new_n86_ & ~new_n119_;
  assign new_n139_ = v5 & ~new_n138_;
  assign new_n140_ = ~v2 & new_n139_;
  assign new_n141_ = ~new_n137_ & ~new_n140_;
  assign new_n142_ = ~v1 & ~new_n141_;
  assign new_n143_ = v1 & new_n132_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = v0 & ~new_n144_;
  assign new_n146_ = ~v4 & new_n55_;
  assign new_n147_ = ~v0 & new_n146_;
  assign new_n148_ = ~new_n145_ & ~new_n147_;
  assign new_n149_ = v7 & ~new_n148_;
  assign new_n150_ = new_n102_ & new_n111_;
  assign new_n151_ = new_n101_ & new_n150_;
  assign new_n152_ = ~new_n149_ & ~new_n151_;
  assign \v8.5  = ~v3 & ~new_n152_;
  assign new_n154_ = ~v0 & v1;
  assign new_n155_ = ~new_n85_ & ~new_n154_;
  assign new_n156_ = v5 & new_n111_;
  assign new_n157_ = ~new_n35_ & ~new_n156_;
  assign new_n158_ = ~v2 & ~new_n157_;
  assign new_n159_ = v2 & ~v5;
  assign new_n160_ = new_n34_ & new_n159_;
  assign new_n161_ = ~new_n158_ & ~new_n160_;
  assign new_n162_ = new_n30_ & new_n161_;
  assign new_n163_ = ~new_n155_ & ~new_n162_;
  assign new_n164_ = v0 & v1;
  assign new_n165_ = ~v0 & ~v1;
  assign new_n166_ = ~new_n164_ & ~new_n165_;
  assign new_n167_ = ~v6 & ~new_n34_;
  assign new_n168_ = ~v5 & ~new_n167_;
  assign new_n169_ = v2 & v5;
  assign new_n170_ = ~v6 & ~v7;
  assign new_n171_ = new_n169_ & new_n170_;
  assign new_n172_ = ~new_n168_ & ~new_n171_;
  assign new_n173_ = ~new_n166_ & ~new_n172_;
  assign new_n174_ = ~new_n163_ & ~new_n173_;
  assign new_n175_ = ~v4 & ~new_n174_;
  assign \v8.6  = ~v3 & new_n175_;
  assign new_n177_ = v1 & v7;
  assign new_n178_ = v5 & ~v7;
  assign new_n179_ = ~v1 & new_n178_;
  assign new_n180_ = ~new_n177_ & ~new_n179_;
  assign new_n181_ = ~v4 & ~new_n180_;
  assign new_n182_ = ~v2 & new_n181_;
  assign new_n183_ = v5 & v7;
  assign new_n184_ = ~v5 & ~v7;
  assign new_n185_ = ~new_n183_ & ~new_n184_;
  assign new_n186_ = v4 & ~new_n185_;
  assign new_n187_ = v2 & new_n186_;
  assign new_n188_ = ~v1 & new_n187_;
  assign new_n189_ = ~new_n182_ & ~new_n188_;
  assign new_n190_ = v6 & ~new_n189_;
  assign new_n191_ = ~v4 & v7;
  assign new_n192_ = v2 & new_n191_;
  assign new_n193_ = v4 & ~v7;
  assign new_n194_ = ~v2 & new_n193_;
  assign new_n195_ = ~new_n192_ & ~new_n194_;
  assign new_n196_ = ~v1 & ~new_n195_;
  assign new_n197_ = v1 & v2;
  assign new_n198_ = ~v4 & ~v7;
  assign new_n199_ = new_n197_ & new_n198_;
  assign new_n200_ = ~new_n196_ & ~new_n199_;
  assign new_n201_ = ~v6 & ~new_n200_;
  assign new_n202_ = v5 & new_n201_;
  assign new_n203_ = ~new_n190_ & ~new_n202_;
  assign new_n204_ = v0 & ~new_n203_;
  assign new_n205_ = v2 & new_n34_;
  assign new_n206_ = ~v2 & new_n111_;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = v1 & ~new_n207_;
  assign new_n209_ = new_n100_ & new_n170_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = v5 & ~new_n210_;
  assign new_n212_ = new_n72_ & new_n126_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~v4 & ~new_n213_;
  assign new_n215_ = ~v0 & new_n214_;
  assign new_n216_ = ~new_n204_ & ~new_n215_;
  assign new_n217_ = ~v3 & ~new_n216_;
  assign \v8.7  = new_n113_ | new_n217_;
  assign new_n219_ = ~v1 & v4;
  assign new_n220_ = v1 & ~v4;
  assign new_n221_ = ~new_n219_ & ~new_n220_;
  assign new_n222_ = v6 & ~new_n221_;
  assign new_n223_ = v0 & new_n222_;
  assign new_n224_ = new_n132_ & new_n154_;
  assign new_n225_ = ~new_n223_ & ~new_n224_;
  assign new_n226_ = v2 & new_n86_;
  assign new_n227_ = new_n85_ & new_n226_;
  assign new_n228_ = new_n225_ & ~new_n227_;
  assign new_n229_ = v5 & ~new_n228_;
  assign new_n230_ = ~v4 & new_n28_;
  assign new_n231_ = ~v0 & new_n230_;
  assign new_n232_ = ~new_n229_ & ~new_n231_;
  assign new_n233_ = ~v3 & ~new_n232_;
  assign new_n234_ = ~new_n76_ & ~new_n233_;
  assign new_n235_ = ~v5 & v7;
  assign new_n236_ = v4 & new_n235_;
  assign new_n237_ = new_n101_ & new_n236_;
  assign new_n238_ = ~v0 & new_n118_;
  assign new_n239_ = ~v4 & new_n178_;
  assign new_n240_ = new_n238_ & new_n239_;
  assign new_n241_ = ~new_n237_ & ~new_n240_;
  assign new_n242_ = v6 & ~new_n241_;
  assign new_n243_ = ~v4 & new_n183_;
  assign new_n244_ = v4 & new_n184_;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = v2 & ~new_n245_;
  assign new_n247_ = ~v2 & ~v4;
  assign new_n248_ = new_n183_ & new_n247_;
  assign new_n249_ = ~new_n246_ & ~new_n248_;
  assign new_n250_ = v1 & ~new_n249_;
  assign new_n251_ = v4 & new_n183_;
  assign new_n252_ = new_n72_ & new_n251_;
  assign new_n253_ = ~new_n250_ & ~new_n252_;
  assign new_n254_ = v0 & ~new_n253_;
  assign new_n255_ = new_n100_ & new_n178_;
  assign new_n256_ = ~new_n235_ & ~new_n255_;
  assign new_n257_ = ~v4 & ~new_n256_;
  assign new_n258_ = ~v0 & new_n257_;
  assign new_n259_ = ~new_n254_ & ~new_n258_;
  assign new_n260_ = ~v6 & ~new_n259_;
  assign new_n261_ = ~new_n242_ & ~new_n260_;
  assign new_n262_ = ~v3 & ~new_n261_;
  assign new_n263_ = ~new_n113_ & ~new_n262_;
  assign \v8.8  = ~new_n234_ | ~new_n263_;
  assign new_n265_ = v4 & new_n28_;
  assign new_n266_ = ~v4 & new_n29_;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = ~new_n140_ & new_n267_;
  assign new_n269_ = ~v1 & ~new_n268_;
  assign new_n270_ = new_n197_ & new_n266_;
  assign new_n271_ = ~new_n269_ & ~new_n270_;
  assign new_n272_ = v4 & ~v5;
  assign new_n273_ = new_n34_ & new_n272_;
  assign new_n274_ = ~new_n150_ & ~new_n273_;
  assign new_n275_ = v2 & ~new_n274_;
  assign new_n276_ = ~v1 & new_n275_;
  assign new_n277_ = v1 & new_n247_;
  assign new_n278_ = v5 & new_n170_;
  assign new_n279_ = new_n277_ & new_n278_;
  assign new_n280_ = ~new_n276_ & ~new_n279_;
  assign new_n281_ = new_n271_ & new_n280_;
  assign new_n282_ = ~v3 & ~new_n281_;
  assign \v8.9  = v0 & new_n282_;
  assign new_n284_ = ~v2 & new_n34_;
  assign new_n285_ = v2 & new_n111_;
  assign new_n286_ = ~new_n284_ & ~new_n285_;
  assign new_n287_ = v1 & ~new_n286_;
  assign new_n288_ = new_n100_ & new_n103_;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign new_n290_ = ~v4 & ~new_n289_;
  assign new_n291_ = ~new_n37_ & ~new_n39_;
  assign new_n292_ = ~v7 & ~new_n291_;
  assign new_n293_ = v4 & new_n292_;
  assign new_n294_ = ~v1 & new_n293_;
  assign new_n295_ = ~new_n290_ & ~new_n294_;
  assign new_n296_ = v5 & ~new_n295_;
  assign new_n297_ = ~v2 & v4;
  assign new_n298_ = ~v1 & new_n297_;
  assign new_n299_ = ~v5 & new_n170_;
  assign new_n300_ = new_n298_ & new_n299_;
  assign new_n301_ = ~new_n296_ & ~new_n300_;
  assign new_n302_ = ~v3 & ~new_n301_;
  assign \v8.10  = v0 & new_n302_;
  assign new_n304_ = v2 & v7;
  assign new_n305_ = ~v2 & ~v7;
  assign new_n306_ = ~new_n304_ & ~new_n305_;
  assign new_n307_ = ~v4 & ~new_n306_;
  assign new_n308_ = v1 & new_n307_;
  assign new_n309_ = v4 & v7;
  assign new_n310_ = new_n72_ & new_n309_;
  assign new_n311_ = ~new_n308_ & ~new_n310_;
  assign new_n312_ = v6 & ~new_n311_;
  assign new_n313_ = v4 & new_n34_;
  assign new_n314_ = new_n100_ & new_n313_;
  assign new_n315_ = ~new_n312_ & ~new_n314_;
  assign new_n316_ = v5 & ~new_n315_;
  assign new_n317_ = ~v2 & v7;
  assign new_n318_ = v2 & ~v7;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = ~v6 & ~new_n319_;
  assign new_n321_ = ~v5 & new_n320_;
  assign new_n322_ = v4 & new_n321_;
  assign new_n323_ = ~v1 & new_n322_;
  assign new_n324_ = ~new_n316_ & ~new_n323_;
  assign new_n325_ = ~v3 & ~new_n324_;
  assign \v8.11  = v0 & new_n325_;
  assign new_n327_ = ~v4 & ~new_n102_;
  assign new_n328_ = ~v3 & ~new_n327_;
  assign new_n329_ = ~v2 & new_n328_;
  assign new_n330_ = ~v1 & new_n329_;
  assign \v8.12  = v0 & new_n330_;
  assign new_n332_ = ~new_n102_ & ~new_n272_;
  assign new_n333_ = v4 & new_n29_;
  assign new_n334_ = new_n332_ & ~new_n333_;
  assign new_n335_ = ~v3 & ~new_n334_;
  assign new_n336_ = v2 & new_n335_;
  assign new_n337_ = ~v1 & new_n336_;
  assign \v8.13  = v0 & new_n337_;
  assign new_n339_ = v2 & ~v3;
  assign new_n340_ = v4 & v5;
  assign new_n341_ = new_n339_ & new_n340_;
  assign new_n342_ = new_n108_ & new_n110_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = ~v1 & ~new_n343_;
  assign new_n345_ = v0 & new_n344_;
  assign new_n346_ = ~v3 & new_n102_;
  assign new_n347_ = new_n238_ & new_n346_;
  assign new_n348_ = ~new_n345_ & ~new_n347_;
  assign new_n349_ = ~new_n72_ & ~new_n197_;
  assign new_n350_ = ~new_n138_ & ~new_n349_;
  assign new_n351_ = ~new_n100_ & ~new_n118_;
  assign new_n352_ = v6 & ~new_n351_;
  assign new_n353_ = ~v4 & new_n352_;
  assign new_n354_ = ~new_n350_ & ~new_n353_;
  assign new_n355_ = ~v5 & ~new_n354_;
  assign new_n356_ = ~new_n220_ & ~new_n298_;
  assign new_n357_ = v6 & ~new_n356_;
  assign new_n358_ = v5 & new_n357_;
  assign new_n359_ = ~new_n355_ & ~new_n358_;
  assign new_n360_ = v0 & ~new_n359_;
  assign new_n361_ = v2 & ~new_n30_;
  assign new_n362_ = ~new_n64_ & ~new_n361_;
  assign new_n363_ = ~v4 & ~new_n362_;
  assign new_n364_ = ~v0 & new_n363_;
  assign new_n365_ = ~new_n360_ & ~new_n364_;
  assign new_n366_ = ~v3 & ~new_n365_;
  assign new_n367_ = new_n348_ & ~new_n366_;
  assign new_n368_ = v2 & v6;
  assign new_n369_ = ~v1 & new_n368_;
  assign new_n370_ = ~v2 & ~v6;
  assign new_n371_ = v1 & new_n370_;
  assign new_n372_ = ~new_n369_ & ~new_n371_;
  assign new_n373_ = v7 & ~new_n372_;
  assign new_n374_ = v0 & new_n373_;
  assign new_n375_ = v1 & new_n368_;
  assign new_n376_ = ~v1 & new_n370_;
  assign new_n377_ = ~new_n375_ & ~new_n376_;
  assign new_n378_ = ~v7 & ~new_n377_;
  assign new_n379_ = ~v0 & new_n378_;
  assign new_n380_ = ~new_n374_ & ~new_n379_;
  assign new_n381_ = v5 & ~new_n380_;
  assign new_n382_ = ~v4 & new_n381_;
  assign new_n383_ = new_n170_ & new_n272_;
  assign new_n384_ = new_n101_ & new_n383_;
  assign new_n385_ = ~new_n382_ & ~new_n384_;
  assign new_n386_ = ~v3 & ~new_n385_;
  assign new_n387_ = v2 & v3;
  assign new_n388_ = new_n85_ & new_n387_;
  assign new_n389_ = new_n110_ & new_n170_;
  assign new_n390_ = new_n388_ & new_n389_;
  assign new_n391_ = ~new_n386_ & ~new_n390_;
  assign \v8.14  = ~new_n367_ | ~new_n391_;
  assign new_n393_ = v2 & new_n235_;
  assign new_n394_ = ~v2 & new_n178_;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign new_n396_ = v3 & ~new_n395_;
  assign new_n397_ = v0 & new_n396_;
  assign new_n398_ = ~v0 & ~v2;
  assign new_n399_ = ~v3 & new_n183_;
  assign new_n400_ = new_n398_ & new_n399_;
  assign new_n401_ = ~new_n397_ & ~new_n400_;
  assign new_n402_ = ~v6 & ~new_n401_;
  assign new_n403_ = ~v0 & new_n339_;
  assign new_n404_ = new_n156_ & new_n403_;
  assign new_n405_ = ~new_n402_ & ~new_n404_;
  assign new_n406_ = ~v1 & ~new_n405_;
  assign new_n407_ = ~v0 & new_n197_;
  assign new_n408_ = ~v3 & v5;
  assign new_n409_ = new_n103_ & new_n408_;
  assign new_n410_ = new_n407_ & new_n409_;
  assign new_n411_ = ~new_n406_ & ~new_n410_;
  assign new_n412_ = ~v4 & ~new_n411_;
  assign new_n413_ = ~new_n368_ & ~new_n370_;
  assign new_n414_ = v0 & ~new_n413_;
  assign new_n415_ = ~v0 & new_n370_;
  assign new_n416_ = ~new_n414_ & ~new_n415_;
  assign new_n417_ = ~v7 & ~new_n416_;
  assign new_n418_ = ~v5 & new_n417_;
  assign new_n419_ = v4 & new_n418_;
  assign new_n420_ = ~v3 & new_n419_;
  assign new_n421_ = v1 & new_n420_;
  assign \v8.15  = new_n412_ | new_n421_;
  assign new_n423_ = v1 & new_n339_;
  assign new_n424_ = new_n265_ & new_n423_;
  assign new_n425_ = ~v1 & new_n108_;
  assign new_n426_ = new_n266_ & new_n425_;
  assign new_n427_ = ~new_n424_ & ~new_n426_;
  assign new_n428_ = v0 & ~new_n427_;
  assign new_n429_ = ~v4 & new_n54_;
  assign new_n430_ = new_n100_ & new_n429_;
  assign new_n431_ = v4 & new_n55_;
  assign new_n432_ = new_n118_ & new_n431_;
  assign new_n433_ = ~new_n430_ & ~new_n432_;
  assign new_n434_ = ~v3 & ~new_n433_;
  assign new_n435_ = ~v0 & new_n434_;
  assign new_n436_ = ~new_n428_ & ~new_n435_;
  assign new_n437_ = v7 & ~new_n436_;
  assign new_n438_ = new_n72_ & new_n429_;
  assign new_n439_ = new_n197_ & new_n431_;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~v7 & ~new_n440_;
  assign new_n442_ = ~v3 & new_n441_;
  assign new_n443_ = ~v0 & new_n442_;
  assign \v8.16  = new_n437_ | new_n443_;
  assign new_n445_ = v7 & ~new_n413_;
  assign new_n446_ = v4 & new_n445_;
  assign new_n447_ = ~v3 & new_n446_;
  assign new_n448_ = v1 & new_n447_;
  assign new_n449_ = ~v1 & new_n387_;
  assign new_n450_ = ~v4 & new_n111_;
  assign new_n451_ = new_n449_ & new_n450_;
  assign new_n452_ = ~new_n448_ & ~new_n451_;
  assign new_n453_ = ~v5 & ~new_n452_;
  assign new_n454_ = new_n34_ & new_n102_;
  assign new_n455_ = new_n425_ & new_n454_;
  assign new_n456_ = ~new_n453_ & ~new_n455_;
  assign new_n457_ = v0 & ~new_n456_;
  assign new_n458_ = v1 & new_n322_;
  assign new_n459_ = v6 & ~new_n306_;
  assign new_n460_ = v5 & new_n459_;
  assign new_n461_ = ~v4 & new_n460_;
  assign new_n462_ = ~v1 & new_n461_;
  assign new_n463_ = ~new_n458_ & ~new_n462_;
  assign new_n464_ = ~v3 & ~new_n463_;
  assign new_n465_ = ~v0 & new_n464_;
  assign \v8.17  = new_n457_ | new_n465_;
  assign \v8.3  = 1'b0;
  assign \v8.4  = 1'b0;
endmodule


