// Benchmark "voter" written by ABC on Thu Sep 14 22:52:17 2023

module voter ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1323_, new_n1324_, new_n1325_, new_n1326_,
    new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_,
    new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_,
    new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_, new_n1344_,
    new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_, new_n1350_,
    new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_, new_n1356_,
    new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_, new_n1362_,
    new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_, new_n1368_,
    new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_, new_n1374_,
    new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_, new_n1380_,
    new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_,
    new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_,
    new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_,
    new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_,
    new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_, new_n1458_,
    new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_, new_n1464_,
    new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_, new_n1470_,
    new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_, new_n1476_,
    new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1500_,
    new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_,
    new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_, new_n1530_,
    new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_,
    new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_, new_n1554_,
    new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_, new_n1560_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_, new_n1644_,
    new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_,
    new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_,
    new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_,
    new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_,
    new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_,
    new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_,
    new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_,
    new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_,
    new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_,
    new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_,
    new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_, new_n1890_,
    new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_, new_n1902_,
    new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_, new_n1908_,
    new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_, new_n1914_,
    new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_, new_n1920_,
    new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_, new_n1926_,
    new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_, new_n1932_,
    new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_, new_n1938_,
    new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_, new_n1944_,
    new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_,
    new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_,
    new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_, new_n1992_,
    new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_, new_n1998_,
    new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_, new_n2004_,
    new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_, new_n2010_,
    new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_, new_n2016_,
    new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_, new_n2022_,
    new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_, new_n2028_,
    new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_, new_n2034_,
    new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_, new_n2040_,
    new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_, new_n2046_,
    new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_, new_n2052_,
    new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_, new_n2058_,
    new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_, new_n2064_,
    new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_, new_n2070_,
    new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_, new_n2076_,
    new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_, new_n2082_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_,
    new_n2120_, new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_,
    new_n2126_, new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_,
    new_n2132_, new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_,
    new_n2138_, new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_,
    new_n2144_, new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_,
    new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_,
    new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_,
    new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_,
    new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_,
    new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_,
    new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_,
    new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_,
    new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_,
    new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_,
    new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_,
    new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_,
    new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_,
    new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_,
    new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_,
    new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_,
    new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_,
    new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_,
    new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_,
    new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_,
    new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_,
    new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_,
    new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_,
    new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_,
    new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_,
    new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_,
    new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_,
    new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_,
    new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_,
    new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_,
    new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_,
    new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_, new_n2509_,
    new_n2510_, new_n2511_, new_n2512_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2621_, new_n2622_, new_n2623_,
    new_n2624_, new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_,
    new_n2630_, new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_,
    new_n2636_, new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_,
    new_n2642_, new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_,
    new_n2648_, new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_,
    new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_,
    new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_,
    new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_,
    new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_,
    new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_,
    new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_,
    new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_,
    new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_,
    new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_,
    new_n2708_, new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_, new_n2779_,
    new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_,
    new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_,
    new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_,
    new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_,
    new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_,
    new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_,
    new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_,
    new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_,
    new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_,
    new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_,
    new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_,
    new_n2846_, new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_, new_n2935_,
    new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_,
    new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_,
    new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_,
    new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_,
    new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_,
    new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_,
    new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_,
    new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_,
    new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_,
    new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_,
    new_n2996_, new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_,
    new_n3140_, new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_,
    new_n3146_, new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_,
    new_n3152_, new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_,
    new_n3158_, new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_,
    new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_,
    new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_,
    new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_,
    new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_,
    new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_,
    new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_,
    new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_,
    new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_,
    new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_,
    new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_,
    new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_,
    new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_,
    new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_,
    new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_,
    new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_,
    new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_,
    new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_,
    new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3271_,
    new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_, new_n3277_,
    new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_, new_n3283_,
    new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_,
    new_n3560_, new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_,
    new_n3566_, new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_,
    new_n3572_, new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_,
    new_n3578_, new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_,
    new_n3584_, new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_,
    new_n3590_, new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_,
    new_n3596_, new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_,
    new_n3602_, new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_,
    new_n3608_, new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_,
    new_n3614_, new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_,
    new_n3620_, new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_,
    new_n3626_, new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_,
    new_n3632_, new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_,
    new_n3638_, new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_,
    new_n3644_, new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_,
    new_n3650_, new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_,
    new_n3656_, new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_,
    new_n3662_, new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_,
    new_n3668_, new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_,
    new_n3674_, new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_,
    new_n3680_, new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_,
    new_n3686_, new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_,
    new_n3692_, new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_,
    new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_,
    new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_, new_n3709_,
    new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_, new_n3715_,
    new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_, new_n3721_,
    new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_, new_n3727_,
    new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_, new_n3733_,
    new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_, new_n3739_,
    new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_, new_n3745_,
    new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_, new_n3751_,
    new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_, new_n3757_,
    new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_, new_n3763_,
    new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_, new_n3769_,
    new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_, new_n3775_,
    new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_, new_n3781_,
    new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_, new_n3787_,
    new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_, new_n3793_,
    new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3853_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_,
    new_n4004_, new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_,
    new_n4010_, new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_,
    new_n4016_, new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_,
    new_n4022_, new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_,
    new_n4028_, new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_,
    new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_,
    new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_,
    new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_,
    new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_,
    new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_,
    new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_,
    new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_,
    new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_,
    new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_,
    new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_,
    new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_,
    new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_,
    new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_,
    new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_,
    new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_,
    new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_,
    new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_,
    new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_,
    new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_,
    new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_,
    new_n4538_, new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_,
    new_n4544_, new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_,
    new_n4550_, new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_,
    new_n4556_, new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_,
    new_n4562_, new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_,
    new_n4568_, new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_,
    new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_,
    new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_,
    new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_,
    new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_,
    new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_, new_n4603_,
    new_n4604_, new_n4605_, new_n4606_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_, new_n4627_,
    new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_,
    new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_, new_n4639_,
    new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_, new_n4645_,
    new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_, new_n4651_,
    new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_, new_n4657_,
    new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_, new_n4663_,
    new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_, new_n4669_,
    new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_, new_n4675_,
    new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_, new_n4681_,
    new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_, new_n4687_,
    new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_, new_n4693_,
    new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_, new_n4699_,
    new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_, new_n4705_,
    new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_, new_n4711_,
    new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_, new_n4717_,
    new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_, new_n4723_,
    new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_, new_n4729_,
    new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_, new_n4735_,
    new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_, new_n4741_,
    new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_, new_n4747_,
    new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_, new_n4753_,
    new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_, new_n4759_,
    new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_, new_n4765_,
    new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_, new_n4771_,
    new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_, new_n4777_,
    new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_,
    new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_,
    new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_,
    new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_,
    new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_,
    new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_,
    new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_,
    new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_, new_n5131_,
    new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_, new_n5137_,
    new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_, new_n5143_,
    new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_, new_n5149_,
    new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_, new_n5155_,
    new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_, new_n5161_,
    new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_, new_n5167_,
    new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_, new_n5173_,
    new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_, new_n5179_,
    new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_, new_n5185_,
    new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_, new_n5191_,
    new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_, new_n5197_,
    new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_, new_n5203_,
    new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_, new_n5209_,
    new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_,
    new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_,
    new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_,
    new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_,
    new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_,
    new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_,
    new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_,
    new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_,
    new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_,
    new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_,
    new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_,
    new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_,
    new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_,
    new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_,
    new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_,
    new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_, new_n5635_,
    new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_, new_n5641_,
    new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_, new_n5647_,
    new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_, new_n5653_,
    new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_, new_n5659_,
    new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_, new_n5665_,
    new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_, new_n5671_,
    new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_, new_n5677_,
    new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_, new_n5683_,
    new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_, new_n5689_,
    new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_, new_n5695_,
    new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_, new_n5701_,
    new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_, new_n5707_,
    new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_, new_n5713_,
    new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_, new_n5719_,
    new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_, new_n5725_,
    new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_, new_n5731_,
    new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_, new_n5737_,
    new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_, new_n5743_,
    new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_, new_n5749_,
    new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_, new_n5755_,
    new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_, new_n5761_,
    new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_, new_n5767_,
    new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_, new_n5773_,
    new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_, new_n5821_,
    new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_, new_n5827_,
    new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_, new_n5833_,
    new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_, new_n5839_,
    new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_, new_n5845_,
    new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_, new_n5851_,
    new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_, new_n5857_,
    new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_,
    new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_,
    new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_,
    new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_,
    new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_,
    new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_,
    new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_,
    new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_,
    new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_,
    new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_,
    new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_,
    new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_,
    new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_,
    new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_,
    new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_,
    new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_,
    new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_,
    new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_,
    new_n7377_, new_n7378_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_,
    new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_,
    new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_,
    new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_,
    new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_,
    new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_,
    new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_,
    new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_,
    new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_,
    new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_,
    new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_,
    new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_,
    new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_,
    new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_,
    new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_,
    new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_,
    new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_,
    new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_,
    new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_,
    new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_,
    new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_,
    new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_,
    new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_,
    new_n8440_, new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_,
    new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_,
    new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_,
    new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_,
    new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_,
    new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_,
    new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_,
    new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_,
    new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_,
    new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_,
    new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_,
    new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_,
    new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_,
    new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_,
    new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_,
    new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_,
    new_n8878_, new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_,
    new_n8884_, new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_,
    new_n8890_, new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_,
    new_n8896_, new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_,
    new_n8914_, new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_,
    new_n8920_, new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_,
    new_n8926_, new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_,
    new_n8932_, new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_,
    new_n8938_, new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_,
    new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_,
    new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_,
    new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_,
    new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_,
    new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11073_, new_n11074_, new_n11075_, new_n11076_,
    new_n11077_, new_n11078_, new_n11079_, new_n11080_, new_n11081_,
    new_n11082_, new_n11083_, new_n11084_, new_n11085_, new_n11086_,
    new_n11087_, new_n11088_, new_n11089_, new_n11090_, new_n11091_,
    new_n11092_, new_n11093_, new_n11094_, new_n11095_, new_n11096_,
    new_n11097_, new_n11098_, new_n11099_, new_n11100_, new_n11101_,
    new_n11102_, new_n11103_, new_n11104_, new_n11105_, new_n11106_,
    new_n11107_, new_n11108_, new_n11109_, new_n11110_, new_n11111_,
    new_n11112_, new_n11113_, new_n11114_, new_n11115_, new_n11116_,
    new_n11117_, new_n11118_, new_n11119_, new_n11120_, new_n11121_,
    new_n11122_, new_n11123_, new_n11124_, new_n11125_, new_n11126_,
    new_n11127_, new_n11128_, new_n11129_, new_n11130_, new_n11131_,
    new_n11132_, new_n11133_, new_n11134_, new_n11135_, new_n11136_,
    new_n11137_, new_n11138_, new_n11139_, new_n11140_, new_n11141_,
    new_n11142_, new_n11143_, new_n11144_, new_n11145_, new_n11146_,
    new_n11147_, new_n11148_, new_n11149_, new_n11150_, new_n11151_,
    new_n11152_, new_n11153_, new_n11154_, new_n11155_, new_n11156_,
    new_n11157_, new_n11158_, new_n11159_, new_n11160_, new_n11161_,
    new_n11162_, new_n11163_, new_n11164_, new_n11165_, new_n11166_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11182_, new_n11183_, new_n11184_, new_n11185_, new_n11186_,
    new_n11187_, new_n11188_, new_n11189_, new_n11190_, new_n11191_,
    new_n11192_, new_n11193_, new_n11194_, new_n11195_, new_n11196_,
    new_n11197_, new_n11198_, new_n11199_, new_n11200_, new_n11201_,
    new_n11202_, new_n11203_, new_n11204_, new_n11205_, new_n11206_,
    new_n11207_, new_n11208_, new_n11209_, new_n11210_, new_n11211_,
    new_n11212_, new_n11213_, new_n11214_, new_n11215_, new_n11216_,
    new_n11217_, new_n11218_, new_n11219_, new_n11220_, new_n11221_,
    new_n11222_, new_n11223_, new_n11224_, new_n11225_, new_n11226_,
    new_n11227_, new_n11228_, new_n11229_, new_n11230_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11300_, new_n11301_, new_n11302_,
    new_n11303_, new_n11304_, new_n11305_, new_n11306_, new_n11307_,
    new_n11308_, new_n11309_, new_n11310_, new_n11311_, new_n11312_,
    new_n11313_, new_n11314_, new_n11315_, new_n11316_, new_n11317_,
    new_n11318_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11395_, new_n11396_, new_n11397_,
    new_n11398_, new_n11399_, new_n11400_, new_n11401_, new_n11402_,
    new_n11403_, new_n11404_, new_n11405_, new_n11406_, new_n11407_,
    new_n11408_, new_n11409_, new_n11410_, new_n11411_, new_n11412_,
    new_n11414_, new_n11415_, new_n11416_, new_n11417_, new_n11418_,
    new_n11419_, new_n11420_, new_n11421_, new_n11422_, new_n11423_,
    new_n11424_, new_n11425_, new_n11426_, new_n11427_, new_n11428_,
    new_n11429_, new_n11430_, new_n11431_, new_n11432_, new_n11433_,
    new_n11434_, new_n11435_, new_n11436_, new_n11437_, new_n11438_,
    new_n11439_, new_n11440_, new_n11441_, new_n11442_, new_n11443_,
    new_n11444_, new_n11445_, new_n11446_, new_n11447_, new_n11448_,
    new_n11449_, new_n11450_, new_n11451_, new_n11452_, new_n11453_,
    new_n11454_, new_n11455_, new_n11456_, new_n11457_, new_n11458_,
    new_n11459_, new_n11460_, new_n11461_, new_n11462_, new_n11463_,
    new_n11464_, new_n11465_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11534_,
    new_n11535_, new_n11536_, new_n11537_, new_n11538_, new_n11539_,
    new_n11540_, new_n11541_, new_n11542_, new_n11543_, new_n11544_,
    new_n11545_, new_n11546_, new_n11547_, new_n11548_, new_n11549_,
    new_n11550_, new_n11551_, new_n11552_, new_n11553_, new_n11554_,
    new_n11555_, new_n11556_, new_n11557_, new_n11558_, new_n11559_,
    new_n11560_, new_n11561_, new_n11562_, new_n11563_, new_n11564_,
    new_n11565_, new_n11566_, new_n11567_, new_n11568_, new_n11569_,
    new_n11570_, new_n11571_, new_n11572_, new_n11573_, new_n11574_,
    new_n11575_, new_n11576_, new_n11577_, new_n11578_, new_n11579_,
    new_n11580_, new_n11581_, new_n11582_, new_n11583_, new_n11584_,
    new_n11585_, new_n11586_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11612_, new_n11613_, new_n11614_,
    new_n11615_, new_n11616_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11690_, new_n11691_,
    new_n11692_, new_n11693_, new_n11694_, new_n11695_, new_n11696_,
    new_n11697_, new_n11698_, new_n11699_, new_n11700_, new_n11701_,
    new_n11702_, new_n11703_, new_n11704_, new_n11705_, new_n11706_,
    new_n11707_, new_n11708_, new_n11709_, new_n11710_, new_n11711_,
    new_n11712_, new_n11713_, new_n11714_, new_n11715_, new_n11716_,
    new_n11717_, new_n11718_, new_n11719_, new_n11720_, new_n11721_,
    new_n11722_, new_n11723_, new_n11724_, new_n11725_, new_n11726_,
    new_n11727_, new_n11728_, new_n11729_, new_n11730_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11761_,
    new_n11762_, new_n11763_, new_n11764_, new_n11765_, new_n11766_,
    new_n11767_, new_n11768_, new_n11769_, new_n11770_, new_n11771_,
    new_n11772_, new_n11773_, new_n11774_, new_n11775_, new_n11776_,
    new_n11777_, new_n11778_, new_n11779_, new_n11780_, new_n11781_,
    new_n11782_, new_n11783_, new_n11784_, new_n11785_, new_n11786_,
    new_n11787_, new_n11788_, new_n11789_, new_n11790_, new_n11791_,
    new_n11792_, new_n11793_, new_n11794_, new_n11795_, new_n11796_,
    new_n11797_, new_n11798_, new_n11799_, new_n11800_, new_n11801_,
    new_n11802_, new_n11803_, new_n11804_, new_n11805_, new_n11806_,
    new_n11807_, new_n11808_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11874_, new_n11875_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11906_, new_n11907_, new_n11908_,
    new_n11909_, new_n11910_, new_n11911_, new_n11912_, new_n11913_,
    new_n11914_, new_n11915_, new_n11916_, new_n11917_, new_n11918_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12484_, new_n12485_, new_n12486_, new_n12487_, new_n12488_,
    new_n12489_, new_n12490_, new_n12491_, new_n12492_, new_n12493_,
    new_n12494_, new_n12495_, new_n12496_, new_n12497_, new_n12498_,
    new_n12499_, new_n12500_, new_n12501_, new_n12502_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14445_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14456_,
    new_n14457_, new_n14458_, new_n14459_, new_n14460_, new_n14461_,
    new_n14462_, new_n14463_, new_n14464_, new_n14465_, new_n14466_,
    new_n14467_, new_n14468_, new_n14469_, new_n14470_, new_n14471_,
    new_n14472_, new_n14473_, new_n14474_, new_n14475_, new_n14476_,
    new_n14477_, new_n14478_, new_n14479_, new_n14480_, new_n14481_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14487_, new_n14488_, new_n14489_, new_n14490_, new_n14491_,
    new_n14492_, new_n14493_, new_n14494_, new_n14495_, new_n14496_,
    new_n14497_, new_n14498_, new_n14499_, new_n14500_, new_n14501_,
    new_n14502_, new_n14503_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14522_, new_n14523_, new_n14524_, new_n14525_, new_n14526_,
    new_n14527_, new_n14528_, new_n14529_, new_n14530_, new_n14531_,
    new_n14532_, new_n14533_, new_n14534_, new_n14535_, new_n14536_,
    new_n14537_, new_n14538_, new_n14539_, new_n14540_, new_n14541_,
    new_n14542_, new_n14543_, new_n14544_, new_n14545_, new_n14546_,
    new_n14547_, new_n14548_, new_n14549_, new_n14550_, new_n14551_,
    new_n14552_, new_n14553_, new_n14554_, new_n14555_, new_n14556_,
    new_n14557_, new_n14558_, new_n14559_, new_n14560_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14575_, new_n14576_,
    new_n14577_, new_n14578_, new_n14579_, new_n14580_, new_n14581_,
    new_n14582_, new_n14583_, new_n14584_, new_n14585_, new_n14586_,
    new_n14587_, new_n14588_, new_n14589_, new_n14590_, new_n14591_,
    new_n14592_, new_n14593_, new_n14594_, new_n14595_, new_n14596_,
    new_n14597_, new_n14598_, new_n14599_, new_n14600_, new_n14601_,
    new_n14602_, new_n14603_, new_n14604_, new_n14605_, new_n14606_,
    new_n14607_, new_n14608_, new_n14609_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14620_, new_n14621_,
    new_n14622_, new_n14623_, new_n14624_, new_n14625_, new_n14626_,
    new_n14627_, new_n14628_, new_n14629_, new_n14630_, new_n14631_,
    new_n14632_, new_n14633_, new_n14634_, new_n14635_, new_n14636_,
    new_n14637_, new_n14638_, new_n14639_, new_n14640_, new_n14641_,
    new_n14642_, new_n14643_, new_n14644_, new_n14645_, new_n14646_,
    new_n14647_, new_n14648_, new_n14649_, new_n14650_, new_n14651_,
    new_n14652_, new_n14653_, new_n14654_, new_n14655_, new_n14656_,
    new_n14657_, new_n14658_, new_n14659_, new_n14660_, new_n14661_,
    new_n14662_, new_n14663_, new_n14664_, new_n14665_, new_n14666_,
    new_n14667_, new_n14668_, new_n14669_, new_n14670_, new_n14671_,
    new_n14672_, new_n14673_, new_n14674_, new_n14675_, new_n14676_,
    new_n14677_, new_n14678_, new_n14679_, new_n14680_, new_n14681_,
    new_n14682_, new_n14683_, new_n14684_, new_n14685_, new_n14686_,
    new_n14687_, new_n14688_, new_n14689_, new_n14690_, new_n14691_,
    new_n14692_, new_n14693_, new_n14694_, new_n14695_, new_n14696_,
    new_n14697_, new_n14698_, new_n14699_, new_n14700_, new_n14701_,
    new_n14702_, new_n14703_, new_n14704_, new_n14705_, new_n14706_,
    new_n14707_, new_n14708_, new_n14709_, new_n14710_, new_n14711_,
    new_n14712_, new_n14713_, new_n14714_, new_n14715_, new_n14716_,
    new_n14717_, new_n14718_, new_n14719_, new_n14720_, new_n14721_,
    new_n14722_, new_n14723_, new_n14724_, new_n14725_, new_n14726_,
    new_n14727_, new_n14728_, new_n14729_, new_n14730_, new_n14731_,
    new_n14732_, new_n14733_, new_n14734_, new_n14735_, new_n14736_,
    new_n14737_, new_n14738_, new_n14739_, new_n14740_, new_n14741_,
    new_n14742_, new_n14743_, new_n14744_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14781_,
    new_n14782_, new_n14783_, new_n14784_, new_n14785_, new_n14786_,
    new_n14787_, new_n14788_, new_n14789_, new_n14790_, new_n14791_,
    new_n14792_, new_n14793_, new_n14794_, new_n14795_, new_n14796_,
    new_n14797_, new_n14798_, new_n14799_, new_n14800_, new_n14801_,
    new_n14802_, new_n14803_, new_n14804_, new_n14805_, new_n14806_,
    new_n14807_, new_n14808_, new_n14809_, new_n14810_, new_n14811_,
    new_n14812_, new_n14813_, new_n14814_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14958_, new_n14959_, new_n14960_, new_n14961_,
    new_n14962_, new_n14963_, new_n14964_, new_n14965_, new_n14966_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14976_,
    new_n14977_, new_n14978_, new_n14979_, new_n14980_, new_n14981_,
    new_n14982_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15113_, new_n15114_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15127_, new_n15128_, new_n15129_, new_n15130_, new_n15131_,
    new_n15132_, new_n15133_, new_n15134_, new_n15135_, new_n15136_,
    new_n15137_, new_n15138_, new_n15139_, new_n15140_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15179_, new_n15180_, new_n15181_,
    new_n15182_, new_n15183_, new_n15184_, new_n15185_, new_n15186_,
    new_n15187_, new_n15188_, new_n15189_, new_n15190_, new_n15191_,
    new_n15192_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15206_,
    new_n15207_, new_n15208_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15213_, new_n15214_, new_n15215_, new_n15216_,
    new_n15217_, new_n15218_, new_n15219_, new_n15220_, new_n15221_,
    new_n15222_, new_n15223_, new_n15224_, new_n15225_, new_n15226_,
    new_n15227_, new_n15228_, new_n15229_, new_n15230_, new_n15231_,
    new_n15232_, new_n15233_, new_n15234_, new_n15235_, new_n15236_,
    new_n15237_, new_n15238_, new_n15239_, new_n15240_, new_n15241_,
    new_n15242_, new_n15243_, new_n15244_, new_n15245_, new_n15246_,
    new_n15247_, new_n15248_, new_n15249_, new_n15250_, new_n15251_,
    new_n15252_, new_n15253_, new_n15254_, new_n15255_, new_n15256_,
    new_n15257_, new_n15258_, new_n15259_, new_n15260_, new_n15261_,
    new_n15262_, new_n15263_, new_n15264_, new_n15265_, new_n15266_,
    new_n15267_, new_n15268_, new_n15269_, new_n15270_, new_n15271_,
    new_n15272_, new_n15273_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15280_, new_n15281_,
    new_n15282_, new_n15283_, new_n15284_, new_n15285_, new_n15286_,
    new_n15287_, new_n15288_, new_n15289_, new_n15290_, new_n15291_,
    new_n15292_, new_n15293_, new_n15294_, new_n15295_, new_n15296_,
    new_n15297_, new_n15298_, new_n15299_, new_n15300_, new_n15301_,
    new_n15302_, new_n15303_, new_n15304_, new_n15305_, new_n15306_,
    new_n15307_, new_n15308_, new_n15309_, new_n15310_, new_n15311_,
    new_n15312_, new_n15313_, new_n15314_, new_n15315_, new_n15316_,
    new_n15317_, new_n15318_, new_n15319_, new_n15320_, new_n15321_,
    new_n15322_, new_n15323_, new_n15324_, new_n15325_, new_n15326_,
    new_n15327_, new_n15328_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15434_, new_n15435_, new_n15436_,
    new_n15437_, new_n15438_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15470_, new_n15471_,
    new_n15472_, new_n15473_, new_n15474_, new_n15475_, new_n15476_,
    new_n15477_, new_n15478_, new_n15479_, new_n15480_, new_n15481_,
    new_n15482_, new_n15483_, new_n15484_, new_n15485_, new_n15486_,
    new_n15487_, new_n15488_, new_n15489_, new_n15490_, new_n15491_,
    new_n15492_, new_n15493_, new_n15494_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15544_, new_n15545_, new_n15546_,
    new_n15547_, new_n15548_, new_n15549_, new_n15550_, new_n15551_,
    new_n15552_, new_n15553_, new_n15554_, new_n15555_, new_n15556_,
    new_n15557_, new_n15558_, new_n15559_, new_n15560_, new_n15561_,
    new_n15562_, new_n15563_, new_n15564_, new_n15565_, new_n15566_,
    new_n15567_, new_n15568_, new_n15569_, new_n15570_, new_n15571_,
    new_n15572_, new_n15573_, new_n15574_, new_n15575_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15580_, new_n15581_,
    new_n15582_, new_n15583_, new_n15584_, new_n15585_, new_n15586_,
    new_n15587_, new_n15588_, new_n15589_, new_n15590_, new_n15591_,
    new_n15592_, new_n15593_, new_n15594_, new_n15595_, new_n15596_,
    new_n15597_, new_n15598_, new_n15599_, new_n15600_, new_n15601_,
    new_n15602_, new_n15603_, new_n15604_, new_n15605_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15611_,
    new_n15612_, new_n15613_, new_n15614_, new_n15615_, new_n15616_,
    new_n15617_, new_n15618_, new_n15619_, new_n15620_, new_n15621_,
    new_n15622_, new_n15623_, new_n15624_, new_n15625_, new_n15626_,
    new_n15627_, new_n15628_, new_n15629_, new_n15630_, new_n15631_,
    new_n15632_, new_n15633_, new_n15634_, new_n15635_, new_n15636_,
    new_n15637_, new_n15638_, new_n15639_, new_n15640_, new_n15641_,
    new_n15642_, new_n15643_, new_n15644_, new_n15645_, new_n15646_,
    new_n15647_, new_n15648_, new_n15649_, new_n15650_, new_n15651_,
    new_n15652_, new_n15653_, new_n15654_, new_n15655_, new_n15656_,
    new_n15657_, new_n15658_, new_n15659_, new_n15660_, new_n15661_,
    new_n15662_, new_n15663_, new_n15664_, new_n15665_, new_n15666_,
    new_n15667_, new_n15668_, new_n15669_, new_n15670_, new_n15671_,
    new_n15672_, new_n15673_, new_n15674_, new_n15675_, new_n15676_,
    new_n15677_, new_n15678_, new_n15679_, new_n15680_, new_n15681_,
    new_n15682_, new_n15683_, new_n15684_, new_n15685_, new_n15686_,
    new_n15687_, new_n15688_, new_n15689_, new_n15690_, new_n15691_,
    new_n15692_, new_n15693_, new_n15694_, new_n15695_, new_n15696_,
    new_n15697_, new_n15698_, new_n15699_, new_n15700_, new_n15701_,
    new_n15702_, new_n15703_, new_n15704_, new_n15705_, new_n15706_,
    new_n15707_, new_n15708_, new_n15709_, new_n15710_, new_n15711_,
    new_n15712_, new_n15713_, new_n15714_, new_n15715_, new_n15716_,
    new_n15717_, new_n15718_, new_n15719_, new_n15720_, new_n15721_,
    new_n15722_, new_n15723_, new_n15724_, new_n15725_, new_n15726_,
    new_n15727_, new_n15728_, new_n15729_, new_n15730_, new_n15731_,
    new_n15732_, new_n15733_, new_n15734_, new_n15735_, new_n15736_,
    new_n15737_, new_n15738_, new_n15739_, new_n15740_, new_n15741_,
    new_n15742_, new_n15743_, new_n15744_, new_n15745_, new_n15746_,
    new_n15747_, new_n15748_, new_n15749_, new_n15750_, new_n15751_,
    new_n15752_, new_n15753_, new_n15754_, new_n15755_, new_n15756_,
    new_n15757_, new_n15758_, new_n15759_, new_n15760_, new_n15761_,
    new_n15762_, new_n15763_, new_n15764_, new_n15765_, new_n15766_,
    new_n15767_, new_n15768_, new_n15769_, new_n15770_, new_n15771_,
    new_n15772_, new_n15773_, new_n15774_, new_n15775_, new_n15776_,
    new_n15777_, new_n15778_, new_n15779_, new_n15780_, new_n15781_,
    new_n15782_, new_n15783_, new_n15784_, new_n15785_, new_n15786_,
    new_n15787_, new_n15788_, new_n15789_, new_n15790_, new_n15791_,
    new_n15792_, new_n15793_, new_n15794_, new_n15795_, new_n15796_,
    new_n15797_, new_n15798_, new_n15799_, new_n15800_, new_n15801_,
    new_n15802_, new_n15803_, new_n15804_, new_n15805_, new_n15806_,
    new_n15807_, new_n15808_, new_n15809_, new_n15810_, new_n15811_,
    new_n15812_, new_n15813_, new_n15814_, new_n15815_, new_n15816_,
    new_n15817_, new_n15818_, new_n15819_, new_n15820_, new_n15821_,
    new_n15822_, new_n15823_, new_n15824_, new_n15825_, new_n15826_,
    new_n15827_, new_n15828_, new_n15829_, new_n15830_, new_n15831_,
    new_n15832_, new_n15833_, new_n15834_, new_n15835_, new_n15836_,
    new_n15837_, new_n15838_, new_n15839_, new_n15840_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15850_, new_n15851_,
    new_n15852_, new_n15853_, new_n15854_, new_n15855_, new_n15856_,
    new_n15857_, new_n15858_, new_n15859_, new_n15860_, new_n15861_,
    new_n15862_, new_n15863_, new_n15864_, new_n15865_, new_n15866_,
    new_n15867_, new_n15868_, new_n15869_, new_n15870_, new_n15871_,
    new_n15872_, new_n15873_, new_n15874_, new_n15875_, new_n15876_,
    new_n15877_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15889_, new_n15890_, new_n15891_,
    new_n15892_, new_n15893_, new_n15894_, new_n15895_, new_n15896_,
    new_n15897_, new_n15898_, new_n15899_, new_n15900_, new_n15901_,
    new_n15902_, new_n15903_, new_n15904_, new_n15905_, new_n15906_,
    new_n15907_, new_n15908_, new_n15909_, new_n15910_, new_n15911_,
    new_n15912_, new_n15913_, new_n15914_, new_n15915_, new_n15916_,
    new_n15917_, new_n15918_, new_n15919_, new_n15920_, new_n15921_,
    new_n15922_, new_n15923_, new_n15924_, new_n15925_, new_n15926_,
    new_n15927_, new_n15928_, new_n15929_, new_n15930_, new_n15931_,
    new_n15932_, new_n15933_, new_n15934_, new_n15935_, new_n15936_,
    new_n15937_, new_n15938_, new_n15939_, new_n15940_, new_n15941_,
    new_n15942_, new_n15943_, new_n15944_, new_n15945_, new_n15946_,
    new_n15947_, new_n15948_, new_n15949_, new_n15950_, new_n15951_,
    new_n15952_, new_n15953_, new_n15954_, new_n15955_, new_n15956_,
    new_n15957_, new_n15958_, new_n15959_, new_n15960_, new_n15961_,
    new_n15962_, new_n15963_, new_n15964_, new_n15965_, new_n15966_,
    new_n15967_, new_n15968_, new_n15969_, new_n15970_, new_n15971_,
    new_n15972_, new_n15973_, new_n15974_, new_n15975_, new_n15976_,
    new_n15977_, new_n15978_, new_n15979_, new_n15980_, new_n15981_,
    new_n15982_, new_n15983_, new_n15984_, new_n15985_, new_n15986_,
    new_n15987_, new_n15988_, new_n15989_, new_n15990_, new_n15991_,
    new_n15992_, new_n15993_, new_n15994_, new_n15995_, new_n15996_,
    new_n15997_, new_n15998_, new_n15999_, new_n16000_, new_n16001_,
    new_n16002_, new_n16003_, new_n16004_, new_n16005_, new_n16006_,
    new_n16007_, new_n16008_, new_n16009_, new_n16010_, new_n16011_,
    new_n16012_, new_n16013_, new_n16014_, new_n16015_, new_n16016_,
    new_n16017_, new_n16018_, new_n16019_, new_n16020_, new_n16021_,
    new_n16022_, new_n16023_, new_n16024_, new_n16025_, new_n16026_,
    new_n16027_, new_n16028_, new_n16029_, new_n16030_, new_n16031_,
    new_n16032_, new_n16033_, new_n16034_, new_n16035_, new_n16036_,
    new_n16037_, new_n16038_, new_n16039_, new_n16040_, new_n16041_,
    new_n16042_, new_n16043_, new_n16044_, new_n16045_, new_n16046_,
    new_n16047_, new_n16048_, new_n16049_, new_n16050_, new_n16051_,
    new_n16052_, new_n16053_, new_n16054_, new_n16055_, new_n16056_,
    new_n16057_, new_n16058_, new_n16059_, new_n16060_, new_n16061_,
    new_n16062_, new_n16063_, new_n16064_, new_n16065_, new_n16066_,
    new_n16067_, new_n16068_, new_n16069_, new_n16070_, new_n16071_,
    new_n16072_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_, new_n16078_, new_n16079_, new_n16080_, new_n16081_,
    new_n16082_, new_n16083_, new_n16084_, new_n16085_, new_n16086_,
    new_n16087_, new_n16088_, new_n16089_, new_n16090_, new_n16091_,
    new_n16092_, new_n16093_, new_n16094_, new_n16095_, new_n16096_,
    new_n16097_, new_n16098_, new_n16099_, new_n16100_, new_n16101_,
    new_n16102_, new_n16103_, new_n16104_, new_n16105_, new_n16106_,
    new_n16107_, new_n16108_, new_n16109_, new_n16110_, new_n16111_,
    new_n16112_, new_n16113_, new_n16114_, new_n16115_, new_n16116_,
    new_n16117_, new_n16118_, new_n16119_, new_n16120_, new_n16121_,
    new_n16122_, new_n16123_, new_n16124_, new_n16125_, new_n16126_,
    new_n16127_, new_n16128_, new_n16129_, new_n16130_, new_n16131_,
    new_n16132_, new_n16133_, new_n16134_, new_n16135_, new_n16136_,
    new_n16137_, new_n16138_, new_n16139_, new_n16140_, new_n16141_,
    new_n16142_, new_n16143_, new_n16144_, new_n16145_, new_n16146_,
    new_n16147_, new_n16148_, new_n16149_, new_n16150_, new_n16151_,
    new_n16152_, new_n16153_, new_n16154_, new_n16155_, new_n16156_,
    new_n16157_, new_n16158_, new_n16159_, new_n16160_, new_n16161_,
    new_n16162_, new_n16163_, new_n16164_, new_n16165_, new_n16166_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16274_, new_n16275_, new_n16276_,
    new_n16277_, new_n16278_, new_n16279_, new_n16280_, new_n16281_,
    new_n16282_, new_n16283_, new_n16284_, new_n16285_, new_n16286_,
    new_n16287_, new_n16288_, new_n16289_, new_n16290_, new_n16291_,
    new_n16292_, new_n16293_, new_n16294_, new_n16295_, new_n16296_,
    new_n16297_, new_n16298_, new_n16299_, new_n16300_, new_n16301_,
    new_n16302_, new_n16303_, new_n16304_, new_n16305_, new_n16306_,
    new_n16307_, new_n16308_, new_n16309_, new_n16310_, new_n16311_,
    new_n16312_, new_n16313_, new_n16314_, new_n16315_, new_n16316_,
    new_n16317_, new_n16318_, new_n16319_, new_n16320_, new_n16321_,
    new_n16322_, new_n16323_, new_n16324_, new_n16325_, new_n16326_,
    new_n16327_, new_n16328_, new_n16329_, new_n16330_, new_n16331_,
    new_n16332_, new_n16333_, new_n16334_, new_n16335_, new_n16336_,
    new_n16337_, new_n16338_, new_n16339_, new_n16340_, new_n16341_,
    new_n16342_, new_n16343_, new_n16344_, new_n16345_, new_n16346_,
    new_n16347_, new_n16348_, new_n16349_, new_n16350_, new_n16351_,
    new_n16352_, new_n16353_, new_n16354_, new_n16355_, new_n16356_,
    new_n16357_, new_n16358_, new_n16359_, new_n16360_, new_n16361_,
    new_n16362_, new_n16363_, new_n16364_, new_n16365_, new_n16366_,
    new_n16367_, new_n16368_, new_n16369_, new_n16370_, new_n16371_,
    new_n16372_, new_n16373_, new_n16374_, new_n16375_, new_n16376_,
    new_n16377_, new_n16378_, new_n16379_, new_n16380_, new_n16381_,
    new_n16382_, new_n16383_, new_n16384_, new_n16385_, new_n16386_,
    new_n16387_, new_n16388_, new_n16389_, new_n16390_, new_n16391_,
    new_n16392_, new_n16393_, new_n16394_, new_n16395_, new_n16396_,
    new_n16397_, new_n16398_, new_n16399_, new_n16400_, new_n16401_,
    new_n16402_, new_n16403_, new_n16404_, new_n16405_, new_n16406_,
    new_n16407_, new_n16408_, new_n16409_, new_n16410_, new_n16411_,
    new_n16412_, new_n16413_, new_n16414_, new_n16415_, new_n16416_,
    new_n16417_, new_n16418_, new_n16419_, new_n16420_, new_n16421_,
    new_n16422_, new_n16423_, new_n16424_, new_n16425_, new_n16426_,
    new_n16427_, new_n16428_, new_n16429_, new_n16430_, new_n16431_,
    new_n16432_, new_n16433_, new_n16434_, new_n16435_, new_n16436_,
    new_n16437_, new_n16438_, new_n16439_, new_n16440_, new_n16441_,
    new_n16442_, new_n16443_, new_n16444_, new_n16445_, new_n16446_,
    new_n16447_, new_n16448_, new_n16449_, new_n16450_, new_n16451_,
    new_n16452_, new_n16453_, new_n16454_, new_n16455_, new_n16456_,
    new_n16457_, new_n16458_, new_n16459_, new_n16460_, new_n16461_,
    new_n16462_, new_n16463_, new_n16464_, new_n16465_, new_n16466_,
    new_n16467_, new_n16468_, new_n16469_, new_n16470_, new_n16471_,
    new_n16472_, new_n16473_, new_n16474_, new_n16475_, new_n16476_,
    new_n16477_, new_n16478_, new_n16479_, new_n16480_, new_n16481_,
    new_n16482_, new_n16483_, new_n16484_, new_n16485_, new_n16486_,
    new_n16487_, new_n16488_, new_n16489_, new_n16490_, new_n16491_,
    new_n16492_, new_n16493_, new_n16494_, new_n16495_, new_n16496_,
    new_n16497_, new_n16498_, new_n16499_, new_n16500_, new_n16501_,
    new_n16502_, new_n16503_, new_n16504_, new_n16505_, new_n16506_,
    new_n16507_, new_n16508_, new_n16509_, new_n16510_, new_n16511_,
    new_n16512_, new_n16513_, new_n16514_, new_n16515_, new_n16516_,
    new_n16517_, new_n16518_, new_n16519_, new_n16520_, new_n16521_,
    new_n16522_, new_n16523_, new_n16524_, new_n16525_, new_n16526_,
    new_n16527_, new_n16528_, new_n16529_, new_n16530_, new_n16531_,
    new_n16532_, new_n16533_, new_n16534_, new_n16535_, new_n16536_,
    new_n16537_, new_n16538_, new_n16539_, new_n16540_, new_n16541_,
    new_n16542_, new_n16543_, new_n16544_, new_n16545_, new_n16546_,
    new_n16547_, new_n16548_, new_n16549_, new_n16550_, new_n16551_,
    new_n16552_, new_n16553_, new_n16554_, new_n16555_, new_n16556_,
    new_n16557_, new_n16558_, new_n16559_, new_n16560_, new_n16561_,
    new_n16562_, new_n16563_, new_n16564_, new_n16565_, new_n16566_,
    new_n16567_, new_n16568_, new_n16569_, new_n16570_, new_n16571_,
    new_n16572_, new_n16573_, new_n16574_, new_n16575_, new_n16576_,
    new_n16577_, new_n16578_, new_n16579_, new_n16580_, new_n16581_,
    new_n16582_, new_n16583_, new_n16584_, new_n16585_, new_n16586_,
    new_n16587_, new_n16588_, new_n16589_, new_n16590_, new_n16591_,
    new_n16592_, new_n16593_, new_n16594_, new_n16595_, new_n16596_,
    new_n16597_, new_n16598_, new_n16599_, new_n16600_, new_n16601_,
    new_n16602_, new_n16603_, new_n16604_, new_n16605_, new_n16606_,
    new_n16607_, new_n16608_, new_n16609_, new_n16610_, new_n16611_,
    new_n16612_, new_n16613_, new_n16614_, new_n16615_, new_n16616_,
    new_n16617_, new_n16618_, new_n16619_, new_n16620_, new_n16621_,
    new_n16622_, new_n16623_, new_n16624_, new_n16625_, new_n16626_,
    new_n16627_, new_n16628_, new_n16629_, new_n16630_, new_n16631_,
    new_n16632_, new_n16633_, new_n16634_, new_n16635_, new_n16636_,
    new_n16637_, new_n16638_, new_n16639_, new_n16640_, new_n16641_,
    new_n16642_, new_n16643_, new_n16644_, new_n16645_, new_n16646_,
    new_n16647_, new_n16648_, new_n16649_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16727_, new_n16728_, new_n16729_, new_n16730_, new_n16731_,
    new_n16732_, new_n16733_, new_n16734_, new_n16735_, new_n16736_,
    new_n16737_, new_n16738_, new_n16739_, new_n16740_, new_n16741_,
    new_n16742_, new_n16743_, new_n16744_, new_n16745_, new_n16746_,
    new_n16747_, new_n16748_, new_n16749_, new_n16750_, new_n16751_,
    new_n16752_, new_n16753_, new_n16754_, new_n16755_, new_n16756_,
    new_n16757_, new_n16758_, new_n16759_, new_n16760_, new_n16761_,
    new_n16762_, new_n16763_, new_n16764_, new_n16765_, new_n16766_,
    new_n16767_, new_n16768_, new_n16769_, new_n16770_, new_n16771_,
    new_n16772_, new_n16773_, new_n16774_, new_n16775_, new_n16776_,
    new_n16777_, new_n16778_, new_n16779_, new_n16780_, new_n16781_,
    new_n16782_, new_n16783_, new_n16784_, new_n16785_, new_n16786_,
    new_n16787_, new_n16788_, new_n16789_, new_n16790_, new_n16791_,
    new_n16792_, new_n16793_, new_n16794_, new_n16795_, new_n16796_,
    new_n16797_, new_n16798_, new_n16799_, new_n16800_, new_n16801_,
    new_n16802_, new_n16803_, new_n16804_, new_n16805_, new_n16806_,
    new_n16807_, new_n16808_, new_n16809_, new_n16810_, new_n16811_,
    new_n16812_, new_n16813_, new_n16814_, new_n16815_, new_n16816_,
    new_n16817_, new_n16818_, new_n16819_, new_n16820_, new_n16821_,
    new_n16822_, new_n16823_, new_n16824_, new_n16825_, new_n16826_,
    new_n16827_, new_n16828_, new_n16829_, new_n16830_, new_n16831_,
    new_n16832_, new_n16833_, new_n16834_, new_n16835_, new_n16836_,
    new_n16837_, new_n16838_, new_n16839_, new_n16840_, new_n16841_,
    new_n16842_, new_n16843_, new_n16844_, new_n16845_, new_n16846_,
    new_n16847_, new_n16848_, new_n16849_, new_n16850_, new_n16851_,
    new_n16852_, new_n16853_, new_n16854_, new_n16855_, new_n16856_,
    new_n16857_, new_n16858_, new_n16859_, new_n16860_, new_n16861_,
    new_n16862_, new_n16864_, new_n16865_, new_n16866_, new_n16867_,
    new_n16868_, new_n16869_, new_n16870_, new_n16871_, new_n16872_,
    new_n16873_, new_n16874_, new_n16875_, new_n16876_, new_n16877_,
    new_n16878_, new_n16879_, new_n16880_, new_n16881_, new_n16882_,
    new_n16883_, new_n16884_, new_n16885_, new_n16886_, new_n16887_,
    new_n16888_, new_n16889_, new_n16890_, new_n16891_, new_n16892_,
    new_n16893_, new_n16894_, new_n16895_, new_n16896_, new_n16897_,
    new_n16898_, new_n16899_, new_n16900_, new_n16901_, new_n16902_,
    new_n16903_, new_n16904_, new_n16905_, new_n16906_, new_n16907_,
    new_n16908_, new_n16909_, new_n16910_, new_n16911_, new_n16912_,
    new_n16913_, new_n16914_, new_n16915_, new_n16916_, new_n16917_,
    new_n16918_, new_n16919_, new_n16920_, new_n16921_, new_n16922_,
    new_n16923_, new_n16924_, new_n16925_, new_n16926_, new_n16927_,
    new_n16928_, new_n16929_, new_n16930_, new_n16931_, new_n16932_,
    new_n16933_, new_n16934_, new_n16935_, new_n16936_, new_n16937_,
    new_n16938_, new_n16939_, new_n16940_, new_n16941_, new_n16942_,
    new_n16943_, new_n16944_, new_n16945_, new_n16946_, new_n16947_,
    new_n16948_, new_n16949_, new_n16950_, new_n16951_, new_n16952_,
    new_n16953_, new_n16954_, new_n16955_, new_n16956_, new_n16957_,
    new_n16958_, new_n16959_, new_n16960_, new_n16961_, new_n16962_,
    new_n16963_, new_n16964_, new_n16965_, new_n16966_, new_n16967_,
    new_n16968_, new_n16969_, new_n16970_, new_n16971_, new_n16972_,
    new_n16973_, new_n16974_, new_n16975_, new_n16976_, new_n16977_,
    new_n16978_, new_n16979_, new_n16980_, new_n16981_, new_n16982_,
    new_n16984_, new_n16985_, new_n16986_, new_n16987_, new_n16988_,
    new_n16989_, new_n16990_, new_n16991_, new_n16992_, new_n16993_,
    new_n16994_, new_n16995_, new_n16996_, new_n16997_, new_n16998_,
    new_n16999_, new_n17000_, new_n17001_, new_n17002_, new_n17003_,
    new_n17004_, new_n17005_, new_n17006_, new_n17007_, new_n17008_,
    new_n17009_, new_n17010_, new_n17011_, new_n17012_, new_n17013_,
    new_n17014_, new_n17015_, new_n17016_, new_n17017_, new_n17018_,
    new_n17019_, new_n17020_, new_n17021_, new_n17022_, new_n17023_,
    new_n17024_, new_n17025_, new_n17026_, new_n17027_, new_n17028_,
    new_n17029_, new_n17030_, new_n17031_, new_n17032_, new_n17033_,
    new_n17034_, new_n17035_, new_n17036_, new_n17037_, new_n17038_,
    new_n17039_, new_n17040_, new_n17041_, new_n17042_, new_n17043_,
    new_n17044_, new_n17045_, new_n17046_, new_n17047_, new_n17048_,
    new_n17049_, new_n17050_, new_n17051_, new_n17052_, new_n17053_,
    new_n17054_, new_n17055_, new_n17056_, new_n17057_, new_n17058_,
    new_n17059_, new_n17060_, new_n17061_, new_n17062_, new_n17063_,
    new_n17064_, new_n17065_, new_n17066_, new_n17067_, new_n17068_,
    new_n17069_, new_n17070_, new_n17071_, new_n17072_, new_n17073_,
    new_n17074_, new_n17075_, new_n17076_, new_n17077_, new_n17078_,
    new_n17079_, new_n17080_, new_n17081_, new_n17082_, new_n17083_,
    new_n17084_, new_n17085_, new_n17086_, new_n17087_, new_n17088_,
    new_n17089_, new_n17090_, new_n17091_, new_n17092_, new_n17093_,
    new_n17094_, new_n17095_, new_n17096_, new_n17097_, new_n17098_,
    new_n17099_, new_n17100_, new_n17101_, new_n17102_, new_n17103_,
    new_n17104_, new_n17105_, new_n17106_, new_n17107_, new_n17108_,
    new_n17109_, new_n17110_, new_n17111_, new_n17112_, new_n17113_,
    new_n17114_, new_n17115_, new_n17116_, new_n17117_, new_n17118_,
    new_n17119_, new_n17120_, new_n17121_, new_n17122_, new_n17123_,
    new_n17124_, new_n17125_, new_n17126_, new_n17127_, new_n17128_,
    new_n17129_, new_n17130_, new_n17131_, new_n17132_, new_n17133_,
    new_n17134_, new_n17135_, new_n17136_, new_n17137_, new_n17138_,
    new_n17139_, new_n17140_, new_n17141_, new_n17142_, new_n17143_,
    new_n17144_, new_n17145_, new_n17146_, new_n17147_, new_n17148_,
    new_n17149_, new_n17150_, new_n17151_, new_n17152_, new_n17153_,
    new_n17154_, new_n17155_, new_n17156_, new_n17157_, new_n17158_,
    new_n17159_, new_n17160_, new_n17161_, new_n17162_, new_n17163_,
    new_n17164_, new_n17165_, new_n17166_, new_n17167_, new_n17168_,
    new_n17169_, new_n17170_, new_n17171_, new_n17172_, new_n17173_,
    new_n17174_, new_n17175_, new_n17176_, new_n17177_, new_n17178_,
    new_n17179_, new_n17180_, new_n17181_, new_n17182_, new_n17183_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17229_, new_n17230_, new_n17231_, new_n17232_, new_n17233_,
    new_n17234_, new_n17235_, new_n17236_, new_n17237_, new_n17238_,
    new_n17239_, new_n17240_, new_n17241_, new_n17242_, new_n17243_,
    new_n17244_, new_n17245_, new_n17246_, new_n17247_, new_n17248_,
    new_n17249_, new_n17250_, new_n17251_, new_n17252_, new_n17253_,
    new_n17254_, new_n17255_, new_n17256_, new_n17257_, new_n17258_,
    new_n17259_, new_n17260_, new_n17261_, new_n17262_, new_n17263_,
    new_n17264_, new_n17265_, new_n17266_, new_n17267_, new_n17268_,
    new_n17269_, new_n17270_, new_n17271_, new_n17272_, new_n17273_,
    new_n17274_, new_n17275_, new_n17276_, new_n17277_, new_n17278_,
    new_n17279_, new_n17280_, new_n17281_, new_n17282_, new_n17283_,
    new_n17284_, new_n17285_, new_n17286_, new_n17287_, new_n17288_,
    new_n17289_, new_n17290_, new_n17291_, new_n17292_, new_n17293_,
    new_n17294_, new_n17295_, new_n17296_, new_n17297_, new_n17298_,
    new_n17299_, new_n17300_, new_n17301_, new_n17302_, new_n17303_,
    new_n17304_, new_n17305_, new_n17306_, new_n17307_, new_n17308_,
    new_n17309_, new_n17310_, new_n17311_, new_n17312_, new_n17313_,
    new_n17314_, new_n17315_, new_n17316_, new_n17317_, new_n17318_,
    new_n17319_, new_n17320_, new_n17321_, new_n17322_, new_n17323_,
    new_n17324_, new_n17325_, new_n17326_, new_n17327_, new_n17328_,
    new_n17329_, new_n17330_, new_n17331_, new_n17332_, new_n17333_,
    new_n17334_, new_n17335_, new_n17336_, new_n17337_, new_n17338_,
    new_n17339_, new_n17340_, new_n17341_, new_n17342_, new_n17343_,
    new_n17344_, new_n17345_, new_n17346_, new_n17347_, new_n17348_,
    new_n17349_, new_n17350_, new_n17351_, new_n17352_, new_n17353_,
    new_n17354_, new_n17355_, new_n17356_, new_n17357_, new_n17358_,
    new_n17359_, new_n17360_, new_n17361_, new_n17362_, new_n17363_,
    new_n17364_, new_n17365_, new_n17366_, new_n17367_, new_n17368_,
    new_n17369_, new_n17370_, new_n17371_, new_n17372_, new_n17373_,
    new_n17374_, new_n17375_, new_n17376_, new_n17377_, new_n17378_,
    new_n17379_, new_n17380_, new_n17381_, new_n17382_, new_n17383_,
    new_n17384_, new_n17385_, new_n17386_, new_n17387_, new_n17388_,
    new_n17389_, new_n17390_, new_n17391_, new_n17392_, new_n17393_,
    new_n17394_, new_n17395_, new_n17396_, new_n17397_, new_n17398_,
    new_n17399_, new_n17400_, new_n17401_, new_n17402_, new_n17403_,
    new_n17404_, new_n17405_, new_n17406_, new_n17407_, new_n17408_,
    new_n17409_, new_n17410_, new_n17411_, new_n17412_, new_n17413_,
    new_n17414_, new_n17415_, new_n17416_, new_n17417_, new_n17418_,
    new_n17419_, new_n17420_, new_n17421_, new_n17422_, new_n17423_,
    new_n17424_, new_n17425_, new_n17426_, new_n17427_, new_n17428_,
    new_n17429_, new_n17430_, new_n17431_, new_n17432_, new_n17433_,
    new_n17434_, new_n17435_, new_n17436_, new_n17437_, new_n17438_,
    new_n17439_, new_n17440_, new_n17441_, new_n17442_, new_n17443_,
    new_n17444_, new_n17445_, new_n17446_, new_n17447_, new_n17448_,
    new_n17449_, new_n17450_, new_n17451_, new_n17452_, new_n17453_,
    new_n17454_, new_n17455_, new_n17456_, new_n17457_, new_n17458_,
    new_n17459_, new_n17460_, new_n17461_, new_n17462_, new_n17463_,
    new_n17464_, new_n17465_, new_n17466_, new_n17467_, new_n17468_,
    new_n17469_, new_n17470_, new_n17471_, new_n17472_, new_n17473_,
    new_n17474_, new_n17475_, new_n17476_, new_n17477_, new_n17478_,
    new_n17479_, new_n17480_, new_n17481_, new_n17482_, new_n17483_,
    new_n17484_, new_n17485_, new_n17486_, new_n17487_, new_n17488_,
    new_n17489_, new_n17490_, new_n17491_, new_n17492_, new_n17493_,
    new_n17494_, new_n17495_, new_n17496_, new_n17497_, new_n17498_,
    new_n17499_, new_n17500_, new_n17501_, new_n17502_, new_n17503_,
    new_n17504_, new_n17505_, new_n17506_, new_n17507_, new_n17508_,
    new_n17509_, new_n17510_, new_n17511_, new_n17512_, new_n17513_,
    new_n17514_, new_n17515_, new_n17516_, new_n17517_, new_n17518_,
    new_n17519_, new_n17520_, new_n17521_, new_n17522_, new_n17523_,
    new_n17524_, new_n17525_, new_n17526_, new_n17527_, new_n17528_,
    new_n17529_, new_n17530_, new_n17531_, new_n17532_, new_n17533_,
    new_n17534_, new_n17535_, new_n17536_, new_n17537_, new_n17538_,
    new_n17539_, new_n17540_, new_n17541_, new_n17542_, new_n17543_,
    new_n17544_, new_n17545_, new_n17546_, new_n17547_, new_n17548_,
    new_n17549_, new_n17550_, new_n17551_, new_n17552_, new_n17553_,
    new_n17554_, new_n17555_, new_n17556_, new_n17557_, new_n17558_,
    new_n17559_, new_n17560_, new_n17561_, new_n17562_, new_n17563_,
    new_n17564_, new_n17565_, new_n17566_, new_n17567_, new_n17568_,
    new_n17569_, new_n17570_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17576_, new_n17577_, new_n17578_,
    new_n17579_, new_n17580_, new_n17581_, new_n17582_, new_n17583_,
    new_n17584_, new_n17585_, new_n17586_, new_n17587_, new_n17588_,
    new_n17589_, new_n17590_, new_n17591_, new_n17592_, new_n17593_,
    new_n17594_, new_n17595_, new_n17596_, new_n17597_, new_n17598_,
    new_n17599_, new_n17600_, new_n17601_, new_n17602_, new_n17603_,
    new_n17604_, new_n17605_, new_n17606_, new_n17607_, new_n17608_,
    new_n17609_, new_n17612_, new_n17613_, new_n17614_, new_n17615_,
    new_n17616_, new_n17617_, new_n17618_, new_n17619_, new_n17620_,
    new_n17621_, new_n17622_, new_n17623_, new_n17624_, new_n17625_,
    new_n17626_, new_n17627_, new_n17628_, new_n17629_, new_n17630_,
    new_n17631_, new_n17632_, new_n17633_, new_n17634_, new_n17635_,
    new_n17636_, new_n17637_, new_n17638_, new_n17639_, new_n17640_,
    new_n17641_, new_n17642_, new_n17643_, new_n17644_, new_n17645_,
    new_n17646_, new_n17647_, new_n17648_, new_n17649_, new_n17650_,
    new_n17651_, new_n17652_, new_n17653_, new_n17654_, new_n17655_,
    new_n17656_, new_n17657_, new_n17658_, new_n17659_, new_n17660_,
    new_n17661_, new_n17662_, new_n17663_, new_n17664_, new_n17665_,
    new_n17666_, new_n17667_, new_n17668_, new_n17669_, new_n17670_,
    new_n17671_, new_n17672_, new_n17673_, new_n17674_, new_n17675_,
    new_n17676_, new_n17677_, new_n17678_, new_n17679_, new_n17680_,
    new_n17681_, new_n17682_, new_n17683_, new_n17684_, new_n17685_,
    new_n17686_, new_n17687_, new_n17688_, new_n17689_, new_n17690_,
    new_n17691_, new_n17692_, new_n17693_, new_n17694_, new_n17695_,
    new_n17696_, new_n17697_, new_n17698_, new_n17699_, new_n17700_,
    new_n17701_, new_n17702_, new_n17703_, new_n17704_, new_n17705_,
    new_n17706_, new_n17707_, new_n17708_, new_n17709_, new_n17710_,
    new_n17711_, new_n17712_, new_n17713_, new_n17714_, new_n17715_,
    new_n17716_, new_n17717_, new_n17718_, new_n17719_, new_n17720_,
    new_n17721_, new_n17722_, new_n17723_, new_n17724_, new_n17725_,
    new_n17726_, new_n17727_, new_n17728_, new_n17729_, new_n17730_,
    new_n17731_, new_n17732_, new_n17733_, new_n17734_, new_n17735_,
    new_n17736_, new_n17737_, new_n17738_, new_n17739_, new_n17740_,
    new_n17741_, new_n17742_, new_n17743_, new_n17744_, new_n17745_,
    new_n17746_, new_n17751_, new_n17752_, new_n17753_, new_n17754_,
    new_n17755_, new_n17756_, new_n17757_, new_n17758_, new_n17759_,
    new_n17760_, new_n17761_, new_n17762_, new_n17763_, new_n17764_,
    new_n17765_, new_n17766_, new_n17767_, new_n17768_, new_n17769_,
    new_n17770_, new_n17771_, new_n17772_, new_n17773_, new_n17774_,
    new_n17775_, new_n17776_, new_n17777_, new_n17778_, new_n17779_,
    new_n17780_, new_n17781_, new_n17782_, new_n17783_, new_n17784_,
    new_n17785_, new_n17786_, new_n17787_, new_n17788_, new_n17789_,
    new_n17790_, new_n17791_, new_n17792_, new_n17793_, new_n17794_,
    new_n17795_, new_n17796_, new_n17797_, new_n17798_, new_n17799_,
    new_n17800_, new_n17801_, new_n17802_, new_n17803_, new_n17804_,
    new_n17805_, new_n17806_, new_n17807_, new_n17808_, new_n17809_,
    new_n17810_, new_n17811_, new_n17812_, new_n17813_, new_n17814_,
    new_n17815_, new_n17816_, new_n17817_, new_n17818_, new_n17819_,
    new_n17820_, new_n17821_, new_n17822_, new_n17823_, new_n17824_,
    new_n17825_;
  INV_X1     g00000(.I(\A[835] ), .ZN(new_n1003_));
  INV_X1     g00001(.I(\A[836] ), .ZN(new_n1004_));
  NAND2_X1   g00002(.A1(new_n1004_), .A2(\A[837] ), .ZN(new_n1005_));
  INV_X1     g00003(.I(\A[837] ), .ZN(new_n1006_));
  NAND2_X1   g00004(.A1(new_n1006_), .A2(\A[836] ), .ZN(new_n1007_));
  AOI21_X1   g00005(.A1(new_n1005_), .A2(new_n1007_), .B(new_n1003_), .ZN(new_n1008_));
  NAND2_X1   g00006(.A1(\A[836] ), .A2(\A[837] ), .ZN(new_n1009_));
  NAND2_X1   g00007(.A1(new_n1004_), .A2(new_n1006_), .ZN(new_n1010_));
  AOI21_X1   g00008(.A1(new_n1010_), .A2(new_n1009_), .B(\A[835] ), .ZN(new_n1011_));
  NOR2_X1    g00009(.A1(new_n1011_), .A2(new_n1008_), .ZN(new_n1012_));
  INV_X1     g00010(.I(\A[838] ), .ZN(new_n1013_));
  INV_X1     g00011(.I(\A[839] ), .ZN(new_n1014_));
  NAND2_X1   g00012(.A1(new_n1014_), .A2(\A[840] ), .ZN(new_n1015_));
  INV_X1     g00013(.I(\A[840] ), .ZN(new_n1016_));
  NAND2_X1   g00014(.A1(new_n1016_), .A2(\A[839] ), .ZN(new_n1017_));
  AOI21_X1   g00015(.A1(new_n1015_), .A2(new_n1017_), .B(new_n1013_), .ZN(new_n1018_));
  NAND2_X1   g00016(.A1(\A[839] ), .A2(\A[840] ), .ZN(new_n1019_));
  NAND2_X1   g00017(.A1(new_n1014_), .A2(new_n1016_), .ZN(new_n1020_));
  AOI21_X1   g00018(.A1(new_n1020_), .A2(new_n1019_), .B(\A[838] ), .ZN(new_n1021_));
  NOR2_X1    g00019(.A1(new_n1021_), .A2(new_n1018_), .ZN(new_n1022_));
  NAND2_X1   g00020(.A1(new_n1009_), .A2(new_n1003_), .ZN(new_n1023_));
  NAND2_X1   g00021(.A1(new_n1023_), .A2(new_n1010_), .ZN(new_n1024_));
  NAND2_X1   g00022(.A1(new_n1019_), .A2(new_n1013_), .ZN(new_n1025_));
  NAND2_X1   g00023(.A1(new_n1025_), .A2(new_n1020_), .ZN(new_n1026_));
  NAND2_X1   g00024(.A1(new_n1024_), .A2(new_n1026_), .ZN(new_n1027_));
  NOR3_X1    g00025(.A1(new_n1012_), .A2(new_n1022_), .A3(new_n1027_), .ZN(new_n1028_));
  INV_X1     g00026(.I(\A[844] ), .ZN(new_n1029_));
  INV_X1     g00027(.I(\A[845] ), .ZN(new_n1030_));
  NAND2_X1   g00028(.A1(new_n1030_), .A2(\A[846] ), .ZN(new_n1031_));
  INV_X1     g00029(.I(\A[846] ), .ZN(new_n1032_));
  NAND2_X1   g00030(.A1(new_n1032_), .A2(\A[845] ), .ZN(new_n1033_));
  AOI21_X1   g00031(.A1(new_n1031_), .A2(new_n1033_), .B(new_n1029_), .ZN(new_n1034_));
  NAND2_X1   g00032(.A1(\A[845] ), .A2(\A[846] ), .ZN(new_n1035_));
  NOR2_X1    g00033(.A1(\A[845] ), .A2(\A[846] ), .ZN(new_n1036_));
  INV_X1     g00034(.I(new_n1036_), .ZN(new_n1037_));
  AOI21_X1   g00035(.A1(new_n1037_), .A2(new_n1035_), .B(\A[844] ), .ZN(new_n1038_));
  NOR2_X1    g00036(.A1(new_n1038_), .A2(new_n1034_), .ZN(new_n1039_));
  INV_X1     g00037(.I(\A[841] ), .ZN(new_n1040_));
  INV_X1     g00038(.I(\A[842] ), .ZN(new_n1041_));
  NAND2_X1   g00039(.A1(new_n1041_), .A2(\A[843] ), .ZN(new_n1042_));
  INV_X1     g00040(.I(\A[843] ), .ZN(new_n1043_));
  NAND2_X1   g00041(.A1(new_n1043_), .A2(\A[842] ), .ZN(new_n1044_));
  AOI21_X1   g00042(.A1(new_n1042_), .A2(new_n1044_), .B(new_n1040_), .ZN(new_n1045_));
  NAND2_X1   g00043(.A1(new_n1041_), .A2(new_n1043_), .ZN(new_n1046_));
  NAND2_X1   g00044(.A1(\A[842] ), .A2(\A[843] ), .ZN(new_n1047_));
  AOI21_X1   g00045(.A1(new_n1046_), .A2(new_n1047_), .B(\A[841] ), .ZN(new_n1048_));
  NOR2_X1    g00046(.A1(new_n1048_), .A2(new_n1045_), .ZN(new_n1049_));
  NAND2_X1   g00047(.A1(new_n1047_), .A2(new_n1040_), .ZN(new_n1050_));
  NAND2_X1   g00048(.A1(new_n1050_), .A2(new_n1046_), .ZN(new_n1051_));
  AOI21_X1   g00049(.A1(new_n1029_), .A2(new_n1035_), .B(new_n1036_), .ZN(new_n1052_));
  INV_X1     g00050(.I(new_n1052_), .ZN(new_n1053_));
  NAND2_X1   g00051(.A1(new_n1053_), .A2(new_n1051_), .ZN(new_n1054_));
  NOR3_X1    g00052(.A1(new_n1039_), .A2(new_n1054_), .A3(new_n1049_), .ZN(new_n1055_));
  NAND2_X1   g00053(.A1(new_n1055_), .A2(new_n1028_), .ZN(new_n1056_));
  INV_X1     g00054(.I(new_n1049_), .ZN(new_n1057_));
  NOR2_X1    g00055(.A1(new_n1057_), .A2(new_n1054_), .ZN(new_n1058_));
  INV_X1     g00056(.I(new_n1051_), .ZN(new_n1059_));
  NOR2_X1    g00057(.A1(new_n1059_), .A2(new_n1052_), .ZN(new_n1060_));
  NOR2_X1    g00058(.A1(new_n1060_), .A2(new_n1049_), .ZN(new_n1061_));
  OAI21_X1   g00059(.A1(new_n1058_), .A2(new_n1061_), .B(new_n1039_), .ZN(new_n1062_));
  INV_X1     g00060(.I(new_n1039_), .ZN(new_n1063_));
  NAND2_X1   g00061(.A1(new_n1060_), .A2(new_n1049_), .ZN(new_n1064_));
  NAND2_X1   g00062(.A1(new_n1057_), .A2(new_n1054_), .ZN(new_n1065_));
  NAND3_X1   g00063(.A1(new_n1065_), .A2(new_n1064_), .A3(new_n1063_), .ZN(new_n1066_));
  INV_X1     g00064(.I(new_n1028_), .ZN(new_n1067_));
  NAND2_X1   g00065(.A1(new_n1059_), .A2(new_n1052_), .ZN(new_n1068_));
  NAND3_X1   g00066(.A1(new_n1063_), .A2(new_n1057_), .A3(new_n1068_), .ZN(new_n1069_));
  NOR2_X1    g00067(.A1(new_n1067_), .A2(new_n1069_), .ZN(new_n1070_));
  INV_X1     g00068(.I(new_n1022_), .ZN(new_n1071_));
  XNOR2_X1   g00069(.A1(new_n1012_), .A2(new_n1027_), .ZN(new_n1072_));
  NOR2_X1    g00070(.A1(new_n1072_), .A2(new_n1071_), .ZN(new_n1073_));
  XOR2_X1    g00071(.A1(new_n1012_), .A2(new_n1027_), .Z(new_n1074_));
  NOR2_X1    g00072(.A1(new_n1074_), .A2(new_n1022_), .ZN(new_n1075_));
  NOR2_X1    g00073(.A1(new_n1073_), .A2(new_n1075_), .ZN(new_n1076_));
  AND2_X2    g00074(.A1(new_n1062_), .A2(new_n1066_), .Z(new_n1077_));
  NOR2_X1    g00075(.A1(new_n1077_), .A2(new_n1056_), .ZN(new_n1078_));
  INV_X1     g00076(.I(new_n1056_), .ZN(new_n1079_));
  NAND2_X1   g00077(.A1(new_n1062_), .A2(new_n1066_), .ZN(new_n1080_));
  INV_X1     g00078(.I(new_n1080_), .ZN(new_n1081_));
  NOR2_X1    g00079(.A1(new_n1081_), .A2(new_n1079_), .ZN(new_n1082_));
  NOR2_X1    g00080(.A1(new_n1080_), .A2(new_n1056_), .ZN(new_n1083_));
  OAI21_X1   g00081(.A1(new_n1082_), .A2(new_n1083_), .B(new_n1076_), .ZN(new_n1084_));
  XNOR2_X1   g00082(.A1(new_n1055_), .A2(new_n1028_), .ZN(new_n1085_));
  INV_X1     g00083(.I(\A[823] ), .ZN(new_n1086_));
  INV_X1     g00084(.I(\A[824] ), .ZN(new_n1087_));
  NAND2_X1   g00085(.A1(new_n1087_), .A2(\A[825] ), .ZN(new_n1088_));
  INV_X1     g00086(.I(\A[825] ), .ZN(new_n1089_));
  NAND2_X1   g00087(.A1(new_n1089_), .A2(\A[824] ), .ZN(new_n1090_));
  AOI21_X1   g00088(.A1(new_n1088_), .A2(new_n1090_), .B(new_n1086_), .ZN(new_n1091_));
  NAND2_X1   g00089(.A1(\A[824] ), .A2(\A[825] ), .ZN(new_n1092_));
  NAND2_X1   g00090(.A1(new_n1087_), .A2(new_n1089_), .ZN(new_n1093_));
  AOI21_X1   g00091(.A1(new_n1093_), .A2(new_n1092_), .B(\A[823] ), .ZN(new_n1094_));
  NOR2_X1    g00092(.A1(new_n1094_), .A2(new_n1091_), .ZN(new_n1095_));
  INV_X1     g00093(.I(\A[826] ), .ZN(new_n1096_));
  INV_X1     g00094(.I(\A[827] ), .ZN(new_n1097_));
  NAND2_X1   g00095(.A1(new_n1097_), .A2(\A[828] ), .ZN(new_n1098_));
  INV_X1     g00096(.I(\A[828] ), .ZN(new_n1099_));
  NAND2_X1   g00097(.A1(new_n1099_), .A2(\A[827] ), .ZN(new_n1100_));
  AOI21_X1   g00098(.A1(new_n1098_), .A2(new_n1100_), .B(new_n1096_), .ZN(new_n1101_));
  NAND2_X1   g00099(.A1(\A[827] ), .A2(\A[828] ), .ZN(new_n1102_));
  NOR2_X1    g00100(.A1(\A[827] ), .A2(\A[828] ), .ZN(new_n1103_));
  INV_X1     g00101(.I(new_n1103_), .ZN(new_n1104_));
  AOI21_X1   g00102(.A1(new_n1104_), .A2(new_n1102_), .B(\A[826] ), .ZN(new_n1105_));
  NOR2_X1    g00103(.A1(new_n1105_), .A2(new_n1101_), .ZN(new_n1106_));
  NAND2_X1   g00104(.A1(new_n1092_), .A2(new_n1086_), .ZN(new_n1107_));
  NAND2_X1   g00105(.A1(new_n1107_), .A2(new_n1093_), .ZN(new_n1108_));
  NAND2_X1   g00106(.A1(new_n1102_), .A2(new_n1096_), .ZN(new_n1109_));
  NAND2_X1   g00107(.A1(new_n1109_), .A2(new_n1104_), .ZN(new_n1110_));
  NAND2_X1   g00108(.A1(new_n1110_), .A2(new_n1108_), .ZN(new_n1111_));
  NOR3_X1    g00109(.A1(new_n1095_), .A2(new_n1106_), .A3(new_n1111_), .ZN(new_n1112_));
  INV_X1     g00110(.I(\A[829] ), .ZN(new_n1113_));
  INV_X1     g00111(.I(\A[830] ), .ZN(new_n1114_));
  NAND2_X1   g00112(.A1(new_n1114_), .A2(\A[831] ), .ZN(new_n1115_));
  INV_X1     g00113(.I(\A[831] ), .ZN(new_n1116_));
  NAND2_X1   g00114(.A1(new_n1116_), .A2(\A[830] ), .ZN(new_n1117_));
  AOI21_X1   g00115(.A1(new_n1115_), .A2(new_n1117_), .B(new_n1113_), .ZN(new_n1118_));
  NOR2_X1    g00116(.A1(\A[830] ), .A2(\A[831] ), .ZN(new_n1119_));
  INV_X1     g00117(.I(new_n1119_), .ZN(new_n1120_));
  NAND2_X1   g00118(.A1(\A[830] ), .A2(\A[831] ), .ZN(new_n1121_));
  AOI21_X1   g00119(.A1(new_n1120_), .A2(new_n1121_), .B(\A[829] ), .ZN(new_n1122_));
  NOR2_X1    g00120(.A1(new_n1122_), .A2(new_n1118_), .ZN(new_n1123_));
  INV_X1     g00121(.I(\A[832] ), .ZN(new_n1124_));
  INV_X1     g00122(.I(\A[833] ), .ZN(new_n1125_));
  NAND2_X1   g00123(.A1(new_n1125_), .A2(\A[834] ), .ZN(new_n1126_));
  INV_X1     g00124(.I(\A[834] ), .ZN(new_n1127_));
  NAND2_X1   g00125(.A1(new_n1127_), .A2(\A[833] ), .ZN(new_n1128_));
  AOI21_X1   g00126(.A1(new_n1126_), .A2(new_n1128_), .B(new_n1124_), .ZN(new_n1129_));
  NAND2_X1   g00127(.A1(\A[833] ), .A2(\A[834] ), .ZN(new_n1130_));
  NOR2_X1    g00128(.A1(\A[833] ), .A2(\A[834] ), .ZN(new_n1131_));
  INV_X1     g00129(.I(new_n1131_), .ZN(new_n1132_));
  AOI21_X1   g00130(.A1(new_n1132_), .A2(new_n1130_), .B(\A[832] ), .ZN(new_n1133_));
  NOR2_X1    g00131(.A1(new_n1133_), .A2(new_n1129_), .ZN(new_n1134_));
  AOI21_X1   g00132(.A1(new_n1113_), .A2(new_n1121_), .B(new_n1119_), .ZN(new_n1135_));
  AOI21_X1   g00133(.A1(new_n1124_), .A2(new_n1130_), .B(new_n1131_), .ZN(new_n1136_));
  NOR2_X1    g00134(.A1(new_n1135_), .A2(new_n1136_), .ZN(new_n1137_));
  INV_X1     g00135(.I(new_n1137_), .ZN(new_n1138_));
  NOR3_X1    g00136(.A1(new_n1138_), .A2(new_n1123_), .A3(new_n1134_), .ZN(new_n1139_));
  XNOR2_X1   g00137(.A1(new_n1139_), .A2(new_n1112_), .ZN(new_n1140_));
  NOR2_X1    g00138(.A1(new_n1116_), .A2(\A[830] ), .ZN(new_n1141_));
  NOR2_X1    g00139(.A1(new_n1114_), .A2(\A[831] ), .ZN(new_n1142_));
  OAI21_X1   g00140(.A1(new_n1141_), .A2(new_n1142_), .B(\A[829] ), .ZN(new_n1143_));
  INV_X1     g00141(.I(new_n1121_), .ZN(new_n1144_));
  OAI21_X1   g00142(.A1(new_n1144_), .A2(new_n1119_), .B(new_n1113_), .ZN(new_n1145_));
  NAND2_X1   g00143(.A1(new_n1143_), .A2(new_n1145_), .ZN(new_n1146_));
  NOR2_X1    g00144(.A1(new_n1138_), .A2(new_n1146_), .ZN(new_n1147_));
  NOR2_X1    g00145(.A1(new_n1123_), .A2(new_n1137_), .ZN(new_n1148_));
  OAI21_X1   g00146(.A1(new_n1147_), .A2(new_n1148_), .B(new_n1134_), .ZN(new_n1149_));
  INV_X1     g00147(.I(new_n1134_), .ZN(new_n1150_));
  NAND2_X1   g00148(.A1(new_n1123_), .A2(new_n1137_), .ZN(new_n1151_));
  NAND2_X1   g00149(.A1(new_n1138_), .A2(new_n1146_), .ZN(new_n1152_));
  NAND3_X1   g00150(.A1(new_n1152_), .A2(new_n1151_), .A3(new_n1150_), .ZN(new_n1153_));
  NAND2_X1   g00151(.A1(new_n1149_), .A2(new_n1153_), .ZN(new_n1154_));
  NAND2_X1   g00152(.A1(new_n1139_), .A2(new_n1112_), .ZN(new_n1155_));
  INV_X1     g00153(.I(new_n1155_), .ZN(new_n1156_));
  INV_X1     g00154(.I(new_n1106_), .ZN(new_n1157_));
  INV_X1     g00155(.I(new_n1108_), .ZN(new_n1158_));
  AOI21_X1   g00156(.A1(new_n1096_), .A2(new_n1102_), .B(new_n1103_), .ZN(new_n1159_));
  NOR2_X1    g00157(.A1(new_n1158_), .A2(new_n1159_), .ZN(new_n1160_));
  NAND2_X1   g00158(.A1(new_n1160_), .A2(new_n1095_), .ZN(new_n1161_));
  INV_X1     g00159(.I(new_n1095_), .ZN(new_n1162_));
  NAND2_X1   g00160(.A1(new_n1162_), .A2(new_n1111_), .ZN(new_n1163_));
  AOI21_X1   g00161(.A1(new_n1163_), .A2(new_n1161_), .B(new_n1157_), .ZN(new_n1164_));
  NOR2_X1    g00162(.A1(new_n1162_), .A2(new_n1111_), .ZN(new_n1165_));
  NOR2_X1    g00163(.A1(new_n1160_), .A2(new_n1095_), .ZN(new_n1166_));
  NOR3_X1    g00164(.A1(new_n1165_), .A2(new_n1166_), .A3(new_n1106_), .ZN(new_n1167_));
  NOR2_X1    g00165(.A1(new_n1167_), .A2(new_n1164_), .ZN(new_n1168_));
  AND2_X2    g00166(.A1(new_n1135_), .A2(new_n1136_), .Z(new_n1169_));
  NOR3_X1    g00167(.A1(new_n1169_), .A2(new_n1123_), .A3(new_n1134_), .ZN(new_n1170_));
  AND2_X2    g00168(.A1(new_n1170_), .A2(new_n1112_), .Z(new_n1171_));
  NOR3_X1    g00169(.A1(new_n1168_), .A2(new_n1154_), .A3(new_n1156_), .ZN(new_n1172_));
  NAND3_X1   g00170(.A1(new_n1172_), .A2(new_n1085_), .A3(new_n1140_), .ZN(new_n1173_));
  XOR2_X1    g00171(.A1(new_n1084_), .A2(new_n1173_), .Z(new_n1174_));
  NAND2_X1   g00172(.A1(new_n1174_), .A2(new_n1078_), .ZN(new_n1175_));
  NAND2_X1   g00173(.A1(new_n1085_), .A2(new_n1140_), .ZN(new_n1176_));
  INV_X1     g00174(.I(new_n1176_), .ZN(new_n1177_));
  NOR2_X1    g00175(.A1(new_n1085_), .A2(new_n1140_), .ZN(new_n1178_));
  INV_X1     g00176(.I(\A[811] ), .ZN(new_n1179_));
  INV_X1     g00177(.I(\A[812] ), .ZN(new_n1180_));
  NAND2_X1   g00178(.A1(new_n1180_), .A2(\A[813] ), .ZN(new_n1181_));
  INV_X1     g00179(.I(\A[813] ), .ZN(new_n1182_));
  NAND2_X1   g00180(.A1(new_n1182_), .A2(\A[812] ), .ZN(new_n1183_));
  AOI21_X1   g00181(.A1(new_n1181_), .A2(new_n1183_), .B(new_n1179_), .ZN(new_n1184_));
  NAND2_X1   g00182(.A1(\A[812] ), .A2(\A[813] ), .ZN(new_n1185_));
  NAND2_X1   g00183(.A1(new_n1180_), .A2(new_n1182_), .ZN(new_n1186_));
  AOI21_X1   g00184(.A1(new_n1186_), .A2(new_n1185_), .B(\A[811] ), .ZN(new_n1187_));
  NOR2_X1    g00185(.A1(new_n1187_), .A2(new_n1184_), .ZN(new_n1188_));
  INV_X1     g00186(.I(\A[814] ), .ZN(new_n1189_));
  INV_X1     g00187(.I(\A[815] ), .ZN(new_n1190_));
  NAND2_X1   g00188(.A1(new_n1190_), .A2(\A[816] ), .ZN(new_n1191_));
  INV_X1     g00189(.I(\A[816] ), .ZN(new_n1192_));
  NAND2_X1   g00190(.A1(new_n1192_), .A2(\A[815] ), .ZN(new_n1193_));
  AOI21_X1   g00191(.A1(new_n1191_), .A2(new_n1193_), .B(new_n1189_), .ZN(new_n1194_));
  NAND2_X1   g00192(.A1(\A[815] ), .A2(\A[816] ), .ZN(new_n1195_));
  NAND2_X1   g00193(.A1(new_n1190_), .A2(new_n1192_), .ZN(new_n1196_));
  AOI21_X1   g00194(.A1(new_n1196_), .A2(new_n1195_), .B(\A[814] ), .ZN(new_n1197_));
  NOR2_X1    g00195(.A1(new_n1197_), .A2(new_n1194_), .ZN(new_n1198_));
  NAND2_X1   g00196(.A1(new_n1185_), .A2(new_n1179_), .ZN(new_n1199_));
  NAND2_X1   g00197(.A1(new_n1199_), .A2(new_n1186_), .ZN(new_n1200_));
  NAND2_X1   g00198(.A1(new_n1195_), .A2(new_n1189_), .ZN(new_n1201_));
  NAND2_X1   g00199(.A1(new_n1201_), .A2(new_n1196_), .ZN(new_n1202_));
  NAND2_X1   g00200(.A1(new_n1200_), .A2(new_n1202_), .ZN(new_n1203_));
  NOR3_X1    g00201(.A1(new_n1188_), .A2(new_n1198_), .A3(new_n1203_), .ZN(new_n1204_));
  INV_X1     g00202(.I(\A[817] ), .ZN(new_n1205_));
  INV_X1     g00203(.I(\A[818] ), .ZN(new_n1206_));
  NAND2_X1   g00204(.A1(new_n1206_), .A2(\A[819] ), .ZN(new_n1207_));
  INV_X1     g00205(.I(\A[819] ), .ZN(new_n1208_));
  NAND2_X1   g00206(.A1(new_n1208_), .A2(\A[818] ), .ZN(new_n1209_));
  AOI21_X1   g00207(.A1(new_n1207_), .A2(new_n1209_), .B(new_n1205_), .ZN(new_n1210_));
  NOR2_X1    g00208(.A1(\A[818] ), .A2(\A[819] ), .ZN(new_n1211_));
  INV_X1     g00209(.I(new_n1211_), .ZN(new_n1212_));
  NAND2_X1   g00210(.A1(\A[818] ), .A2(\A[819] ), .ZN(new_n1213_));
  AOI21_X1   g00211(.A1(new_n1212_), .A2(new_n1213_), .B(\A[817] ), .ZN(new_n1214_));
  NOR2_X1    g00212(.A1(new_n1214_), .A2(new_n1210_), .ZN(new_n1215_));
  INV_X1     g00213(.I(\A[820] ), .ZN(new_n1216_));
  INV_X1     g00214(.I(\A[821] ), .ZN(new_n1217_));
  NAND2_X1   g00215(.A1(new_n1217_), .A2(\A[822] ), .ZN(new_n1218_));
  INV_X1     g00216(.I(\A[822] ), .ZN(new_n1219_));
  NAND2_X1   g00217(.A1(new_n1219_), .A2(\A[821] ), .ZN(new_n1220_));
  AOI21_X1   g00218(.A1(new_n1218_), .A2(new_n1220_), .B(new_n1216_), .ZN(new_n1221_));
  NAND2_X1   g00219(.A1(\A[821] ), .A2(\A[822] ), .ZN(new_n1222_));
  NOR2_X1    g00220(.A1(\A[821] ), .A2(\A[822] ), .ZN(new_n1223_));
  INV_X1     g00221(.I(new_n1223_), .ZN(new_n1224_));
  AOI21_X1   g00222(.A1(new_n1224_), .A2(new_n1222_), .B(\A[820] ), .ZN(new_n1225_));
  NOR2_X1    g00223(.A1(new_n1225_), .A2(new_n1221_), .ZN(new_n1226_));
  AOI21_X1   g00224(.A1(new_n1205_), .A2(new_n1213_), .B(new_n1211_), .ZN(new_n1227_));
  AOI21_X1   g00225(.A1(new_n1216_), .A2(new_n1222_), .B(new_n1223_), .ZN(new_n1228_));
  OR2_X2     g00226(.A1(new_n1227_), .A2(new_n1228_), .Z(new_n1229_));
  NOR3_X1    g00227(.A1(new_n1229_), .A2(new_n1215_), .A3(new_n1226_), .ZN(new_n1230_));
  XOR2_X1    g00228(.A1(new_n1230_), .A2(new_n1204_), .Z(new_n1231_));
  INV_X1     g00229(.I(\A[807] ), .ZN(new_n1232_));
  NOR2_X1    g00230(.A1(new_n1232_), .A2(\A[806] ), .ZN(new_n1233_));
  INV_X1     g00231(.I(\A[806] ), .ZN(new_n1234_));
  NOR2_X1    g00232(.A1(new_n1234_), .A2(\A[807] ), .ZN(new_n1235_));
  OAI21_X1   g00233(.A1(new_n1233_), .A2(new_n1235_), .B(\A[805] ), .ZN(new_n1236_));
  INV_X1     g00234(.I(\A[805] ), .ZN(new_n1237_));
  NAND2_X1   g00235(.A1(\A[806] ), .A2(\A[807] ), .ZN(new_n1238_));
  INV_X1     g00236(.I(new_n1238_), .ZN(new_n1239_));
  NOR2_X1    g00237(.A1(\A[806] ), .A2(\A[807] ), .ZN(new_n1240_));
  OAI21_X1   g00238(.A1(new_n1239_), .A2(new_n1240_), .B(new_n1237_), .ZN(new_n1241_));
  NAND2_X1   g00239(.A1(new_n1236_), .A2(new_n1241_), .ZN(new_n1242_));
  INV_X1     g00240(.I(\A[810] ), .ZN(new_n1243_));
  NOR2_X1    g00241(.A1(new_n1243_), .A2(\A[809] ), .ZN(new_n1244_));
  INV_X1     g00242(.I(\A[809] ), .ZN(new_n1245_));
  NOR2_X1    g00243(.A1(new_n1245_), .A2(\A[810] ), .ZN(new_n1246_));
  OAI21_X1   g00244(.A1(new_n1244_), .A2(new_n1246_), .B(\A[808] ), .ZN(new_n1247_));
  INV_X1     g00245(.I(\A[808] ), .ZN(new_n1248_));
  NAND2_X1   g00246(.A1(\A[809] ), .A2(\A[810] ), .ZN(new_n1249_));
  INV_X1     g00247(.I(new_n1249_), .ZN(new_n1250_));
  NOR2_X1    g00248(.A1(\A[809] ), .A2(\A[810] ), .ZN(new_n1251_));
  OAI21_X1   g00249(.A1(new_n1250_), .A2(new_n1251_), .B(new_n1248_), .ZN(new_n1252_));
  NAND2_X1   g00250(.A1(new_n1247_), .A2(new_n1252_), .ZN(new_n1253_));
  AOI21_X1   g00251(.A1(new_n1237_), .A2(new_n1238_), .B(new_n1240_), .ZN(new_n1254_));
  AOI21_X1   g00252(.A1(new_n1248_), .A2(new_n1249_), .B(new_n1251_), .ZN(new_n1255_));
  NOR2_X1    g00253(.A1(new_n1254_), .A2(new_n1255_), .ZN(new_n1256_));
  NAND3_X1   g00254(.A1(new_n1242_), .A2(new_n1253_), .A3(new_n1256_), .ZN(new_n1257_));
  INV_X1     g00255(.I(\A[799] ), .ZN(new_n1258_));
  INV_X1     g00256(.I(\A[800] ), .ZN(new_n1259_));
  NAND2_X1   g00257(.A1(new_n1259_), .A2(\A[801] ), .ZN(new_n1260_));
  INV_X1     g00258(.I(\A[801] ), .ZN(new_n1261_));
  NAND2_X1   g00259(.A1(new_n1261_), .A2(\A[800] ), .ZN(new_n1262_));
  AOI21_X1   g00260(.A1(new_n1260_), .A2(new_n1262_), .B(new_n1258_), .ZN(new_n1263_));
  NAND2_X1   g00261(.A1(\A[800] ), .A2(\A[801] ), .ZN(new_n1264_));
  NAND2_X1   g00262(.A1(new_n1259_), .A2(new_n1261_), .ZN(new_n1265_));
  AOI21_X1   g00263(.A1(new_n1265_), .A2(new_n1264_), .B(\A[799] ), .ZN(new_n1266_));
  NOR2_X1    g00264(.A1(new_n1266_), .A2(new_n1263_), .ZN(new_n1267_));
  INV_X1     g00265(.I(\A[802] ), .ZN(new_n1268_));
  INV_X1     g00266(.I(\A[803] ), .ZN(new_n1269_));
  NAND2_X1   g00267(.A1(new_n1269_), .A2(\A[804] ), .ZN(new_n1270_));
  INV_X1     g00268(.I(\A[804] ), .ZN(new_n1271_));
  NAND2_X1   g00269(.A1(new_n1271_), .A2(\A[803] ), .ZN(new_n1272_));
  AOI21_X1   g00270(.A1(new_n1270_), .A2(new_n1272_), .B(new_n1268_), .ZN(new_n1273_));
  NAND2_X1   g00271(.A1(\A[803] ), .A2(\A[804] ), .ZN(new_n1274_));
  NAND2_X1   g00272(.A1(new_n1269_), .A2(new_n1271_), .ZN(new_n1275_));
  AOI21_X1   g00273(.A1(new_n1275_), .A2(new_n1274_), .B(\A[802] ), .ZN(new_n1276_));
  NOR2_X1    g00274(.A1(new_n1276_), .A2(new_n1273_), .ZN(new_n1277_));
  NAND2_X1   g00275(.A1(new_n1264_), .A2(new_n1258_), .ZN(new_n1278_));
  NAND2_X1   g00276(.A1(new_n1278_), .A2(new_n1265_), .ZN(new_n1279_));
  NAND2_X1   g00277(.A1(new_n1274_), .A2(new_n1268_), .ZN(new_n1280_));
  NAND2_X1   g00278(.A1(new_n1280_), .A2(new_n1275_), .ZN(new_n1281_));
  NAND2_X1   g00279(.A1(new_n1279_), .A2(new_n1281_), .ZN(new_n1282_));
  NOR3_X1    g00280(.A1(new_n1267_), .A2(new_n1277_), .A3(new_n1282_), .ZN(new_n1283_));
  XNOR2_X1   g00281(.A1(new_n1283_), .A2(new_n1257_), .ZN(new_n1284_));
  NAND2_X1   g00282(.A1(new_n1231_), .A2(new_n1284_), .ZN(new_n1285_));
  XNOR2_X1   g00283(.A1(new_n1230_), .A2(new_n1204_), .ZN(new_n1286_));
  XOR2_X1    g00284(.A1(new_n1283_), .A2(new_n1257_), .Z(new_n1287_));
  NAND2_X1   g00285(.A1(new_n1286_), .A2(new_n1287_), .ZN(new_n1288_));
  NAND2_X1   g00286(.A1(new_n1285_), .A2(new_n1288_), .ZN(new_n1289_));
  NOR3_X1    g00287(.A1(new_n1289_), .A2(new_n1177_), .A3(new_n1178_), .ZN(new_n1290_));
  INV_X1     g00288(.I(new_n1290_), .ZN(new_n1291_));
  INV_X1     g00289(.I(new_n1198_), .ZN(new_n1292_));
  NAND3_X1   g00290(.A1(new_n1188_), .A2(new_n1200_), .A3(new_n1202_), .ZN(new_n1293_));
  INV_X1     g00291(.I(new_n1188_), .ZN(new_n1294_));
  NAND2_X1   g00292(.A1(new_n1294_), .A2(new_n1203_), .ZN(new_n1295_));
  AOI21_X1   g00293(.A1(new_n1295_), .A2(new_n1293_), .B(new_n1292_), .ZN(new_n1296_));
  AND3_X2    g00294(.A1(new_n1293_), .A2(new_n1295_), .A3(new_n1292_), .Z(new_n1297_));
  NOR2_X1    g00295(.A1(new_n1297_), .A2(new_n1296_), .ZN(new_n1298_));
  AND2_X2    g00296(.A1(new_n1230_), .A2(new_n1204_), .Z(new_n1299_));
  NOR2_X1    g00297(.A1(new_n1208_), .A2(\A[818] ), .ZN(new_n1300_));
  NOR2_X1    g00298(.A1(new_n1206_), .A2(\A[819] ), .ZN(new_n1301_));
  OAI21_X1   g00299(.A1(new_n1300_), .A2(new_n1301_), .B(\A[817] ), .ZN(new_n1302_));
  INV_X1     g00300(.I(new_n1213_), .ZN(new_n1303_));
  OAI21_X1   g00301(.A1(new_n1303_), .A2(new_n1211_), .B(new_n1205_), .ZN(new_n1304_));
  NAND2_X1   g00302(.A1(new_n1302_), .A2(new_n1304_), .ZN(new_n1305_));
  NOR2_X1    g00303(.A1(new_n1229_), .A2(new_n1305_), .ZN(new_n1306_));
  NOR2_X1    g00304(.A1(new_n1227_), .A2(new_n1228_), .ZN(new_n1307_));
  NOR2_X1    g00305(.A1(new_n1215_), .A2(new_n1307_), .ZN(new_n1308_));
  OAI21_X1   g00306(.A1(new_n1306_), .A2(new_n1308_), .B(new_n1226_), .ZN(new_n1309_));
  INV_X1     g00307(.I(new_n1226_), .ZN(new_n1310_));
  NAND2_X1   g00308(.A1(new_n1215_), .A2(new_n1307_), .ZN(new_n1311_));
  NAND2_X1   g00309(.A1(new_n1229_), .A2(new_n1305_), .ZN(new_n1312_));
  NAND3_X1   g00310(.A1(new_n1312_), .A2(new_n1311_), .A3(new_n1310_), .ZN(new_n1313_));
  NAND2_X1   g00311(.A1(new_n1309_), .A2(new_n1313_), .ZN(new_n1314_));
  XOR2_X1    g00312(.A1(new_n1314_), .A2(new_n1299_), .Z(new_n1315_));
  NAND2_X1   g00313(.A1(new_n1315_), .A2(new_n1298_), .ZN(new_n1316_));
  INV_X1     g00314(.I(new_n1314_), .ZN(new_n1317_));
  NAND2_X1   g00315(.A1(new_n1227_), .A2(new_n1228_), .ZN(new_n1318_));
  NAND4_X1   g00316(.A1(new_n1204_), .A2(new_n1305_), .A3(new_n1310_), .A4(new_n1318_), .ZN(new_n1319_));
  NOR2_X1    g00317(.A1(new_n1317_), .A2(new_n1319_), .ZN(new_n1320_));
  INV_X1     g00318(.I(new_n1320_), .ZN(new_n1321_));
  NAND4_X1   g00319(.A1(new_n1204_), .A2(new_n1305_), .A3(new_n1310_), .A4(new_n1307_), .ZN(new_n1323_));
  INV_X1     g00320(.I(new_n1323_), .ZN(new_n1324_));
  NOR2_X1    g00321(.A1(new_n1231_), .A2(new_n1284_), .ZN(new_n1325_));
  NOR4_X1    g00322(.A1(new_n1257_), .A2(new_n1267_), .A3(new_n1277_), .A4(new_n1282_), .ZN(new_n1326_));
  INV_X1     g00323(.I(new_n1326_), .ZN(new_n1327_));
  INV_X1     g00324(.I(new_n1253_), .ZN(new_n1328_));
  INV_X1     g00325(.I(new_n1256_), .ZN(new_n1329_));
  NOR2_X1    g00326(.A1(new_n1329_), .A2(new_n1242_), .ZN(new_n1330_));
  AND2_X2    g00327(.A1(new_n1236_), .A2(new_n1241_), .Z(new_n1331_));
  NOR2_X1    g00328(.A1(new_n1331_), .A2(new_n1256_), .ZN(new_n1332_));
  OAI21_X1   g00329(.A1(new_n1332_), .A2(new_n1330_), .B(new_n1328_), .ZN(new_n1333_));
  OR3_X2     g00330(.A1(new_n1332_), .A2(new_n1328_), .A3(new_n1330_), .Z(new_n1334_));
  XOR2_X1    g00331(.A1(new_n1242_), .A2(new_n1253_), .Z(new_n1335_));
  NAND2_X1   g00332(.A1(new_n1335_), .A2(new_n1256_), .ZN(new_n1336_));
  NAND4_X1   g00333(.A1(new_n1336_), .A2(new_n1334_), .A3(new_n1327_), .A4(new_n1333_), .ZN(new_n1337_));
  INV_X1     g00334(.I(new_n1277_), .ZN(new_n1338_));
  NAND3_X1   g00335(.A1(new_n1267_), .A2(new_n1279_), .A3(new_n1281_), .ZN(new_n1339_));
  OAI21_X1   g00336(.A1(new_n1263_), .A2(new_n1266_), .B(new_n1282_), .ZN(new_n1340_));
  AOI21_X1   g00337(.A1(new_n1340_), .A2(new_n1339_), .B(new_n1338_), .ZN(new_n1341_));
  INV_X1     g00338(.I(new_n1341_), .ZN(new_n1342_));
  NAND3_X1   g00339(.A1(new_n1340_), .A2(new_n1339_), .A3(new_n1338_), .ZN(new_n1343_));
  NAND2_X1   g00340(.A1(new_n1342_), .A2(new_n1343_), .ZN(new_n1344_));
  XNOR2_X1   g00341(.A1(new_n1267_), .A2(new_n1277_), .ZN(new_n1345_));
  NOR3_X1    g00342(.A1(new_n1267_), .A2(new_n1277_), .A3(new_n1282_), .ZN(new_n1346_));
  NAND4_X1   g00343(.A1(new_n1345_), .A2(new_n1242_), .A3(new_n1253_), .A4(new_n1256_), .ZN(new_n1347_));
  NAND4_X1   g00344(.A1(new_n1325_), .A2(new_n1337_), .A3(new_n1344_), .A4(new_n1347_), .ZN(new_n1348_));
  NOR2_X1    g00345(.A1(new_n1348_), .A2(new_n1324_), .ZN(new_n1349_));
  INV_X1     g00346(.I(new_n1333_), .ZN(new_n1350_));
  NOR3_X1    g00347(.A1(new_n1332_), .A2(new_n1328_), .A3(new_n1330_), .ZN(new_n1351_));
  XNOR2_X1   g00348(.A1(new_n1242_), .A2(new_n1253_), .ZN(new_n1352_));
  NOR2_X1    g00349(.A1(new_n1352_), .A2(new_n1329_), .ZN(new_n1353_));
  NOR4_X1    g00350(.A1(new_n1353_), .A2(new_n1350_), .A3(new_n1326_), .A4(new_n1351_), .ZN(new_n1354_));
  INV_X1     g00351(.I(new_n1343_), .ZN(new_n1355_));
  NOR2_X1    g00352(.A1(new_n1355_), .A2(new_n1341_), .ZN(new_n1356_));
  INV_X1     g00353(.I(new_n1347_), .ZN(new_n1357_));
  NOR4_X1    g00354(.A1(new_n1288_), .A2(new_n1354_), .A3(new_n1356_), .A4(new_n1357_), .ZN(new_n1358_));
  NOR2_X1    g00355(.A1(new_n1358_), .A2(new_n1323_), .ZN(new_n1359_));
  OAI21_X1   g00356(.A1(new_n1359_), .A2(new_n1349_), .B(new_n1316_), .ZN(new_n1360_));
  INV_X1     g00357(.I(new_n1316_), .ZN(new_n1361_));
  NAND2_X1   g00358(.A1(new_n1358_), .A2(new_n1323_), .ZN(new_n1362_));
  NAND2_X1   g00359(.A1(new_n1348_), .A2(new_n1324_), .ZN(new_n1363_));
  NAND3_X1   g00360(.A1(new_n1361_), .A2(new_n1362_), .A3(new_n1363_), .ZN(new_n1364_));
  AOI21_X1   g00361(.A1(new_n1364_), .A2(new_n1360_), .B(new_n1291_), .ZN(new_n1365_));
  INV_X1     g00362(.I(\A[790] ), .ZN(new_n1366_));
  INV_X1     g00363(.I(\A[791] ), .ZN(new_n1367_));
  NAND2_X1   g00364(.A1(new_n1367_), .A2(\A[792] ), .ZN(new_n1368_));
  INV_X1     g00365(.I(\A[792] ), .ZN(new_n1369_));
  NAND2_X1   g00366(.A1(new_n1369_), .A2(\A[791] ), .ZN(new_n1370_));
  AOI21_X1   g00367(.A1(new_n1368_), .A2(new_n1370_), .B(new_n1366_), .ZN(new_n1371_));
  NOR2_X1    g00368(.A1(\A[791] ), .A2(\A[792] ), .ZN(new_n1372_));
  INV_X1     g00369(.I(new_n1372_), .ZN(new_n1373_));
  NAND2_X1   g00370(.A1(\A[791] ), .A2(\A[792] ), .ZN(new_n1374_));
  AOI21_X1   g00371(.A1(new_n1373_), .A2(new_n1374_), .B(\A[790] ), .ZN(new_n1375_));
  NOR2_X1    g00372(.A1(new_n1375_), .A2(new_n1371_), .ZN(new_n1376_));
  AOI21_X1   g00373(.A1(new_n1366_), .A2(new_n1374_), .B(new_n1372_), .ZN(new_n1377_));
  INV_X1     g00374(.I(\A[787] ), .ZN(new_n1378_));
  NOR2_X1    g00375(.A1(\A[788] ), .A2(\A[789] ), .ZN(new_n1379_));
  NAND2_X1   g00376(.A1(\A[788] ), .A2(\A[789] ), .ZN(new_n1380_));
  AOI21_X1   g00377(.A1(new_n1378_), .A2(new_n1380_), .B(new_n1379_), .ZN(new_n1381_));
  NOR2_X1    g00378(.A1(new_n1377_), .A2(new_n1381_), .ZN(new_n1382_));
  INV_X1     g00379(.I(\A[788] ), .ZN(new_n1383_));
  NAND2_X1   g00380(.A1(new_n1383_), .A2(\A[789] ), .ZN(new_n1384_));
  INV_X1     g00381(.I(\A[789] ), .ZN(new_n1385_));
  NAND2_X1   g00382(.A1(new_n1385_), .A2(\A[788] ), .ZN(new_n1386_));
  AOI21_X1   g00383(.A1(new_n1384_), .A2(new_n1386_), .B(new_n1378_), .ZN(new_n1387_));
  INV_X1     g00384(.I(new_n1379_), .ZN(new_n1388_));
  AOI21_X1   g00385(.A1(new_n1388_), .A2(new_n1380_), .B(\A[787] ), .ZN(new_n1389_));
  NOR2_X1    g00386(.A1(new_n1389_), .A2(new_n1387_), .ZN(new_n1390_));
  NAND2_X1   g00387(.A1(new_n1390_), .A2(new_n1382_), .ZN(new_n1391_));
  INV_X1     g00388(.I(new_n1382_), .ZN(new_n1392_));
  NOR2_X1    g00389(.A1(new_n1385_), .A2(\A[788] ), .ZN(new_n1393_));
  NOR2_X1    g00390(.A1(new_n1383_), .A2(\A[789] ), .ZN(new_n1394_));
  OAI21_X1   g00391(.A1(new_n1393_), .A2(new_n1394_), .B(\A[787] ), .ZN(new_n1395_));
  INV_X1     g00392(.I(new_n1380_), .ZN(new_n1396_));
  OAI21_X1   g00393(.A1(new_n1396_), .A2(new_n1379_), .B(new_n1378_), .ZN(new_n1397_));
  NAND2_X1   g00394(.A1(new_n1395_), .A2(new_n1397_), .ZN(new_n1398_));
  NAND2_X1   g00395(.A1(new_n1392_), .A2(new_n1398_), .ZN(new_n1399_));
  NAND2_X1   g00396(.A1(new_n1399_), .A2(new_n1391_), .ZN(new_n1400_));
  NAND2_X1   g00397(.A1(new_n1400_), .A2(new_n1376_), .ZN(new_n1401_));
  NOR2_X1    g00398(.A1(new_n1369_), .A2(\A[791] ), .ZN(new_n1402_));
  NOR2_X1    g00399(.A1(new_n1367_), .A2(\A[792] ), .ZN(new_n1403_));
  OAI21_X1   g00400(.A1(new_n1402_), .A2(new_n1403_), .B(\A[790] ), .ZN(new_n1404_));
  INV_X1     g00401(.I(new_n1374_), .ZN(new_n1405_));
  OAI21_X1   g00402(.A1(new_n1405_), .A2(new_n1372_), .B(new_n1366_), .ZN(new_n1406_));
  NAND2_X1   g00403(.A1(new_n1404_), .A2(new_n1406_), .ZN(new_n1407_));
  NAND3_X1   g00404(.A1(new_n1399_), .A2(new_n1391_), .A3(new_n1407_), .ZN(new_n1408_));
  NAND2_X1   g00405(.A1(new_n1401_), .A2(new_n1408_), .ZN(new_n1409_));
  INV_X1     g00406(.I(new_n1409_), .ZN(new_n1410_));
  INV_X1     g00407(.I(\A[798] ), .ZN(new_n1411_));
  NOR2_X1    g00408(.A1(new_n1411_), .A2(\A[797] ), .ZN(new_n1412_));
  INV_X1     g00409(.I(\A[797] ), .ZN(new_n1413_));
  NOR2_X1    g00410(.A1(new_n1413_), .A2(\A[798] ), .ZN(new_n1414_));
  OAI21_X1   g00411(.A1(new_n1412_), .A2(new_n1414_), .B(\A[796] ), .ZN(new_n1415_));
  INV_X1     g00412(.I(\A[796] ), .ZN(new_n1416_));
  NOR2_X1    g00413(.A1(\A[797] ), .A2(\A[798] ), .ZN(new_n1417_));
  NAND2_X1   g00414(.A1(\A[797] ), .A2(\A[798] ), .ZN(new_n1418_));
  INV_X1     g00415(.I(new_n1418_), .ZN(new_n1419_));
  OAI21_X1   g00416(.A1(new_n1419_), .A2(new_n1417_), .B(new_n1416_), .ZN(new_n1420_));
  NAND2_X1   g00417(.A1(new_n1415_), .A2(new_n1420_), .ZN(new_n1421_));
  AOI21_X1   g00418(.A1(new_n1416_), .A2(new_n1418_), .B(new_n1417_), .ZN(new_n1422_));
  INV_X1     g00419(.I(\A[793] ), .ZN(new_n1423_));
  NOR2_X1    g00420(.A1(\A[794] ), .A2(\A[795] ), .ZN(new_n1424_));
  NAND2_X1   g00421(.A1(\A[794] ), .A2(\A[795] ), .ZN(new_n1425_));
  AOI21_X1   g00422(.A1(new_n1423_), .A2(new_n1425_), .B(new_n1424_), .ZN(new_n1426_));
  NOR2_X1    g00423(.A1(new_n1422_), .A2(new_n1426_), .ZN(new_n1427_));
  INV_X1     g00424(.I(\A[794] ), .ZN(new_n1428_));
  NAND2_X1   g00425(.A1(new_n1428_), .A2(\A[795] ), .ZN(new_n1429_));
  INV_X1     g00426(.I(\A[795] ), .ZN(new_n1430_));
  NAND2_X1   g00427(.A1(new_n1430_), .A2(\A[794] ), .ZN(new_n1431_));
  AOI21_X1   g00428(.A1(new_n1429_), .A2(new_n1431_), .B(new_n1423_), .ZN(new_n1432_));
  INV_X1     g00429(.I(new_n1424_), .ZN(new_n1433_));
  AOI21_X1   g00430(.A1(new_n1433_), .A2(new_n1425_), .B(\A[793] ), .ZN(new_n1434_));
  NOR2_X1    g00431(.A1(new_n1434_), .A2(new_n1432_), .ZN(new_n1435_));
  NAND2_X1   g00432(.A1(new_n1435_), .A2(new_n1427_), .ZN(new_n1436_));
  INV_X1     g00433(.I(new_n1427_), .ZN(new_n1437_));
  NOR2_X1    g00434(.A1(new_n1430_), .A2(\A[794] ), .ZN(new_n1438_));
  NOR2_X1    g00435(.A1(new_n1428_), .A2(\A[795] ), .ZN(new_n1439_));
  OAI21_X1   g00436(.A1(new_n1438_), .A2(new_n1439_), .B(\A[793] ), .ZN(new_n1440_));
  INV_X1     g00437(.I(new_n1425_), .ZN(new_n1441_));
  OAI21_X1   g00438(.A1(new_n1441_), .A2(new_n1424_), .B(new_n1423_), .ZN(new_n1442_));
  NAND2_X1   g00439(.A1(new_n1440_), .A2(new_n1442_), .ZN(new_n1443_));
  NAND2_X1   g00440(.A1(new_n1437_), .A2(new_n1443_), .ZN(new_n1444_));
  AOI21_X1   g00441(.A1(new_n1444_), .A2(new_n1436_), .B(new_n1421_), .ZN(new_n1445_));
  NAND2_X1   g00442(.A1(new_n1413_), .A2(\A[798] ), .ZN(new_n1446_));
  NAND2_X1   g00443(.A1(new_n1411_), .A2(\A[797] ), .ZN(new_n1447_));
  AOI21_X1   g00444(.A1(new_n1446_), .A2(new_n1447_), .B(new_n1416_), .ZN(new_n1448_));
  INV_X1     g00445(.I(new_n1417_), .ZN(new_n1449_));
  AOI21_X1   g00446(.A1(new_n1449_), .A2(new_n1418_), .B(\A[796] ), .ZN(new_n1450_));
  NOR2_X1    g00447(.A1(new_n1450_), .A2(new_n1448_), .ZN(new_n1451_));
  NOR2_X1    g00448(.A1(new_n1437_), .A2(new_n1443_), .ZN(new_n1452_));
  NOR2_X1    g00449(.A1(new_n1435_), .A2(new_n1427_), .ZN(new_n1453_));
  NOR3_X1    g00450(.A1(new_n1452_), .A2(new_n1453_), .A3(new_n1451_), .ZN(new_n1454_));
  NOR2_X1    g00451(.A1(new_n1454_), .A2(new_n1445_), .ZN(new_n1455_));
  NOR2_X1    g00452(.A1(new_n1376_), .A2(new_n1390_), .ZN(new_n1456_));
  NOR2_X1    g00453(.A1(new_n1407_), .A2(new_n1398_), .ZN(new_n1457_));
  NOR2_X1    g00454(.A1(new_n1421_), .A2(new_n1443_), .ZN(new_n1458_));
  NOR2_X1    g00455(.A1(new_n1451_), .A2(new_n1435_), .ZN(new_n1459_));
  NOR4_X1    g00456(.A1(new_n1456_), .A2(new_n1457_), .A3(new_n1459_), .A4(new_n1458_), .ZN(new_n1460_));
  NAND2_X1   g00457(.A1(new_n1422_), .A2(new_n1426_), .ZN(new_n1461_));
  INV_X1     g00458(.I(new_n1461_), .ZN(new_n1462_));
  NAND2_X1   g00459(.A1(new_n1458_), .A2(new_n1462_), .ZN(new_n1463_));
  NAND3_X1   g00460(.A1(new_n1407_), .A2(new_n1398_), .A3(new_n1382_), .ZN(new_n1464_));
  NAND3_X1   g00461(.A1(new_n1460_), .A2(new_n1463_), .A3(new_n1464_), .ZN(new_n1465_));
  XOR2_X1    g00462(.A1(new_n1465_), .A2(new_n1455_), .Z(new_n1466_));
  NAND2_X1   g00463(.A1(new_n1466_), .A2(new_n1410_), .ZN(new_n1467_));
  INV_X1     g00464(.I(new_n1467_), .ZN(new_n1468_));
  INV_X1     g00465(.I(\A[775] ), .ZN(new_n1469_));
  INV_X1     g00466(.I(\A[776] ), .ZN(new_n1470_));
  NAND2_X1   g00467(.A1(new_n1470_), .A2(\A[777] ), .ZN(new_n1471_));
  INV_X1     g00468(.I(\A[777] ), .ZN(new_n1472_));
  NAND2_X1   g00469(.A1(new_n1472_), .A2(\A[776] ), .ZN(new_n1473_));
  AOI21_X1   g00470(.A1(new_n1471_), .A2(new_n1473_), .B(new_n1469_), .ZN(new_n1474_));
  NOR2_X1    g00471(.A1(\A[776] ), .A2(\A[777] ), .ZN(new_n1475_));
  INV_X1     g00472(.I(new_n1475_), .ZN(new_n1476_));
  NAND2_X1   g00473(.A1(\A[776] ), .A2(\A[777] ), .ZN(new_n1477_));
  AOI21_X1   g00474(.A1(new_n1476_), .A2(new_n1477_), .B(\A[775] ), .ZN(new_n1478_));
  NOR2_X1    g00475(.A1(new_n1478_), .A2(new_n1474_), .ZN(new_n1479_));
  INV_X1     g00476(.I(\A[778] ), .ZN(new_n1480_));
  INV_X1     g00477(.I(\A[779] ), .ZN(new_n1481_));
  NAND2_X1   g00478(.A1(new_n1481_), .A2(\A[780] ), .ZN(new_n1482_));
  INV_X1     g00479(.I(\A[780] ), .ZN(new_n1483_));
  NAND2_X1   g00480(.A1(new_n1483_), .A2(\A[779] ), .ZN(new_n1484_));
  AOI21_X1   g00481(.A1(new_n1482_), .A2(new_n1484_), .B(new_n1480_), .ZN(new_n1485_));
  NOR2_X1    g00482(.A1(\A[779] ), .A2(\A[780] ), .ZN(new_n1486_));
  INV_X1     g00483(.I(new_n1486_), .ZN(new_n1487_));
  NAND2_X1   g00484(.A1(\A[779] ), .A2(\A[780] ), .ZN(new_n1488_));
  AOI21_X1   g00485(.A1(new_n1487_), .A2(new_n1488_), .B(\A[778] ), .ZN(new_n1489_));
  NOR2_X1    g00486(.A1(new_n1489_), .A2(new_n1485_), .ZN(new_n1490_));
  NOR2_X1    g00487(.A1(new_n1479_), .A2(new_n1490_), .ZN(new_n1491_));
  NOR2_X1    g00488(.A1(new_n1472_), .A2(\A[776] ), .ZN(new_n1492_));
  NOR2_X1    g00489(.A1(new_n1470_), .A2(\A[777] ), .ZN(new_n1493_));
  OAI21_X1   g00490(.A1(new_n1492_), .A2(new_n1493_), .B(\A[775] ), .ZN(new_n1494_));
  INV_X1     g00491(.I(new_n1477_), .ZN(new_n1495_));
  OAI21_X1   g00492(.A1(new_n1495_), .A2(new_n1475_), .B(new_n1469_), .ZN(new_n1496_));
  NAND2_X1   g00493(.A1(new_n1494_), .A2(new_n1496_), .ZN(new_n1497_));
  NOR2_X1    g00494(.A1(new_n1483_), .A2(\A[779] ), .ZN(new_n1498_));
  NOR2_X1    g00495(.A1(new_n1481_), .A2(\A[780] ), .ZN(new_n1499_));
  OAI21_X1   g00496(.A1(new_n1498_), .A2(new_n1499_), .B(\A[778] ), .ZN(new_n1500_));
  INV_X1     g00497(.I(new_n1488_), .ZN(new_n1501_));
  OAI21_X1   g00498(.A1(new_n1501_), .A2(new_n1486_), .B(new_n1480_), .ZN(new_n1502_));
  NAND2_X1   g00499(.A1(new_n1500_), .A2(new_n1502_), .ZN(new_n1503_));
  NOR2_X1    g00500(.A1(new_n1497_), .A2(new_n1503_), .ZN(new_n1504_));
  NOR2_X1    g00501(.A1(new_n1491_), .A2(new_n1504_), .ZN(new_n1505_));
  INV_X1     g00502(.I(\A[781] ), .ZN(new_n1506_));
  INV_X1     g00503(.I(\A[782] ), .ZN(new_n1507_));
  NAND2_X1   g00504(.A1(new_n1507_), .A2(\A[783] ), .ZN(new_n1508_));
  INV_X1     g00505(.I(\A[783] ), .ZN(new_n1509_));
  NAND2_X1   g00506(.A1(new_n1509_), .A2(\A[782] ), .ZN(new_n1510_));
  AOI21_X1   g00507(.A1(new_n1508_), .A2(new_n1510_), .B(new_n1506_), .ZN(new_n1511_));
  NOR2_X1    g00508(.A1(\A[782] ), .A2(\A[783] ), .ZN(new_n1512_));
  INV_X1     g00509(.I(new_n1512_), .ZN(new_n1513_));
  NAND2_X1   g00510(.A1(\A[782] ), .A2(\A[783] ), .ZN(new_n1514_));
  AOI21_X1   g00511(.A1(new_n1513_), .A2(new_n1514_), .B(\A[781] ), .ZN(new_n1515_));
  NOR2_X1    g00512(.A1(new_n1515_), .A2(new_n1511_), .ZN(new_n1516_));
  INV_X1     g00513(.I(\A[784] ), .ZN(new_n1517_));
  INV_X1     g00514(.I(\A[785] ), .ZN(new_n1518_));
  NAND2_X1   g00515(.A1(new_n1518_), .A2(\A[786] ), .ZN(new_n1519_));
  INV_X1     g00516(.I(\A[786] ), .ZN(new_n1520_));
  NAND2_X1   g00517(.A1(new_n1520_), .A2(\A[785] ), .ZN(new_n1521_));
  AOI21_X1   g00518(.A1(new_n1519_), .A2(new_n1521_), .B(new_n1517_), .ZN(new_n1522_));
  NOR2_X1    g00519(.A1(\A[785] ), .A2(\A[786] ), .ZN(new_n1523_));
  INV_X1     g00520(.I(new_n1523_), .ZN(new_n1524_));
  NAND2_X1   g00521(.A1(\A[785] ), .A2(\A[786] ), .ZN(new_n1525_));
  AOI21_X1   g00522(.A1(new_n1524_), .A2(new_n1525_), .B(\A[784] ), .ZN(new_n1526_));
  NOR2_X1    g00523(.A1(new_n1526_), .A2(new_n1522_), .ZN(new_n1527_));
  NAND2_X1   g00524(.A1(new_n1516_), .A2(new_n1527_), .ZN(new_n1528_));
  NOR2_X1    g00525(.A1(new_n1509_), .A2(\A[782] ), .ZN(new_n1529_));
  NOR2_X1    g00526(.A1(new_n1507_), .A2(\A[783] ), .ZN(new_n1530_));
  OAI21_X1   g00527(.A1(new_n1529_), .A2(new_n1530_), .B(\A[781] ), .ZN(new_n1531_));
  INV_X1     g00528(.I(new_n1514_), .ZN(new_n1532_));
  OAI21_X1   g00529(.A1(new_n1532_), .A2(new_n1512_), .B(new_n1506_), .ZN(new_n1533_));
  NAND2_X1   g00530(.A1(new_n1531_), .A2(new_n1533_), .ZN(new_n1534_));
  NOR2_X1    g00531(.A1(new_n1520_), .A2(\A[785] ), .ZN(new_n1535_));
  NOR2_X1    g00532(.A1(new_n1518_), .A2(\A[786] ), .ZN(new_n1536_));
  OAI21_X1   g00533(.A1(new_n1535_), .A2(new_n1536_), .B(\A[784] ), .ZN(new_n1537_));
  INV_X1     g00534(.I(new_n1525_), .ZN(new_n1538_));
  OAI21_X1   g00535(.A1(new_n1538_), .A2(new_n1523_), .B(new_n1517_), .ZN(new_n1539_));
  NAND2_X1   g00536(.A1(new_n1537_), .A2(new_n1539_), .ZN(new_n1540_));
  NAND2_X1   g00537(.A1(new_n1534_), .A2(new_n1540_), .ZN(new_n1541_));
  INV_X1     g00538(.I(new_n1528_), .ZN(new_n1542_));
  AOI21_X1   g00539(.A1(new_n1517_), .A2(new_n1525_), .B(new_n1523_), .ZN(new_n1543_));
  INV_X1     g00540(.I(new_n1543_), .ZN(new_n1544_));
  AOI21_X1   g00541(.A1(new_n1506_), .A2(new_n1514_), .B(new_n1512_), .ZN(new_n1545_));
  INV_X1     g00542(.I(new_n1545_), .ZN(new_n1546_));
  NOR2_X1    g00543(.A1(new_n1544_), .A2(new_n1546_), .ZN(new_n1547_));
  AOI21_X1   g00544(.A1(new_n1469_), .A2(new_n1477_), .B(new_n1475_), .ZN(new_n1548_));
  AOI21_X1   g00545(.A1(new_n1480_), .A2(new_n1488_), .B(new_n1486_), .ZN(new_n1549_));
  NOR2_X1    g00546(.A1(new_n1548_), .A2(new_n1549_), .ZN(new_n1550_));
  INV_X1     g00547(.I(new_n1550_), .ZN(new_n1551_));
  NOR3_X1    g00548(.A1(new_n1551_), .A2(new_n1479_), .A3(new_n1490_), .ZN(new_n1552_));
  AOI21_X1   g00549(.A1(new_n1542_), .A2(new_n1547_), .B(new_n1552_), .ZN(new_n1553_));
  NAND4_X1   g00550(.A1(new_n1553_), .A2(new_n1505_), .A3(new_n1528_), .A4(new_n1541_), .ZN(new_n1554_));
  NOR2_X1    g00551(.A1(new_n1543_), .A2(new_n1545_), .ZN(new_n1555_));
  NAND2_X1   g00552(.A1(new_n1516_), .A2(new_n1555_), .ZN(new_n1556_));
  INV_X1     g00553(.I(new_n1555_), .ZN(new_n1557_));
  NAND2_X1   g00554(.A1(new_n1557_), .A2(new_n1534_), .ZN(new_n1558_));
  AOI21_X1   g00555(.A1(new_n1558_), .A2(new_n1556_), .B(new_n1540_), .ZN(new_n1559_));
  NAND3_X1   g00556(.A1(new_n1558_), .A2(new_n1556_), .A3(new_n1540_), .ZN(new_n1560_));
  INV_X1     g00557(.I(new_n1560_), .ZN(new_n1561_));
  NOR2_X1    g00558(.A1(new_n1561_), .A2(new_n1559_), .ZN(new_n1562_));
  NAND2_X1   g00559(.A1(new_n1479_), .A2(new_n1550_), .ZN(new_n1563_));
  NAND2_X1   g00560(.A1(new_n1551_), .A2(new_n1497_), .ZN(new_n1564_));
  NAND2_X1   g00561(.A1(new_n1564_), .A2(new_n1563_), .ZN(new_n1565_));
  NAND2_X1   g00562(.A1(new_n1565_), .A2(new_n1490_), .ZN(new_n1566_));
  NAND3_X1   g00563(.A1(new_n1564_), .A2(new_n1563_), .A3(new_n1503_), .ZN(new_n1567_));
  NAND2_X1   g00564(.A1(new_n1566_), .A2(new_n1567_), .ZN(new_n1568_));
  XNOR2_X1   g00565(.A1(new_n1543_), .A2(new_n1545_), .ZN(new_n1569_));
  OAI21_X1   g00566(.A1(new_n1547_), .A2(new_n1555_), .B(new_n1528_), .ZN(new_n1570_));
  OAI21_X1   g00567(.A1(new_n1528_), .A2(new_n1569_), .B(new_n1570_), .ZN(new_n1571_));
  NAND3_X1   g00568(.A1(new_n1505_), .A2(new_n1528_), .A3(new_n1541_), .ZN(new_n1572_));
  INV_X1     g00569(.I(new_n1547_), .ZN(new_n1573_));
  NAND4_X1   g00570(.A1(new_n1552_), .A2(new_n1534_), .A3(new_n1540_), .A4(new_n1573_), .ZN(new_n1574_));
  NOR2_X1    g00571(.A1(new_n1572_), .A2(new_n1574_), .ZN(new_n1575_));
  NAND2_X1   g00572(.A1(new_n1575_), .A2(new_n1571_), .ZN(new_n1576_));
  NAND4_X1   g00573(.A1(new_n1576_), .A2(new_n1554_), .A3(new_n1562_), .A4(new_n1568_), .ZN(new_n1577_));
  NAND3_X1   g00574(.A1(new_n1497_), .A2(new_n1503_), .A3(new_n1550_), .ZN(new_n1578_));
  NAND2_X1   g00575(.A1(new_n1505_), .A2(new_n1578_), .ZN(new_n1579_));
  NOR2_X1    g00576(.A1(new_n1456_), .A2(new_n1457_), .ZN(new_n1580_));
  NAND2_X1   g00577(.A1(new_n1580_), .A2(new_n1464_), .ZN(new_n1581_));
  XOR2_X1    g00578(.A1(new_n1579_), .A2(new_n1581_), .Z(new_n1582_));
  NOR2_X1    g00579(.A1(new_n1459_), .A2(new_n1458_), .ZN(new_n1583_));
  NAND2_X1   g00580(.A1(new_n1528_), .A2(new_n1541_), .ZN(new_n1584_));
  XOR2_X1    g00581(.A1(new_n1583_), .A2(new_n1584_), .Z(new_n1585_));
  INV_X1     g00582(.I(new_n1585_), .ZN(new_n1586_));
  NAND2_X1   g00583(.A1(new_n1582_), .A2(new_n1586_), .ZN(new_n1587_));
  NOR2_X1    g00584(.A1(new_n1587_), .A2(new_n1577_), .ZN(new_n1588_));
  OR2_X2     g00585(.A1(new_n1454_), .A2(new_n1445_), .Z(new_n1589_));
  NOR2_X1    g00586(.A1(new_n1459_), .A2(new_n1458_), .ZN(new_n1590_));
  AND4_X2    g00587(.A1(new_n1580_), .A2(new_n1590_), .A3(new_n1463_), .A4(new_n1464_), .Z(new_n1591_));
  XOR2_X1    g00588(.A1(new_n1422_), .A2(new_n1426_), .Z(new_n1592_));
  NAND2_X1   g00589(.A1(new_n1458_), .A2(new_n1592_), .ZN(new_n1593_));
  NOR2_X1    g00590(.A1(new_n1462_), .A2(new_n1427_), .ZN(new_n1594_));
  OAI21_X1   g00591(.A1(new_n1458_), .A2(new_n1594_), .B(new_n1593_), .ZN(new_n1595_));
  NAND2_X1   g00592(.A1(new_n1459_), .A2(new_n1461_), .ZN(new_n1596_));
  NOR2_X1    g00593(.A1(new_n1596_), .A2(new_n1464_), .ZN(new_n1597_));
  NAND3_X1   g00594(.A1(new_n1595_), .A2(new_n1460_), .A3(new_n1597_), .ZN(new_n1598_));
  NOR2_X1    g00595(.A1(new_n1410_), .A2(new_n1598_), .ZN(new_n1599_));
  OAI21_X1   g00596(.A1(new_n1599_), .A2(new_n1589_), .B(new_n1591_), .ZN(new_n1600_));
  NAND2_X1   g00597(.A1(new_n1588_), .A2(new_n1600_), .ZN(new_n1601_));
  INV_X1     g00598(.I(new_n1601_), .ZN(new_n1602_));
  NOR2_X1    g00599(.A1(new_n1588_), .A2(new_n1600_), .ZN(new_n1603_));
  OAI21_X1   g00600(.A1(new_n1602_), .A2(new_n1603_), .B(new_n1468_), .ZN(new_n1604_));
  INV_X1     g00601(.I(new_n1579_), .ZN(new_n1605_));
  XNOR2_X1   g00602(.A1(new_n1581_), .A2(new_n1583_), .ZN(new_n1606_));
  NAND2_X1   g00603(.A1(new_n1606_), .A2(new_n1584_), .ZN(new_n1607_));
  INV_X1     g00604(.I(new_n1584_), .ZN(new_n1608_));
  XOR2_X1    g00605(.A1(new_n1581_), .A2(new_n1583_), .Z(new_n1609_));
  NAND2_X1   g00606(.A1(new_n1609_), .A2(new_n1608_), .ZN(new_n1610_));
  AOI21_X1   g00607(.A1(new_n1607_), .A2(new_n1610_), .B(new_n1605_), .ZN(new_n1611_));
  NAND3_X1   g00608(.A1(new_n1607_), .A2(new_n1610_), .A3(new_n1605_), .ZN(new_n1612_));
  INV_X1     g00609(.I(new_n1612_), .ZN(new_n1613_));
  INV_X1     g00610(.I(\A[771] ), .ZN(new_n1614_));
  NOR2_X1    g00611(.A1(new_n1614_), .A2(\A[770] ), .ZN(new_n1615_));
  INV_X1     g00612(.I(\A[770] ), .ZN(new_n1616_));
  NOR2_X1    g00613(.A1(new_n1616_), .A2(\A[771] ), .ZN(new_n1617_));
  OAI21_X1   g00614(.A1(new_n1615_), .A2(new_n1617_), .B(\A[769] ), .ZN(new_n1618_));
  INV_X1     g00615(.I(\A[769] ), .ZN(new_n1619_));
  NAND2_X1   g00616(.A1(\A[770] ), .A2(\A[771] ), .ZN(new_n1620_));
  INV_X1     g00617(.I(new_n1620_), .ZN(new_n1621_));
  NOR2_X1    g00618(.A1(\A[770] ), .A2(\A[771] ), .ZN(new_n1622_));
  OAI21_X1   g00619(.A1(new_n1621_), .A2(new_n1622_), .B(new_n1619_), .ZN(new_n1623_));
  NAND2_X1   g00620(.A1(new_n1618_), .A2(new_n1623_), .ZN(new_n1624_));
  INV_X1     g00621(.I(\A[774] ), .ZN(new_n1625_));
  NOR2_X1    g00622(.A1(new_n1625_), .A2(\A[773] ), .ZN(new_n1626_));
  INV_X1     g00623(.I(\A[773] ), .ZN(new_n1627_));
  NOR2_X1    g00624(.A1(new_n1627_), .A2(\A[774] ), .ZN(new_n1628_));
  OAI21_X1   g00625(.A1(new_n1626_), .A2(new_n1628_), .B(\A[772] ), .ZN(new_n1629_));
  INV_X1     g00626(.I(\A[772] ), .ZN(new_n1630_));
  NAND2_X1   g00627(.A1(\A[773] ), .A2(\A[774] ), .ZN(new_n1631_));
  INV_X1     g00628(.I(new_n1631_), .ZN(new_n1632_));
  NOR2_X1    g00629(.A1(\A[773] ), .A2(\A[774] ), .ZN(new_n1633_));
  OAI21_X1   g00630(.A1(new_n1632_), .A2(new_n1633_), .B(new_n1630_), .ZN(new_n1634_));
  NAND2_X1   g00631(.A1(new_n1629_), .A2(new_n1634_), .ZN(new_n1635_));
  AOI21_X1   g00632(.A1(new_n1619_), .A2(new_n1620_), .B(new_n1622_), .ZN(new_n1636_));
  AOI21_X1   g00633(.A1(new_n1630_), .A2(new_n1631_), .B(new_n1633_), .ZN(new_n1637_));
  NOR2_X1    g00634(.A1(new_n1636_), .A2(new_n1637_), .ZN(new_n1638_));
  NAND3_X1   g00635(.A1(new_n1624_), .A2(new_n1635_), .A3(new_n1638_), .ZN(new_n1639_));
  INV_X1     g00636(.I(\A[763] ), .ZN(new_n1640_));
  INV_X1     g00637(.I(\A[764] ), .ZN(new_n1641_));
  NAND2_X1   g00638(.A1(new_n1641_), .A2(\A[765] ), .ZN(new_n1642_));
  INV_X1     g00639(.I(\A[765] ), .ZN(new_n1643_));
  NAND2_X1   g00640(.A1(new_n1643_), .A2(\A[764] ), .ZN(new_n1644_));
  AOI21_X1   g00641(.A1(new_n1642_), .A2(new_n1644_), .B(new_n1640_), .ZN(new_n1645_));
  NAND2_X1   g00642(.A1(\A[764] ), .A2(\A[765] ), .ZN(new_n1646_));
  NAND2_X1   g00643(.A1(new_n1641_), .A2(new_n1643_), .ZN(new_n1647_));
  AOI21_X1   g00644(.A1(new_n1647_), .A2(new_n1646_), .B(\A[763] ), .ZN(new_n1648_));
  NOR2_X1    g00645(.A1(new_n1648_), .A2(new_n1645_), .ZN(new_n1649_));
  INV_X1     g00646(.I(\A[766] ), .ZN(new_n1650_));
  INV_X1     g00647(.I(\A[767] ), .ZN(new_n1651_));
  NAND2_X1   g00648(.A1(new_n1651_), .A2(\A[768] ), .ZN(new_n1652_));
  INV_X1     g00649(.I(\A[768] ), .ZN(new_n1653_));
  NAND2_X1   g00650(.A1(new_n1653_), .A2(\A[767] ), .ZN(new_n1654_));
  AOI21_X1   g00651(.A1(new_n1652_), .A2(new_n1654_), .B(new_n1650_), .ZN(new_n1655_));
  NAND2_X1   g00652(.A1(\A[767] ), .A2(\A[768] ), .ZN(new_n1656_));
  NAND2_X1   g00653(.A1(new_n1651_), .A2(new_n1653_), .ZN(new_n1657_));
  AOI21_X1   g00654(.A1(new_n1657_), .A2(new_n1656_), .B(\A[766] ), .ZN(new_n1658_));
  NOR2_X1    g00655(.A1(new_n1658_), .A2(new_n1655_), .ZN(new_n1659_));
  NAND2_X1   g00656(.A1(new_n1646_), .A2(new_n1640_), .ZN(new_n1660_));
  NAND2_X1   g00657(.A1(new_n1660_), .A2(new_n1647_), .ZN(new_n1661_));
  NAND2_X1   g00658(.A1(new_n1656_), .A2(new_n1650_), .ZN(new_n1662_));
  NAND2_X1   g00659(.A1(new_n1662_), .A2(new_n1657_), .ZN(new_n1663_));
  NAND2_X1   g00660(.A1(new_n1661_), .A2(new_n1663_), .ZN(new_n1664_));
  NOR3_X1    g00661(.A1(new_n1649_), .A2(new_n1659_), .A3(new_n1664_), .ZN(new_n1665_));
  XOR2_X1    g00662(.A1(new_n1665_), .A2(new_n1639_), .Z(new_n1666_));
  INV_X1     g00663(.I(\A[759] ), .ZN(new_n1667_));
  NOR2_X1    g00664(.A1(new_n1667_), .A2(\A[758] ), .ZN(new_n1668_));
  INV_X1     g00665(.I(\A[758] ), .ZN(new_n1669_));
  NOR2_X1    g00666(.A1(new_n1669_), .A2(\A[759] ), .ZN(new_n1670_));
  OAI21_X1   g00667(.A1(new_n1668_), .A2(new_n1670_), .B(\A[757] ), .ZN(new_n1671_));
  INV_X1     g00668(.I(\A[757] ), .ZN(new_n1672_));
  NOR2_X1    g00669(.A1(new_n1669_), .A2(new_n1667_), .ZN(new_n1673_));
  NOR2_X1    g00670(.A1(\A[758] ), .A2(\A[759] ), .ZN(new_n1674_));
  OAI21_X1   g00671(.A1(new_n1673_), .A2(new_n1674_), .B(new_n1672_), .ZN(new_n1675_));
  NAND2_X1   g00672(.A1(new_n1675_), .A2(new_n1671_), .ZN(new_n1676_));
  INV_X1     g00673(.I(\A[762] ), .ZN(new_n1677_));
  NOR2_X1    g00674(.A1(new_n1677_), .A2(\A[761] ), .ZN(new_n1678_));
  INV_X1     g00675(.I(\A[761] ), .ZN(new_n1679_));
  NOR2_X1    g00676(.A1(new_n1679_), .A2(\A[762] ), .ZN(new_n1680_));
  OAI21_X1   g00677(.A1(new_n1678_), .A2(new_n1680_), .B(\A[760] ), .ZN(new_n1681_));
  INV_X1     g00678(.I(\A[760] ), .ZN(new_n1682_));
  NOR2_X1    g00679(.A1(new_n1679_), .A2(new_n1677_), .ZN(new_n1683_));
  NOR2_X1    g00680(.A1(\A[761] ), .A2(\A[762] ), .ZN(new_n1684_));
  OAI21_X1   g00681(.A1(new_n1683_), .A2(new_n1684_), .B(new_n1682_), .ZN(new_n1685_));
  NAND2_X1   g00682(.A1(new_n1685_), .A2(new_n1681_), .ZN(new_n1686_));
  INV_X1     g00683(.I(new_n1674_), .ZN(new_n1687_));
  OAI21_X1   g00684(.A1(\A[757] ), .A2(new_n1673_), .B(new_n1687_), .ZN(new_n1688_));
  INV_X1     g00685(.I(new_n1684_), .ZN(new_n1689_));
  OAI21_X1   g00686(.A1(\A[760] ), .A2(new_n1683_), .B(new_n1689_), .ZN(new_n1690_));
  NAND2_X1   g00687(.A1(new_n1688_), .A2(new_n1690_), .ZN(new_n1691_));
  INV_X1     g00688(.I(new_n1691_), .ZN(new_n1692_));
  NAND3_X1   g00689(.A1(new_n1692_), .A2(new_n1676_), .A3(new_n1686_), .ZN(new_n1693_));
  INV_X1     g00690(.I(\A[751] ), .ZN(new_n1694_));
  INV_X1     g00691(.I(\A[752] ), .ZN(new_n1695_));
  NAND2_X1   g00692(.A1(new_n1695_), .A2(\A[753] ), .ZN(new_n1696_));
  INV_X1     g00693(.I(\A[753] ), .ZN(new_n1697_));
  NAND2_X1   g00694(.A1(new_n1697_), .A2(\A[752] ), .ZN(new_n1698_));
  AOI21_X1   g00695(.A1(new_n1696_), .A2(new_n1698_), .B(new_n1694_), .ZN(new_n1699_));
  NAND2_X1   g00696(.A1(\A[752] ), .A2(\A[753] ), .ZN(new_n1700_));
  NAND2_X1   g00697(.A1(new_n1695_), .A2(new_n1697_), .ZN(new_n1701_));
  AOI21_X1   g00698(.A1(new_n1701_), .A2(new_n1700_), .B(\A[751] ), .ZN(new_n1702_));
  NOR2_X1    g00699(.A1(new_n1702_), .A2(new_n1699_), .ZN(new_n1703_));
  INV_X1     g00700(.I(\A[754] ), .ZN(new_n1704_));
  INV_X1     g00701(.I(\A[755] ), .ZN(new_n1705_));
  NAND2_X1   g00702(.A1(new_n1705_), .A2(\A[756] ), .ZN(new_n1706_));
  INV_X1     g00703(.I(\A[756] ), .ZN(new_n1707_));
  NAND2_X1   g00704(.A1(new_n1707_), .A2(\A[755] ), .ZN(new_n1708_));
  AOI21_X1   g00705(.A1(new_n1706_), .A2(new_n1708_), .B(new_n1704_), .ZN(new_n1709_));
  NAND2_X1   g00706(.A1(\A[755] ), .A2(\A[756] ), .ZN(new_n1710_));
  NAND2_X1   g00707(.A1(new_n1705_), .A2(new_n1707_), .ZN(new_n1711_));
  AOI21_X1   g00708(.A1(new_n1711_), .A2(new_n1710_), .B(\A[754] ), .ZN(new_n1712_));
  NOR2_X1    g00709(.A1(new_n1712_), .A2(new_n1709_), .ZN(new_n1713_));
  NAND2_X1   g00710(.A1(new_n1700_), .A2(new_n1694_), .ZN(new_n1714_));
  NAND2_X1   g00711(.A1(new_n1714_), .A2(new_n1701_), .ZN(new_n1715_));
  NAND2_X1   g00712(.A1(new_n1710_), .A2(new_n1704_), .ZN(new_n1716_));
  NAND2_X1   g00713(.A1(new_n1716_), .A2(new_n1711_), .ZN(new_n1717_));
  NAND2_X1   g00714(.A1(new_n1715_), .A2(new_n1717_), .ZN(new_n1718_));
  NOR3_X1    g00715(.A1(new_n1703_), .A2(new_n1713_), .A3(new_n1718_), .ZN(new_n1719_));
  XOR2_X1    g00716(.A1(new_n1693_), .A2(new_n1719_), .Z(new_n1720_));
  NOR2_X1    g00717(.A1(new_n1720_), .A2(new_n1666_), .ZN(new_n1721_));
  NAND2_X1   g00718(.A1(new_n1720_), .A2(new_n1666_), .ZN(new_n1722_));
  INV_X1     g00719(.I(new_n1722_), .ZN(new_n1723_));
  NOR4_X1    g00720(.A1(new_n1613_), .A2(new_n1611_), .A3(new_n1721_), .A4(new_n1723_), .ZN(new_n1724_));
  NAND3_X1   g00721(.A1(new_n1649_), .A2(new_n1661_), .A3(new_n1663_), .ZN(new_n1725_));
  OR2_X2     g00722(.A1(new_n1648_), .A2(new_n1645_), .Z(new_n1726_));
  NAND2_X1   g00723(.A1(new_n1726_), .A2(new_n1664_), .ZN(new_n1727_));
  NAND2_X1   g00724(.A1(new_n1727_), .A2(new_n1725_), .ZN(new_n1728_));
  NAND2_X1   g00725(.A1(new_n1728_), .A2(new_n1659_), .ZN(new_n1729_));
  OR2_X2     g00726(.A1(new_n1658_), .A2(new_n1655_), .Z(new_n1730_));
  NAND3_X1   g00727(.A1(new_n1727_), .A2(new_n1730_), .A3(new_n1725_), .ZN(new_n1731_));
  NAND2_X1   g00728(.A1(new_n1729_), .A2(new_n1731_), .ZN(new_n1732_));
  INV_X1     g00729(.I(new_n1732_), .ZN(new_n1733_));
  NOR4_X1    g00730(.A1(new_n1639_), .A2(new_n1649_), .A3(new_n1659_), .A4(new_n1664_), .ZN(new_n1734_));
  INV_X1     g00731(.I(new_n1635_), .ZN(new_n1735_));
  INV_X1     g00732(.I(new_n1638_), .ZN(new_n1736_));
  NOR2_X1    g00733(.A1(new_n1736_), .A2(new_n1624_), .ZN(new_n1737_));
  NAND2_X1   g00734(.A1(new_n1616_), .A2(\A[771] ), .ZN(new_n1738_));
  NAND2_X1   g00735(.A1(new_n1614_), .A2(\A[770] ), .ZN(new_n1739_));
  AOI21_X1   g00736(.A1(new_n1738_), .A2(new_n1739_), .B(new_n1619_), .ZN(new_n1740_));
  INV_X1     g00737(.I(new_n1622_), .ZN(new_n1741_));
  AOI21_X1   g00738(.A1(new_n1741_), .A2(new_n1620_), .B(\A[769] ), .ZN(new_n1742_));
  NOR2_X1    g00739(.A1(new_n1742_), .A2(new_n1740_), .ZN(new_n1743_));
  NOR2_X1    g00740(.A1(new_n1743_), .A2(new_n1638_), .ZN(new_n1744_));
  OAI21_X1   g00741(.A1(new_n1737_), .A2(new_n1744_), .B(new_n1735_), .ZN(new_n1745_));
  NAND2_X1   g00742(.A1(new_n1743_), .A2(new_n1638_), .ZN(new_n1746_));
  NAND2_X1   g00743(.A1(new_n1736_), .A2(new_n1624_), .ZN(new_n1747_));
  NAND3_X1   g00744(.A1(new_n1747_), .A2(new_n1746_), .A3(new_n1635_), .ZN(new_n1748_));
  NAND2_X1   g00745(.A1(new_n1745_), .A2(new_n1748_), .ZN(new_n1749_));
  XOR2_X1    g00746(.A1(new_n1743_), .A2(new_n1635_), .Z(new_n1750_));
  NOR2_X1    g00747(.A1(new_n1750_), .A2(new_n1736_), .ZN(new_n1751_));
  NOR2_X1    g00748(.A1(new_n1751_), .A2(new_n1749_), .ZN(new_n1752_));
  XOR2_X1    g00749(.A1(new_n1752_), .A2(new_n1734_), .Z(new_n1753_));
  NAND2_X1   g00750(.A1(new_n1753_), .A2(new_n1733_), .ZN(new_n1754_));
  INV_X1     g00751(.I(new_n1752_), .ZN(new_n1755_));
  NOR2_X1    g00752(.A1(new_n1649_), .A2(new_n1659_), .ZN(new_n1756_));
  NOR2_X1    g00753(.A1(new_n1726_), .A2(new_n1730_), .ZN(new_n1757_));
  NOR2_X1    g00754(.A1(new_n1757_), .A2(new_n1756_), .ZN(new_n1758_));
  NOR3_X1    g00755(.A1(new_n1649_), .A2(new_n1659_), .A3(new_n1664_), .ZN(new_n1759_));
  NOR4_X1    g00756(.A1(new_n1751_), .A2(new_n1639_), .A3(new_n1758_), .A4(new_n1759_), .ZN(new_n1760_));
  NAND3_X1   g00757(.A1(new_n1760_), .A2(new_n1732_), .A3(new_n1749_), .ZN(new_n1761_));
  NAND2_X1   g00758(.A1(new_n1761_), .A2(new_n1755_), .ZN(new_n1762_));
  NOR4_X1    g00759(.A1(new_n1693_), .A2(new_n1703_), .A3(new_n1713_), .A4(new_n1718_), .ZN(new_n1763_));
  XOR2_X1    g00760(.A1(new_n1691_), .A2(new_n1676_), .Z(new_n1764_));
  NOR2_X1    g00761(.A1(new_n1764_), .A2(new_n1686_), .ZN(new_n1765_));
  INV_X1     g00762(.I(new_n1686_), .ZN(new_n1766_));
  XNOR2_X1   g00763(.A1(new_n1691_), .A2(new_n1676_), .ZN(new_n1767_));
  NOR2_X1    g00764(.A1(new_n1767_), .A2(new_n1766_), .ZN(new_n1768_));
  XNOR2_X1   g00765(.A1(new_n1676_), .A2(new_n1686_), .ZN(new_n1769_));
  NOR2_X1    g00766(.A1(new_n1769_), .A2(new_n1691_), .ZN(new_n1770_));
  NOR3_X1    g00767(.A1(new_n1768_), .A2(new_n1770_), .A3(new_n1765_), .ZN(new_n1771_));
  XOR2_X1    g00768(.A1(new_n1703_), .A2(new_n1718_), .Z(new_n1772_));
  XOR2_X1    g00769(.A1(new_n1772_), .A2(new_n1713_), .Z(new_n1773_));
  INV_X1     g00770(.I(new_n1676_), .ZN(new_n1774_));
  NOR2_X1    g00771(.A1(new_n1703_), .A2(new_n1713_), .ZN(new_n1775_));
  OR2_X2     g00772(.A1(new_n1702_), .A2(new_n1699_), .Z(new_n1776_));
  OR2_X2     g00773(.A1(new_n1712_), .A2(new_n1709_), .Z(new_n1777_));
  NOR2_X1    g00774(.A1(new_n1776_), .A2(new_n1777_), .ZN(new_n1778_));
  NAND3_X1   g00775(.A1(new_n1776_), .A2(new_n1715_), .A3(new_n1717_), .ZN(new_n1779_));
  OAI22_X1   g00776(.A1(new_n1775_), .A2(new_n1778_), .B1(new_n1779_), .B2(new_n1713_), .ZN(new_n1780_));
  NOR4_X1    g00777(.A1(new_n1780_), .A2(new_n1774_), .A3(new_n1766_), .A4(new_n1691_), .ZN(new_n1781_));
  NOR4_X1    g00778(.A1(new_n1771_), .A2(new_n1773_), .A3(new_n1763_), .A4(new_n1781_), .ZN(new_n1782_));
  NAND2_X1   g00779(.A1(new_n1782_), .A2(new_n1723_), .ZN(new_n1783_));
  AOI21_X1   g00780(.A1(new_n1734_), .A2(new_n1762_), .B(new_n1783_), .ZN(new_n1784_));
  NOR2_X1    g00781(.A1(new_n1758_), .A2(new_n1759_), .ZN(new_n1785_));
  NAND4_X1   g00782(.A1(new_n1785_), .A2(new_n1624_), .A3(new_n1635_), .A4(new_n1638_), .ZN(new_n1786_));
  NOR2_X1    g00783(.A1(new_n1733_), .A2(new_n1786_), .ZN(new_n1787_));
  OAI21_X1   g00784(.A1(new_n1787_), .A2(new_n1752_), .B(new_n1734_), .ZN(new_n1788_));
  INV_X1     g00785(.I(new_n1763_), .ZN(new_n1789_));
  NAND2_X1   g00786(.A1(new_n1767_), .A2(new_n1766_), .ZN(new_n1790_));
  NAND2_X1   g00787(.A1(new_n1764_), .A2(new_n1686_), .ZN(new_n1791_));
  XOR2_X1    g00788(.A1(new_n1676_), .A2(new_n1686_), .Z(new_n1792_));
  NAND2_X1   g00789(.A1(new_n1792_), .A2(new_n1692_), .ZN(new_n1793_));
  NAND3_X1   g00790(.A1(new_n1790_), .A2(new_n1791_), .A3(new_n1793_), .ZN(new_n1794_));
  NAND2_X1   g00791(.A1(new_n1772_), .A2(new_n1713_), .ZN(new_n1795_));
  XNOR2_X1   g00792(.A1(new_n1703_), .A2(new_n1718_), .ZN(new_n1796_));
  NAND2_X1   g00793(.A1(new_n1796_), .A2(new_n1777_), .ZN(new_n1797_));
  NAND2_X1   g00794(.A1(new_n1797_), .A2(new_n1795_), .ZN(new_n1798_));
  NOR2_X1    g00795(.A1(new_n1778_), .A2(new_n1775_), .ZN(new_n1799_));
  NOR3_X1    g00796(.A1(new_n1703_), .A2(new_n1713_), .A3(new_n1718_), .ZN(new_n1800_));
  NOR2_X1    g00797(.A1(new_n1799_), .A2(new_n1800_), .ZN(new_n1801_));
  NAND4_X1   g00798(.A1(new_n1801_), .A2(new_n1676_), .A3(new_n1686_), .A4(new_n1692_), .ZN(new_n1802_));
  NAND4_X1   g00799(.A1(new_n1802_), .A2(new_n1794_), .A3(new_n1789_), .A4(new_n1798_), .ZN(new_n1803_));
  NOR2_X1    g00800(.A1(new_n1803_), .A2(new_n1722_), .ZN(new_n1804_));
  NOR2_X1    g00801(.A1(new_n1804_), .A2(new_n1788_), .ZN(new_n1805_));
  OAI21_X1   g00802(.A1(new_n1784_), .A2(new_n1805_), .B(new_n1754_), .ZN(new_n1806_));
  INV_X1     g00803(.I(new_n1754_), .ZN(new_n1807_));
  NAND2_X1   g00804(.A1(new_n1804_), .A2(new_n1788_), .ZN(new_n1808_));
  NAND3_X1   g00805(.A1(new_n1783_), .A2(new_n1734_), .A3(new_n1762_), .ZN(new_n1809_));
  NAND3_X1   g00806(.A1(new_n1807_), .A2(new_n1809_), .A3(new_n1808_), .ZN(new_n1810_));
  NAND2_X1   g00807(.A1(new_n1806_), .A2(new_n1810_), .ZN(new_n1811_));
  NAND3_X1   g00808(.A1(new_n1811_), .A2(new_n1604_), .A3(new_n1724_), .ZN(new_n1812_));
  INV_X1     g00809(.I(new_n1603_), .ZN(new_n1813_));
  AOI21_X1   g00810(.A1(new_n1813_), .A2(new_n1601_), .B(new_n1467_), .ZN(new_n1814_));
  NAND3_X1   g00811(.A1(new_n1811_), .A2(new_n1814_), .A3(new_n1724_), .ZN(new_n1815_));
  INV_X1     g00812(.I(new_n1611_), .ZN(new_n1816_));
  NOR2_X1    g00813(.A1(new_n1723_), .A2(new_n1721_), .ZN(new_n1817_));
  AOI21_X1   g00814(.A1(new_n1816_), .A2(new_n1612_), .B(new_n1817_), .ZN(new_n1818_));
  NOR2_X1    g00815(.A1(new_n1177_), .A2(new_n1178_), .ZN(new_n1819_));
  XOR2_X1    g00816(.A1(new_n1819_), .A2(new_n1289_), .Z(new_n1820_));
  NOR3_X1    g00817(.A1(new_n1724_), .A2(new_n1818_), .A3(new_n1820_), .ZN(new_n1821_));
  INV_X1     g00818(.I(new_n1821_), .ZN(new_n1822_));
  AOI21_X1   g00819(.A1(new_n1812_), .A2(new_n1815_), .B(new_n1822_), .ZN(new_n1823_));
  NOR3_X1    g00820(.A1(new_n1823_), .A2(new_n1175_), .A3(new_n1365_), .ZN(new_n1824_));
  INV_X1     g00821(.I(new_n1824_), .ZN(new_n1825_));
  INV_X1     g00822(.I(\A[739] ), .ZN(new_n1826_));
  INV_X1     g00823(.I(\A[740] ), .ZN(new_n1827_));
  NAND2_X1   g00824(.A1(new_n1827_), .A2(\A[741] ), .ZN(new_n1828_));
  INV_X1     g00825(.I(\A[741] ), .ZN(new_n1829_));
  NAND2_X1   g00826(.A1(new_n1829_), .A2(\A[740] ), .ZN(new_n1830_));
  AOI21_X1   g00827(.A1(new_n1828_), .A2(new_n1830_), .B(new_n1826_), .ZN(new_n1831_));
  NAND2_X1   g00828(.A1(\A[740] ), .A2(\A[741] ), .ZN(new_n1832_));
  NAND2_X1   g00829(.A1(new_n1827_), .A2(new_n1829_), .ZN(new_n1833_));
  AOI21_X1   g00830(.A1(new_n1833_), .A2(new_n1832_), .B(\A[739] ), .ZN(new_n1834_));
  NOR2_X1    g00831(.A1(new_n1834_), .A2(new_n1831_), .ZN(new_n1835_));
  INV_X1     g00832(.I(\A[742] ), .ZN(new_n1836_));
  INV_X1     g00833(.I(\A[743] ), .ZN(new_n1837_));
  NAND2_X1   g00834(.A1(new_n1837_), .A2(\A[744] ), .ZN(new_n1838_));
  INV_X1     g00835(.I(\A[744] ), .ZN(new_n1839_));
  NAND2_X1   g00836(.A1(new_n1839_), .A2(\A[743] ), .ZN(new_n1840_));
  AOI21_X1   g00837(.A1(new_n1838_), .A2(new_n1840_), .B(new_n1836_), .ZN(new_n1841_));
  NAND2_X1   g00838(.A1(\A[743] ), .A2(\A[744] ), .ZN(new_n1842_));
  NAND2_X1   g00839(.A1(new_n1837_), .A2(new_n1839_), .ZN(new_n1843_));
  AOI21_X1   g00840(.A1(new_n1843_), .A2(new_n1842_), .B(\A[742] ), .ZN(new_n1844_));
  NOR2_X1    g00841(.A1(new_n1844_), .A2(new_n1841_), .ZN(new_n1845_));
  NAND2_X1   g00842(.A1(new_n1832_), .A2(new_n1826_), .ZN(new_n1846_));
  NAND2_X1   g00843(.A1(new_n1846_), .A2(new_n1833_), .ZN(new_n1847_));
  NAND2_X1   g00844(.A1(new_n1842_), .A2(new_n1836_), .ZN(new_n1848_));
  NAND2_X1   g00845(.A1(new_n1848_), .A2(new_n1843_), .ZN(new_n1849_));
  NAND2_X1   g00846(.A1(new_n1847_), .A2(new_n1849_), .ZN(new_n1850_));
  NOR3_X1    g00847(.A1(new_n1835_), .A2(new_n1845_), .A3(new_n1850_), .ZN(new_n1851_));
  INV_X1     g00848(.I(\A[745] ), .ZN(new_n1852_));
  INV_X1     g00849(.I(\A[746] ), .ZN(new_n1853_));
  NAND2_X1   g00850(.A1(new_n1853_), .A2(\A[747] ), .ZN(new_n1854_));
  INV_X1     g00851(.I(\A[747] ), .ZN(new_n1855_));
  NAND2_X1   g00852(.A1(new_n1855_), .A2(\A[746] ), .ZN(new_n1856_));
  AOI21_X1   g00853(.A1(new_n1854_), .A2(new_n1856_), .B(new_n1852_), .ZN(new_n1857_));
  NAND2_X1   g00854(.A1(\A[746] ), .A2(\A[747] ), .ZN(new_n1858_));
  NOR2_X1    g00855(.A1(\A[746] ), .A2(\A[747] ), .ZN(new_n1859_));
  INV_X1     g00856(.I(new_n1859_), .ZN(new_n1860_));
  AOI21_X1   g00857(.A1(new_n1860_), .A2(new_n1858_), .B(\A[745] ), .ZN(new_n1861_));
  NOR2_X1    g00858(.A1(new_n1861_), .A2(new_n1857_), .ZN(new_n1862_));
  INV_X1     g00859(.I(\A[748] ), .ZN(new_n1863_));
  INV_X1     g00860(.I(\A[749] ), .ZN(new_n1864_));
  NAND2_X1   g00861(.A1(new_n1864_), .A2(\A[750] ), .ZN(new_n1865_));
  INV_X1     g00862(.I(\A[750] ), .ZN(new_n1866_));
  NAND2_X1   g00863(.A1(new_n1866_), .A2(\A[749] ), .ZN(new_n1867_));
  AOI21_X1   g00864(.A1(new_n1865_), .A2(new_n1867_), .B(new_n1863_), .ZN(new_n1868_));
  NAND2_X1   g00865(.A1(\A[749] ), .A2(\A[750] ), .ZN(new_n1869_));
  NOR2_X1    g00866(.A1(\A[749] ), .A2(\A[750] ), .ZN(new_n1870_));
  INV_X1     g00867(.I(new_n1870_), .ZN(new_n1871_));
  AOI21_X1   g00868(.A1(new_n1871_), .A2(new_n1869_), .B(\A[748] ), .ZN(new_n1872_));
  NOR2_X1    g00869(.A1(new_n1872_), .A2(new_n1868_), .ZN(new_n1873_));
  AOI21_X1   g00870(.A1(new_n1852_), .A2(new_n1858_), .B(new_n1859_), .ZN(new_n1874_));
  AOI21_X1   g00871(.A1(new_n1863_), .A2(new_n1869_), .B(new_n1870_), .ZN(new_n1875_));
  OR2_X2     g00872(.A1(new_n1874_), .A2(new_n1875_), .Z(new_n1876_));
  NOR3_X1    g00873(.A1(new_n1876_), .A2(new_n1862_), .A3(new_n1873_), .ZN(new_n1877_));
  NAND2_X1   g00874(.A1(new_n1877_), .A2(new_n1851_), .ZN(new_n1878_));
  NOR2_X1    g00875(.A1(new_n1855_), .A2(\A[746] ), .ZN(new_n1879_));
  NOR2_X1    g00876(.A1(new_n1853_), .A2(\A[747] ), .ZN(new_n1880_));
  OAI21_X1   g00877(.A1(new_n1879_), .A2(new_n1880_), .B(\A[745] ), .ZN(new_n1881_));
  INV_X1     g00878(.I(new_n1858_), .ZN(new_n1882_));
  OAI21_X1   g00879(.A1(new_n1882_), .A2(new_n1859_), .B(new_n1852_), .ZN(new_n1883_));
  NAND2_X1   g00880(.A1(new_n1881_), .A2(new_n1883_), .ZN(new_n1884_));
  NOR2_X1    g00881(.A1(new_n1876_), .A2(new_n1884_), .ZN(new_n1885_));
  NOR2_X1    g00882(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1886_));
  NOR2_X1    g00883(.A1(new_n1862_), .A2(new_n1886_), .ZN(new_n1887_));
  OAI21_X1   g00884(.A1(new_n1885_), .A2(new_n1887_), .B(new_n1873_), .ZN(new_n1888_));
  INV_X1     g00885(.I(new_n1873_), .ZN(new_n1889_));
  NAND2_X1   g00886(.A1(new_n1862_), .A2(new_n1886_), .ZN(new_n1890_));
  NAND2_X1   g00887(.A1(new_n1876_), .A2(new_n1884_), .ZN(new_n1891_));
  NAND3_X1   g00888(.A1(new_n1891_), .A2(new_n1890_), .A3(new_n1889_), .ZN(new_n1892_));
  NAND2_X1   g00889(.A1(new_n1874_), .A2(new_n1875_), .ZN(new_n1893_));
  AND4_X2    g00890(.A1(new_n1851_), .A2(new_n1884_), .A3(new_n1889_), .A4(new_n1893_), .Z(new_n1894_));
  INV_X1     g00891(.I(new_n1845_), .ZN(new_n1895_));
  XNOR2_X1   g00892(.A1(new_n1835_), .A2(new_n1850_), .ZN(new_n1896_));
  NOR2_X1    g00893(.A1(new_n1896_), .A2(new_n1895_), .ZN(new_n1897_));
  XOR2_X1    g00894(.A1(new_n1835_), .A2(new_n1850_), .Z(new_n1898_));
  NOR2_X1    g00895(.A1(new_n1898_), .A2(new_n1845_), .ZN(new_n1899_));
  NOR2_X1    g00896(.A1(new_n1897_), .A2(new_n1899_), .ZN(new_n1900_));
  AND2_X2    g00897(.A1(new_n1888_), .A2(new_n1892_), .Z(new_n1901_));
  NOR2_X1    g00898(.A1(new_n1901_), .A2(new_n1878_), .ZN(new_n1902_));
  INV_X1     g00899(.I(new_n1902_), .ZN(new_n1903_));
  NAND2_X1   g00900(.A1(new_n1898_), .A2(new_n1845_), .ZN(new_n1904_));
  NAND2_X1   g00901(.A1(new_n1896_), .A2(new_n1895_), .ZN(new_n1905_));
  NAND2_X1   g00902(.A1(new_n1905_), .A2(new_n1904_), .ZN(new_n1906_));
  NAND2_X1   g00903(.A1(new_n1888_), .A2(new_n1892_), .ZN(new_n1907_));
  XOR2_X1    g00904(.A1(new_n1907_), .A2(new_n1878_), .Z(new_n1908_));
  XNOR2_X1   g00905(.A1(new_n1877_), .A2(new_n1851_), .ZN(new_n1909_));
  INV_X1     g00906(.I(\A[727] ), .ZN(new_n1910_));
  INV_X1     g00907(.I(\A[728] ), .ZN(new_n1911_));
  NAND2_X1   g00908(.A1(new_n1911_), .A2(\A[729] ), .ZN(new_n1912_));
  INV_X1     g00909(.I(\A[729] ), .ZN(new_n1913_));
  NAND2_X1   g00910(.A1(new_n1913_), .A2(\A[728] ), .ZN(new_n1914_));
  AOI21_X1   g00911(.A1(new_n1912_), .A2(new_n1914_), .B(new_n1910_), .ZN(new_n1915_));
  NAND2_X1   g00912(.A1(\A[728] ), .A2(\A[729] ), .ZN(new_n1916_));
  NAND2_X1   g00913(.A1(new_n1911_), .A2(new_n1913_), .ZN(new_n1917_));
  AOI21_X1   g00914(.A1(new_n1917_), .A2(new_n1916_), .B(\A[727] ), .ZN(new_n1918_));
  NOR2_X1    g00915(.A1(new_n1918_), .A2(new_n1915_), .ZN(new_n1919_));
  INV_X1     g00916(.I(\A[730] ), .ZN(new_n1920_));
  INV_X1     g00917(.I(\A[731] ), .ZN(new_n1921_));
  NAND2_X1   g00918(.A1(new_n1921_), .A2(\A[732] ), .ZN(new_n1922_));
  INV_X1     g00919(.I(\A[732] ), .ZN(new_n1923_));
  NAND2_X1   g00920(.A1(new_n1923_), .A2(\A[731] ), .ZN(new_n1924_));
  AOI21_X1   g00921(.A1(new_n1922_), .A2(new_n1924_), .B(new_n1920_), .ZN(new_n1925_));
  NAND2_X1   g00922(.A1(\A[731] ), .A2(\A[732] ), .ZN(new_n1926_));
  NOR2_X1    g00923(.A1(\A[731] ), .A2(\A[732] ), .ZN(new_n1927_));
  INV_X1     g00924(.I(new_n1927_), .ZN(new_n1928_));
  AOI21_X1   g00925(.A1(new_n1928_), .A2(new_n1926_), .B(\A[730] ), .ZN(new_n1929_));
  NOR2_X1    g00926(.A1(new_n1929_), .A2(new_n1925_), .ZN(new_n1930_));
  NAND2_X1   g00927(.A1(new_n1916_), .A2(new_n1910_), .ZN(new_n1931_));
  NAND2_X1   g00928(.A1(new_n1931_), .A2(new_n1917_), .ZN(new_n1932_));
  NAND2_X1   g00929(.A1(new_n1926_), .A2(new_n1920_), .ZN(new_n1933_));
  NAND2_X1   g00930(.A1(new_n1933_), .A2(new_n1928_), .ZN(new_n1934_));
  NAND2_X1   g00931(.A1(new_n1934_), .A2(new_n1932_), .ZN(new_n1935_));
  NOR3_X1    g00932(.A1(new_n1919_), .A2(new_n1930_), .A3(new_n1935_), .ZN(new_n1936_));
  INV_X1     g00933(.I(\A[735] ), .ZN(new_n1937_));
  NOR2_X1    g00934(.A1(new_n1937_), .A2(\A[734] ), .ZN(new_n1938_));
  INV_X1     g00935(.I(\A[734] ), .ZN(new_n1939_));
  NOR2_X1    g00936(.A1(new_n1939_), .A2(\A[735] ), .ZN(new_n1940_));
  OAI21_X1   g00937(.A1(new_n1938_), .A2(new_n1940_), .B(\A[733] ), .ZN(new_n1941_));
  INV_X1     g00938(.I(\A[733] ), .ZN(new_n1942_));
  NOR2_X1    g00939(.A1(\A[734] ), .A2(\A[735] ), .ZN(new_n1943_));
  NAND2_X1   g00940(.A1(\A[734] ), .A2(\A[735] ), .ZN(new_n1944_));
  INV_X1     g00941(.I(new_n1944_), .ZN(new_n1945_));
  OAI21_X1   g00942(.A1(new_n1945_), .A2(new_n1943_), .B(new_n1942_), .ZN(new_n1946_));
  NAND2_X1   g00943(.A1(new_n1941_), .A2(new_n1946_), .ZN(new_n1947_));
  INV_X1     g00944(.I(\A[738] ), .ZN(new_n1948_));
  NOR2_X1    g00945(.A1(new_n1948_), .A2(\A[737] ), .ZN(new_n1949_));
  INV_X1     g00946(.I(\A[737] ), .ZN(new_n1950_));
  NOR2_X1    g00947(.A1(new_n1950_), .A2(\A[738] ), .ZN(new_n1951_));
  OAI21_X1   g00948(.A1(new_n1949_), .A2(new_n1951_), .B(\A[736] ), .ZN(new_n1952_));
  INV_X1     g00949(.I(\A[736] ), .ZN(new_n1953_));
  NAND2_X1   g00950(.A1(\A[737] ), .A2(\A[738] ), .ZN(new_n1954_));
  INV_X1     g00951(.I(new_n1954_), .ZN(new_n1955_));
  NOR2_X1    g00952(.A1(\A[737] ), .A2(\A[738] ), .ZN(new_n1956_));
  OAI21_X1   g00953(.A1(new_n1955_), .A2(new_n1956_), .B(new_n1953_), .ZN(new_n1957_));
  NAND2_X1   g00954(.A1(new_n1952_), .A2(new_n1957_), .ZN(new_n1958_));
  AOI21_X1   g00955(.A1(new_n1942_), .A2(new_n1944_), .B(new_n1943_), .ZN(new_n1959_));
  AOI21_X1   g00956(.A1(new_n1953_), .A2(new_n1954_), .B(new_n1956_), .ZN(new_n1960_));
  NOR2_X1    g00957(.A1(new_n1959_), .A2(new_n1960_), .ZN(new_n1961_));
  NAND3_X1   g00958(.A1(new_n1947_), .A2(new_n1958_), .A3(new_n1961_), .ZN(new_n1962_));
  XOR2_X1    g00959(.A1(new_n1936_), .A2(new_n1962_), .Z(new_n1963_));
  NAND2_X1   g00960(.A1(new_n1909_), .A2(new_n1963_), .ZN(new_n1964_));
  NAND2_X1   g00961(.A1(new_n1950_), .A2(\A[738] ), .ZN(new_n1965_));
  NAND2_X1   g00962(.A1(new_n1948_), .A2(\A[737] ), .ZN(new_n1966_));
  AOI21_X1   g00963(.A1(new_n1965_), .A2(new_n1966_), .B(new_n1953_), .ZN(new_n1967_));
  INV_X1     g00964(.I(new_n1956_), .ZN(new_n1968_));
  AOI21_X1   g00965(.A1(new_n1968_), .A2(new_n1954_), .B(\A[736] ), .ZN(new_n1969_));
  NOR2_X1    g00966(.A1(new_n1969_), .A2(new_n1967_), .ZN(new_n1970_));
  INV_X1     g00967(.I(new_n1961_), .ZN(new_n1971_));
  NOR2_X1    g00968(.A1(new_n1971_), .A2(new_n1947_), .ZN(new_n1972_));
  NAND2_X1   g00969(.A1(new_n1939_), .A2(\A[735] ), .ZN(new_n1973_));
  NAND2_X1   g00970(.A1(new_n1937_), .A2(\A[734] ), .ZN(new_n1974_));
  AOI21_X1   g00971(.A1(new_n1973_), .A2(new_n1974_), .B(new_n1942_), .ZN(new_n1975_));
  INV_X1     g00972(.I(new_n1943_), .ZN(new_n1976_));
  AOI21_X1   g00973(.A1(new_n1976_), .A2(new_n1944_), .B(\A[733] ), .ZN(new_n1977_));
  NOR2_X1    g00974(.A1(new_n1977_), .A2(new_n1975_), .ZN(new_n1978_));
  NOR2_X1    g00975(.A1(new_n1978_), .A2(new_n1961_), .ZN(new_n1979_));
  OAI21_X1   g00976(.A1(new_n1972_), .A2(new_n1979_), .B(new_n1970_), .ZN(new_n1980_));
  NAND2_X1   g00977(.A1(new_n1978_), .A2(new_n1961_), .ZN(new_n1981_));
  NAND2_X1   g00978(.A1(new_n1971_), .A2(new_n1947_), .ZN(new_n1982_));
  NAND3_X1   g00979(.A1(new_n1982_), .A2(new_n1981_), .A3(new_n1958_), .ZN(new_n1983_));
  AND2_X2    g00980(.A1(new_n1980_), .A2(new_n1983_), .Z(new_n1984_));
  INV_X1     g00981(.I(new_n1936_), .ZN(new_n1985_));
  NOR2_X1    g00982(.A1(new_n1985_), .A2(new_n1962_), .ZN(new_n1986_));
  INV_X1     g00983(.I(new_n1986_), .ZN(new_n1987_));
  INV_X1     g00984(.I(new_n1919_), .ZN(new_n1988_));
  NOR2_X1    g00985(.A1(new_n1988_), .A2(new_n1935_), .ZN(new_n1989_));
  INV_X1     g00986(.I(new_n1935_), .ZN(new_n1990_));
  NOR2_X1    g00987(.A1(new_n1990_), .A2(new_n1919_), .ZN(new_n1991_));
  OAI21_X1   g00988(.A1(new_n1989_), .A2(new_n1991_), .B(new_n1930_), .ZN(new_n1992_));
  OR2_X2     g00989(.A1(new_n1929_), .A2(new_n1925_), .Z(new_n1993_));
  NAND2_X1   g00990(.A1(new_n1990_), .A2(new_n1919_), .ZN(new_n1994_));
  NAND2_X1   g00991(.A1(new_n1988_), .A2(new_n1935_), .ZN(new_n1995_));
  NAND3_X1   g00992(.A1(new_n1995_), .A2(new_n1994_), .A3(new_n1993_), .ZN(new_n1996_));
  NAND2_X1   g00993(.A1(new_n1992_), .A2(new_n1996_), .ZN(new_n1997_));
  AND2_X2    g00994(.A1(new_n1959_), .A2(new_n1960_), .Z(new_n1998_));
  NOR4_X1    g00995(.A1(new_n1985_), .A2(new_n1978_), .A3(new_n1970_), .A4(new_n1998_), .ZN(new_n1999_));
  NAND3_X1   g00996(.A1(new_n1984_), .A2(new_n1997_), .A3(new_n1987_), .ZN(new_n2000_));
  NOR2_X1    g00997(.A1(new_n2000_), .A2(new_n1964_), .ZN(new_n2001_));
  OAI21_X1   g00998(.A1(new_n1906_), .A2(new_n1908_), .B(new_n2001_), .ZN(new_n2002_));
  OR3_X2     g00999(.A1(new_n2001_), .A2(new_n1906_), .A3(new_n1908_), .Z(new_n2003_));
  AOI21_X1   g01000(.A1(new_n2003_), .A2(new_n2002_), .B(new_n1903_), .ZN(new_n2004_));
  INV_X1     g01001(.I(new_n2004_), .ZN(new_n2005_));
  INV_X1     g01002(.I(\A[718] ), .ZN(new_n2006_));
  INV_X1     g01003(.I(\A[719] ), .ZN(new_n2007_));
  NAND2_X1   g01004(.A1(new_n2007_), .A2(\A[720] ), .ZN(new_n2008_));
  INV_X1     g01005(.I(\A[720] ), .ZN(new_n2009_));
  NAND2_X1   g01006(.A1(new_n2009_), .A2(\A[719] ), .ZN(new_n2010_));
  AOI21_X1   g01007(.A1(new_n2008_), .A2(new_n2010_), .B(new_n2006_), .ZN(new_n2011_));
  NAND2_X1   g01008(.A1(\A[719] ), .A2(\A[720] ), .ZN(new_n2012_));
  NAND2_X1   g01009(.A1(new_n2007_), .A2(new_n2009_), .ZN(new_n2013_));
  AOI21_X1   g01010(.A1(new_n2013_), .A2(new_n2012_), .B(\A[718] ), .ZN(new_n2014_));
  NOR2_X1    g01011(.A1(new_n2014_), .A2(new_n2011_), .ZN(new_n2015_));
  INV_X1     g01012(.I(\A[715] ), .ZN(new_n2016_));
  INV_X1     g01013(.I(\A[716] ), .ZN(new_n2017_));
  NAND2_X1   g01014(.A1(new_n2017_), .A2(\A[717] ), .ZN(new_n2018_));
  INV_X1     g01015(.I(\A[717] ), .ZN(new_n2019_));
  NAND2_X1   g01016(.A1(new_n2019_), .A2(\A[716] ), .ZN(new_n2020_));
  AOI21_X1   g01017(.A1(new_n2018_), .A2(new_n2020_), .B(new_n2016_), .ZN(new_n2021_));
  NAND2_X1   g01018(.A1(\A[716] ), .A2(\A[717] ), .ZN(new_n2022_));
  NAND2_X1   g01019(.A1(new_n2017_), .A2(new_n2019_), .ZN(new_n2023_));
  AOI21_X1   g01020(.A1(new_n2023_), .A2(new_n2022_), .B(\A[715] ), .ZN(new_n2024_));
  NOR2_X1    g01021(.A1(new_n2024_), .A2(new_n2021_), .ZN(new_n2025_));
  INV_X1     g01022(.I(new_n2025_), .ZN(new_n2026_));
  NAND2_X1   g01023(.A1(new_n2012_), .A2(new_n2006_), .ZN(new_n2027_));
  NAND2_X1   g01024(.A1(new_n2027_), .A2(new_n2013_), .ZN(new_n2028_));
  NAND2_X1   g01025(.A1(new_n2022_), .A2(new_n2016_), .ZN(new_n2029_));
  NAND2_X1   g01026(.A1(new_n2029_), .A2(new_n2023_), .ZN(new_n2030_));
  NAND2_X1   g01027(.A1(new_n2028_), .A2(new_n2030_), .ZN(new_n2031_));
  NOR2_X1    g01028(.A1(new_n2026_), .A2(new_n2031_), .ZN(new_n2032_));
  INV_X1     g01029(.I(new_n2031_), .ZN(new_n2033_));
  NOR2_X1    g01030(.A1(new_n2033_), .A2(new_n2025_), .ZN(new_n2034_));
  OAI21_X1   g01031(.A1(new_n2032_), .A2(new_n2034_), .B(new_n2015_), .ZN(new_n2035_));
  INV_X1     g01032(.I(new_n2015_), .ZN(new_n2036_));
  NAND2_X1   g01033(.A1(new_n2033_), .A2(new_n2025_), .ZN(new_n2037_));
  NAND2_X1   g01034(.A1(new_n2026_), .A2(new_n2031_), .ZN(new_n2038_));
  NAND3_X1   g01035(.A1(new_n2038_), .A2(new_n2037_), .A3(new_n2036_), .ZN(new_n2039_));
  NAND2_X1   g01036(.A1(new_n2035_), .A2(new_n2039_), .ZN(new_n2040_));
  INV_X1     g01037(.I(new_n2040_), .ZN(new_n2041_));
  NOR3_X1    g01038(.A1(new_n2015_), .A2(new_n2025_), .A3(new_n2031_), .ZN(new_n2042_));
  INV_X1     g01039(.I(\A[721] ), .ZN(new_n2043_));
  INV_X1     g01040(.I(\A[722] ), .ZN(new_n2044_));
  NAND2_X1   g01041(.A1(new_n2044_), .A2(\A[723] ), .ZN(new_n2045_));
  INV_X1     g01042(.I(\A[723] ), .ZN(new_n2046_));
  NAND2_X1   g01043(.A1(new_n2046_), .A2(\A[722] ), .ZN(new_n2047_));
  AOI21_X1   g01044(.A1(new_n2045_), .A2(new_n2047_), .B(new_n2043_), .ZN(new_n2048_));
  NAND2_X1   g01045(.A1(\A[722] ), .A2(\A[723] ), .ZN(new_n2049_));
  NOR2_X1    g01046(.A1(\A[722] ), .A2(\A[723] ), .ZN(new_n2050_));
  INV_X1     g01047(.I(new_n2050_), .ZN(new_n2051_));
  AOI21_X1   g01048(.A1(new_n2051_), .A2(new_n2049_), .B(\A[721] ), .ZN(new_n2052_));
  NOR2_X1    g01049(.A1(new_n2052_), .A2(new_n2048_), .ZN(new_n2053_));
  INV_X1     g01050(.I(\A[724] ), .ZN(new_n2054_));
  INV_X1     g01051(.I(\A[725] ), .ZN(new_n2055_));
  NAND2_X1   g01052(.A1(new_n2055_), .A2(\A[726] ), .ZN(new_n2056_));
  INV_X1     g01053(.I(\A[726] ), .ZN(new_n2057_));
  NAND2_X1   g01054(.A1(new_n2057_), .A2(\A[725] ), .ZN(new_n2058_));
  AOI21_X1   g01055(.A1(new_n2056_), .A2(new_n2058_), .B(new_n2054_), .ZN(new_n2059_));
  NAND2_X1   g01056(.A1(\A[725] ), .A2(\A[726] ), .ZN(new_n2060_));
  NOR2_X1    g01057(.A1(\A[725] ), .A2(\A[726] ), .ZN(new_n2061_));
  INV_X1     g01058(.I(new_n2061_), .ZN(new_n2062_));
  AOI21_X1   g01059(.A1(new_n2062_), .A2(new_n2060_), .B(\A[724] ), .ZN(new_n2063_));
  NOR2_X1    g01060(.A1(new_n2063_), .A2(new_n2059_), .ZN(new_n2064_));
  AOI21_X1   g01061(.A1(new_n2043_), .A2(new_n2049_), .B(new_n2050_), .ZN(new_n2065_));
  AOI21_X1   g01062(.A1(new_n2054_), .A2(new_n2060_), .B(new_n2061_), .ZN(new_n2066_));
  NOR2_X1    g01063(.A1(new_n2065_), .A2(new_n2066_), .ZN(new_n2067_));
  INV_X1     g01064(.I(new_n2067_), .ZN(new_n2068_));
  NOR3_X1    g01065(.A1(new_n2068_), .A2(new_n2053_), .A3(new_n2064_), .ZN(new_n2069_));
  NAND2_X1   g01066(.A1(new_n2069_), .A2(new_n2042_), .ZN(new_n2070_));
  INV_X1     g01067(.I(new_n2070_), .ZN(new_n2071_));
  NOR2_X1    g01068(.A1(new_n2046_), .A2(\A[722] ), .ZN(new_n2072_));
  NOR2_X1    g01069(.A1(new_n2044_), .A2(\A[723] ), .ZN(new_n2073_));
  OAI21_X1   g01070(.A1(new_n2072_), .A2(new_n2073_), .B(\A[721] ), .ZN(new_n2074_));
  INV_X1     g01071(.I(new_n2049_), .ZN(new_n2075_));
  OAI21_X1   g01072(.A1(new_n2075_), .A2(new_n2050_), .B(new_n2043_), .ZN(new_n2076_));
  NAND2_X1   g01073(.A1(new_n2074_), .A2(new_n2076_), .ZN(new_n2077_));
  NOR2_X1    g01074(.A1(new_n2068_), .A2(new_n2077_), .ZN(new_n2078_));
  NOR2_X1    g01075(.A1(new_n2053_), .A2(new_n2067_), .ZN(new_n2079_));
  OAI21_X1   g01076(.A1(new_n2078_), .A2(new_n2079_), .B(new_n2064_), .ZN(new_n2080_));
  INV_X1     g01077(.I(new_n2064_), .ZN(new_n2081_));
  NAND2_X1   g01078(.A1(new_n2053_), .A2(new_n2067_), .ZN(new_n2082_));
  NAND2_X1   g01079(.A1(new_n2068_), .A2(new_n2077_), .ZN(new_n2083_));
  NAND3_X1   g01080(.A1(new_n2083_), .A2(new_n2082_), .A3(new_n2081_), .ZN(new_n2084_));
  NAND2_X1   g01081(.A1(new_n2080_), .A2(new_n2084_), .ZN(new_n2085_));
  XOR2_X1    g01082(.A1(new_n2085_), .A2(new_n2071_), .Z(new_n2086_));
  NAND2_X1   g01083(.A1(new_n2086_), .A2(new_n2041_), .ZN(new_n2087_));
  INV_X1     g01084(.I(new_n2085_), .ZN(new_n2088_));
  NAND2_X1   g01085(.A1(new_n2065_), .A2(new_n2066_), .ZN(new_n2089_));
  NAND4_X1   g01086(.A1(new_n2042_), .A2(new_n2077_), .A3(new_n2081_), .A4(new_n2089_), .ZN(new_n2090_));
  NOR2_X1    g01087(.A1(new_n2088_), .A2(new_n2090_), .ZN(new_n2091_));
  INV_X1     g01088(.I(new_n2091_), .ZN(new_n2092_));
  NAND4_X1   g01089(.A1(new_n2042_), .A2(new_n2077_), .A3(new_n2081_), .A4(new_n2067_), .ZN(new_n2094_));
  INV_X1     g01090(.I(new_n2094_), .ZN(new_n2095_));
  INV_X1     g01091(.I(\A[706] ), .ZN(new_n2096_));
  INV_X1     g01092(.I(\A[707] ), .ZN(new_n2097_));
  NAND2_X1   g01093(.A1(new_n2097_), .A2(\A[708] ), .ZN(new_n2098_));
  INV_X1     g01094(.I(\A[708] ), .ZN(new_n2099_));
  NAND2_X1   g01095(.A1(new_n2099_), .A2(\A[707] ), .ZN(new_n2100_));
  AOI21_X1   g01096(.A1(new_n2098_), .A2(new_n2100_), .B(new_n2096_), .ZN(new_n2101_));
  NAND2_X1   g01097(.A1(\A[707] ), .A2(\A[708] ), .ZN(new_n2102_));
  NOR2_X1    g01098(.A1(\A[707] ), .A2(\A[708] ), .ZN(new_n2103_));
  INV_X1     g01099(.I(new_n2103_), .ZN(new_n2104_));
  AOI21_X1   g01100(.A1(new_n2104_), .A2(new_n2102_), .B(\A[706] ), .ZN(new_n2105_));
  NOR2_X1    g01101(.A1(new_n2105_), .A2(new_n2101_), .ZN(new_n2106_));
  INV_X1     g01102(.I(\A[703] ), .ZN(new_n2107_));
  INV_X1     g01103(.I(\A[704] ), .ZN(new_n2108_));
  NAND2_X1   g01104(.A1(new_n2108_), .A2(\A[705] ), .ZN(new_n2109_));
  INV_X1     g01105(.I(\A[705] ), .ZN(new_n2110_));
  NAND2_X1   g01106(.A1(new_n2110_), .A2(\A[704] ), .ZN(new_n2111_));
  AOI21_X1   g01107(.A1(new_n2109_), .A2(new_n2111_), .B(new_n2107_), .ZN(new_n2112_));
  NOR2_X1    g01108(.A1(\A[704] ), .A2(\A[705] ), .ZN(new_n2113_));
  INV_X1     g01109(.I(new_n2113_), .ZN(new_n2114_));
  NAND2_X1   g01110(.A1(\A[704] ), .A2(\A[705] ), .ZN(new_n2115_));
  AOI21_X1   g01111(.A1(new_n2114_), .A2(new_n2115_), .B(\A[703] ), .ZN(new_n2116_));
  NOR2_X1    g01112(.A1(new_n2116_), .A2(new_n2112_), .ZN(new_n2117_));
  NOR2_X1    g01113(.A1(new_n2106_), .A2(new_n2117_), .ZN(new_n2118_));
  NOR2_X1    g01114(.A1(new_n2099_), .A2(\A[707] ), .ZN(new_n2119_));
  NOR2_X1    g01115(.A1(new_n2097_), .A2(\A[708] ), .ZN(new_n2120_));
  OAI21_X1   g01116(.A1(new_n2119_), .A2(new_n2120_), .B(\A[706] ), .ZN(new_n2121_));
  INV_X1     g01117(.I(new_n2102_), .ZN(new_n2122_));
  OAI21_X1   g01118(.A1(new_n2122_), .A2(new_n2103_), .B(new_n2096_), .ZN(new_n2123_));
  NAND2_X1   g01119(.A1(new_n2121_), .A2(new_n2123_), .ZN(new_n2124_));
  NOR2_X1    g01120(.A1(new_n2110_), .A2(\A[704] ), .ZN(new_n2125_));
  NOR2_X1    g01121(.A1(new_n2108_), .A2(\A[705] ), .ZN(new_n2126_));
  OAI21_X1   g01122(.A1(new_n2125_), .A2(new_n2126_), .B(\A[703] ), .ZN(new_n2127_));
  INV_X1     g01123(.I(new_n2115_), .ZN(new_n2128_));
  OAI21_X1   g01124(.A1(new_n2128_), .A2(new_n2113_), .B(new_n2107_), .ZN(new_n2129_));
  NAND2_X1   g01125(.A1(new_n2127_), .A2(new_n2129_), .ZN(new_n2130_));
  NOR2_X1    g01126(.A1(new_n2124_), .A2(new_n2130_), .ZN(new_n2131_));
  NOR2_X1    g01127(.A1(new_n2118_), .A2(new_n2131_), .ZN(new_n2132_));
  INV_X1     g01128(.I(\A[712] ), .ZN(new_n2133_));
  INV_X1     g01129(.I(\A[713] ), .ZN(new_n2134_));
  NAND2_X1   g01130(.A1(new_n2134_), .A2(\A[714] ), .ZN(new_n2135_));
  INV_X1     g01131(.I(\A[714] ), .ZN(new_n2136_));
  NAND2_X1   g01132(.A1(new_n2136_), .A2(\A[713] ), .ZN(new_n2137_));
  AOI21_X1   g01133(.A1(new_n2135_), .A2(new_n2137_), .B(new_n2133_), .ZN(new_n2138_));
  NOR2_X1    g01134(.A1(\A[713] ), .A2(\A[714] ), .ZN(new_n2139_));
  INV_X1     g01135(.I(new_n2139_), .ZN(new_n2140_));
  NAND2_X1   g01136(.A1(\A[713] ), .A2(\A[714] ), .ZN(new_n2141_));
  AOI21_X1   g01137(.A1(new_n2140_), .A2(new_n2141_), .B(\A[712] ), .ZN(new_n2142_));
  NOR2_X1    g01138(.A1(new_n2142_), .A2(new_n2138_), .ZN(new_n2143_));
  INV_X1     g01139(.I(\A[709] ), .ZN(new_n2144_));
  INV_X1     g01140(.I(\A[710] ), .ZN(new_n2145_));
  NAND2_X1   g01141(.A1(new_n2145_), .A2(\A[711] ), .ZN(new_n2146_));
  INV_X1     g01142(.I(\A[711] ), .ZN(new_n2147_));
  NAND2_X1   g01143(.A1(new_n2147_), .A2(\A[710] ), .ZN(new_n2148_));
  AOI21_X1   g01144(.A1(new_n2146_), .A2(new_n2148_), .B(new_n2144_), .ZN(new_n2149_));
  NOR2_X1    g01145(.A1(\A[710] ), .A2(\A[711] ), .ZN(new_n2150_));
  INV_X1     g01146(.I(new_n2150_), .ZN(new_n2151_));
  NAND2_X1   g01147(.A1(\A[710] ), .A2(\A[711] ), .ZN(new_n2152_));
  AOI21_X1   g01148(.A1(new_n2151_), .A2(new_n2152_), .B(\A[709] ), .ZN(new_n2153_));
  NOR2_X1    g01149(.A1(new_n2153_), .A2(new_n2149_), .ZN(new_n2154_));
  NOR2_X1    g01150(.A1(new_n2143_), .A2(new_n2154_), .ZN(new_n2155_));
  NOR2_X1    g01151(.A1(new_n2136_), .A2(\A[713] ), .ZN(new_n2156_));
  NOR2_X1    g01152(.A1(new_n2134_), .A2(\A[714] ), .ZN(new_n2157_));
  OAI21_X1   g01153(.A1(new_n2156_), .A2(new_n2157_), .B(\A[712] ), .ZN(new_n2158_));
  INV_X1     g01154(.I(new_n2141_), .ZN(new_n2159_));
  OAI21_X1   g01155(.A1(new_n2159_), .A2(new_n2139_), .B(new_n2133_), .ZN(new_n2160_));
  NAND2_X1   g01156(.A1(new_n2158_), .A2(new_n2160_), .ZN(new_n2161_));
  NOR2_X1    g01157(.A1(new_n2147_), .A2(\A[710] ), .ZN(new_n2162_));
  NOR2_X1    g01158(.A1(new_n2145_), .A2(\A[711] ), .ZN(new_n2163_));
  OAI21_X1   g01159(.A1(new_n2162_), .A2(new_n2163_), .B(\A[709] ), .ZN(new_n2164_));
  INV_X1     g01160(.I(new_n2152_), .ZN(new_n2165_));
  OAI21_X1   g01161(.A1(new_n2165_), .A2(new_n2150_), .B(new_n2144_), .ZN(new_n2166_));
  NAND2_X1   g01162(.A1(new_n2164_), .A2(new_n2166_), .ZN(new_n2167_));
  NOR2_X1    g01163(.A1(new_n2161_), .A2(new_n2167_), .ZN(new_n2168_));
  NOR2_X1    g01164(.A1(new_n2155_), .A2(new_n2168_), .ZN(new_n2169_));
  AOI21_X1   g01165(.A1(new_n2144_), .A2(new_n2152_), .B(new_n2150_), .ZN(new_n2170_));
  AOI21_X1   g01166(.A1(new_n2133_), .A2(new_n2141_), .B(new_n2139_), .ZN(new_n2171_));
  NOR2_X1    g01167(.A1(new_n2170_), .A2(new_n2171_), .ZN(new_n2172_));
  INV_X1     g01168(.I(new_n2172_), .ZN(new_n2173_));
  NOR2_X1    g01169(.A1(new_n2173_), .A2(new_n2143_), .ZN(new_n2174_));
  AOI21_X1   g01170(.A1(new_n2107_), .A2(new_n2115_), .B(new_n2113_), .ZN(new_n2175_));
  AOI21_X1   g01171(.A1(new_n2096_), .A2(new_n2102_), .B(new_n2103_), .ZN(new_n2176_));
  OR2_X2     g01172(.A1(new_n2175_), .A2(new_n2176_), .Z(new_n2177_));
  NOR3_X1    g01173(.A1(new_n2106_), .A2(new_n2177_), .A3(new_n2117_), .ZN(new_n2178_));
  NAND3_X1   g01174(.A1(new_n2178_), .A2(new_n2174_), .A3(new_n2167_), .ZN(new_n2179_));
  NOR3_X1    g01175(.A1(new_n2179_), .A2(new_n2132_), .A3(new_n2169_), .ZN(new_n2180_));
  INV_X1     g01176(.I(new_n2180_), .ZN(new_n2181_));
  NOR2_X1    g01177(.A1(new_n2173_), .A2(new_n2167_), .ZN(new_n2182_));
  NOR2_X1    g01178(.A1(new_n2154_), .A2(new_n2172_), .ZN(new_n2183_));
  OAI21_X1   g01179(.A1(new_n2182_), .A2(new_n2183_), .B(new_n2143_), .ZN(new_n2184_));
  NAND2_X1   g01180(.A1(new_n2154_), .A2(new_n2172_), .ZN(new_n2185_));
  NAND2_X1   g01181(.A1(new_n2173_), .A2(new_n2167_), .ZN(new_n2186_));
  NAND3_X1   g01182(.A1(new_n2186_), .A2(new_n2185_), .A3(new_n2161_), .ZN(new_n2187_));
  XOR2_X1    g01183(.A1(new_n2161_), .A2(new_n2167_), .Z(new_n2188_));
  NAND2_X1   g01184(.A1(new_n2188_), .A2(new_n2172_), .ZN(new_n2189_));
  NAND3_X1   g01185(.A1(new_n2189_), .A2(new_n2184_), .A3(new_n2187_), .ZN(new_n2190_));
  NOR2_X1    g01186(.A1(new_n2175_), .A2(new_n2176_), .ZN(new_n2191_));
  NAND2_X1   g01187(.A1(new_n2117_), .A2(new_n2191_), .ZN(new_n2192_));
  NAND2_X1   g01188(.A1(new_n2177_), .A2(new_n2130_), .ZN(new_n2193_));
  NAND2_X1   g01189(.A1(new_n2193_), .A2(new_n2192_), .ZN(new_n2194_));
  XOR2_X1    g01190(.A1(new_n2194_), .A2(new_n2124_), .Z(new_n2195_));
  NAND2_X1   g01191(.A1(new_n2124_), .A2(new_n2191_), .ZN(new_n2196_));
  OAI22_X1   g01192(.A1(new_n2118_), .A2(new_n2131_), .B1(new_n2196_), .B2(new_n2117_), .ZN(new_n2197_));
  NOR4_X1    g01193(.A1(new_n2197_), .A2(new_n2143_), .A3(new_n2154_), .A4(new_n2173_), .ZN(new_n2198_));
  INV_X1     g01194(.I(new_n2198_), .ZN(new_n2199_));
  NAND4_X1   g01195(.A1(new_n2199_), .A2(new_n2190_), .A3(new_n2195_), .A4(new_n2181_), .ZN(new_n2200_));
  XNOR2_X1   g01196(.A1(new_n2069_), .A2(new_n2042_), .ZN(new_n2201_));
  NAND3_X1   g01197(.A1(new_n2161_), .A2(new_n2167_), .A3(new_n2172_), .ZN(new_n2202_));
  NOR3_X1    g01198(.A1(new_n2177_), .A2(new_n2106_), .A3(new_n2117_), .ZN(new_n2203_));
  XOR2_X1    g01199(.A1(new_n2203_), .A2(new_n2202_), .Z(new_n2204_));
  NAND2_X1   g01200(.A1(new_n2201_), .A2(new_n2204_), .ZN(new_n2205_));
  NOR3_X1    g01201(.A1(new_n2200_), .A2(new_n2095_), .A3(new_n2205_), .ZN(new_n2206_));
  NAND2_X1   g01202(.A1(new_n2184_), .A2(new_n2187_), .ZN(new_n2207_));
  XOR2_X1    g01203(.A1(new_n2143_), .A2(new_n2167_), .Z(new_n2208_));
  NOR2_X1    g01204(.A1(new_n2208_), .A2(new_n2173_), .ZN(new_n2209_));
  NOR2_X1    g01205(.A1(new_n2209_), .A2(new_n2207_), .ZN(new_n2210_));
  XOR2_X1    g01206(.A1(new_n2194_), .A2(new_n2106_), .Z(new_n2211_));
  NOR4_X1    g01207(.A1(new_n2210_), .A2(new_n2211_), .A3(new_n2180_), .A4(new_n2198_), .ZN(new_n2212_));
  INV_X1     g01208(.I(new_n2205_), .ZN(new_n2213_));
  AOI21_X1   g01209(.A1(new_n2212_), .A2(new_n2213_), .B(new_n2094_), .ZN(new_n2214_));
  OAI21_X1   g01210(.A1(new_n2206_), .A2(new_n2214_), .B(new_n2087_), .ZN(new_n2215_));
  XOR2_X1    g01211(.A1(new_n2085_), .A2(new_n2070_), .Z(new_n2216_));
  NOR2_X1    g01212(.A1(new_n2216_), .A2(new_n2040_), .ZN(new_n2217_));
  NAND3_X1   g01213(.A1(new_n2212_), .A2(new_n2213_), .A3(new_n2094_), .ZN(new_n2218_));
  OAI21_X1   g01214(.A1(new_n2200_), .A2(new_n2205_), .B(new_n2095_), .ZN(new_n2219_));
  NAND3_X1   g01215(.A1(new_n2219_), .A2(new_n2218_), .A3(new_n2217_), .ZN(new_n2220_));
  XOR2_X1    g01216(.A1(new_n1877_), .A2(new_n1851_), .Z(new_n2221_));
  XNOR2_X1   g01217(.A1(new_n1936_), .A2(new_n1962_), .ZN(new_n2222_));
  NOR2_X1    g01218(.A1(new_n2221_), .A2(new_n2222_), .ZN(new_n2223_));
  NOR2_X1    g01219(.A1(new_n1909_), .A2(new_n1963_), .ZN(new_n2224_));
  NOR2_X1    g01220(.A1(new_n2223_), .A2(new_n2224_), .ZN(new_n2225_));
  NOR2_X1    g01221(.A1(new_n2201_), .A2(new_n2204_), .ZN(new_n2226_));
  NOR2_X1    g01222(.A1(new_n2213_), .A2(new_n2226_), .ZN(new_n2227_));
  NAND2_X1   g01223(.A1(new_n2227_), .A2(new_n2225_), .ZN(new_n2228_));
  AOI21_X1   g01224(.A1(new_n2215_), .A2(new_n2220_), .B(new_n2228_), .ZN(new_n2229_));
  NOR2_X1    g01225(.A1(new_n2005_), .A2(new_n2229_), .ZN(new_n2230_));
  INV_X1     g01226(.I(new_n2230_), .ZN(new_n2231_));
  INV_X1     g01227(.I(\A[691] ), .ZN(new_n2232_));
  INV_X1     g01228(.I(\A[692] ), .ZN(new_n2233_));
  NAND2_X1   g01229(.A1(new_n2233_), .A2(\A[693] ), .ZN(new_n2234_));
  INV_X1     g01230(.I(\A[693] ), .ZN(new_n2235_));
  NAND2_X1   g01231(.A1(new_n2235_), .A2(\A[692] ), .ZN(new_n2236_));
  AOI21_X1   g01232(.A1(new_n2234_), .A2(new_n2236_), .B(new_n2232_), .ZN(new_n2237_));
  NAND2_X1   g01233(.A1(new_n2233_), .A2(new_n2235_), .ZN(new_n2238_));
  NAND2_X1   g01234(.A1(\A[692] ), .A2(\A[693] ), .ZN(new_n2239_));
  AOI21_X1   g01235(.A1(new_n2238_), .A2(new_n2239_), .B(\A[691] ), .ZN(new_n2240_));
  NOR2_X1    g01236(.A1(new_n2240_), .A2(new_n2237_), .ZN(new_n2241_));
  INV_X1     g01237(.I(\A[694] ), .ZN(new_n2242_));
  INV_X1     g01238(.I(\A[695] ), .ZN(new_n2243_));
  INV_X1     g01239(.I(\A[696] ), .ZN(new_n2244_));
  NAND2_X1   g01240(.A1(new_n2239_), .A2(new_n2232_), .ZN(new_n2245_));
  NAND2_X1   g01241(.A1(new_n2245_), .A2(new_n2238_), .ZN(new_n2246_));
  NAND4_X1   g01242(.A1(new_n2246_), .A2(new_n2242_), .A3(new_n2243_), .A4(new_n2244_), .ZN(new_n2247_));
  NOR2_X1    g01243(.A1(new_n2247_), .A2(new_n2241_), .ZN(new_n2248_));
  INV_X1     g01244(.I(\A[699] ), .ZN(new_n2249_));
  NOR2_X1    g01245(.A1(new_n2249_), .A2(\A[698] ), .ZN(new_n2250_));
  INV_X1     g01246(.I(\A[698] ), .ZN(new_n2251_));
  NOR2_X1    g01247(.A1(new_n2251_), .A2(\A[699] ), .ZN(new_n2252_));
  OAI21_X1   g01248(.A1(new_n2250_), .A2(new_n2252_), .B(\A[697] ), .ZN(new_n2253_));
  INV_X1     g01249(.I(\A[697] ), .ZN(new_n2254_));
  NOR2_X1    g01250(.A1(\A[698] ), .A2(\A[699] ), .ZN(new_n2255_));
  NOR2_X1    g01251(.A1(new_n2251_), .A2(new_n2249_), .ZN(new_n2256_));
  OAI21_X1   g01252(.A1(new_n2256_), .A2(new_n2255_), .B(new_n2254_), .ZN(new_n2257_));
  NAND2_X1   g01253(.A1(new_n2257_), .A2(new_n2253_), .ZN(new_n2258_));
  INV_X1     g01254(.I(\A[702] ), .ZN(new_n2259_));
  NOR2_X1    g01255(.A1(new_n2259_), .A2(\A[701] ), .ZN(new_n2260_));
  INV_X1     g01256(.I(\A[701] ), .ZN(new_n2261_));
  NOR2_X1    g01257(.A1(new_n2261_), .A2(\A[702] ), .ZN(new_n2262_));
  OAI21_X1   g01258(.A1(new_n2260_), .A2(new_n2262_), .B(\A[700] ), .ZN(new_n2263_));
  INV_X1     g01259(.I(\A[700] ), .ZN(new_n2264_));
  NOR2_X1    g01260(.A1(new_n2261_), .A2(new_n2259_), .ZN(new_n2265_));
  NOR2_X1    g01261(.A1(\A[701] ), .A2(\A[702] ), .ZN(new_n2266_));
  OAI21_X1   g01262(.A1(new_n2265_), .A2(new_n2266_), .B(new_n2264_), .ZN(new_n2267_));
  NAND2_X1   g01263(.A1(new_n2267_), .A2(new_n2263_), .ZN(new_n2268_));
  NOR2_X1    g01264(.A1(new_n2256_), .A2(\A[697] ), .ZN(new_n2269_));
  NOR2_X1    g01265(.A1(new_n2265_), .A2(\A[700] ), .ZN(new_n2270_));
  OAI22_X1   g01266(.A1(new_n2255_), .A2(new_n2269_), .B1(new_n2270_), .B2(new_n2266_), .ZN(new_n2271_));
  INV_X1     g01267(.I(new_n2271_), .ZN(new_n2272_));
  NAND4_X1   g01268(.A1(new_n2248_), .A2(new_n2272_), .A3(new_n2258_), .A4(new_n2268_), .ZN(new_n2273_));
  INV_X1     g01269(.I(new_n2258_), .ZN(new_n2274_));
  INV_X1     g01270(.I(new_n2268_), .ZN(new_n2275_));
  NOR2_X1    g01271(.A1(new_n2274_), .A2(new_n2275_), .ZN(new_n2276_));
  NOR2_X1    g01272(.A1(new_n2258_), .A2(new_n2268_), .ZN(new_n2277_));
  NOR2_X1    g01273(.A1(new_n2276_), .A2(new_n2277_), .ZN(new_n2278_));
  NOR2_X1    g01274(.A1(new_n2244_), .A2(\A[695] ), .ZN(new_n2279_));
  NOR2_X1    g01275(.A1(new_n2243_), .A2(\A[696] ), .ZN(new_n2280_));
  OAI21_X1   g01276(.A1(new_n2279_), .A2(new_n2280_), .B(\A[694] ), .ZN(new_n2281_));
  NOR2_X1    g01277(.A1(new_n2243_), .A2(new_n2244_), .ZN(new_n2282_));
  NOR2_X1    g01278(.A1(\A[695] ), .A2(\A[696] ), .ZN(new_n2283_));
  OAI21_X1   g01279(.A1(new_n2282_), .A2(new_n2283_), .B(new_n2242_), .ZN(new_n2284_));
  NAND2_X1   g01280(.A1(new_n2284_), .A2(new_n2281_), .ZN(new_n2285_));
  INV_X1     g01281(.I(new_n2285_), .ZN(new_n2286_));
  NOR2_X1    g01282(.A1(new_n2286_), .A2(new_n2241_), .ZN(new_n2287_));
  NOR3_X1    g01283(.A1(new_n2285_), .A2(new_n2237_), .A3(new_n2240_), .ZN(new_n2288_));
  NOR2_X1    g01284(.A1(new_n2287_), .A2(new_n2288_), .ZN(new_n2289_));
  NOR3_X1    g01285(.A1(new_n2278_), .A2(new_n2289_), .A3(new_n2273_), .ZN(new_n2290_));
  INV_X1     g01286(.I(new_n2290_), .ZN(new_n2291_));
  XNOR2_X1   g01287(.A1(new_n2271_), .A2(new_n2258_), .ZN(new_n2292_));
  NAND2_X1   g01288(.A1(new_n2292_), .A2(new_n2275_), .ZN(new_n2293_));
  XOR2_X1    g01289(.A1(new_n2271_), .A2(new_n2258_), .Z(new_n2294_));
  NAND2_X1   g01290(.A1(new_n2294_), .A2(new_n2268_), .ZN(new_n2295_));
  XOR2_X1    g01291(.A1(new_n2258_), .A2(new_n2268_), .Z(new_n2296_));
  NAND2_X1   g01292(.A1(new_n2296_), .A2(new_n2272_), .ZN(new_n2297_));
  NAND3_X1   g01293(.A1(new_n2293_), .A2(new_n2295_), .A3(new_n2297_), .ZN(new_n2298_));
  OAI22_X1   g01294(.A1(new_n2287_), .A2(new_n2288_), .B1(new_n2241_), .B2(new_n2247_), .ZN(new_n2299_));
  NOR4_X1    g01295(.A1(new_n2299_), .A2(new_n2274_), .A3(new_n2275_), .A4(new_n2271_), .ZN(new_n2300_));
  NOR2_X1    g01296(.A1(new_n2282_), .A2(\A[694] ), .ZN(new_n2301_));
  OAI21_X1   g01297(.A1(new_n2283_), .A2(new_n2301_), .B(new_n2246_), .ZN(new_n2302_));
  XOR2_X1    g01298(.A1(new_n2302_), .A2(new_n2241_), .Z(new_n2303_));
  XOR2_X1    g01299(.A1(new_n2303_), .A2(new_n2285_), .Z(new_n2304_));
  NAND2_X1   g01300(.A1(new_n2304_), .A2(new_n2300_), .ZN(new_n2305_));
  AOI21_X1   g01301(.A1(new_n2305_), .A2(new_n2298_), .B(new_n2291_), .ZN(new_n2306_));
  XOR2_X1    g01302(.A1(new_n2298_), .A2(new_n2290_), .Z(new_n2307_));
  NOR2_X1    g01303(.A1(new_n2307_), .A2(new_n2304_), .ZN(new_n2308_));
  INV_X1     g01304(.I(\A[682] ), .ZN(new_n2309_));
  INV_X1     g01305(.I(\A[683] ), .ZN(new_n2310_));
  NAND2_X1   g01306(.A1(new_n2310_), .A2(\A[684] ), .ZN(new_n2311_));
  INV_X1     g01307(.I(\A[684] ), .ZN(new_n2312_));
  NAND2_X1   g01308(.A1(new_n2312_), .A2(\A[683] ), .ZN(new_n2313_));
  AOI21_X1   g01309(.A1(new_n2311_), .A2(new_n2313_), .B(new_n2309_), .ZN(new_n2314_));
  NAND2_X1   g01310(.A1(\A[683] ), .A2(\A[684] ), .ZN(new_n2315_));
  NOR2_X1    g01311(.A1(\A[683] ), .A2(\A[684] ), .ZN(new_n2316_));
  INV_X1     g01312(.I(new_n2316_), .ZN(new_n2317_));
  AOI21_X1   g01313(.A1(new_n2317_), .A2(new_n2315_), .B(\A[682] ), .ZN(new_n2318_));
  NOR2_X1    g01314(.A1(new_n2318_), .A2(new_n2314_), .ZN(new_n2319_));
  INV_X1     g01315(.I(\A[679] ), .ZN(new_n2320_));
  INV_X1     g01316(.I(\A[680] ), .ZN(new_n2321_));
  NAND2_X1   g01317(.A1(new_n2321_), .A2(\A[681] ), .ZN(new_n2322_));
  INV_X1     g01318(.I(\A[681] ), .ZN(new_n2323_));
  NAND2_X1   g01319(.A1(new_n2323_), .A2(\A[680] ), .ZN(new_n2324_));
  AOI21_X1   g01320(.A1(new_n2322_), .A2(new_n2324_), .B(new_n2320_), .ZN(new_n2325_));
  NOR2_X1    g01321(.A1(\A[680] ), .A2(\A[681] ), .ZN(new_n2326_));
  INV_X1     g01322(.I(new_n2326_), .ZN(new_n2327_));
  NAND2_X1   g01323(.A1(\A[680] ), .A2(\A[681] ), .ZN(new_n2328_));
  AOI21_X1   g01324(.A1(new_n2327_), .A2(new_n2328_), .B(\A[679] ), .ZN(new_n2329_));
  NOR2_X1    g01325(.A1(new_n2329_), .A2(new_n2325_), .ZN(new_n2330_));
  NOR2_X1    g01326(.A1(new_n2319_), .A2(new_n2330_), .ZN(new_n2331_));
  NOR2_X1    g01327(.A1(new_n2312_), .A2(\A[683] ), .ZN(new_n2332_));
  NOR2_X1    g01328(.A1(new_n2310_), .A2(\A[684] ), .ZN(new_n2333_));
  OAI21_X1   g01329(.A1(new_n2332_), .A2(new_n2333_), .B(\A[682] ), .ZN(new_n2334_));
  INV_X1     g01330(.I(new_n2315_), .ZN(new_n2335_));
  OAI21_X1   g01331(.A1(new_n2335_), .A2(new_n2316_), .B(new_n2309_), .ZN(new_n2336_));
  NAND2_X1   g01332(.A1(new_n2334_), .A2(new_n2336_), .ZN(new_n2337_));
  NOR2_X1    g01333(.A1(new_n2323_), .A2(\A[680] ), .ZN(new_n2338_));
  NOR2_X1    g01334(.A1(new_n2321_), .A2(\A[681] ), .ZN(new_n2339_));
  OAI21_X1   g01335(.A1(new_n2338_), .A2(new_n2339_), .B(\A[679] ), .ZN(new_n2340_));
  INV_X1     g01336(.I(new_n2328_), .ZN(new_n2341_));
  OAI21_X1   g01337(.A1(new_n2341_), .A2(new_n2326_), .B(new_n2320_), .ZN(new_n2342_));
  NAND2_X1   g01338(.A1(new_n2340_), .A2(new_n2342_), .ZN(new_n2343_));
  NOR2_X1    g01339(.A1(new_n2337_), .A2(new_n2343_), .ZN(new_n2344_));
  NOR2_X1    g01340(.A1(new_n2331_), .A2(new_n2344_), .ZN(new_n2345_));
  INV_X1     g01341(.I(\A[690] ), .ZN(new_n2346_));
  NOR2_X1    g01342(.A1(new_n2346_), .A2(\A[689] ), .ZN(new_n2347_));
  INV_X1     g01343(.I(\A[689] ), .ZN(new_n2348_));
  NOR2_X1    g01344(.A1(new_n2348_), .A2(\A[690] ), .ZN(new_n2349_));
  OAI21_X1   g01345(.A1(new_n2347_), .A2(new_n2349_), .B(\A[688] ), .ZN(new_n2350_));
  INV_X1     g01346(.I(\A[688] ), .ZN(new_n2351_));
  NOR2_X1    g01347(.A1(\A[689] ), .A2(\A[690] ), .ZN(new_n2352_));
  NAND2_X1   g01348(.A1(\A[689] ), .A2(\A[690] ), .ZN(new_n2353_));
  INV_X1     g01349(.I(new_n2353_), .ZN(new_n2354_));
  OAI21_X1   g01350(.A1(new_n2354_), .A2(new_n2352_), .B(new_n2351_), .ZN(new_n2355_));
  NAND2_X1   g01351(.A1(new_n2350_), .A2(new_n2355_), .ZN(new_n2356_));
  INV_X1     g01352(.I(new_n2356_), .ZN(new_n2357_));
  INV_X1     g01353(.I(\A[687] ), .ZN(new_n2358_));
  NOR2_X1    g01354(.A1(new_n2358_), .A2(\A[686] ), .ZN(new_n2359_));
  INV_X1     g01355(.I(\A[686] ), .ZN(new_n2360_));
  NOR2_X1    g01356(.A1(new_n2360_), .A2(\A[687] ), .ZN(new_n2361_));
  OAI21_X1   g01357(.A1(new_n2359_), .A2(new_n2361_), .B(\A[685] ), .ZN(new_n2362_));
  INV_X1     g01358(.I(\A[685] ), .ZN(new_n2363_));
  NOR2_X1    g01359(.A1(\A[686] ), .A2(\A[687] ), .ZN(new_n2364_));
  NAND2_X1   g01360(.A1(\A[686] ), .A2(\A[687] ), .ZN(new_n2365_));
  INV_X1     g01361(.I(new_n2365_), .ZN(new_n2366_));
  OAI21_X1   g01362(.A1(new_n2366_), .A2(new_n2364_), .B(new_n2363_), .ZN(new_n2367_));
  AND2_X2    g01363(.A1(new_n2362_), .A2(new_n2367_), .Z(new_n2368_));
  NOR2_X1    g01364(.A1(new_n2357_), .A2(new_n2368_), .ZN(new_n2369_));
  NAND2_X1   g01365(.A1(new_n2362_), .A2(new_n2367_), .ZN(new_n2370_));
  NOR2_X1    g01366(.A1(new_n2356_), .A2(new_n2370_), .ZN(new_n2371_));
  NOR2_X1    g01367(.A1(new_n2369_), .A2(new_n2371_), .ZN(new_n2372_));
  AOI21_X1   g01368(.A1(new_n2363_), .A2(new_n2365_), .B(new_n2364_), .ZN(new_n2373_));
  AOI21_X1   g01369(.A1(new_n2351_), .A2(new_n2353_), .B(new_n2352_), .ZN(new_n2374_));
  NOR2_X1    g01370(.A1(new_n2373_), .A2(new_n2374_), .ZN(new_n2375_));
  AOI21_X1   g01371(.A1(new_n2320_), .A2(new_n2328_), .B(new_n2326_), .ZN(new_n2376_));
  AOI21_X1   g01372(.A1(new_n2309_), .A2(new_n2315_), .B(new_n2316_), .ZN(new_n2377_));
  NOR2_X1    g01373(.A1(new_n2376_), .A2(new_n2377_), .ZN(new_n2378_));
  INV_X1     g01374(.I(new_n2378_), .ZN(new_n2379_));
  NOR3_X1    g01375(.A1(new_n2379_), .A2(new_n2319_), .A3(new_n2330_), .ZN(new_n2380_));
  NAND4_X1   g01376(.A1(new_n2380_), .A2(new_n2356_), .A3(new_n2370_), .A4(new_n2375_), .ZN(new_n2381_));
  NOR3_X1    g01377(.A1(new_n2381_), .A2(new_n2372_), .A3(new_n2345_), .ZN(new_n2382_));
  XNOR2_X1   g01378(.A1(new_n2370_), .A2(new_n2375_), .ZN(new_n2383_));
  NOR2_X1    g01379(.A1(new_n2383_), .A2(new_n2356_), .ZN(new_n2384_));
  XOR2_X1    g01380(.A1(new_n2370_), .A2(new_n2375_), .Z(new_n2385_));
  NOR2_X1    g01381(.A1(new_n2385_), .A2(new_n2357_), .ZN(new_n2386_));
  INV_X1     g01382(.I(new_n2375_), .ZN(new_n2387_));
  XNOR2_X1   g01383(.A1(new_n2356_), .A2(new_n2370_), .ZN(new_n2388_));
  NOR2_X1    g01384(.A1(new_n2388_), .A2(new_n2387_), .ZN(new_n2389_));
  NOR3_X1    g01385(.A1(new_n2389_), .A2(new_n2384_), .A3(new_n2386_), .ZN(new_n2390_));
  NAND2_X1   g01386(.A1(new_n2330_), .A2(new_n2378_), .ZN(new_n2391_));
  NAND2_X1   g01387(.A1(new_n2379_), .A2(new_n2343_), .ZN(new_n2392_));
  AOI21_X1   g01388(.A1(new_n2392_), .A2(new_n2391_), .B(new_n2337_), .ZN(new_n2393_));
  AND3_X2    g01389(.A1(new_n2392_), .A2(new_n2337_), .A3(new_n2391_), .Z(new_n2394_));
  NOR2_X1    g01390(.A1(new_n2394_), .A2(new_n2393_), .ZN(new_n2395_));
  NAND2_X1   g01391(.A1(new_n2337_), .A2(new_n2378_), .ZN(new_n2396_));
  OAI22_X1   g01392(.A1(new_n2331_), .A2(new_n2344_), .B1(new_n2396_), .B2(new_n2330_), .ZN(new_n2397_));
  NOR4_X1    g01393(.A1(new_n2397_), .A2(new_n2357_), .A3(new_n2368_), .A4(new_n2387_), .ZN(new_n2398_));
  NOR4_X1    g01394(.A1(new_n2390_), .A2(new_n2382_), .A3(new_n2395_), .A4(new_n2398_), .ZN(new_n2399_));
  NAND3_X1   g01395(.A1(new_n2272_), .A2(new_n2258_), .A3(new_n2268_), .ZN(new_n2400_));
  NOR3_X1    g01396(.A1(new_n2286_), .A2(new_n2241_), .A3(new_n2302_), .ZN(new_n2401_));
  XNOR2_X1   g01397(.A1(new_n2400_), .A2(new_n2401_), .ZN(new_n2402_));
  NAND3_X1   g01398(.A1(new_n2356_), .A2(new_n2370_), .A3(new_n2375_), .ZN(new_n2403_));
  NOR3_X1    g01399(.A1(new_n2379_), .A2(new_n2319_), .A3(new_n2330_), .ZN(new_n2404_));
  XOR2_X1    g01400(.A1(new_n2404_), .A2(new_n2403_), .Z(new_n2405_));
  INV_X1     g01401(.I(new_n2405_), .ZN(new_n2406_));
  NOR2_X1    g01402(.A1(new_n2402_), .A2(new_n2406_), .ZN(new_n2407_));
  NAND2_X1   g01403(.A1(new_n2399_), .A2(new_n2407_), .ZN(new_n2408_));
  NOR2_X1    g01404(.A1(new_n2308_), .A2(new_n2408_), .ZN(new_n2409_));
  XOR2_X1    g01405(.A1(new_n2303_), .A2(new_n2286_), .Z(new_n2410_));
  XOR2_X1    g01406(.A1(new_n2298_), .A2(new_n2291_), .Z(new_n2411_));
  NAND2_X1   g01407(.A1(new_n2411_), .A2(new_n2410_), .ZN(new_n2412_));
  INV_X1     g01408(.I(new_n2382_), .ZN(new_n2413_));
  NAND2_X1   g01409(.A1(new_n2385_), .A2(new_n2357_), .ZN(new_n2414_));
  NAND2_X1   g01410(.A1(new_n2383_), .A2(new_n2356_), .ZN(new_n2415_));
  XOR2_X1    g01411(.A1(new_n2356_), .A2(new_n2370_), .Z(new_n2416_));
  NAND2_X1   g01412(.A1(new_n2416_), .A2(new_n2375_), .ZN(new_n2417_));
  NAND3_X1   g01413(.A1(new_n2417_), .A2(new_n2415_), .A3(new_n2414_), .ZN(new_n2418_));
  INV_X1     g01414(.I(new_n2395_), .ZN(new_n2419_));
  INV_X1     g01415(.I(new_n2398_), .ZN(new_n2420_));
  NAND4_X1   g01416(.A1(new_n2413_), .A2(new_n2419_), .A3(new_n2420_), .A4(new_n2418_), .ZN(new_n2421_));
  XOR2_X1    g01417(.A1(new_n2400_), .A2(new_n2401_), .Z(new_n2422_));
  NAND2_X1   g01418(.A1(new_n2422_), .A2(new_n2405_), .ZN(new_n2423_));
  NOR2_X1    g01419(.A1(new_n2421_), .A2(new_n2423_), .ZN(new_n2424_));
  NOR2_X1    g01420(.A1(new_n2412_), .A2(new_n2424_), .ZN(new_n2425_));
  OAI21_X1   g01421(.A1(new_n2409_), .A2(new_n2425_), .B(new_n2306_), .ZN(new_n2426_));
  INV_X1     g01422(.I(\A[672] ), .ZN(new_n2427_));
  NOR2_X1    g01423(.A1(new_n2427_), .A2(\A[671] ), .ZN(new_n2428_));
  INV_X1     g01424(.I(\A[671] ), .ZN(new_n2429_));
  NOR2_X1    g01425(.A1(new_n2429_), .A2(\A[672] ), .ZN(new_n2430_));
  OAI21_X1   g01426(.A1(new_n2428_), .A2(new_n2430_), .B(\A[670] ), .ZN(new_n2431_));
  INV_X1     g01427(.I(\A[670] ), .ZN(new_n2432_));
  NAND2_X1   g01428(.A1(\A[671] ), .A2(\A[672] ), .ZN(new_n2433_));
  INV_X1     g01429(.I(new_n2433_), .ZN(new_n2434_));
  NOR2_X1    g01430(.A1(\A[671] ), .A2(\A[672] ), .ZN(new_n2435_));
  OAI21_X1   g01431(.A1(new_n2434_), .A2(new_n2435_), .B(new_n2432_), .ZN(new_n2436_));
  NAND2_X1   g01432(.A1(new_n2431_), .A2(new_n2436_), .ZN(new_n2437_));
  INV_X1     g01433(.I(\A[669] ), .ZN(new_n2438_));
  NOR2_X1    g01434(.A1(new_n2438_), .A2(\A[668] ), .ZN(new_n2439_));
  INV_X1     g01435(.I(\A[668] ), .ZN(new_n2440_));
  NOR2_X1    g01436(.A1(new_n2440_), .A2(\A[669] ), .ZN(new_n2441_));
  OAI21_X1   g01437(.A1(new_n2439_), .A2(new_n2441_), .B(\A[667] ), .ZN(new_n2442_));
  INV_X1     g01438(.I(\A[667] ), .ZN(new_n2443_));
  NAND2_X1   g01439(.A1(\A[668] ), .A2(\A[669] ), .ZN(new_n2444_));
  INV_X1     g01440(.I(new_n2444_), .ZN(new_n2445_));
  NOR2_X1    g01441(.A1(\A[668] ), .A2(\A[669] ), .ZN(new_n2446_));
  OAI21_X1   g01442(.A1(new_n2445_), .A2(new_n2446_), .B(new_n2443_), .ZN(new_n2447_));
  NAND2_X1   g01443(.A1(new_n2442_), .A2(new_n2447_), .ZN(new_n2448_));
  AOI21_X1   g01444(.A1(new_n2432_), .A2(new_n2433_), .B(new_n2435_), .ZN(new_n2449_));
  AOI21_X1   g01445(.A1(new_n2443_), .A2(new_n2444_), .B(new_n2446_), .ZN(new_n2450_));
  NOR2_X1    g01446(.A1(new_n2449_), .A2(new_n2450_), .ZN(new_n2451_));
  XOR2_X1    g01447(.A1(new_n2448_), .A2(new_n2451_), .Z(new_n2452_));
  XOR2_X1    g01448(.A1(new_n2452_), .A2(new_n2437_), .Z(new_n2453_));
  NAND2_X1   g01449(.A1(new_n2440_), .A2(\A[669] ), .ZN(new_n2454_));
  NAND2_X1   g01450(.A1(new_n2438_), .A2(\A[668] ), .ZN(new_n2455_));
  AOI21_X1   g01451(.A1(new_n2454_), .A2(new_n2455_), .B(new_n2443_), .ZN(new_n2456_));
  INV_X1     g01452(.I(new_n2446_), .ZN(new_n2457_));
  AOI21_X1   g01453(.A1(new_n2457_), .A2(new_n2444_), .B(\A[667] ), .ZN(new_n2458_));
  NOR2_X1    g01454(.A1(new_n2458_), .A2(new_n2456_), .ZN(new_n2459_));
  NAND2_X1   g01455(.A1(new_n2437_), .A2(new_n2451_), .ZN(new_n2460_));
  NOR2_X1    g01456(.A1(new_n2460_), .A2(new_n2459_), .ZN(new_n2461_));
  INV_X1     g01457(.I(\A[675] ), .ZN(new_n2462_));
  NOR2_X1    g01458(.A1(new_n2462_), .A2(\A[674] ), .ZN(new_n2463_));
  INV_X1     g01459(.I(\A[674] ), .ZN(new_n2464_));
  NOR2_X1    g01460(.A1(new_n2464_), .A2(\A[675] ), .ZN(new_n2465_));
  OAI21_X1   g01461(.A1(new_n2463_), .A2(new_n2465_), .B(\A[673] ), .ZN(new_n2466_));
  INV_X1     g01462(.I(\A[673] ), .ZN(new_n2467_));
  NOR2_X1    g01463(.A1(\A[674] ), .A2(\A[675] ), .ZN(new_n2468_));
  NAND2_X1   g01464(.A1(\A[674] ), .A2(\A[675] ), .ZN(new_n2469_));
  INV_X1     g01465(.I(new_n2469_), .ZN(new_n2470_));
  OAI21_X1   g01466(.A1(new_n2470_), .A2(new_n2468_), .B(new_n2467_), .ZN(new_n2471_));
  NAND2_X1   g01467(.A1(new_n2466_), .A2(new_n2471_), .ZN(new_n2472_));
  INV_X1     g01468(.I(\A[678] ), .ZN(new_n2473_));
  NOR2_X1    g01469(.A1(new_n2473_), .A2(\A[677] ), .ZN(new_n2474_));
  INV_X1     g01470(.I(\A[677] ), .ZN(new_n2475_));
  NOR2_X1    g01471(.A1(new_n2475_), .A2(\A[678] ), .ZN(new_n2476_));
  OAI21_X1   g01472(.A1(new_n2474_), .A2(new_n2476_), .B(\A[676] ), .ZN(new_n2477_));
  INV_X1     g01473(.I(\A[676] ), .ZN(new_n2478_));
  NAND2_X1   g01474(.A1(\A[677] ), .A2(\A[678] ), .ZN(new_n2479_));
  INV_X1     g01475(.I(new_n2479_), .ZN(new_n2480_));
  NOR2_X1    g01476(.A1(\A[677] ), .A2(\A[678] ), .ZN(new_n2481_));
  OAI21_X1   g01477(.A1(new_n2480_), .A2(new_n2481_), .B(new_n2478_), .ZN(new_n2482_));
  NAND2_X1   g01478(.A1(new_n2477_), .A2(new_n2482_), .ZN(new_n2483_));
  AOI21_X1   g01479(.A1(new_n2467_), .A2(new_n2469_), .B(new_n2468_), .ZN(new_n2484_));
  AOI21_X1   g01480(.A1(new_n2478_), .A2(new_n2479_), .B(new_n2481_), .ZN(new_n2485_));
  NOR2_X1    g01481(.A1(new_n2484_), .A2(new_n2485_), .ZN(new_n2486_));
  NAND4_X1   g01482(.A1(new_n2461_), .A2(new_n2472_), .A3(new_n2483_), .A4(new_n2486_), .ZN(new_n2487_));
  INV_X1     g01483(.I(new_n2472_), .ZN(new_n2488_));
  AND2_X2    g01484(.A1(new_n2477_), .A2(new_n2482_), .Z(new_n2489_));
  NOR2_X1    g01485(.A1(new_n2488_), .A2(new_n2489_), .ZN(new_n2490_));
  NOR2_X1    g01486(.A1(new_n2472_), .A2(new_n2483_), .ZN(new_n2491_));
  NOR2_X1    g01487(.A1(new_n2490_), .A2(new_n2491_), .ZN(new_n2492_));
  NAND2_X1   g01488(.A1(new_n2429_), .A2(\A[672] ), .ZN(new_n2493_));
  NAND2_X1   g01489(.A1(new_n2427_), .A2(\A[671] ), .ZN(new_n2494_));
  AOI21_X1   g01490(.A1(new_n2493_), .A2(new_n2494_), .B(new_n2432_), .ZN(new_n2495_));
  INV_X1     g01491(.I(new_n2435_), .ZN(new_n2496_));
  AOI21_X1   g01492(.A1(new_n2496_), .A2(new_n2433_), .B(\A[670] ), .ZN(new_n2497_));
  NOR2_X1    g01493(.A1(new_n2497_), .A2(new_n2495_), .ZN(new_n2498_));
  NOR2_X1    g01494(.A1(new_n2498_), .A2(new_n2459_), .ZN(new_n2499_));
  NOR2_X1    g01495(.A1(new_n2437_), .A2(new_n2448_), .ZN(new_n2500_));
  NOR2_X1    g01496(.A1(new_n2499_), .A2(new_n2500_), .ZN(new_n2501_));
  OR3_X2     g01497(.A1(new_n2487_), .A2(new_n2492_), .A3(new_n2501_), .Z(new_n2502_));
  XNOR2_X1   g01498(.A1(new_n2472_), .A2(new_n2486_), .ZN(new_n2503_));
  NOR2_X1    g01499(.A1(new_n2503_), .A2(new_n2483_), .ZN(new_n2504_));
  XOR2_X1    g01500(.A1(new_n2472_), .A2(new_n2486_), .Z(new_n2505_));
  NOR2_X1    g01501(.A1(new_n2505_), .A2(new_n2489_), .ZN(new_n2506_));
  INV_X1     g01502(.I(new_n2486_), .ZN(new_n2507_));
  XNOR2_X1   g01503(.A1(new_n2472_), .A2(new_n2483_), .ZN(new_n2508_));
  NOR2_X1    g01504(.A1(new_n2508_), .A2(new_n2507_), .ZN(new_n2509_));
  NOR3_X1    g01505(.A1(new_n2509_), .A2(new_n2504_), .A3(new_n2506_), .ZN(new_n2510_));
  NAND2_X1   g01506(.A1(new_n2502_), .A2(new_n2510_), .ZN(new_n2511_));
  NOR3_X1    g01507(.A1(new_n2487_), .A2(new_n2492_), .A3(new_n2501_), .ZN(new_n2512_));
  NAND2_X1   g01508(.A1(new_n2505_), .A2(new_n2489_), .ZN(new_n2513_));
  NAND2_X1   g01509(.A1(new_n2503_), .A2(new_n2483_), .ZN(new_n2514_));
  XOR2_X1    g01510(.A1(new_n2472_), .A2(new_n2483_), .Z(new_n2515_));
  NAND2_X1   g01511(.A1(new_n2515_), .A2(new_n2486_), .ZN(new_n2516_));
  NAND3_X1   g01512(.A1(new_n2516_), .A2(new_n2514_), .A3(new_n2513_), .ZN(new_n2517_));
  NAND2_X1   g01513(.A1(new_n2517_), .A2(new_n2512_), .ZN(new_n2518_));
  AOI21_X1   g01514(.A1(new_n2511_), .A2(new_n2518_), .B(new_n2453_), .ZN(new_n2519_));
  INV_X1     g01515(.I(new_n2519_), .ZN(new_n2520_));
  OAI22_X1   g01516(.A1(new_n2499_), .A2(new_n2500_), .B1(new_n2460_), .B2(new_n2459_), .ZN(new_n2521_));
  NOR4_X1    g01517(.A1(new_n2521_), .A2(new_n2488_), .A3(new_n2489_), .A4(new_n2507_), .ZN(new_n2522_));
  NAND2_X1   g01518(.A1(new_n2453_), .A2(new_n2522_), .ZN(new_n2523_));
  AOI21_X1   g01519(.A1(new_n2523_), .A2(new_n2517_), .B(new_n2502_), .ZN(new_n2524_));
  INV_X1     g01520(.I(\A[658] ), .ZN(new_n2525_));
  INV_X1     g01521(.I(\A[659] ), .ZN(new_n2526_));
  NAND2_X1   g01522(.A1(new_n2526_), .A2(\A[660] ), .ZN(new_n2527_));
  INV_X1     g01523(.I(\A[660] ), .ZN(new_n2528_));
  NAND2_X1   g01524(.A1(new_n2528_), .A2(\A[659] ), .ZN(new_n2529_));
  AOI21_X1   g01525(.A1(new_n2527_), .A2(new_n2529_), .B(new_n2525_), .ZN(new_n2530_));
  NAND2_X1   g01526(.A1(\A[659] ), .A2(\A[660] ), .ZN(new_n2531_));
  NOR2_X1    g01527(.A1(\A[659] ), .A2(\A[660] ), .ZN(new_n2532_));
  INV_X1     g01528(.I(new_n2532_), .ZN(new_n2533_));
  AOI21_X1   g01529(.A1(new_n2533_), .A2(new_n2531_), .B(\A[658] ), .ZN(new_n2534_));
  NOR2_X1    g01530(.A1(new_n2534_), .A2(new_n2530_), .ZN(new_n2535_));
  INV_X1     g01531(.I(\A[655] ), .ZN(new_n2536_));
  INV_X1     g01532(.I(\A[656] ), .ZN(new_n2537_));
  NAND2_X1   g01533(.A1(new_n2537_), .A2(\A[657] ), .ZN(new_n2538_));
  INV_X1     g01534(.I(\A[657] ), .ZN(new_n2539_));
  NAND2_X1   g01535(.A1(new_n2539_), .A2(\A[656] ), .ZN(new_n2540_));
  AOI21_X1   g01536(.A1(new_n2538_), .A2(new_n2540_), .B(new_n2536_), .ZN(new_n2541_));
  NOR2_X1    g01537(.A1(\A[656] ), .A2(\A[657] ), .ZN(new_n2542_));
  INV_X1     g01538(.I(new_n2542_), .ZN(new_n2543_));
  NAND2_X1   g01539(.A1(\A[656] ), .A2(\A[657] ), .ZN(new_n2544_));
  AOI21_X1   g01540(.A1(new_n2543_), .A2(new_n2544_), .B(\A[655] ), .ZN(new_n2545_));
  NOR2_X1    g01541(.A1(new_n2545_), .A2(new_n2541_), .ZN(new_n2546_));
  NOR2_X1    g01542(.A1(new_n2535_), .A2(new_n2546_), .ZN(new_n2547_));
  NOR2_X1    g01543(.A1(new_n2528_), .A2(\A[659] ), .ZN(new_n2548_));
  NOR2_X1    g01544(.A1(new_n2526_), .A2(\A[660] ), .ZN(new_n2549_));
  OAI21_X1   g01545(.A1(new_n2548_), .A2(new_n2549_), .B(\A[658] ), .ZN(new_n2550_));
  INV_X1     g01546(.I(new_n2531_), .ZN(new_n2551_));
  OAI21_X1   g01547(.A1(new_n2551_), .A2(new_n2532_), .B(new_n2525_), .ZN(new_n2552_));
  NAND2_X1   g01548(.A1(new_n2550_), .A2(new_n2552_), .ZN(new_n2553_));
  NOR2_X1    g01549(.A1(new_n2539_), .A2(\A[656] ), .ZN(new_n2554_));
  NOR2_X1    g01550(.A1(new_n2537_), .A2(\A[657] ), .ZN(new_n2555_));
  OAI21_X1   g01551(.A1(new_n2554_), .A2(new_n2555_), .B(\A[655] ), .ZN(new_n2556_));
  INV_X1     g01552(.I(new_n2544_), .ZN(new_n2557_));
  OAI21_X1   g01553(.A1(new_n2557_), .A2(new_n2542_), .B(new_n2536_), .ZN(new_n2558_));
  NAND2_X1   g01554(.A1(new_n2556_), .A2(new_n2558_), .ZN(new_n2559_));
  NOR2_X1    g01555(.A1(new_n2553_), .A2(new_n2559_), .ZN(new_n2560_));
  NOR2_X1    g01556(.A1(new_n2547_), .A2(new_n2560_), .ZN(new_n2561_));
  INV_X1     g01557(.I(\A[666] ), .ZN(new_n2562_));
  NOR2_X1    g01558(.A1(new_n2562_), .A2(\A[665] ), .ZN(new_n2563_));
  INV_X1     g01559(.I(\A[665] ), .ZN(new_n2564_));
  NOR2_X1    g01560(.A1(new_n2564_), .A2(\A[666] ), .ZN(new_n2565_));
  OAI21_X1   g01561(.A1(new_n2563_), .A2(new_n2565_), .B(\A[664] ), .ZN(new_n2566_));
  INV_X1     g01562(.I(\A[664] ), .ZN(new_n2567_));
  NOR2_X1    g01563(.A1(\A[665] ), .A2(\A[666] ), .ZN(new_n2568_));
  NAND2_X1   g01564(.A1(\A[665] ), .A2(\A[666] ), .ZN(new_n2569_));
  INV_X1     g01565(.I(new_n2569_), .ZN(new_n2570_));
  OAI21_X1   g01566(.A1(new_n2570_), .A2(new_n2568_), .B(new_n2567_), .ZN(new_n2571_));
  AND2_X2    g01567(.A1(new_n2566_), .A2(new_n2571_), .Z(new_n2572_));
  INV_X1     g01568(.I(\A[661] ), .ZN(new_n2573_));
  INV_X1     g01569(.I(\A[662] ), .ZN(new_n2574_));
  NAND2_X1   g01570(.A1(new_n2574_), .A2(\A[663] ), .ZN(new_n2575_));
  INV_X1     g01571(.I(\A[663] ), .ZN(new_n2576_));
  NAND2_X1   g01572(.A1(new_n2576_), .A2(\A[662] ), .ZN(new_n2577_));
  AOI21_X1   g01573(.A1(new_n2575_), .A2(new_n2577_), .B(new_n2573_), .ZN(new_n2578_));
  NOR2_X1    g01574(.A1(\A[662] ), .A2(\A[663] ), .ZN(new_n2579_));
  INV_X1     g01575(.I(new_n2579_), .ZN(new_n2580_));
  NAND2_X1   g01576(.A1(\A[662] ), .A2(\A[663] ), .ZN(new_n2581_));
  AOI21_X1   g01577(.A1(new_n2580_), .A2(new_n2581_), .B(\A[661] ), .ZN(new_n2582_));
  NOR2_X1    g01578(.A1(new_n2582_), .A2(new_n2578_), .ZN(new_n2583_));
  NOR2_X1    g01579(.A1(new_n2572_), .A2(new_n2583_), .ZN(new_n2584_));
  NAND2_X1   g01580(.A1(new_n2566_), .A2(new_n2571_), .ZN(new_n2585_));
  NOR2_X1    g01581(.A1(new_n2576_), .A2(\A[662] ), .ZN(new_n2586_));
  NOR2_X1    g01582(.A1(new_n2574_), .A2(\A[663] ), .ZN(new_n2587_));
  OAI21_X1   g01583(.A1(new_n2586_), .A2(new_n2587_), .B(\A[661] ), .ZN(new_n2588_));
  INV_X1     g01584(.I(new_n2581_), .ZN(new_n2589_));
  OAI21_X1   g01585(.A1(new_n2589_), .A2(new_n2579_), .B(new_n2573_), .ZN(new_n2590_));
  NAND2_X1   g01586(.A1(new_n2588_), .A2(new_n2590_), .ZN(new_n2591_));
  NOR2_X1    g01587(.A1(new_n2585_), .A2(new_n2591_), .ZN(new_n2592_));
  NOR2_X1    g01588(.A1(new_n2584_), .A2(new_n2592_), .ZN(new_n2593_));
  NOR2_X1    g01589(.A1(new_n2593_), .A2(new_n2561_), .ZN(new_n2594_));
  AOI21_X1   g01590(.A1(new_n2573_), .A2(new_n2581_), .B(new_n2579_), .ZN(new_n2595_));
  AOI21_X1   g01591(.A1(new_n2567_), .A2(new_n2569_), .B(new_n2568_), .ZN(new_n2596_));
  NOR2_X1    g01592(.A1(new_n2595_), .A2(new_n2596_), .ZN(new_n2597_));
  NAND3_X1   g01593(.A1(new_n2585_), .A2(new_n2591_), .A3(new_n2597_), .ZN(new_n2598_));
  AOI21_X1   g01594(.A1(new_n2536_), .A2(new_n2544_), .B(new_n2542_), .ZN(new_n2599_));
  AOI21_X1   g01595(.A1(new_n2525_), .A2(new_n2531_), .B(new_n2532_), .ZN(new_n2600_));
  NOR2_X1    g01596(.A1(new_n2599_), .A2(new_n2600_), .ZN(new_n2601_));
  NAND3_X1   g01597(.A1(new_n2553_), .A2(new_n2559_), .A3(new_n2601_), .ZN(new_n2602_));
  NOR2_X1    g01598(.A1(new_n2598_), .A2(new_n2602_), .ZN(new_n2603_));
  NAND2_X1   g01599(.A1(new_n2594_), .A2(new_n2603_), .ZN(new_n2604_));
  INV_X1     g01600(.I(new_n2597_), .ZN(new_n2605_));
  NOR2_X1    g01601(.A1(new_n2605_), .A2(new_n2591_), .ZN(new_n2606_));
  NOR2_X1    g01602(.A1(new_n2583_), .A2(new_n2597_), .ZN(new_n2607_));
  OAI21_X1   g01603(.A1(new_n2606_), .A2(new_n2607_), .B(new_n2572_), .ZN(new_n2608_));
  NAND2_X1   g01604(.A1(new_n2583_), .A2(new_n2597_), .ZN(new_n2609_));
  NAND2_X1   g01605(.A1(new_n2605_), .A2(new_n2591_), .ZN(new_n2610_));
  NAND3_X1   g01606(.A1(new_n2610_), .A2(new_n2609_), .A3(new_n2585_), .ZN(new_n2611_));
  NAND2_X1   g01607(.A1(new_n2608_), .A2(new_n2611_), .ZN(new_n2612_));
  XOR2_X1    g01608(.A1(new_n2583_), .A2(new_n2585_), .Z(new_n2613_));
  NOR2_X1    g01609(.A1(new_n2613_), .A2(new_n2605_), .ZN(new_n2614_));
  NOR2_X1    g01610(.A1(new_n2614_), .A2(new_n2612_), .ZN(new_n2615_));
  NAND2_X1   g01611(.A1(new_n2615_), .A2(new_n2604_), .ZN(new_n2616_));
  NAND2_X1   g01612(.A1(new_n2546_), .A2(new_n2601_), .ZN(new_n2617_));
  INV_X1     g01613(.I(new_n2601_), .ZN(new_n2618_));
  NAND2_X1   g01614(.A1(new_n2618_), .A2(new_n2559_), .ZN(new_n2619_));
  AOI21_X1   g01615(.A1(new_n2619_), .A2(new_n2617_), .B(new_n2553_), .ZN(new_n2620_));
  AND3_X2    g01616(.A1(new_n2619_), .A2(new_n2553_), .A3(new_n2617_), .Z(new_n2621_));
  NOR2_X1    g01617(.A1(new_n2621_), .A2(new_n2620_), .ZN(new_n2622_));
  INV_X1     g01618(.I(new_n2622_), .ZN(new_n2623_));
  XOR2_X1    g01619(.A1(new_n2535_), .A2(new_n2559_), .Z(new_n2624_));
  INV_X1     g01620(.I(new_n2602_), .ZN(new_n2625_));
  NAND4_X1   g01621(.A1(new_n2624_), .A2(new_n2585_), .A3(new_n2591_), .A4(new_n2597_), .ZN(new_n2626_));
  NAND3_X1   g01622(.A1(new_n2472_), .A2(new_n2483_), .A3(new_n2486_), .ZN(new_n2627_));
  OR2_X2     g01623(.A1(new_n2449_), .A2(new_n2450_), .Z(new_n2628_));
  NOR3_X1    g01624(.A1(new_n2628_), .A2(new_n2498_), .A3(new_n2459_), .ZN(new_n2629_));
  XNOR2_X1   g01625(.A1(new_n2629_), .A2(new_n2627_), .ZN(new_n2630_));
  NAND3_X1   g01626(.A1(new_n2585_), .A2(new_n2591_), .A3(new_n2597_), .ZN(new_n2631_));
  NOR3_X1    g01627(.A1(new_n2618_), .A2(new_n2535_), .A3(new_n2546_), .ZN(new_n2632_));
  XNOR2_X1   g01628(.A1(new_n2632_), .A2(new_n2631_), .ZN(new_n2633_));
  NOR2_X1    g01629(.A1(new_n2633_), .A2(new_n2630_), .ZN(new_n2634_));
  NAND4_X1   g01630(.A1(new_n2616_), .A2(new_n2623_), .A3(new_n2626_), .A4(new_n2634_), .ZN(new_n2635_));
  NOR2_X1    g01631(.A1(new_n2524_), .A2(new_n2635_), .ZN(new_n2636_));
  XOR2_X1    g01632(.A1(new_n2459_), .A2(new_n2451_), .Z(new_n2637_));
  NOR2_X1    g01633(.A1(new_n2637_), .A2(new_n2437_), .ZN(new_n2638_));
  NOR2_X1    g01634(.A1(new_n2452_), .A2(new_n2498_), .ZN(new_n2639_));
  NOR2_X1    g01635(.A1(new_n2638_), .A2(new_n2639_), .ZN(new_n2640_));
  INV_X1     g01636(.I(new_n2522_), .ZN(new_n2641_));
  NOR2_X1    g01637(.A1(new_n2641_), .A2(new_n2640_), .ZN(new_n2642_));
  OAI21_X1   g01638(.A1(new_n2642_), .A2(new_n2510_), .B(new_n2512_), .ZN(new_n2643_));
  XOR2_X1    g01639(.A1(new_n2585_), .A2(new_n2591_), .Z(new_n2644_));
  NAND2_X1   g01640(.A1(new_n2644_), .A2(new_n2597_), .ZN(new_n2645_));
  NAND3_X1   g01641(.A1(new_n2645_), .A2(new_n2608_), .A3(new_n2611_), .ZN(new_n2646_));
  NOR2_X1    g01642(.A1(new_n2561_), .A2(new_n2625_), .ZN(new_n2647_));
  NAND4_X1   g01643(.A1(new_n2647_), .A2(new_n2585_), .A3(new_n2591_), .A4(new_n2597_), .ZN(new_n2648_));
  NAND4_X1   g01644(.A1(new_n2623_), .A2(new_n2646_), .A3(new_n2648_), .A4(new_n2604_), .ZN(new_n2649_));
  OR2_X2     g01645(.A1(new_n2633_), .A2(new_n2630_), .Z(new_n2650_));
  NOR2_X1    g01646(.A1(new_n2649_), .A2(new_n2650_), .ZN(new_n2651_));
  NOR2_X1    g01647(.A1(new_n2651_), .A2(new_n2643_), .ZN(new_n2652_));
  OAI21_X1   g01648(.A1(new_n2652_), .A2(new_n2636_), .B(new_n2520_), .ZN(new_n2653_));
  NAND2_X1   g01649(.A1(new_n2651_), .A2(new_n2643_), .ZN(new_n2654_));
  NAND2_X1   g01650(.A1(new_n2524_), .A2(new_n2635_), .ZN(new_n2655_));
  NAND3_X1   g01651(.A1(new_n2654_), .A2(new_n2655_), .A3(new_n2519_), .ZN(new_n2656_));
  NOR2_X1    g01652(.A1(new_n2422_), .A2(new_n2405_), .ZN(new_n2657_));
  NOR2_X1    g01653(.A1(new_n2407_), .A2(new_n2657_), .ZN(new_n2658_));
  AND2_X2    g01654(.A1(new_n2633_), .A2(new_n2630_), .Z(new_n2659_));
  NOR2_X1    g01655(.A1(new_n2659_), .A2(new_n2634_), .ZN(new_n2660_));
  NAND2_X1   g01656(.A1(new_n2658_), .A2(new_n2660_), .ZN(new_n2661_));
  AOI21_X1   g01657(.A1(new_n2653_), .A2(new_n2656_), .B(new_n2661_), .ZN(new_n2662_));
  NAND2_X1   g01658(.A1(new_n2426_), .A2(new_n2662_), .ZN(new_n2663_));
  INV_X1     g01659(.I(new_n2306_), .ZN(new_n2664_));
  NAND2_X1   g01660(.A1(new_n2412_), .A2(new_n2424_), .ZN(new_n2665_));
  NAND2_X1   g01661(.A1(new_n2308_), .A2(new_n2408_), .ZN(new_n2666_));
  AOI21_X1   g01662(.A1(new_n2666_), .A2(new_n2665_), .B(new_n2664_), .ZN(new_n2667_));
  NAND2_X1   g01663(.A1(new_n2667_), .A2(new_n2662_), .ZN(new_n2668_));
  INV_X1     g01664(.I(new_n2228_), .ZN(new_n2669_));
  NOR2_X1    g01665(.A1(new_n2227_), .A2(new_n2225_), .ZN(new_n2670_));
  NOR2_X1    g01666(.A1(new_n2669_), .A2(new_n2670_), .ZN(new_n2671_));
  INV_X1     g01667(.I(new_n2661_), .ZN(new_n2672_));
  NOR2_X1    g01668(.A1(new_n2658_), .A2(new_n2660_), .ZN(new_n2673_));
  NOR2_X1    g01669(.A1(new_n2672_), .A2(new_n2673_), .ZN(new_n2674_));
  NAND2_X1   g01670(.A1(new_n2674_), .A2(new_n2671_), .ZN(new_n2675_));
  AOI21_X1   g01671(.A1(new_n2663_), .A2(new_n2668_), .B(new_n2675_), .ZN(new_n2676_));
  NAND2_X1   g01672(.A1(new_n2676_), .A2(new_n2231_), .ZN(new_n2677_));
  NAND2_X1   g01673(.A1(new_n2676_), .A2(new_n2230_), .ZN(new_n2678_));
  AND2_X2    g01674(.A1(new_n2677_), .A2(new_n2678_), .Z(new_n2679_));
  OAI21_X1   g01675(.A1(new_n1724_), .A2(new_n1818_), .B(new_n1820_), .ZN(new_n2680_));
  INV_X1     g01676(.I(new_n2675_), .ZN(new_n2681_));
  NOR2_X1    g01677(.A1(new_n2674_), .A2(new_n2671_), .ZN(new_n2682_));
  NOR2_X1    g01678(.A1(new_n2681_), .A2(new_n2682_), .ZN(new_n2683_));
  NAND3_X1   g01679(.A1(new_n2683_), .A2(new_n1822_), .A3(new_n2680_), .ZN(new_n2684_));
  NOR2_X1    g01680(.A1(new_n2679_), .A2(new_n2684_), .ZN(new_n2685_));
  NOR2_X1    g01681(.A1(new_n2685_), .A2(new_n1825_), .ZN(new_n2686_));
  NAND2_X1   g01682(.A1(new_n1822_), .A2(new_n2680_), .ZN(new_n2687_));
  OAI21_X1   g01683(.A1(new_n2681_), .A2(new_n2682_), .B(new_n2687_), .ZN(new_n2688_));
  NAND2_X1   g01684(.A1(new_n2688_), .A2(new_n2684_), .ZN(new_n2689_));
  INV_X1     g01685(.I(\A[471] ), .ZN(new_n2690_));
  NOR2_X1    g01686(.A1(new_n2690_), .A2(\A[470] ), .ZN(new_n2691_));
  INV_X1     g01687(.I(\A[470] ), .ZN(new_n2692_));
  NOR2_X1    g01688(.A1(new_n2692_), .A2(\A[471] ), .ZN(new_n2693_));
  OAI21_X1   g01689(.A1(new_n2691_), .A2(new_n2693_), .B(\A[469] ), .ZN(new_n2694_));
  INV_X1     g01690(.I(\A[469] ), .ZN(new_n2695_));
  NOR2_X1    g01691(.A1(\A[470] ), .A2(\A[471] ), .ZN(new_n2696_));
  NOR2_X1    g01692(.A1(new_n2692_), .A2(new_n2690_), .ZN(new_n2697_));
  OAI21_X1   g01693(.A1(new_n2697_), .A2(new_n2696_), .B(new_n2695_), .ZN(new_n2698_));
  NAND2_X1   g01694(.A1(new_n2698_), .A2(new_n2694_), .ZN(new_n2699_));
  INV_X1     g01695(.I(\A[474] ), .ZN(new_n2700_));
  NOR2_X1    g01696(.A1(new_n2700_), .A2(\A[473] ), .ZN(new_n2701_));
  INV_X1     g01697(.I(\A[473] ), .ZN(new_n2702_));
  NOR2_X1    g01698(.A1(new_n2702_), .A2(\A[474] ), .ZN(new_n2703_));
  OAI21_X1   g01699(.A1(new_n2701_), .A2(new_n2703_), .B(\A[472] ), .ZN(new_n2704_));
  INV_X1     g01700(.I(\A[472] ), .ZN(new_n2705_));
  NOR2_X1    g01701(.A1(\A[473] ), .A2(\A[474] ), .ZN(new_n2706_));
  NOR2_X1    g01702(.A1(new_n2702_), .A2(new_n2700_), .ZN(new_n2707_));
  OAI21_X1   g01703(.A1(new_n2707_), .A2(new_n2706_), .B(new_n2705_), .ZN(new_n2708_));
  NAND2_X1   g01704(.A1(new_n2708_), .A2(new_n2704_), .ZN(new_n2709_));
  NOR2_X1    g01705(.A1(new_n2697_), .A2(\A[469] ), .ZN(new_n2710_));
  NOR2_X1    g01706(.A1(new_n2710_), .A2(new_n2696_), .ZN(new_n2711_));
  NOR2_X1    g01707(.A1(new_n2707_), .A2(\A[472] ), .ZN(new_n2712_));
  NOR2_X1    g01708(.A1(new_n2712_), .A2(new_n2706_), .ZN(new_n2713_));
  NOR2_X1    g01709(.A1(new_n2711_), .A2(new_n2713_), .ZN(new_n2714_));
  NAND3_X1   g01710(.A1(new_n2714_), .A2(new_n2699_), .A3(new_n2709_), .ZN(new_n2715_));
  INV_X1     g01711(.I(\A[466] ), .ZN(new_n2716_));
  INV_X1     g01712(.I(\A[467] ), .ZN(new_n2717_));
  NAND2_X1   g01713(.A1(new_n2717_), .A2(\A[468] ), .ZN(new_n2718_));
  INV_X1     g01714(.I(\A[468] ), .ZN(new_n2719_));
  NAND2_X1   g01715(.A1(new_n2719_), .A2(\A[467] ), .ZN(new_n2720_));
  AOI21_X1   g01716(.A1(new_n2718_), .A2(new_n2720_), .B(new_n2716_), .ZN(new_n2721_));
  NAND2_X1   g01717(.A1(\A[467] ), .A2(\A[468] ), .ZN(new_n2722_));
  NAND2_X1   g01718(.A1(new_n2717_), .A2(new_n2719_), .ZN(new_n2723_));
  AOI21_X1   g01719(.A1(new_n2723_), .A2(new_n2722_), .B(\A[466] ), .ZN(new_n2724_));
  NOR2_X1    g01720(.A1(new_n2724_), .A2(new_n2721_), .ZN(new_n2725_));
  INV_X1     g01721(.I(\A[463] ), .ZN(new_n2726_));
  INV_X1     g01722(.I(\A[464] ), .ZN(new_n2727_));
  NAND2_X1   g01723(.A1(new_n2727_), .A2(\A[465] ), .ZN(new_n2728_));
  INV_X1     g01724(.I(\A[465] ), .ZN(new_n2729_));
  NAND2_X1   g01725(.A1(new_n2729_), .A2(\A[464] ), .ZN(new_n2730_));
  AOI21_X1   g01726(.A1(new_n2728_), .A2(new_n2730_), .B(new_n2726_), .ZN(new_n2731_));
  NAND2_X1   g01727(.A1(new_n2727_), .A2(new_n2729_), .ZN(new_n2732_));
  NAND2_X1   g01728(.A1(\A[464] ), .A2(\A[465] ), .ZN(new_n2733_));
  AOI21_X1   g01729(.A1(new_n2732_), .A2(new_n2733_), .B(\A[463] ), .ZN(new_n2734_));
  NOR2_X1    g01730(.A1(new_n2734_), .A2(new_n2731_), .ZN(new_n2735_));
  NAND2_X1   g01731(.A1(new_n2733_), .A2(new_n2726_), .ZN(new_n2736_));
  NAND2_X1   g01732(.A1(new_n2736_), .A2(new_n2732_), .ZN(new_n2737_));
  NAND2_X1   g01733(.A1(new_n2722_), .A2(new_n2716_), .ZN(new_n2738_));
  NAND2_X1   g01734(.A1(new_n2738_), .A2(new_n2723_), .ZN(new_n2739_));
  NAND2_X1   g01735(.A1(new_n2737_), .A2(new_n2739_), .ZN(new_n2740_));
  NOR3_X1    g01736(.A1(new_n2725_), .A2(new_n2735_), .A3(new_n2740_), .ZN(new_n2741_));
  XOR2_X1    g01737(.A1(new_n2715_), .A2(new_n2741_), .Z(new_n2742_));
  INV_X1     g01738(.I(\A[483] ), .ZN(new_n2743_));
  NOR2_X1    g01739(.A1(new_n2743_), .A2(\A[482] ), .ZN(new_n2744_));
  INV_X1     g01740(.I(\A[482] ), .ZN(new_n2745_));
  NOR2_X1    g01741(.A1(new_n2745_), .A2(\A[483] ), .ZN(new_n2746_));
  OAI21_X1   g01742(.A1(new_n2744_), .A2(new_n2746_), .B(\A[481] ), .ZN(new_n2747_));
  INV_X1     g01743(.I(\A[481] ), .ZN(new_n2748_));
  NOR2_X1    g01744(.A1(\A[482] ), .A2(\A[483] ), .ZN(new_n2749_));
  NAND2_X1   g01745(.A1(\A[482] ), .A2(\A[483] ), .ZN(new_n2750_));
  INV_X1     g01746(.I(new_n2750_), .ZN(new_n2751_));
  OAI21_X1   g01747(.A1(new_n2751_), .A2(new_n2749_), .B(new_n2748_), .ZN(new_n2752_));
  NAND2_X1   g01748(.A1(new_n2747_), .A2(new_n2752_), .ZN(new_n2753_));
  INV_X1     g01749(.I(\A[486] ), .ZN(new_n2754_));
  NOR2_X1    g01750(.A1(new_n2754_), .A2(\A[485] ), .ZN(new_n2755_));
  INV_X1     g01751(.I(\A[485] ), .ZN(new_n2756_));
  NOR2_X1    g01752(.A1(new_n2756_), .A2(\A[486] ), .ZN(new_n2757_));
  OAI21_X1   g01753(.A1(new_n2755_), .A2(new_n2757_), .B(\A[484] ), .ZN(new_n2758_));
  INV_X1     g01754(.I(\A[484] ), .ZN(new_n2759_));
  NAND2_X1   g01755(.A1(\A[485] ), .A2(\A[486] ), .ZN(new_n2760_));
  INV_X1     g01756(.I(new_n2760_), .ZN(new_n2761_));
  NOR2_X1    g01757(.A1(\A[485] ), .A2(\A[486] ), .ZN(new_n2762_));
  OAI21_X1   g01758(.A1(new_n2761_), .A2(new_n2762_), .B(new_n2759_), .ZN(new_n2763_));
  NAND2_X1   g01759(.A1(new_n2758_), .A2(new_n2763_), .ZN(new_n2764_));
  AOI21_X1   g01760(.A1(new_n2748_), .A2(new_n2750_), .B(new_n2749_), .ZN(new_n2765_));
  AOI21_X1   g01761(.A1(new_n2759_), .A2(new_n2760_), .B(new_n2762_), .ZN(new_n2766_));
  NOR2_X1    g01762(.A1(new_n2765_), .A2(new_n2766_), .ZN(new_n2767_));
  NAND3_X1   g01763(.A1(new_n2753_), .A2(new_n2764_), .A3(new_n2767_), .ZN(new_n2768_));
  INV_X1     g01764(.I(\A[475] ), .ZN(new_n2769_));
  INV_X1     g01765(.I(\A[476] ), .ZN(new_n2770_));
  NAND2_X1   g01766(.A1(new_n2770_), .A2(\A[477] ), .ZN(new_n2771_));
  INV_X1     g01767(.I(\A[477] ), .ZN(new_n2772_));
  NAND2_X1   g01768(.A1(new_n2772_), .A2(\A[476] ), .ZN(new_n2773_));
  AOI21_X1   g01769(.A1(new_n2771_), .A2(new_n2773_), .B(new_n2769_), .ZN(new_n2774_));
  NAND2_X1   g01770(.A1(new_n2770_), .A2(new_n2772_), .ZN(new_n2775_));
  NAND2_X1   g01771(.A1(\A[476] ), .A2(\A[477] ), .ZN(new_n2776_));
  AOI21_X1   g01772(.A1(new_n2775_), .A2(new_n2776_), .B(\A[475] ), .ZN(new_n2777_));
  NOR2_X1    g01773(.A1(new_n2777_), .A2(new_n2774_), .ZN(new_n2778_));
  INV_X1     g01774(.I(\A[478] ), .ZN(new_n2779_));
  INV_X1     g01775(.I(\A[479] ), .ZN(new_n2780_));
  NAND2_X1   g01776(.A1(new_n2780_), .A2(\A[480] ), .ZN(new_n2781_));
  INV_X1     g01777(.I(\A[480] ), .ZN(new_n2782_));
  NAND2_X1   g01778(.A1(new_n2782_), .A2(\A[479] ), .ZN(new_n2783_));
  AOI21_X1   g01779(.A1(new_n2781_), .A2(new_n2783_), .B(new_n2779_), .ZN(new_n2784_));
  NAND2_X1   g01780(.A1(\A[479] ), .A2(\A[480] ), .ZN(new_n2785_));
  NAND2_X1   g01781(.A1(new_n2780_), .A2(new_n2782_), .ZN(new_n2786_));
  AOI21_X1   g01782(.A1(new_n2786_), .A2(new_n2785_), .B(\A[478] ), .ZN(new_n2787_));
  NOR2_X1    g01783(.A1(new_n2787_), .A2(new_n2784_), .ZN(new_n2788_));
  NAND2_X1   g01784(.A1(new_n2776_), .A2(new_n2769_), .ZN(new_n2789_));
  NAND2_X1   g01785(.A1(new_n2789_), .A2(new_n2775_), .ZN(new_n2790_));
  NAND2_X1   g01786(.A1(new_n2785_), .A2(new_n2779_), .ZN(new_n2791_));
  NAND2_X1   g01787(.A1(new_n2791_), .A2(new_n2786_), .ZN(new_n2792_));
  NAND2_X1   g01788(.A1(new_n2790_), .A2(new_n2792_), .ZN(new_n2793_));
  NOR3_X1    g01789(.A1(new_n2778_), .A2(new_n2788_), .A3(new_n2793_), .ZN(new_n2794_));
  XOR2_X1    g01790(.A1(new_n2794_), .A2(new_n2768_), .Z(new_n2795_));
  NAND2_X1   g01791(.A1(new_n2742_), .A2(new_n2795_), .ZN(new_n2796_));
  INV_X1     g01792(.I(new_n2796_), .ZN(new_n2797_));
  NOR2_X1    g01793(.A1(new_n2742_), .A2(new_n2795_), .ZN(new_n2798_));
  NOR2_X1    g01794(.A1(new_n2797_), .A2(new_n2798_), .ZN(new_n2799_));
  INV_X1     g01795(.I(\A[507] ), .ZN(new_n2800_));
  NOR2_X1    g01796(.A1(new_n2800_), .A2(\A[506] ), .ZN(new_n2801_));
  INV_X1     g01797(.I(\A[506] ), .ZN(new_n2802_));
  NOR2_X1    g01798(.A1(new_n2802_), .A2(\A[507] ), .ZN(new_n2803_));
  OAI21_X1   g01799(.A1(new_n2801_), .A2(new_n2803_), .B(\A[505] ), .ZN(new_n2804_));
  NOR2_X1    g01800(.A1(\A[506] ), .A2(\A[507] ), .ZN(new_n2805_));
  NOR2_X1    g01801(.A1(new_n2802_), .A2(new_n2800_), .ZN(new_n2806_));
  NOR2_X1    g01802(.A1(new_n2806_), .A2(new_n2805_), .ZN(new_n2807_));
  OAI21_X1   g01803(.A1(\A[505] ), .A2(new_n2807_), .B(new_n2804_), .ZN(new_n2808_));
  INV_X1     g01804(.I(\A[510] ), .ZN(new_n2809_));
  NOR2_X1    g01805(.A1(new_n2809_), .A2(\A[509] ), .ZN(new_n2810_));
  INV_X1     g01806(.I(\A[509] ), .ZN(new_n2811_));
  NOR2_X1    g01807(.A1(new_n2811_), .A2(\A[510] ), .ZN(new_n2812_));
  OAI21_X1   g01808(.A1(new_n2810_), .A2(new_n2812_), .B(\A[508] ), .ZN(new_n2813_));
  INV_X1     g01809(.I(\A[508] ), .ZN(new_n2814_));
  NOR2_X1    g01810(.A1(new_n2811_), .A2(new_n2809_), .ZN(new_n2815_));
  NOR2_X1    g01811(.A1(\A[509] ), .A2(\A[510] ), .ZN(new_n2816_));
  OAI21_X1   g01812(.A1(new_n2815_), .A2(new_n2816_), .B(new_n2814_), .ZN(new_n2817_));
  NAND2_X1   g01813(.A1(new_n2817_), .A2(new_n2813_), .ZN(new_n2818_));
  NOR2_X1    g01814(.A1(new_n2806_), .A2(\A[505] ), .ZN(new_n2819_));
  NOR2_X1    g01815(.A1(new_n2815_), .A2(\A[508] ), .ZN(new_n2820_));
  OAI22_X1   g01816(.A1(new_n2805_), .A2(new_n2819_), .B1(new_n2820_), .B2(new_n2816_), .ZN(new_n2821_));
  INV_X1     g01817(.I(new_n2821_), .ZN(new_n2822_));
  NAND3_X1   g01818(.A1(new_n2822_), .A2(new_n2808_), .A3(new_n2818_), .ZN(new_n2823_));
  INV_X1     g01819(.I(\A[499] ), .ZN(new_n2824_));
  INV_X1     g01820(.I(\A[500] ), .ZN(new_n2825_));
  NAND2_X1   g01821(.A1(new_n2825_), .A2(\A[501] ), .ZN(new_n2826_));
  INV_X1     g01822(.I(\A[501] ), .ZN(new_n2827_));
  NAND2_X1   g01823(.A1(new_n2827_), .A2(\A[500] ), .ZN(new_n2828_));
  AOI21_X1   g01824(.A1(new_n2826_), .A2(new_n2828_), .B(new_n2824_), .ZN(new_n2829_));
  NAND2_X1   g01825(.A1(new_n2825_), .A2(new_n2827_), .ZN(new_n2830_));
  NAND2_X1   g01826(.A1(\A[500] ), .A2(\A[501] ), .ZN(new_n2831_));
  AOI21_X1   g01827(.A1(new_n2830_), .A2(new_n2831_), .B(\A[499] ), .ZN(new_n2832_));
  NOR2_X1    g01828(.A1(new_n2832_), .A2(new_n2829_), .ZN(new_n2833_));
  INV_X1     g01829(.I(\A[502] ), .ZN(new_n2834_));
  INV_X1     g01830(.I(\A[503] ), .ZN(new_n2835_));
  NAND2_X1   g01831(.A1(new_n2835_), .A2(\A[504] ), .ZN(new_n2836_));
  INV_X1     g01832(.I(\A[504] ), .ZN(new_n2837_));
  NAND2_X1   g01833(.A1(new_n2837_), .A2(\A[503] ), .ZN(new_n2838_));
  AOI21_X1   g01834(.A1(new_n2836_), .A2(new_n2838_), .B(new_n2834_), .ZN(new_n2839_));
  NAND2_X1   g01835(.A1(\A[503] ), .A2(\A[504] ), .ZN(new_n2840_));
  NAND2_X1   g01836(.A1(new_n2835_), .A2(new_n2837_), .ZN(new_n2841_));
  AOI21_X1   g01837(.A1(new_n2841_), .A2(new_n2840_), .B(\A[502] ), .ZN(new_n2842_));
  NOR2_X1    g01838(.A1(new_n2842_), .A2(new_n2839_), .ZN(new_n2843_));
  NAND2_X1   g01839(.A1(new_n2831_), .A2(new_n2824_), .ZN(new_n2844_));
  NAND2_X1   g01840(.A1(new_n2844_), .A2(new_n2830_), .ZN(new_n2845_));
  NAND2_X1   g01841(.A1(new_n2840_), .A2(new_n2834_), .ZN(new_n2846_));
  NAND2_X1   g01842(.A1(new_n2846_), .A2(new_n2841_), .ZN(new_n2847_));
  NAND2_X1   g01843(.A1(new_n2845_), .A2(new_n2847_), .ZN(new_n2848_));
  NOR3_X1    g01844(.A1(new_n2833_), .A2(new_n2843_), .A3(new_n2848_), .ZN(new_n2849_));
  XOR2_X1    g01845(.A1(new_n2823_), .A2(new_n2849_), .Z(new_n2850_));
  INV_X1     g01846(.I(\A[495] ), .ZN(new_n2851_));
  NOR2_X1    g01847(.A1(new_n2851_), .A2(\A[494] ), .ZN(new_n2852_));
  INV_X1     g01848(.I(\A[494] ), .ZN(new_n2853_));
  NOR2_X1    g01849(.A1(new_n2853_), .A2(\A[495] ), .ZN(new_n2854_));
  OAI21_X1   g01850(.A1(new_n2852_), .A2(new_n2854_), .B(\A[493] ), .ZN(new_n2855_));
  INV_X1     g01851(.I(\A[493] ), .ZN(new_n2856_));
  NOR2_X1    g01852(.A1(\A[494] ), .A2(\A[495] ), .ZN(new_n2857_));
  NOR2_X1    g01853(.A1(new_n2853_), .A2(new_n2851_), .ZN(new_n2858_));
  OAI21_X1   g01854(.A1(new_n2858_), .A2(new_n2857_), .B(new_n2856_), .ZN(new_n2859_));
  NAND2_X1   g01855(.A1(new_n2859_), .A2(new_n2855_), .ZN(new_n2860_));
  INV_X1     g01856(.I(\A[498] ), .ZN(new_n2861_));
  NOR2_X1    g01857(.A1(new_n2861_), .A2(\A[497] ), .ZN(new_n2862_));
  INV_X1     g01858(.I(\A[497] ), .ZN(new_n2863_));
  NOR2_X1    g01859(.A1(new_n2863_), .A2(\A[498] ), .ZN(new_n2864_));
  OAI21_X1   g01860(.A1(new_n2862_), .A2(new_n2864_), .B(\A[496] ), .ZN(new_n2865_));
  INV_X1     g01861(.I(\A[496] ), .ZN(new_n2866_));
  NOR2_X1    g01862(.A1(\A[497] ), .A2(\A[498] ), .ZN(new_n2867_));
  NOR2_X1    g01863(.A1(new_n2863_), .A2(new_n2861_), .ZN(new_n2868_));
  OAI21_X1   g01864(.A1(new_n2868_), .A2(new_n2867_), .B(new_n2866_), .ZN(new_n2869_));
  NAND2_X1   g01865(.A1(new_n2869_), .A2(new_n2865_), .ZN(new_n2870_));
  NOR2_X1    g01866(.A1(new_n2858_), .A2(\A[493] ), .ZN(new_n2871_));
  NOR2_X1    g01867(.A1(new_n2868_), .A2(\A[496] ), .ZN(new_n2872_));
  OAI22_X1   g01868(.A1(new_n2857_), .A2(new_n2871_), .B1(new_n2872_), .B2(new_n2867_), .ZN(new_n2873_));
  INV_X1     g01869(.I(new_n2873_), .ZN(new_n2874_));
  NAND3_X1   g01870(.A1(new_n2874_), .A2(new_n2860_), .A3(new_n2870_), .ZN(new_n2875_));
  INV_X1     g01871(.I(\A[487] ), .ZN(new_n2876_));
  INV_X1     g01872(.I(\A[488] ), .ZN(new_n2877_));
  NAND2_X1   g01873(.A1(new_n2877_), .A2(\A[489] ), .ZN(new_n2878_));
  INV_X1     g01874(.I(\A[489] ), .ZN(new_n2879_));
  NAND2_X1   g01875(.A1(new_n2879_), .A2(\A[488] ), .ZN(new_n2880_));
  AOI21_X1   g01876(.A1(new_n2878_), .A2(new_n2880_), .B(new_n2876_), .ZN(new_n2881_));
  NAND2_X1   g01877(.A1(new_n2877_), .A2(new_n2879_), .ZN(new_n2882_));
  NAND2_X1   g01878(.A1(\A[488] ), .A2(\A[489] ), .ZN(new_n2883_));
  AOI21_X1   g01879(.A1(new_n2882_), .A2(new_n2883_), .B(\A[487] ), .ZN(new_n2884_));
  NOR2_X1    g01880(.A1(new_n2884_), .A2(new_n2881_), .ZN(new_n2885_));
  INV_X1     g01881(.I(\A[490] ), .ZN(new_n2886_));
  INV_X1     g01882(.I(\A[491] ), .ZN(new_n2887_));
  NAND2_X1   g01883(.A1(new_n2887_), .A2(\A[492] ), .ZN(new_n2888_));
  INV_X1     g01884(.I(\A[492] ), .ZN(new_n2889_));
  NAND2_X1   g01885(.A1(new_n2889_), .A2(\A[491] ), .ZN(new_n2890_));
  AOI21_X1   g01886(.A1(new_n2888_), .A2(new_n2890_), .B(new_n2886_), .ZN(new_n2891_));
  NAND2_X1   g01887(.A1(\A[491] ), .A2(\A[492] ), .ZN(new_n2892_));
  NAND2_X1   g01888(.A1(new_n2887_), .A2(new_n2889_), .ZN(new_n2893_));
  AOI21_X1   g01889(.A1(new_n2893_), .A2(new_n2892_), .B(\A[490] ), .ZN(new_n2894_));
  NOR2_X1    g01890(.A1(new_n2894_), .A2(new_n2891_), .ZN(new_n2895_));
  NAND2_X1   g01891(.A1(new_n2883_), .A2(new_n2876_), .ZN(new_n2896_));
  NAND2_X1   g01892(.A1(new_n2896_), .A2(new_n2882_), .ZN(new_n2897_));
  NAND2_X1   g01893(.A1(new_n2892_), .A2(new_n2886_), .ZN(new_n2898_));
  NAND2_X1   g01894(.A1(new_n2898_), .A2(new_n2893_), .ZN(new_n2899_));
  NAND2_X1   g01895(.A1(new_n2897_), .A2(new_n2899_), .ZN(new_n2900_));
  NOR3_X1    g01896(.A1(new_n2885_), .A2(new_n2895_), .A3(new_n2900_), .ZN(new_n2901_));
  XOR2_X1    g01897(.A1(new_n2875_), .A2(new_n2901_), .Z(new_n2902_));
  AND2_X2    g01898(.A1(new_n2850_), .A2(new_n2902_), .Z(new_n2903_));
  NOR2_X1    g01899(.A1(new_n2850_), .A2(new_n2902_), .ZN(new_n2904_));
  NOR2_X1    g01900(.A1(new_n2903_), .A2(new_n2904_), .ZN(new_n2905_));
  NAND2_X1   g01901(.A1(new_n2905_), .A2(new_n2799_), .ZN(new_n2906_));
  INV_X1     g01902(.I(new_n2906_), .ZN(new_n2907_));
  NOR2_X1    g01903(.A1(new_n2905_), .A2(new_n2799_), .ZN(new_n2908_));
  NOR2_X1    g01904(.A1(new_n2907_), .A2(new_n2908_), .ZN(new_n2909_));
  INV_X1     g01905(.I(\A[555] ), .ZN(new_n2910_));
  NOR2_X1    g01906(.A1(new_n2910_), .A2(\A[554] ), .ZN(new_n2911_));
  INV_X1     g01907(.I(\A[554] ), .ZN(new_n2912_));
  NOR2_X1    g01908(.A1(new_n2912_), .A2(\A[555] ), .ZN(new_n2913_));
  OAI21_X1   g01909(.A1(new_n2911_), .A2(new_n2913_), .B(\A[553] ), .ZN(new_n2914_));
  INV_X1     g01910(.I(\A[553] ), .ZN(new_n2915_));
  NOR2_X1    g01911(.A1(\A[554] ), .A2(\A[555] ), .ZN(new_n2916_));
  NAND2_X1   g01912(.A1(\A[554] ), .A2(\A[555] ), .ZN(new_n2917_));
  INV_X1     g01913(.I(new_n2917_), .ZN(new_n2918_));
  OAI21_X1   g01914(.A1(new_n2918_), .A2(new_n2916_), .B(new_n2915_), .ZN(new_n2919_));
  NAND2_X1   g01915(.A1(new_n2914_), .A2(new_n2919_), .ZN(new_n2920_));
  INV_X1     g01916(.I(\A[558] ), .ZN(new_n2921_));
  NOR2_X1    g01917(.A1(new_n2921_), .A2(\A[557] ), .ZN(new_n2922_));
  INV_X1     g01918(.I(\A[557] ), .ZN(new_n2923_));
  NOR2_X1    g01919(.A1(new_n2923_), .A2(\A[558] ), .ZN(new_n2924_));
  OAI21_X1   g01920(.A1(new_n2922_), .A2(new_n2924_), .B(\A[556] ), .ZN(new_n2925_));
  INV_X1     g01921(.I(\A[556] ), .ZN(new_n2926_));
  NAND2_X1   g01922(.A1(\A[557] ), .A2(\A[558] ), .ZN(new_n2927_));
  INV_X1     g01923(.I(new_n2927_), .ZN(new_n2928_));
  NOR2_X1    g01924(.A1(\A[557] ), .A2(\A[558] ), .ZN(new_n2929_));
  OAI21_X1   g01925(.A1(new_n2928_), .A2(new_n2929_), .B(new_n2926_), .ZN(new_n2930_));
  NAND2_X1   g01926(.A1(new_n2925_), .A2(new_n2930_), .ZN(new_n2931_));
  AOI21_X1   g01927(.A1(new_n2915_), .A2(new_n2917_), .B(new_n2916_), .ZN(new_n2932_));
  AOI21_X1   g01928(.A1(new_n2926_), .A2(new_n2927_), .B(new_n2929_), .ZN(new_n2933_));
  NOR2_X1    g01929(.A1(new_n2932_), .A2(new_n2933_), .ZN(new_n2934_));
  NAND3_X1   g01930(.A1(new_n2920_), .A2(new_n2931_), .A3(new_n2934_), .ZN(new_n2935_));
  INV_X1     g01931(.I(\A[547] ), .ZN(new_n2936_));
  INV_X1     g01932(.I(\A[548] ), .ZN(new_n2937_));
  NAND2_X1   g01933(.A1(new_n2937_), .A2(\A[549] ), .ZN(new_n2938_));
  INV_X1     g01934(.I(\A[549] ), .ZN(new_n2939_));
  NAND2_X1   g01935(.A1(new_n2939_), .A2(\A[548] ), .ZN(new_n2940_));
  AOI21_X1   g01936(.A1(new_n2938_), .A2(new_n2940_), .B(new_n2936_), .ZN(new_n2941_));
  NAND2_X1   g01937(.A1(new_n2937_), .A2(new_n2939_), .ZN(new_n2942_));
  NAND2_X1   g01938(.A1(\A[548] ), .A2(\A[549] ), .ZN(new_n2943_));
  AOI21_X1   g01939(.A1(new_n2942_), .A2(new_n2943_), .B(\A[547] ), .ZN(new_n2944_));
  NOR2_X1    g01940(.A1(new_n2944_), .A2(new_n2941_), .ZN(new_n2945_));
  INV_X1     g01941(.I(\A[550] ), .ZN(new_n2946_));
  INV_X1     g01942(.I(\A[551] ), .ZN(new_n2947_));
  NAND2_X1   g01943(.A1(new_n2947_), .A2(\A[552] ), .ZN(new_n2948_));
  INV_X1     g01944(.I(\A[552] ), .ZN(new_n2949_));
  NAND2_X1   g01945(.A1(new_n2949_), .A2(\A[551] ), .ZN(new_n2950_));
  AOI21_X1   g01946(.A1(new_n2948_), .A2(new_n2950_), .B(new_n2946_), .ZN(new_n2951_));
  NAND2_X1   g01947(.A1(\A[551] ), .A2(\A[552] ), .ZN(new_n2952_));
  NAND2_X1   g01948(.A1(new_n2947_), .A2(new_n2949_), .ZN(new_n2953_));
  AOI21_X1   g01949(.A1(new_n2953_), .A2(new_n2952_), .B(\A[550] ), .ZN(new_n2954_));
  NOR2_X1    g01950(.A1(new_n2954_), .A2(new_n2951_), .ZN(new_n2955_));
  NAND2_X1   g01951(.A1(new_n2943_), .A2(new_n2936_), .ZN(new_n2956_));
  NAND2_X1   g01952(.A1(new_n2956_), .A2(new_n2942_), .ZN(new_n2957_));
  NAND2_X1   g01953(.A1(new_n2952_), .A2(new_n2946_), .ZN(new_n2958_));
  NAND2_X1   g01954(.A1(new_n2958_), .A2(new_n2953_), .ZN(new_n2959_));
  NAND2_X1   g01955(.A1(new_n2957_), .A2(new_n2959_), .ZN(new_n2960_));
  NOR3_X1    g01956(.A1(new_n2945_), .A2(new_n2955_), .A3(new_n2960_), .ZN(new_n2961_));
  XOR2_X1    g01957(.A1(new_n2961_), .A2(new_n2935_), .Z(new_n2962_));
  INV_X1     g01958(.I(\A[543] ), .ZN(new_n2963_));
  NOR2_X1    g01959(.A1(new_n2963_), .A2(\A[542] ), .ZN(new_n2964_));
  INV_X1     g01960(.I(\A[542] ), .ZN(new_n2965_));
  NOR2_X1    g01961(.A1(new_n2965_), .A2(\A[543] ), .ZN(new_n2966_));
  OAI21_X1   g01962(.A1(new_n2964_), .A2(new_n2966_), .B(\A[541] ), .ZN(new_n2967_));
  INV_X1     g01963(.I(\A[541] ), .ZN(new_n2968_));
  NOR2_X1    g01964(.A1(new_n2965_), .A2(new_n2963_), .ZN(new_n2969_));
  NOR2_X1    g01965(.A1(\A[542] ), .A2(\A[543] ), .ZN(new_n2970_));
  OAI21_X1   g01966(.A1(new_n2969_), .A2(new_n2970_), .B(new_n2968_), .ZN(new_n2971_));
  NAND2_X1   g01967(.A1(new_n2971_), .A2(new_n2967_), .ZN(new_n2972_));
  INV_X1     g01968(.I(\A[546] ), .ZN(new_n2973_));
  NOR2_X1    g01969(.A1(new_n2973_), .A2(\A[545] ), .ZN(new_n2974_));
  INV_X1     g01970(.I(\A[545] ), .ZN(new_n2975_));
  NOR2_X1    g01971(.A1(new_n2975_), .A2(\A[546] ), .ZN(new_n2976_));
  OAI21_X1   g01972(.A1(new_n2974_), .A2(new_n2976_), .B(\A[544] ), .ZN(new_n2977_));
  INV_X1     g01973(.I(\A[544] ), .ZN(new_n2978_));
  NOR2_X1    g01974(.A1(new_n2975_), .A2(new_n2973_), .ZN(new_n2979_));
  NOR2_X1    g01975(.A1(\A[545] ), .A2(\A[546] ), .ZN(new_n2980_));
  OAI21_X1   g01976(.A1(new_n2979_), .A2(new_n2980_), .B(new_n2978_), .ZN(new_n2981_));
  NAND2_X1   g01977(.A1(new_n2981_), .A2(new_n2977_), .ZN(new_n2982_));
  NOR2_X1    g01978(.A1(new_n2969_), .A2(\A[541] ), .ZN(new_n2983_));
  NOR2_X1    g01979(.A1(new_n2979_), .A2(\A[544] ), .ZN(new_n2984_));
  OAI22_X1   g01980(.A1(new_n2970_), .A2(new_n2983_), .B1(new_n2984_), .B2(new_n2980_), .ZN(new_n2985_));
  INV_X1     g01981(.I(new_n2985_), .ZN(new_n2986_));
  NAND3_X1   g01982(.A1(new_n2986_), .A2(new_n2972_), .A3(new_n2982_), .ZN(new_n2987_));
  INV_X1     g01983(.I(\A[535] ), .ZN(new_n2988_));
  INV_X1     g01984(.I(\A[536] ), .ZN(new_n2989_));
  NAND2_X1   g01985(.A1(new_n2989_), .A2(\A[537] ), .ZN(new_n2990_));
  INV_X1     g01986(.I(\A[537] ), .ZN(new_n2991_));
  NAND2_X1   g01987(.A1(new_n2991_), .A2(\A[536] ), .ZN(new_n2992_));
  AOI21_X1   g01988(.A1(new_n2990_), .A2(new_n2992_), .B(new_n2988_), .ZN(new_n2993_));
  NAND2_X1   g01989(.A1(\A[536] ), .A2(\A[537] ), .ZN(new_n2994_));
  NAND2_X1   g01990(.A1(new_n2989_), .A2(new_n2991_), .ZN(new_n2995_));
  AOI21_X1   g01991(.A1(new_n2995_), .A2(new_n2994_), .B(\A[535] ), .ZN(new_n2996_));
  NOR2_X1    g01992(.A1(new_n2996_), .A2(new_n2993_), .ZN(new_n2997_));
  INV_X1     g01993(.I(\A[538] ), .ZN(new_n2998_));
  INV_X1     g01994(.I(\A[539] ), .ZN(new_n2999_));
  NAND2_X1   g01995(.A1(new_n2999_), .A2(\A[540] ), .ZN(new_n3000_));
  INV_X1     g01996(.I(\A[540] ), .ZN(new_n3001_));
  NAND2_X1   g01997(.A1(new_n3001_), .A2(\A[539] ), .ZN(new_n3002_));
  AOI21_X1   g01998(.A1(new_n3000_), .A2(new_n3002_), .B(new_n2998_), .ZN(new_n3003_));
  NAND2_X1   g01999(.A1(\A[539] ), .A2(\A[540] ), .ZN(new_n3004_));
  NAND2_X1   g02000(.A1(new_n2999_), .A2(new_n3001_), .ZN(new_n3005_));
  AOI21_X1   g02001(.A1(new_n3005_), .A2(new_n3004_), .B(\A[538] ), .ZN(new_n3006_));
  NOR2_X1    g02002(.A1(new_n3006_), .A2(new_n3003_), .ZN(new_n3007_));
  NAND2_X1   g02003(.A1(new_n2994_), .A2(new_n2988_), .ZN(new_n3008_));
  NAND2_X1   g02004(.A1(new_n3008_), .A2(new_n2995_), .ZN(new_n3009_));
  NAND2_X1   g02005(.A1(new_n3004_), .A2(new_n2998_), .ZN(new_n3010_));
  NAND2_X1   g02006(.A1(new_n3010_), .A2(new_n3005_), .ZN(new_n3011_));
  NAND2_X1   g02007(.A1(new_n3009_), .A2(new_n3011_), .ZN(new_n3012_));
  NOR3_X1    g02008(.A1(new_n2997_), .A2(new_n3007_), .A3(new_n3012_), .ZN(new_n3013_));
  XOR2_X1    g02009(.A1(new_n2987_), .A2(new_n3013_), .Z(new_n3014_));
  NAND2_X1   g02010(.A1(new_n3014_), .A2(new_n2962_), .ZN(new_n3015_));
  INV_X1     g02011(.I(new_n3015_), .ZN(new_n3016_));
  NOR2_X1    g02012(.A1(new_n3014_), .A2(new_n2962_), .ZN(new_n3017_));
  NOR2_X1    g02013(.A1(new_n3016_), .A2(new_n3017_), .ZN(new_n3018_));
  INV_X1     g02014(.I(\A[531] ), .ZN(new_n3019_));
  NOR2_X1    g02015(.A1(new_n3019_), .A2(\A[530] ), .ZN(new_n3020_));
  INV_X1     g02016(.I(\A[530] ), .ZN(new_n3021_));
  NOR2_X1    g02017(.A1(new_n3021_), .A2(\A[531] ), .ZN(new_n3022_));
  OAI21_X1   g02018(.A1(new_n3020_), .A2(new_n3022_), .B(\A[529] ), .ZN(new_n3023_));
  INV_X1     g02019(.I(\A[529] ), .ZN(new_n3024_));
  NOR2_X1    g02020(.A1(\A[530] ), .A2(\A[531] ), .ZN(new_n3025_));
  NAND2_X1   g02021(.A1(\A[530] ), .A2(\A[531] ), .ZN(new_n3026_));
  INV_X1     g02022(.I(new_n3026_), .ZN(new_n3027_));
  OAI21_X1   g02023(.A1(new_n3027_), .A2(new_n3025_), .B(new_n3024_), .ZN(new_n3028_));
  NAND2_X1   g02024(.A1(new_n3023_), .A2(new_n3028_), .ZN(new_n3029_));
  INV_X1     g02025(.I(\A[534] ), .ZN(new_n3030_));
  NOR2_X1    g02026(.A1(new_n3030_), .A2(\A[533] ), .ZN(new_n3031_));
  INV_X1     g02027(.I(\A[533] ), .ZN(new_n3032_));
  NOR2_X1    g02028(.A1(new_n3032_), .A2(\A[534] ), .ZN(new_n3033_));
  OAI21_X1   g02029(.A1(new_n3031_), .A2(new_n3033_), .B(\A[532] ), .ZN(new_n3034_));
  INV_X1     g02030(.I(\A[532] ), .ZN(new_n3035_));
  NAND2_X1   g02031(.A1(\A[533] ), .A2(\A[534] ), .ZN(new_n3036_));
  INV_X1     g02032(.I(new_n3036_), .ZN(new_n3037_));
  NOR2_X1    g02033(.A1(\A[533] ), .A2(\A[534] ), .ZN(new_n3038_));
  OAI21_X1   g02034(.A1(new_n3037_), .A2(new_n3038_), .B(new_n3035_), .ZN(new_n3039_));
  NAND2_X1   g02035(.A1(new_n3034_), .A2(new_n3039_), .ZN(new_n3040_));
  AOI21_X1   g02036(.A1(new_n3024_), .A2(new_n3026_), .B(new_n3025_), .ZN(new_n3041_));
  AOI21_X1   g02037(.A1(new_n3035_), .A2(new_n3036_), .B(new_n3038_), .ZN(new_n3042_));
  NOR2_X1    g02038(.A1(new_n3041_), .A2(new_n3042_), .ZN(new_n3043_));
  NAND3_X1   g02039(.A1(new_n3029_), .A2(new_n3040_), .A3(new_n3043_), .ZN(new_n3044_));
  INV_X1     g02040(.I(\A[523] ), .ZN(new_n3045_));
  INV_X1     g02041(.I(\A[524] ), .ZN(new_n3046_));
  NAND2_X1   g02042(.A1(new_n3046_), .A2(\A[525] ), .ZN(new_n3047_));
  INV_X1     g02043(.I(\A[525] ), .ZN(new_n3048_));
  NAND2_X1   g02044(.A1(new_n3048_), .A2(\A[524] ), .ZN(new_n3049_));
  AOI21_X1   g02045(.A1(new_n3047_), .A2(new_n3049_), .B(new_n3045_), .ZN(new_n3050_));
  NAND2_X1   g02046(.A1(new_n3046_), .A2(new_n3048_), .ZN(new_n3051_));
  NAND2_X1   g02047(.A1(\A[524] ), .A2(\A[525] ), .ZN(new_n3052_));
  AOI21_X1   g02048(.A1(new_n3051_), .A2(new_n3052_), .B(\A[523] ), .ZN(new_n3053_));
  NOR2_X1    g02049(.A1(new_n3053_), .A2(new_n3050_), .ZN(new_n3054_));
  INV_X1     g02050(.I(\A[526] ), .ZN(new_n3055_));
  INV_X1     g02051(.I(\A[527] ), .ZN(new_n3056_));
  NAND2_X1   g02052(.A1(new_n3056_), .A2(\A[528] ), .ZN(new_n3057_));
  INV_X1     g02053(.I(\A[528] ), .ZN(new_n3058_));
  NAND2_X1   g02054(.A1(new_n3058_), .A2(\A[527] ), .ZN(new_n3059_));
  AOI21_X1   g02055(.A1(new_n3057_), .A2(new_n3059_), .B(new_n3055_), .ZN(new_n3060_));
  NAND2_X1   g02056(.A1(\A[527] ), .A2(\A[528] ), .ZN(new_n3061_));
  NAND2_X1   g02057(.A1(new_n3056_), .A2(new_n3058_), .ZN(new_n3062_));
  AOI21_X1   g02058(.A1(new_n3062_), .A2(new_n3061_), .B(\A[526] ), .ZN(new_n3063_));
  NOR2_X1    g02059(.A1(new_n3063_), .A2(new_n3060_), .ZN(new_n3064_));
  NAND2_X1   g02060(.A1(new_n3052_), .A2(new_n3045_), .ZN(new_n3065_));
  NAND2_X1   g02061(.A1(new_n3065_), .A2(new_n3051_), .ZN(new_n3066_));
  NAND2_X1   g02062(.A1(new_n3061_), .A2(new_n3055_), .ZN(new_n3067_));
  NAND2_X1   g02063(.A1(new_n3067_), .A2(new_n3062_), .ZN(new_n3068_));
  NAND2_X1   g02064(.A1(new_n3066_), .A2(new_n3068_), .ZN(new_n3069_));
  NOR3_X1    g02065(.A1(new_n3054_), .A2(new_n3064_), .A3(new_n3069_), .ZN(new_n3070_));
  XOR2_X1    g02066(.A1(new_n3070_), .A2(new_n3044_), .Z(new_n3071_));
  INV_X1     g02067(.I(\A[519] ), .ZN(new_n3072_));
  NOR2_X1    g02068(.A1(new_n3072_), .A2(\A[518] ), .ZN(new_n3073_));
  INV_X1     g02069(.I(\A[518] ), .ZN(new_n3074_));
  NOR2_X1    g02070(.A1(new_n3074_), .A2(\A[519] ), .ZN(new_n3075_));
  OAI21_X1   g02071(.A1(new_n3073_), .A2(new_n3075_), .B(\A[517] ), .ZN(new_n3076_));
  INV_X1     g02072(.I(\A[517] ), .ZN(new_n3077_));
  NOR2_X1    g02073(.A1(\A[518] ), .A2(\A[519] ), .ZN(new_n3078_));
  NOR2_X1    g02074(.A1(new_n3074_), .A2(new_n3072_), .ZN(new_n3079_));
  OAI21_X1   g02075(.A1(new_n3079_), .A2(new_n3078_), .B(new_n3077_), .ZN(new_n3080_));
  NAND2_X1   g02076(.A1(new_n3080_), .A2(new_n3076_), .ZN(new_n3081_));
  INV_X1     g02077(.I(\A[522] ), .ZN(new_n3082_));
  NOR2_X1    g02078(.A1(new_n3082_), .A2(\A[521] ), .ZN(new_n3083_));
  INV_X1     g02079(.I(\A[521] ), .ZN(new_n3084_));
  NOR2_X1    g02080(.A1(new_n3084_), .A2(\A[522] ), .ZN(new_n3085_));
  OAI21_X1   g02081(.A1(new_n3083_), .A2(new_n3085_), .B(\A[520] ), .ZN(new_n3086_));
  INV_X1     g02082(.I(\A[520] ), .ZN(new_n3087_));
  NOR2_X1    g02083(.A1(\A[521] ), .A2(\A[522] ), .ZN(new_n3088_));
  NAND2_X1   g02084(.A1(\A[521] ), .A2(\A[522] ), .ZN(new_n3089_));
  INV_X1     g02085(.I(new_n3089_), .ZN(new_n3090_));
  OAI21_X1   g02086(.A1(new_n3090_), .A2(new_n3088_), .B(new_n3087_), .ZN(new_n3091_));
  NAND2_X1   g02087(.A1(new_n3086_), .A2(new_n3091_), .ZN(new_n3092_));
  NOR2_X1    g02088(.A1(new_n3079_), .A2(\A[517] ), .ZN(new_n3093_));
  NOR2_X1    g02089(.A1(new_n3093_), .A2(new_n3078_), .ZN(new_n3094_));
  NOR2_X1    g02090(.A1(new_n3090_), .A2(\A[520] ), .ZN(new_n3095_));
  NOR2_X1    g02091(.A1(new_n3095_), .A2(new_n3088_), .ZN(new_n3096_));
  NOR2_X1    g02092(.A1(new_n3094_), .A2(new_n3096_), .ZN(new_n3097_));
  NAND3_X1   g02093(.A1(new_n3097_), .A2(new_n3081_), .A3(new_n3092_), .ZN(new_n3098_));
  INV_X1     g02094(.I(\A[511] ), .ZN(new_n3099_));
  INV_X1     g02095(.I(\A[512] ), .ZN(new_n3100_));
  NAND2_X1   g02096(.A1(new_n3100_), .A2(\A[513] ), .ZN(new_n3101_));
  INV_X1     g02097(.I(\A[513] ), .ZN(new_n3102_));
  NAND2_X1   g02098(.A1(new_n3102_), .A2(\A[512] ), .ZN(new_n3103_));
  AOI21_X1   g02099(.A1(new_n3101_), .A2(new_n3103_), .B(new_n3099_), .ZN(new_n3104_));
  NAND2_X1   g02100(.A1(new_n3100_), .A2(new_n3102_), .ZN(new_n3105_));
  NAND2_X1   g02101(.A1(\A[512] ), .A2(\A[513] ), .ZN(new_n3106_));
  AOI21_X1   g02102(.A1(new_n3105_), .A2(new_n3106_), .B(\A[511] ), .ZN(new_n3107_));
  NOR2_X1    g02103(.A1(new_n3107_), .A2(new_n3104_), .ZN(new_n3108_));
  INV_X1     g02104(.I(\A[514] ), .ZN(new_n3109_));
  INV_X1     g02105(.I(\A[515] ), .ZN(new_n3110_));
  NAND2_X1   g02106(.A1(new_n3110_), .A2(\A[516] ), .ZN(new_n3111_));
  INV_X1     g02107(.I(\A[516] ), .ZN(new_n3112_));
  NAND2_X1   g02108(.A1(new_n3112_), .A2(\A[515] ), .ZN(new_n3113_));
  AOI21_X1   g02109(.A1(new_n3111_), .A2(new_n3113_), .B(new_n3109_), .ZN(new_n3114_));
  NAND2_X1   g02110(.A1(\A[515] ), .A2(\A[516] ), .ZN(new_n3115_));
  NAND2_X1   g02111(.A1(new_n3110_), .A2(new_n3112_), .ZN(new_n3116_));
  AOI21_X1   g02112(.A1(new_n3116_), .A2(new_n3115_), .B(\A[514] ), .ZN(new_n3117_));
  NOR2_X1    g02113(.A1(new_n3117_), .A2(new_n3114_), .ZN(new_n3118_));
  NAND2_X1   g02114(.A1(new_n3106_), .A2(new_n3099_), .ZN(new_n3119_));
  NAND2_X1   g02115(.A1(new_n3119_), .A2(new_n3105_), .ZN(new_n3120_));
  NAND2_X1   g02116(.A1(new_n3115_), .A2(new_n3109_), .ZN(new_n3121_));
  NAND2_X1   g02117(.A1(new_n3121_), .A2(new_n3116_), .ZN(new_n3122_));
  NAND2_X1   g02118(.A1(new_n3120_), .A2(new_n3122_), .ZN(new_n3123_));
  NOR3_X1    g02119(.A1(new_n3108_), .A2(new_n3118_), .A3(new_n3123_), .ZN(new_n3124_));
  XOR2_X1    g02120(.A1(new_n3098_), .A2(new_n3124_), .Z(new_n3125_));
  NAND2_X1   g02121(.A1(new_n3125_), .A2(new_n3071_), .ZN(new_n3126_));
  INV_X1     g02122(.I(new_n3126_), .ZN(new_n3127_));
  NOR2_X1    g02123(.A1(new_n3125_), .A2(new_n3071_), .ZN(new_n3128_));
  NOR2_X1    g02124(.A1(new_n3127_), .A2(new_n3128_), .ZN(new_n3129_));
  NAND2_X1   g02125(.A1(new_n3018_), .A2(new_n3129_), .ZN(new_n3130_));
  INV_X1     g02126(.I(new_n3130_), .ZN(new_n3131_));
  NOR2_X1    g02127(.A1(new_n3018_), .A2(new_n3129_), .ZN(new_n3132_));
  NOR2_X1    g02128(.A1(new_n3131_), .A2(new_n3132_), .ZN(new_n3133_));
  NAND2_X1   g02129(.A1(new_n2909_), .A2(new_n3133_), .ZN(new_n3134_));
  INV_X1     g02130(.I(new_n3134_), .ZN(new_n3135_));
  NOR2_X1    g02131(.A1(new_n2909_), .A2(new_n3133_), .ZN(new_n3136_));
  NOR2_X1    g02132(.A1(new_n3135_), .A2(new_n3136_), .ZN(new_n3137_));
  INV_X1     g02133(.I(\A[651] ), .ZN(new_n3138_));
  NOR2_X1    g02134(.A1(new_n3138_), .A2(\A[650] ), .ZN(new_n3139_));
  INV_X1     g02135(.I(\A[650] ), .ZN(new_n3140_));
  NOR2_X1    g02136(.A1(new_n3140_), .A2(\A[651] ), .ZN(new_n3141_));
  OAI21_X1   g02137(.A1(new_n3139_), .A2(new_n3141_), .B(\A[649] ), .ZN(new_n3142_));
  INV_X1     g02138(.I(\A[649] ), .ZN(new_n3143_));
  NAND2_X1   g02139(.A1(\A[650] ), .A2(\A[651] ), .ZN(new_n3144_));
  INV_X1     g02140(.I(new_n3144_), .ZN(new_n3145_));
  NOR2_X1    g02141(.A1(\A[650] ), .A2(\A[651] ), .ZN(new_n3146_));
  OAI21_X1   g02142(.A1(new_n3145_), .A2(new_n3146_), .B(new_n3143_), .ZN(new_n3147_));
  NAND2_X1   g02143(.A1(new_n3142_), .A2(new_n3147_), .ZN(new_n3148_));
  INV_X1     g02144(.I(\A[654] ), .ZN(new_n3149_));
  NOR2_X1    g02145(.A1(new_n3149_), .A2(\A[653] ), .ZN(new_n3150_));
  INV_X1     g02146(.I(\A[653] ), .ZN(new_n3151_));
  NOR2_X1    g02147(.A1(new_n3151_), .A2(\A[654] ), .ZN(new_n3152_));
  OAI21_X1   g02148(.A1(new_n3150_), .A2(new_n3152_), .B(\A[652] ), .ZN(new_n3153_));
  INV_X1     g02149(.I(\A[652] ), .ZN(new_n3154_));
  NAND2_X1   g02150(.A1(\A[653] ), .A2(\A[654] ), .ZN(new_n3155_));
  INV_X1     g02151(.I(new_n3155_), .ZN(new_n3156_));
  NOR2_X1    g02152(.A1(\A[653] ), .A2(\A[654] ), .ZN(new_n3157_));
  OAI21_X1   g02153(.A1(new_n3156_), .A2(new_n3157_), .B(new_n3154_), .ZN(new_n3158_));
  NAND2_X1   g02154(.A1(new_n3153_), .A2(new_n3158_), .ZN(new_n3159_));
  AOI21_X1   g02155(.A1(new_n3143_), .A2(new_n3144_), .B(new_n3146_), .ZN(new_n3160_));
  AOI21_X1   g02156(.A1(new_n3154_), .A2(new_n3155_), .B(new_n3157_), .ZN(new_n3161_));
  NOR2_X1    g02157(.A1(new_n3160_), .A2(new_n3161_), .ZN(new_n3162_));
  NAND3_X1   g02158(.A1(new_n3148_), .A2(new_n3159_), .A3(new_n3162_), .ZN(new_n3163_));
  INV_X1     g02159(.I(\A[643] ), .ZN(new_n3164_));
  INV_X1     g02160(.I(\A[644] ), .ZN(new_n3165_));
  NAND2_X1   g02161(.A1(new_n3165_), .A2(\A[645] ), .ZN(new_n3166_));
  INV_X1     g02162(.I(\A[645] ), .ZN(new_n3167_));
  NAND2_X1   g02163(.A1(new_n3167_), .A2(\A[644] ), .ZN(new_n3168_));
  AOI21_X1   g02164(.A1(new_n3166_), .A2(new_n3168_), .B(new_n3164_), .ZN(new_n3169_));
  NAND2_X1   g02165(.A1(\A[644] ), .A2(\A[645] ), .ZN(new_n3170_));
  NAND2_X1   g02166(.A1(new_n3165_), .A2(new_n3167_), .ZN(new_n3171_));
  AOI21_X1   g02167(.A1(new_n3171_), .A2(new_n3170_), .B(\A[643] ), .ZN(new_n3172_));
  NOR2_X1    g02168(.A1(new_n3172_), .A2(new_n3169_), .ZN(new_n3173_));
  INV_X1     g02169(.I(\A[646] ), .ZN(new_n3174_));
  INV_X1     g02170(.I(\A[647] ), .ZN(new_n3175_));
  NAND2_X1   g02171(.A1(new_n3175_), .A2(\A[648] ), .ZN(new_n3176_));
  INV_X1     g02172(.I(\A[648] ), .ZN(new_n3177_));
  NAND2_X1   g02173(.A1(new_n3177_), .A2(\A[647] ), .ZN(new_n3178_));
  AOI21_X1   g02174(.A1(new_n3176_), .A2(new_n3178_), .B(new_n3174_), .ZN(new_n3179_));
  NAND2_X1   g02175(.A1(\A[647] ), .A2(\A[648] ), .ZN(new_n3180_));
  NOR2_X1    g02176(.A1(\A[647] ), .A2(\A[648] ), .ZN(new_n3181_));
  INV_X1     g02177(.I(new_n3181_), .ZN(new_n3182_));
  AOI21_X1   g02178(.A1(new_n3182_), .A2(new_n3180_), .B(\A[646] ), .ZN(new_n3183_));
  NOR2_X1    g02179(.A1(new_n3183_), .A2(new_n3179_), .ZN(new_n3184_));
  NAND2_X1   g02180(.A1(new_n3170_), .A2(new_n3164_), .ZN(new_n3185_));
  NAND2_X1   g02181(.A1(new_n3185_), .A2(new_n3171_), .ZN(new_n3186_));
  AOI21_X1   g02182(.A1(new_n3174_), .A2(new_n3180_), .B(new_n3181_), .ZN(new_n3187_));
  INV_X1     g02183(.I(new_n3187_), .ZN(new_n3188_));
  NAND2_X1   g02184(.A1(new_n3188_), .A2(new_n3186_), .ZN(new_n3189_));
  NOR3_X1    g02185(.A1(new_n3173_), .A2(new_n3189_), .A3(new_n3184_), .ZN(new_n3190_));
  XOR2_X1    g02186(.A1(new_n3190_), .A2(new_n3163_), .Z(new_n3191_));
  INV_X1     g02187(.I(\A[639] ), .ZN(new_n3192_));
  NOR2_X1    g02188(.A1(new_n3192_), .A2(\A[638] ), .ZN(new_n3193_));
  INV_X1     g02189(.I(\A[638] ), .ZN(new_n3194_));
  NOR2_X1    g02190(.A1(new_n3194_), .A2(\A[639] ), .ZN(new_n3195_));
  OAI21_X1   g02191(.A1(new_n3193_), .A2(new_n3195_), .B(\A[637] ), .ZN(new_n3196_));
  INV_X1     g02192(.I(\A[637] ), .ZN(new_n3197_));
  NAND2_X1   g02193(.A1(\A[638] ), .A2(\A[639] ), .ZN(new_n3198_));
  INV_X1     g02194(.I(new_n3198_), .ZN(new_n3199_));
  NOR2_X1    g02195(.A1(\A[638] ), .A2(\A[639] ), .ZN(new_n3200_));
  OAI21_X1   g02196(.A1(new_n3199_), .A2(new_n3200_), .B(new_n3197_), .ZN(new_n3201_));
  NAND2_X1   g02197(.A1(new_n3196_), .A2(new_n3201_), .ZN(new_n3202_));
  INV_X1     g02198(.I(\A[642] ), .ZN(new_n3203_));
  NOR2_X1    g02199(.A1(new_n3203_), .A2(\A[641] ), .ZN(new_n3204_));
  INV_X1     g02200(.I(\A[641] ), .ZN(new_n3205_));
  NOR2_X1    g02201(.A1(new_n3205_), .A2(\A[642] ), .ZN(new_n3206_));
  OAI21_X1   g02202(.A1(new_n3204_), .A2(new_n3206_), .B(\A[640] ), .ZN(new_n3207_));
  INV_X1     g02203(.I(\A[640] ), .ZN(new_n3208_));
  NAND2_X1   g02204(.A1(\A[641] ), .A2(\A[642] ), .ZN(new_n3209_));
  INV_X1     g02205(.I(new_n3209_), .ZN(new_n3210_));
  NOR2_X1    g02206(.A1(\A[641] ), .A2(\A[642] ), .ZN(new_n3211_));
  OAI21_X1   g02207(.A1(new_n3210_), .A2(new_n3211_), .B(new_n3208_), .ZN(new_n3212_));
  NAND2_X1   g02208(.A1(new_n3207_), .A2(new_n3212_), .ZN(new_n3213_));
  AOI21_X1   g02209(.A1(new_n3197_), .A2(new_n3198_), .B(new_n3200_), .ZN(new_n3214_));
  AOI21_X1   g02210(.A1(new_n3208_), .A2(new_n3209_), .B(new_n3211_), .ZN(new_n3215_));
  NOR2_X1    g02211(.A1(new_n3214_), .A2(new_n3215_), .ZN(new_n3216_));
  NAND3_X1   g02212(.A1(new_n3202_), .A2(new_n3213_), .A3(new_n3216_), .ZN(new_n3217_));
  INV_X1     g02213(.I(\A[631] ), .ZN(new_n3218_));
  INV_X1     g02214(.I(\A[632] ), .ZN(new_n3219_));
  NAND2_X1   g02215(.A1(new_n3219_), .A2(\A[633] ), .ZN(new_n3220_));
  INV_X1     g02216(.I(\A[633] ), .ZN(new_n3221_));
  NAND2_X1   g02217(.A1(new_n3221_), .A2(\A[632] ), .ZN(new_n3222_));
  AOI21_X1   g02218(.A1(new_n3220_), .A2(new_n3222_), .B(new_n3218_), .ZN(new_n3223_));
  NAND2_X1   g02219(.A1(\A[632] ), .A2(\A[633] ), .ZN(new_n3224_));
  NAND2_X1   g02220(.A1(new_n3219_), .A2(new_n3221_), .ZN(new_n3225_));
  AOI21_X1   g02221(.A1(new_n3225_), .A2(new_n3224_), .B(\A[631] ), .ZN(new_n3226_));
  NOR2_X1    g02222(.A1(new_n3226_), .A2(new_n3223_), .ZN(new_n3227_));
  INV_X1     g02223(.I(\A[634] ), .ZN(new_n3228_));
  INV_X1     g02224(.I(\A[635] ), .ZN(new_n3229_));
  NAND2_X1   g02225(.A1(new_n3229_), .A2(\A[636] ), .ZN(new_n3230_));
  INV_X1     g02226(.I(\A[636] ), .ZN(new_n3231_));
  NAND2_X1   g02227(.A1(new_n3231_), .A2(\A[635] ), .ZN(new_n3232_));
  AOI21_X1   g02228(.A1(new_n3230_), .A2(new_n3232_), .B(new_n3228_), .ZN(new_n3233_));
  NAND2_X1   g02229(.A1(\A[635] ), .A2(\A[636] ), .ZN(new_n3234_));
  NAND2_X1   g02230(.A1(new_n3229_), .A2(new_n3231_), .ZN(new_n3235_));
  AOI21_X1   g02231(.A1(new_n3235_), .A2(new_n3234_), .B(\A[634] ), .ZN(new_n3236_));
  NOR2_X1    g02232(.A1(new_n3236_), .A2(new_n3233_), .ZN(new_n3237_));
  NAND2_X1   g02233(.A1(new_n3224_), .A2(new_n3218_), .ZN(new_n3238_));
  NAND2_X1   g02234(.A1(new_n3238_), .A2(new_n3225_), .ZN(new_n3239_));
  NAND2_X1   g02235(.A1(new_n3234_), .A2(new_n3228_), .ZN(new_n3240_));
  NAND2_X1   g02236(.A1(new_n3240_), .A2(new_n3235_), .ZN(new_n3241_));
  NAND2_X1   g02237(.A1(new_n3239_), .A2(new_n3241_), .ZN(new_n3242_));
  NOR3_X1    g02238(.A1(new_n3227_), .A2(new_n3237_), .A3(new_n3242_), .ZN(new_n3243_));
  XOR2_X1    g02239(.A1(new_n3243_), .A2(new_n3217_), .Z(new_n3244_));
  NOR2_X1    g02240(.A1(new_n3191_), .A2(new_n3244_), .ZN(new_n3245_));
  NAND2_X1   g02241(.A1(new_n3191_), .A2(new_n3244_), .ZN(new_n3246_));
  INV_X1     g02242(.I(new_n3246_), .ZN(new_n3247_));
  NOR2_X1    g02243(.A1(new_n3247_), .A2(new_n3245_), .ZN(new_n3248_));
  INV_X1     g02244(.I(\A[627] ), .ZN(new_n3249_));
  NOR2_X1    g02245(.A1(new_n3249_), .A2(\A[626] ), .ZN(new_n3250_));
  INV_X1     g02246(.I(\A[626] ), .ZN(new_n3251_));
  NOR2_X1    g02247(.A1(new_n3251_), .A2(\A[627] ), .ZN(new_n3252_));
  OAI21_X1   g02248(.A1(new_n3250_), .A2(new_n3252_), .B(\A[625] ), .ZN(new_n3253_));
  INV_X1     g02249(.I(\A[625] ), .ZN(new_n3254_));
  NAND2_X1   g02250(.A1(\A[626] ), .A2(\A[627] ), .ZN(new_n3255_));
  INV_X1     g02251(.I(new_n3255_), .ZN(new_n3256_));
  NOR2_X1    g02252(.A1(\A[626] ), .A2(\A[627] ), .ZN(new_n3257_));
  OAI21_X1   g02253(.A1(new_n3256_), .A2(new_n3257_), .B(new_n3254_), .ZN(new_n3258_));
  NAND2_X1   g02254(.A1(new_n3253_), .A2(new_n3258_), .ZN(new_n3259_));
  INV_X1     g02255(.I(\A[630] ), .ZN(new_n3260_));
  NOR2_X1    g02256(.A1(new_n3260_), .A2(\A[629] ), .ZN(new_n3261_));
  INV_X1     g02257(.I(\A[629] ), .ZN(new_n3262_));
  NOR2_X1    g02258(.A1(new_n3262_), .A2(\A[630] ), .ZN(new_n3263_));
  OAI21_X1   g02259(.A1(new_n3261_), .A2(new_n3263_), .B(\A[628] ), .ZN(new_n3264_));
  INV_X1     g02260(.I(\A[628] ), .ZN(new_n3265_));
  NAND2_X1   g02261(.A1(\A[629] ), .A2(\A[630] ), .ZN(new_n3266_));
  INV_X1     g02262(.I(new_n3266_), .ZN(new_n3267_));
  NOR2_X1    g02263(.A1(\A[629] ), .A2(\A[630] ), .ZN(new_n3268_));
  OAI21_X1   g02264(.A1(new_n3267_), .A2(new_n3268_), .B(new_n3265_), .ZN(new_n3269_));
  NAND2_X1   g02265(.A1(new_n3264_), .A2(new_n3269_), .ZN(new_n3270_));
  AOI21_X1   g02266(.A1(new_n3254_), .A2(new_n3255_), .B(new_n3257_), .ZN(new_n3271_));
  AOI21_X1   g02267(.A1(new_n3265_), .A2(new_n3266_), .B(new_n3268_), .ZN(new_n3272_));
  NOR2_X1    g02268(.A1(new_n3271_), .A2(new_n3272_), .ZN(new_n3273_));
  NAND3_X1   g02269(.A1(new_n3259_), .A2(new_n3270_), .A3(new_n3273_), .ZN(new_n3274_));
  INV_X1     g02270(.I(\A[619] ), .ZN(new_n3275_));
  INV_X1     g02271(.I(\A[620] ), .ZN(new_n3276_));
  NAND2_X1   g02272(.A1(new_n3276_), .A2(\A[621] ), .ZN(new_n3277_));
  INV_X1     g02273(.I(\A[621] ), .ZN(new_n3278_));
  NAND2_X1   g02274(.A1(new_n3278_), .A2(\A[620] ), .ZN(new_n3279_));
  AOI21_X1   g02275(.A1(new_n3277_), .A2(new_n3279_), .B(new_n3275_), .ZN(new_n3280_));
  NAND2_X1   g02276(.A1(\A[620] ), .A2(\A[621] ), .ZN(new_n3281_));
  NAND2_X1   g02277(.A1(new_n3276_), .A2(new_n3278_), .ZN(new_n3282_));
  AOI21_X1   g02278(.A1(new_n3282_), .A2(new_n3281_), .B(\A[619] ), .ZN(new_n3283_));
  NOR2_X1    g02279(.A1(new_n3283_), .A2(new_n3280_), .ZN(new_n3284_));
  INV_X1     g02280(.I(\A[622] ), .ZN(new_n3285_));
  INV_X1     g02281(.I(\A[623] ), .ZN(new_n3286_));
  NAND2_X1   g02282(.A1(new_n3286_), .A2(\A[624] ), .ZN(new_n3287_));
  INV_X1     g02283(.I(\A[624] ), .ZN(new_n3288_));
  NAND2_X1   g02284(.A1(new_n3288_), .A2(\A[623] ), .ZN(new_n3289_));
  AOI21_X1   g02285(.A1(new_n3287_), .A2(new_n3289_), .B(new_n3285_), .ZN(new_n3290_));
  NAND2_X1   g02286(.A1(\A[623] ), .A2(\A[624] ), .ZN(new_n3291_));
  NOR2_X1    g02287(.A1(\A[623] ), .A2(\A[624] ), .ZN(new_n3292_));
  INV_X1     g02288(.I(new_n3292_), .ZN(new_n3293_));
  AOI21_X1   g02289(.A1(new_n3293_), .A2(new_n3291_), .B(\A[622] ), .ZN(new_n3294_));
  NOR2_X1    g02290(.A1(new_n3294_), .A2(new_n3290_), .ZN(new_n3295_));
  NAND2_X1   g02291(.A1(new_n3281_), .A2(new_n3275_), .ZN(new_n3296_));
  NAND2_X1   g02292(.A1(new_n3296_), .A2(new_n3282_), .ZN(new_n3297_));
  NAND2_X1   g02293(.A1(new_n3291_), .A2(new_n3285_), .ZN(new_n3298_));
  NAND2_X1   g02294(.A1(new_n3298_), .A2(new_n3293_), .ZN(new_n3299_));
  NAND2_X1   g02295(.A1(new_n3299_), .A2(new_n3297_), .ZN(new_n3300_));
  NOR3_X1    g02296(.A1(new_n3284_), .A2(new_n3295_), .A3(new_n3300_), .ZN(new_n3301_));
  XOR2_X1    g02297(.A1(new_n3301_), .A2(new_n3274_), .Z(new_n3302_));
  INV_X1     g02298(.I(\A[615] ), .ZN(new_n3303_));
  NOR2_X1    g02299(.A1(new_n3303_), .A2(\A[614] ), .ZN(new_n3304_));
  INV_X1     g02300(.I(\A[614] ), .ZN(new_n3305_));
  NOR2_X1    g02301(.A1(new_n3305_), .A2(\A[615] ), .ZN(new_n3306_));
  OAI21_X1   g02302(.A1(new_n3304_), .A2(new_n3306_), .B(\A[613] ), .ZN(new_n3307_));
  INV_X1     g02303(.I(\A[613] ), .ZN(new_n3308_));
  NAND2_X1   g02304(.A1(\A[614] ), .A2(\A[615] ), .ZN(new_n3309_));
  INV_X1     g02305(.I(new_n3309_), .ZN(new_n3310_));
  NOR2_X1    g02306(.A1(\A[614] ), .A2(\A[615] ), .ZN(new_n3311_));
  OAI21_X1   g02307(.A1(new_n3310_), .A2(new_n3311_), .B(new_n3308_), .ZN(new_n3312_));
  NAND2_X1   g02308(.A1(new_n3307_), .A2(new_n3312_), .ZN(new_n3313_));
  INV_X1     g02309(.I(\A[618] ), .ZN(new_n3314_));
  NOR2_X1    g02310(.A1(new_n3314_), .A2(\A[617] ), .ZN(new_n3315_));
  INV_X1     g02311(.I(\A[617] ), .ZN(new_n3316_));
  NOR2_X1    g02312(.A1(new_n3316_), .A2(\A[618] ), .ZN(new_n3317_));
  OAI21_X1   g02313(.A1(new_n3315_), .A2(new_n3317_), .B(\A[616] ), .ZN(new_n3318_));
  INV_X1     g02314(.I(\A[616] ), .ZN(new_n3319_));
  NAND2_X1   g02315(.A1(\A[617] ), .A2(\A[618] ), .ZN(new_n3320_));
  INV_X1     g02316(.I(new_n3320_), .ZN(new_n3321_));
  NOR2_X1    g02317(.A1(\A[617] ), .A2(\A[618] ), .ZN(new_n3322_));
  OAI21_X1   g02318(.A1(new_n3321_), .A2(new_n3322_), .B(new_n3319_), .ZN(new_n3323_));
  NAND2_X1   g02319(.A1(new_n3318_), .A2(new_n3323_), .ZN(new_n3324_));
  AOI21_X1   g02320(.A1(new_n3308_), .A2(new_n3309_), .B(new_n3311_), .ZN(new_n3325_));
  AOI21_X1   g02321(.A1(new_n3319_), .A2(new_n3320_), .B(new_n3322_), .ZN(new_n3326_));
  NOR2_X1    g02322(.A1(new_n3325_), .A2(new_n3326_), .ZN(new_n3327_));
  NAND3_X1   g02323(.A1(new_n3313_), .A2(new_n3324_), .A3(new_n3327_), .ZN(new_n3328_));
  INV_X1     g02324(.I(\A[607] ), .ZN(new_n3329_));
  INV_X1     g02325(.I(\A[608] ), .ZN(new_n3330_));
  NAND2_X1   g02326(.A1(new_n3330_), .A2(\A[609] ), .ZN(new_n3331_));
  INV_X1     g02327(.I(\A[609] ), .ZN(new_n3332_));
  NAND2_X1   g02328(.A1(new_n3332_), .A2(\A[608] ), .ZN(new_n3333_));
  AOI21_X1   g02329(.A1(new_n3331_), .A2(new_n3333_), .B(new_n3329_), .ZN(new_n3334_));
  NAND2_X1   g02330(.A1(\A[608] ), .A2(\A[609] ), .ZN(new_n3335_));
  NAND2_X1   g02331(.A1(new_n3330_), .A2(new_n3332_), .ZN(new_n3336_));
  AOI21_X1   g02332(.A1(new_n3336_), .A2(new_n3335_), .B(\A[607] ), .ZN(new_n3337_));
  NOR2_X1    g02333(.A1(new_n3337_), .A2(new_n3334_), .ZN(new_n3338_));
  INV_X1     g02334(.I(\A[610] ), .ZN(new_n3339_));
  INV_X1     g02335(.I(\A[611] ), .ZN(new_n3340_));
  NAND2_X1   g02336(.A1(new_n3340_), .A2(\A[612] ), .ZN(new_n3341_));
  INV_X1     g02337(.I(\A[612] ), .ZN(new_n3342_));
  NAND2_X1   g02338(.A1(new_n3342_), .A2(\A[611] ), .ZN(new_n3343_));
  AOI21_X1   g02339(.A1(new_n3341_), .A2(new_n3343_), .B(new_n3339_), .ZN(new_n3344_));
  NAND2_X1   g02340(.A1(\A[611] ), .A2(\A[612] ), .ZN(new_n3345_));
  NAND2_X1   g02341(.A1(new_n3340_), .A2(new_n3342_), .ZN(new_n3346_));
  AOI21_X1   g02342(.A1(new_n3346_), .A2(new_n3345_), .B(\A[610] ), .ZN(new_n3347_));
  NOR2_X1    g02343(.A1(new_n3347_), .A2(new_n3344_), .ZN(new_n3348_));
  NAND2_X1   g02344(.A1(new_n3335_), .A2(new_n3329_), .ZN(new_n3349_));
  NAND2_X1   g02345(.A1(new_n3349_), .A2(new_n3336_), .ZN(new_n3350_));
  NAND2_X1   g02346(.A1(new_n3345_), .A2(new_n3339_), .ZN(new_n3351_));
  NAND2_X1   g02347(.A1(new_n3351_), .A2(new_n3346_), .ZN(new_n3352_));
  NAND2_X1   g02348(.A1(new_n3350_), .A2(new_n3352_), .ZN(new_n3353_));
  NOR3_X1    g02349(.A1(new_n3338_), .A2(new_n3348_), .A3(new_n3353_), .ZN(new_n3354_));
  XOR2_X1    g02350(.A1(new_n3354_), .A2(new_n3328_), .Z(new_n3355_));
  NOR2_X1    g02351(.A1(new_n3302_), .A2(new_n3355_), .ZN(new_n3356_));
  AND2_X2    g02352(.A1(new_n3302_), .A2(new_n3355_), .Z(new_n3357_));
  NOR2_X1    g02353(.A1(new_n3357_), .A2(new_n3356_), .ZN(new_n3358_));
  NOR2_X1    g02354(.A1(new_n3248_), .A2(new_n3358_), .ZN(new_n3359_));
  NAND2_X1   g02355(.A1(new_n3248_), .A2(new_n3358_), .ZN(new_n3360_));
  INV_X1     g02356(.I(new_n3360_), .ZN(new_n3361_));
  NOR2_X1    g02357(.A1(new_n3361_), .A2(new_n3359_), .ZN(new_n3362_));
  INV_X1     g02358(.I(\A[603] ), .ZN(new_n3363_));
  NOR2_X1    g02359(.A1(new_n3363_), .A2(\A[602] ), .ZN(new_n3364_));
  INV_X1     g02360(.I(\A[602] ), .ZN(new_n3365_));
  NOR2_X1    g02361(.A1(new_n3365_), .A2(\A[603] ), .ZN(new_n3366_));
  OAI21_X1   g02362(.A1(new_n3364_), .A2(new_n3366_), .B(\A[601] ), .ZN(new_n3367_));
  INV_X1     g02363(.I(\A[601] ), .ZN(new_n3368_));
  NAND2_X1   g02364(.A1(\A[602] ), .A2(\A[603] ), .ZN(new_n3369_));
  INV_X1     g02365(.I(new_n3369_), .ZN(new_n3370_));
  NOR2_X1    g02366(.A1(\A[602] ), .A2(\A[603] ), .ZN(new_n3371_));
  OAI21_X1   g02367(.A1(new_n3370_), .A2(new_n3371_), .B(new_n3368_), .ZN(new_n3372_));
  NAND2_X1   g02368(.A1(new_n3367_), .A2(new_n3372_), .ZN(new_n3373_));
  INV_X1     g02369(.I(\A[606] ), .ZN(new_n3374_));
  NOR2_X1    g02370(.A1(new_n3374_), .A2(\A[605] ), .ZN(new_n3375_));
  INV_X1     g02371(.I(\A[605] ), .ZN(new_n3376_));
  NOR2_X1    g02372(.A1(new_n3376_), .A2(\A[606] ), .ZN(new_n3377_));
  OAI21_X1   g02373(.A1(new_n3375_), .A2(new_n3377_), .B(\A[604] ), .ZN(new_n3378_));
  INV_X1     g02374(.I(\A[604] ), .ZN(new_n3379_));
  NAND2_X1   g02375(.A1(\A[605] ), .A2(\A[606] ), .ZN(new_n3380_));
  INV_X1     g02376(.I(new_n3380_), .ZN(new_n3381_));
  NOR2_X1    g02377(.A1(\A[605] ), .A2(\A[606] ), .ZN(new_n3382_));
  OAI21_X1   g02378(.A1(new_n3381_), .A2(new_n3382_), .B(new_n3379_), .ZN(new_n3383_));
  NAND2_X1   g02379(.A1(new_n3378_), .A2(new_n3383_), .ZN(new_n3384_));
  AOI21_X1   g02380(.A1(new_n3368_), .A2(new_n3369_), .B(new_n3371_), .ZN(new_n3385_));
  AOI21_X1   g02381(.A1(new_n3379_), .A2(new_n3380_), .B(new_n3382_), .ZN(new_n3386_));
  NOR2_X1    g02382(.A1(new_n3385_), .A2(new_n3386_), .ZN(new_n3387_));
  NAND3_X1   g02383(.A1(new_n3373_), .A2(new_n3384_), .A3(new_n3387_), .ZN(new_n3388_));
  INV_X1     g02384(.I(\A[595] ), .ZN(new_n3389_));
  INV_X1     g02385(.I(\A[596] ), .ZN(new_n3390_));
  NAND2_X1   g02386(.A1(new_n3390_), .A2(\A[597] ), .ZN(new_n3391_));
  INV_X1     g02387(.I(\A[597] ), .ZN(new_n3392_));
  NAND2_X1   g02388(.A1(new_n3392_), .A2(\A[596] ), .ZN(new_n3393_));
  AOI21_X1   g02389(.A1(new_n3391_), .A2(new_n3393_), .B(new_n3389_), .ZN(new_n3394_));
  NAND2_X1   g02390(.A1(\A[596] ), .A2(\A[597] ), .ZN(new_n3395_));
  NAND2_X1   g02391(.A1(new_n3390_), .A2(new_n3392_), .ZN(new_n3396_));
  AOI21_X1   g02392(.A1(new_n3396_), .A2(new_n3395_), .B(\A[595] ), .ZN(new_n3397_));
  NOR2_X1    g02393(.A1(new_n3397_), .A2(new_n3394_), .ZN(new_n3398_));
  INV_X1     g02394(.I(\A[598] ), .ZN(new_n3399_));
  INV_X1     g02395(.I(\A[599] ), .ZN(new_n3400_));
  NAND2_X1   g02396(.A1(new_n3400_), .A2(\A[600] ), .ZN(new_n3401_));
  INV_X1     g02397(.I(\A[600] ), .ZN(new_n3402_));
  NAND2_X1   g02398(.A1(new_n3402_), .A2(\A[599] ), .ZN(new_n3403_));
  AOI21_X1   g02399(.A1(new_n3401_), .A2(new_n3403_), .B(new_n3399_), .ZN(new_n3404_));
  NAND2_X1   g02400(.A1(\A[599] ), .A2(\A[600] ), .ZN(new_n3405_));
  NOR2_X1    g02401(.A1(\A[599] ), .A2(\A[600] ), .ZN(new_n3406_));
  INV_X1     g02402(.I(new_n3406_), .ZN(new_n3407_));
  AOI21_X1   g02403(.A1(new_n3407_), .A2(new_n3405_), .B(\A[598] ), .ZN(new_n3408_));
  NOR2_X1    g02404(.A1(new_n3408_), .A2(new_n3404_), .ZN(new_n3409_));
  NAND2_X1   g02405(.A1(new_n3395_), .A2(new_n3389_), .ZN(new_n3410_));
  NAND2_X1   g02406(.A1(new_n3410_), .A2(new_n3396_), .ZN(new_n3411_));
  AOI21_X1   g02407(.A1(new_n3399_), .A2(new_n3405_), .B(new_n3406_), .ZN(new_n3412_));
  INV_X1     g02408(.I(new_n3412_), .ZN(new_n3413_));
  NAND2_X1   g02409(.A1(new_n3413_), .A2(new_n3411_), .ZN(new_n3414_));
  NOR3_X1    g02410(.A1(new_n3398_), .A2(new_n3414_), .A3(new_n3409_), .ZN(new_n3415_));
  XOR2_X1    g02411(.A1(new_n3415_), .A2(new_n3388_), .Z(new_n3416_));
  INV_X1     g02412(.I(\A[591] ), .ZN(new_n3417_));
  NOR2_X1    g02413(.A1(new_n3417_), .A2(\A[590] ), .ZN(new_n3418_));
  INV_X1     g02414(.I(\A[590] ), .ZN(new_n3419_));
  NOR2_X1    g02415(.A1(new_n3419_), .A2(\A[591] ), .ZN(new_n3420_));
  OAI21_X1   g02416(.A1(new_n3418_), .A2(new_n3420_), .B(\A[589] ), .ZN(new_n3421_));
  INV_X1     g02417(.I(\A[589] ), .ZN(new_n3422_));
  NAND2_X1   g02418(.A1(\A[590] ), .A2(\A[591] ), .ZN(new_n3423_));
  INV_X1     g02419(.I(new_n3423_), .ZN(new_n3424_));
  NOR2_X1    g02420(.A1(\A[590] ), .A2(\A[591] ), .ZN(new_n3425_));
  OAI21_X1   g02421(.A1(new_n3424_), .A2(new_n3425_), .B(new_n3422_), .ZN(new_n3426_));
  NAND2_X1   g02422(.A1(new_n3421_), .A2(new_n3426_), .ZN(new_n3427_));
  INV_X1     g02423(.I(\A[594] ), .ZN(new_n3428_));
  NOR2_X1    g02424(.A1(new_n3428_), .A2(\A[593] ), .ZN(new_n3429_));
  INV_X1     g02425(.I(\A[593] ), .ZN(new_n3430_));
  NOR2_X1    g02426(.A1(new_n3430_), .A2(\A[594] ), .ZN(new_n3431_));
  OAI21_X1   g02427(.A1(new_n3429_), .A2(new_n3431_), .B(\A[592] ), .ZN(new_n3432_));
  INV_X1     g02428(.I(\A[592] ), .ZN(new_n3433_));
  NAND2_X1   g02429(.A1(\A[593] ), .A2(\A[594] ), .ZN(new_n3434_));
  INV_X1     g02430(.I(new_n3434_), .ZN(new_n3435_));
  NOR2_X1    g02431(.A1(\A[593] ), .A2(\A[594] ), .ZN(new_n3436_));
  OAI21_X1   g02432(.A1(new_n3435_), .A2(new_n3436_), .B(new_n3433_), .ZN(new_n3437_));
  NAND2_X1   g02433(.A1(new_n3432_), .A2(new_n3437_), .ZN(new_n3438_));
  AOI21_X1   g02434(.A1(new_n3422_), .A2(new_n3423_), .B(new_n3425_), .ZN(new_n3439_));
  AOI21_X1   g02435(.A1(new_n3433_), .A2(new_n3434_), .B(new_n3436_), .ZN(new_n3440_));
  NOR2_X1    g02436(.A1(new_n3439_), .A2(new_n3440_), .ZN(new_n3441_));
  NAND3_X1   g02437(.A1(new_n3427_), .A2(new_n3438_), .A3(new_n3441_), .ZN(new_n3442_));
  INV_X1     g02438(.I(\A[583] ), .ZN(new_n3443_));
  INV_X1     g02439(.I(\A[584] ), .ZN(new_n3444_));
  NAND2_X1   g02440(.A1(new_n3444_), .A2(\A[585] ), .ZN(new_n3445_));
  INV_X1     g02441(.I(\A[585] ), .ZN(new_n3446_));
  NAND2_X1   g02442(.A1(new_n3446_), .A2(\A[584] ), .ZN(new_n3447_));
  AOI21_X1   g02443(.A1(new_n3445_), .A2(new_n3447_), .B(new_n3443_), .ZN(new_n3448_));
  NAND2_X1   g02444(.A1(\A[584] ), .A2(\A[585] ), .ZN(new_n3449_));
  NAND2_X1   g02445(.A1(new_n3444_), .A2(new_n3446_), .ZN(new_n3450_));
  AOI21_X1   g02446(.A1(new_n3450_), .A2(new_n3449_), .B(\A[583] ), .ZN(new_n3451_));
  NOR2_X1    g02447(.A1(new_n3451_), .A2(new_n3448_), .ZN(new_n3452_));
  INV_X1     g02448(.I(\A[586] ), .ZN(new_n3453_));
  INV_X1     g02449(.I(\A[587] ), .ZN(new_n3454_));
  NAND2_X1   g02450(.A1(new_n3454_), .A2(\A[588] ), .ZN(new_n3455_));
  INV_X1     g02451(.I(\A[588] ), .ZN(new_n3456_));
  NAND2_X1   g02452(.A1(new_n3456_), .A2(\A[587] ), .ZN(new_n3457_));
  AOI21_X1   g02453(.A1(new_n3455_), .A2(new_n3457_), .B(new_n3453_), .ZN(new_n3458_));
  NAND2_X1   g02454(.A1(\A[587] ), .A2(\A[588] ), .ZN(new_n3459_));
  NAND2_X1   g02455(.A1(new_n3454_), .A2(new_n3456_), .ZN(new_n3460_));
  AOI21_X1   g02456(.A1(new_n3460_), .A2(new_n3459_), .B(\A[586] ), .ZN(new_n3461_));
  NOR2_X1    g02457(.A1(new_n3461_), .A2(new_n3458_), .ZN(new_n3462_));
  NAND2_X1   g02458(.A1(new_n3449_), .A2(new_n3443_), .ZN(new_n3463_));
  NAND2_X1   g02459(.A1(new_n3463_), .A2(new_n3450_), .ZN(new_n3464_));
  NAND2_X1   g02460(.A1(new_n3459_), .A2(new_n3453_), .ZN(new_n3465_));
  NAND2_X1   g02461(.A1(new_n3465_), .A2(new_n3460_), .ZN(new_n3466_));
  NAND2_X1   g02462(.A1(new_n3464_), .A2(new_n3466_), .ZN(new_n3467_));
  NOR3_X1    g02463(.A1(new_n3452_), .A2(new_n3462_), .A3(new_n3467_), .ZN(new_n3468_));
  XOR2_X1    g02464(.A1(new_n3468_), .A2(new_n3442_), .Z(new_n3469_));
  NOR2_X1    g02465(.A1(new_n3416_), .A2(new_n3469_), .ZN(new_n3470_));
  NAND2_X1   g02466(.A1(new_n3416_), .A2(new_n3469_), .ZN(new_n3471_));
  INV_X1     g02467(.I(new_n3471_), .ZN(new_n3472_));
  NOR2_X1    g02468(.A1(new_n3472_), .A2(new_n3470_), .ZN(new_n3473_));
  INV_X1     g02469(.I(\A[579] ), .ZN(new_n3474_));
  NOR2_X1    g02470(.A1(new_n3474_), .A2(\A[578] ), .ZN(new_n3475_));
  INV_X1     g02471(.I(\A[578] ), .ZN(new_n3476_));
  NOR2_X1    g02472(.A1(new_n3476_), .A2(\A[579] ), .ZN(new_n3477_));
  OAI21_X1   g02473(.A1(new_n3475_), .A2(new_n3477_), .B(\A[577] ), .ZN(new_n3478_));
  INV_X1     g02474(.I(\A[577] ), .ZN(new_n3479_));
  NAND2_X1   g02475(.A1(\A[578] ), .A2(\A[579] ), .ZN(new_n3480_));
  INV_X1     g02476(.I(new_n3480_), .ZN(new_n3481_));
  NOR2_X1    g02477(.A1(\A[578] ), .A2(\A[579] ), .ZN(new_n3482_));
  OAI21_X1   g02478(.A1(new_n3481_), .A2(new_n3482_), .B(new_n3479_), .ZN(new_n3483_));
  NAND2_X1   g02479(.A1(new_n3478_), .A2(new_n3483_), .ZN(new_n3484_));
  INV_X1     g02480(.I(\A[582] ), .ZN(new_n3485_));
  NOR2_X1    g02481(.A1(new_n3485_), .A2(\A[581] ), .ZN(new_n3486_));
  INV_X1     g02482(.I(\A[581] ), .ZN(new_n3487_));
  NOR2_X1    g02483(.A1(new_n3487_), .A2(\A[582] ), .ZN(new_n3488_));
  OAI21_X1   g02484(.A1(new_n3486_), .A2(new_n3488_), .B(\A[580] ), .ZN(new_n3489_));
  INV_X1     g02485(.I(\A[580] ), .ZN(new_n3490_));
  NAND2_X1   g02486(.A1(\A[581] ), .A2(\A[582] ), .ZN(new_n3491_));
  INV_X1     g02487(.I(new_n3491_), .ZN(new_n3492_));
  NOR2_X1    g02488(.A1(\A[581] ), .A2(\A[582] ), .ZN(new_n3493_));
  OAI21_X1   g02489(.A1(new_n3492_), .A2(new_n3493_), .B(new_n3490_), .ZN(new_n3494_));
  NAND2_X1   g02490(.A1(new_n3489_), .A2(new_n3494_), .ZN(new_n3495_));
  AOI21_X1   g02491(.A1(new_n3479_), .A2(new_n3480_), .B(new_n3482_), .ZN(new_n3496_));
  AOI21_X1   g02492(.A1(new_n3490_), .A2(new_n3491_), .B(new_n3493_), .ZN(new_n3497_));
  NOR2_X1    g02493(.A1(new_n3496_), .A2(new_n3497_), .ZN(new_n3498_));
  NAND3_X1   g02494(.A1(new_n3484_), .A2(new_n3495_), .A3(new_n3498_), .ZN(new_n3499_));
  INV_X1     g02495(.I(\A[571] ), .ZN(new_n3500_));
  INV_X1     g02496(.I(\A[572] ), .ZN(new_n3501_));
  NAND2_X1   g02497(.A1(new_n3501_), .A2(\A[573] ), .ZN(new_n3502_));
  INV_X1     g02498(.I(\A[573] ), .ZN(new_n3503_));
  NAND2_X1   g02499(.A1(new_n3503_), .A2(\A[572] ), .ZN(new_n3504_));
  AOI21_X1   g02500(.A1(new_n3502_), .A2(new_n3504_), .B(new_n3500_), .ZN(new_n3505_));
  NAND2_X1   g02501(.A1(\A[572] ), .A2(\A[573] ), .ZN(new_n3506_));
  NOR2_X1    g02502(.A1(\A[572] ), .A2(\A[573] ), .ZN(new_n3507_));
  INV_X1     g02503(.I(new_n3507_), .ZN(new_n3508_));
  AOI21_X1   g02504(.A1(new_n3508_), .A2(new_n3506_), .B(\A[571] ), .ZN(new_n3509_));
  NOR2_X1    g02505(.A1(new_n3509_), .A2(new_n3505_), .ZN(new_n3510_));
  INV_X1     g02506(.I(\A[574] ), .ZN(new_n3511_));
  INV_X1     g02507(.I(\A[575] ), .ZN(new_n3512_));
  NAND2_X1   g02508(.A1(new_n3512_), .A2(\A[576] ), .ZN(new_n3513_));
  INV_X1     g02509(.I(\A[576] ), .ZN(new_n3514_));
  NAND2_X1   g02510(.A1(new_n3514_), .A2(\A[575] ), .ZN(new_n3515_));
  AOI21_X1   g02511(.A1(new_n3513_), .A2(new_n3515_), .B(new_n3511_), .ZN(new_n3516_));
  NAND2_X1   g02512(.A1(\A[575] ), .A2(\A[576] ), .ZN(new_n3517_));
  NOR2_X1    g02513(.A1(\A[575] ), .A2(\A[576] ), .ZN(new_n3518_));
  INV_X1     g02514(.I(new_n3518_), .ZN(new_n3519_));
  AOI21_X1   g02515(.A1(new_n3519_), .A2(new_n3517_), .B(\A[574] ), .ZN(new_n3520_));
  NOR2_X1    g02516(.A1(new_n3520_), .A2(new_n3516_), .ZN(new_n3521_));
  AOI21_X1   g02517(.A1(new_n3500_), .A2(new_n3506_), .B(new_n3507_), .ZN(new_n3522_));
  AOI21_X1   g02518(.A1(new_n3511_), .A2(new_n3517_), .B(new_n3518_), .ZN(new_n3523_));
  NOR2_X1    g02519(.A1(new_n3522_), .A2(new_n3523_), .ZN(new_n3524_));
  INV_X1     g02520(.I(new_n3524_), .ZN(new_n3525_));
  NOR3_X1    g02521(.A1(new_n3525_), .A2(new_n3510_), .A3(new_n3521_), .ZN(new_n3526_));
  XOR2_X1    g02522(.A1(new_n3526_), .A2(new_n3499_), .Z(new_n3527_));
  INV_X1     g02523(.I(\A[567] ), .ZN(new_n3528_));
  NOR2_X1    g02524(.A1(new_n3528_), .A2(\A[566] ), .ZN(new_n3529_));
  INV_X1     g02525(.I(\A[566] ), .ZN(new_n3530_));
  NOR2_X1    g02526(.A1(new_n3530_), .A2(\A[567] ), .ZN(new_n3531_));
  OAI21_X1   g02527(.A1(new_n3529_), .A2(new_n3531_), .B(\A[565] ), .ZN(new_n3532_));
  INV_X1     g02528(.I(\A[565] ), .ZN(new_n3533_));
  NAND2_X1   g02529(.A1(\A[566] ), .A2(\A[567] ), .ZN(new_n3534_));
  INV_X1     g02530(.I(new_n3534_), .ZN(new_n3535_));
  NOR2_X1    g02531(.A1(\A[566] ), .A2(\A[567] ), .ZN(new_n3536_));
  OAI21_X1   g02532(.A1(new_n3535_), .A2(new_n3536_), .B(new_n3533_), .ZN(new_n3537_));
  NAND2_X1   g02533(.A1(new_n3532_), .A2(new_n3537_), .ZN(new_n3538_));
  INV_X1     g02534(.I(\A[570] ), .ZN(new_n3539_));
  NOR2_X1    g02535(.A1(new_n3539_), .A2(\A[569] ), .ZN(new_n3540_));
  INV_X1     g02536(.I(\A[569] ), .ZN(new_n3541_));
  NOR2_X1    g02537(.A1(new_n3541_), .A2(\A[570] ), .ZN(new_n3542_));
  OAI21_X1   g02538(.A1(new_n3540_), .A2(new_n3542_), .B(\A[568] ), .ZN(new_n3543_));
  INV_X1     g02539(.I(\A[568] ), .ZN(new_n3544_));
  NAND2_X1   g02540(.A1(\A[569] ), .A2(\A[570] ), .ZN(new_n3545_));
  INV_X1     g02541(.I(new_n3545_), .ZN(new_n3546_));
  NOR2_X1    g02542(.A1(\A[569] ), .A2(\A[570] ), .ZN(new_n3547_));
  OAI21_X1   g02543(.A1(new_n3546_), .A2(new_n3547_), .B(new_n3544_), .ZN(new_n3548_));
  NAND2_X1   g02544(.A1(new_n3543_), .A2(new_n3548_), .ZN(new_n3549_));
  AOI21_X1   g02545(.A1(new_n3533_), .A2(new_n3534_), .B(new_n3536_), .ZN(new_n3550_));
  AOI21_X1   g02546(.A1(new_n3544_), .A2(new_n3545_), .B(new_n3547_), .ZN(new_n3551_));
  NOR2_X1    g02547(.A1(new_n3550_), .A2(new_n3551_), .ZN(new_n3552_));
  NAND3_X1   g02548(.A1(new_n3538_), .A2(new_n3549_), .A3(new_n3552_), .ZN(new_n3553_));
  INV_X1     g02549(.I(\A[559] ), .ZN(new_n3554_));
  INV_X1     g02550(.I(\A[560] ), .ZN(new_n3555_));
  NAND2_X1   g02551(.A1(new_n3555_), .A2(\A[561] ), .ZN(new_n3556_));
  INV_X1     g02552(.I(\A[561] ), .ZN(new_n3557_));
  NAND2_X1   g02553(.A1(new_n3557_), .A2(\A[560] ), .ZN(new_n3558_));
  AOI21_X1   g02554(.A1(new_n3556_), .A2(new_n3558_), .B(new_n3554_), .ZN(new_n3559_));
  NAND2_X1   g02555(.A1(\A[560] ), .A2(\A[561] ), .ZN(new_n3560_));
  NAND2_X1   g02556(.A1(new_n3555_), .A2(new_n3557_), .ZN(new_n3561_));
  AOI21_X1   g02557(.A1(new_n3561_), .A2(new_n3560_), .B(\A[559] ), .ZN(new_n3562_));
  NOR2_X1    g02558(.A1(new_n3562_), .A2(new_n3559_), .ZN(new_n3563_));
  INV_X1     g02559(.I(\A[562] ), .ZN(new_n3564_));
  INV_X1     g02560(.I(\A[563] ), .ZN(new_n3565_));
  NAND2_X1   g02561(.A1(new_n3565_), .A2(\A[564] ), .ZN(new_n3566_));
  INV_X1     g02562(.I(\A[564] ), .ZN(new_n3567_));
  NAND2_X1   g02563(.A1(new_n3567_), .A2(\A[563] ), .ZN(new_n3568_));
  AOI21_X1   g02564(.A1(new_n3566_), .A2(new_n3568_), .B(new_n3564_), .ZN(new_n3569_));
  NAND2_X1   g02565(.A1(\A[563] ), .A2(\A[564] ), .ZN(new_n3570_));
  NAND2_X1   g02566(.A1(new_n3565_), .A2(new_n3567_), .ZN(new_n3571_));
  AOI21_X1   g02567(.A1(new_n3571_), .A2(new_n3570_), .B(\A[562] ), .ZN(new_n3572_));
  NOR2_X1    g02568(.A1(new_n3572_), .A2(new_n3569_), .ZN(new_n3573_));
  NAND2_X1   g02569(.A1(new_n3560_), .A2(new_n3554_), .ZN(new_n3574_));
  NAND2_X1   g02570(.A1(new_n3574_), .A2(new_n3561_), .ZN(new_n3575_));
  NAND2_X1   g02571(.A1(new_n3570_), .A2(new_n3564_), .ZN(new_n3576_));
  NAND2_X1   g02572(.A1(new_n3576_), .A2(new_n3571_), .ZN(new_n3577_));
  NAND2_X1   g02573(.A1(new_n3575_), .A2(new_n3577_), .ZN(new_n3578_));
  NOR3_X1    g02574(.A1(new_n3563_), .A2(new_n3573_), .A3(new_n3578_), .ZN(new_n3579_));
  XOR2_X1    g02575(.A1(new_n3579_), .A2(new_n3553_), .Z(new_n3580_));
  NOR2_X1    g02576(.A1(new_n3527_), .A2(new_n3580_), .ZN(new_n3581_));
  XNOR2_X1   g02577(.A1(new_n3526_), .A2(new_n3499_), .ZN(new_n3582_));
  XNOR2_X1   g02578(.A1(new_n3579_), .A2(new_n3553_), .ZN(new_n3583_));
  NOR2_X1    g02579(.A1(new_n3582_), .A2(new_n3583_), .ZN(new_n3584_));
  NOR2_X1    g02580(.A1(new_n3584_), .A2(new_n3581_), .ZN(new_n3585_));
  NOR2_X1    g02581(.A1(new_n3473_), .A2(new_n3585_), .ZN(new_n3586_));
  NAND2_X1   g02582(.A1(new_n3473_), .A2(new_n3585_), .ZN(new_n3587_));
  INV_X1     g02583(.I(new_n3587_), .ZN(new_n3588_));
  NOR2_X1    g02584(.A1(new_n3588_), .A2(new_n3586_), .ZN(new_n3589_));
  NOR2_X1    g02585(.A1(new_n3362_), .A2(new_n3589_), .ZN(new_n3590_));
  NAND2_X1   g02586(.A1(new_n3362_), .A2(new_n3589_), .ZN(new_n3591_));
  INV_X1     g02587(.I(new_n3591_), .ZN(new_n3592_));
  NOR2_X1    g02588(.A1(new_n3592_), .A2(new_n3590_), .ZN(new_n3593_));
  NAND2_X1   g02589(.A1(new_n3137_), .A2(new_n3593_), .ZN(new_n3594_));
  INV_X1     g02590(.I(new_n3594_), .ZN(new_n3595_));
  NOR2_X1    g02591(.A1(new_n3137_), .A2(new_n3593_), .ZN(new_n3596_));
  NOR2_X1    g02592(.A1(new_n3595_), .A2(new_n3596_), .ZN(new_n3597_));
  INV_X1     g02593(.I(new_n3597_), .ZN(new_n3598_));
  NOR2_X1    g02594(.A1(new_n3598_), .A2(new_n2689_), .ZN(new_n3599_));
  NOR4_X1    g02595(.A1(new_n3163_), .A2(new_n3173_), .A3(new_n3184_), .A4(new_n3189_), .ZN(new_n3600_));
  INV_X1     g02596(.I(new_n3600_), .ZN(new_n3601_));
  INV_X1     g02597(.I(new_n3159_), .ZN(new_n3602_));
  INV_X1     g02598(.I(new_n3162_), .ZN(new_n3603_));
  NOR2_X1    g02599(.A1(new_n3603_), .A2(new_n3148_), .ZN(new_n3604_));
  NAND2_X1   g02600(.A1(new_n3140_), .A2(\A[651] ), .ZN(new_n3605_));
  NAND2_X1   g02601(.A1(new_n3138_), .A2(\A[650] ), .ZN(new_n3606_));
  AOI21_X1   g02602(.A1(new_n3605_), .A2(new_n3606_), .B(new_n3143_), .ZN(new_n3607_));
  INV_X1     g02603(.I(new_n3146_), .ZN(new_n3608_));
  AOI21_X1   g02604(.A1(new_n3608_), .A2(new_n3144_), .B(\A[649] ), .ZN(new_n3609_));
  NOR2_X1    g02605(.A1(new_n3609_), .A2(new_n3607_), .ZN(new_n3610_));
  NOR2_X1    g02606(.A1(new_n3610_), .A2(new_n3162_), .ZN(new_n3611_));
  OAI21_X1   g02607(.A1(new_n3604_), .A2(new_n3611_), .B(new_n3602_), .ZN(new_n3612_));
  NAND2_X1   g02608(.A1(new_n3610_), .A2(new_n3162_), .ZN(new_n3613_));
  NAND2_X1   g02609(.A1(new_n3603_), .A2(new_n3148_), .ZN(new_n3614_));
  NAND3_X1   g02610(.A1(new_n3614_), .A2(new_n3613_), .A3(new_n3159_), .ZN(new_n3615_));
  XOR2_X1    g02611(.A1(new_n3148_), .A2(new_n3159_), .Z(new_n3616_));
  NAND2_X1   g02612(.A1(new_n3616_), .A2(new_n3162_), .ZN(new_n3617_));
  NAND3_X1   g02613(.A1(new_n3617_), .A2(new_n3612_), .A3(new_n3615_), .ZN(new_n3618_));
  NAND2_X1   g02614(.A1(new_n3612_), .A2(new_n3615_), .ZN(new_n3619_));
  NOR2_X1    g02615(.A1(new_n3173_), .A2(new_n3184_), .ZN(new_n3620_));
  INV_X1     g02616(.I(new_n3173_), .ZN(new_n3621_));
  INV_X1     g02617(.I(new_n3184_), .ZN(new_n3622_));
  NOR2_X1    g02618(.A1(new_n3621_), .A2(new_n3622_), .ZN(new_n3623_));
  NOR2_X1    g02619(.A1(new_n3623_), .A2(new_n3620_), .ZN(new_n3624_));
  NOR3_X1    g02620(.A1(new_n3173_), .A2(new_n3189_), .A3(new_n3184_), .ZN(new_n3625_));
  NOR3_X1    g02621(.A1(new_n3624_), .A2(new_n3163_), .A3(new_n3625_), .ZN(new_n3626_));
  NOR2_X1    g02622(.A1(new_n3621_), .A2(new_n3189_), .ZN(new_n3627_));
  INV_X1     g02623(.I(new_n3186_), .ZN(new_n3628_));
  NOR2_X1    g02624(.A1(new_n3628_), .A2(new_n3187_), .ZN(new_n3629_));
  NOR2_X1    g02625(.A1(new_n3629_), .A2(new_n3173_), .ZN(new_n3630_));
  OAI21_X1   g02626(.A1(new_n3627_), .A2(new_n3630_), .B(new_n3184_), .ZN(new_n3631_));
  NAND2_X1   g02627(.A1(new_n3629_), .A2(new_n3173_), .ZN(new_n3632_));
  NAND2_X1   g02628(.A1(new_n3621_), .A2(new_n3189_), .ZN(new_n3633_));
  NAND3_X1   g02629(.A1(new_n3633_), .A2(new_n3632_), .A3(new_n3622_), .ZN(new_n3634_));
  NAND2_X1   g02630(.A1(new_n3631_), .A2(new_n3634_), .ZN(new_n3635_));
  NAND4_X1   g02631(.A1(new_n3626_), .A2(new_n3635_), .A3(new_n3619_), .A4(new_n3617_), .ZN(new_n3636_));
  AOI21_X1   g02632(.A1(new_n3636_), .A2(new_n3618_), .B(new_n3601_), .ZN(new_n3637_));
  INV_X1     g02633(.I(new_n3637_), .ZN(new_n3638_));
  INV_X1     g02634(.I(new_n3635_), .ZN(new_n3639_));
  XOR2_X1    g02635(.A1(new_n3618_), .A2(new_n3601_), .Z(new_n3640_));
  NAND2_X1   g02636(.A1(new_n3640_), .A2(new_n3639_), .ZN(new_n3641_));
  NAND4_X1   g02637(.A1(new_n3243_), .A2(new_n3202_), .A3(new_n3213_), .A4(new_n3216_), .ZN(new_n3642_));
  INV_X1     g02638(.I(new_n3213_), .ZN(new_n3643_));
  XOR2_X1    g02639(.A1(new_n3202_), .A2(new_n3216_), .Z(new_n3644_));
  NAND2_X1   g02640(.A1(new_n3644_), .A2(new_n3643_), .ZN(new_n3645_));
  XNOR2_X1   g02641(.A1(new_n3202_), .A2(new_n3216_), .ZN(new_n3646_));
  NAND2_X1   g02642(.A1(new_n3646_), .A2(new_n3213_), .ZN(new_n3647_));
  XOR2_X1    g02643(.A1(new_n3202_), .A2(new_n3213_), .Z(new_n3648_));
  NAND2_X1   g02644(.A1(new_n3648_), .A2(new_n3216_), .ZN(new_n3649_));
  NAND4_X1   g02645(.A1(new_n3649_), .A2(new_n3647_), .A3(new_n3645_), .A4(new_n3642_), .ZN(new_n3650_));
  INV_X1     g02646(.I(new_n3237_), .ZN(new_n3651_));
  NAND3_X1   g02647(.A1(new_n3227_), .A2(new_n3239_), .A3(new_n3241_), .ZN(new_n3652_));
  INV_X1     g02648(.I(new_n3227_), .ZN(new_n3653_));
  NAND2_X1   g02649(.A1(new_n3653_), .A2(new_n3242_), .ZN(new_n3654_));
  AOI21_X1   g02650(.A1(new_n3654_), .A2(new_n3652_), .B(new_n3651_), .ZN(new_n3655_));
  INV_X1     g02651(.I(new_n3655_), .ZN(new_n3656_));
  NAND3_X1   g02652(.A1(new_n3654_), .A2(new_n3651_), .A3(new_n3652_), .ZN(new_n3657_));
  NAND2_X1   g02653(.A1(new_n3656_), .A2(new_n3657_), .ZN(new_n3658_));
  INV_X1     g02654(.I(new_n3202_), .ZN(new_n3659_));
  INV_X1     g02655(.I(new_n3216_), .ZN(new_n3660_));
  XOR2_X1    g02656(.A1(new_n3227_), .A2(new_n3237_), .Z(new_n3661_));
  NOR3_X1    g02657(.A1(new_n3227_), .A2(new_n3237_), .A3(new_n3242_), .ZN(new_n3662_));
  NOR4_X1    g02658(.A1(new_n3661_), .A2(new_n3659_), .A3(new_n3643_), .A4(new_n3660_), .ZN(new_n3663_));
  INV_X1     g02659(.I(new_n3663_), .ZN(new_n3664_));
  NAND3_X1   g02660(.A1(new_n3650_), .A2(new_n3664_), .A3(new_n3658_), .ZN(new_n3665_));
  NOR2_X1    g02661(.A1(new_n3665_), .A2(new_n3246_), .ZN(new_n3666_));
  NAND2_X1   g02662(.A1(new_n3641_), .A2(new_n3666_), .ZN(new_n3667_));
  INV_X1     g02663(.I(new_n3642_), .ZN(new_n3668_));
  NOR2_X1    g02664(.A1(new_n3646_), .A2(new_n3213_), .ZN(new_n3669_));
  NOR2_X1    g02665(.A1(new_n3644_), .A2(new_n3643_), .ZN(new_n3670_));
  XNOR2_X1   g02666(.A1(new_n3202_), .A2(new_n3213_), .ZN(new_n3671_));
  NOR2_X1    g02667(.A1(new_n3671_), .A2(new_n3660_), .ZN(new_n3672_));
  NOR4_X1    g02668(.A1(new_n3672_), .A2(new_n3669_), .A3(new_n3668_), .A4(new_n3670_), .ZN(new_n3673_));
  INV_X1     g02669(.I(new_n3657_), .ZN(new_n3674_));
  NOR2_X1    g02670(.A1(new_n3674_), .A2(new_n3655_), .ZN(new_n3675_));
  NOR3_X1    g02671(.A1(new_n3673_), .A2(new_n3675_), .A3(new_n3663_), .ZN(new_n3676_));
  NAND2_X1   g02672(.A1(new_n3676_), .A2(new_n3247_), .ZN(new_n3677_));
  NAND3_X1   g02673(.A1(new_n3640_), .A2(new_n3677_), .A3(new_n3639_), .ZN(new_n3678_));
  AOI21_X1   g02674(.A1(new_n3667_), .A2(new_n3678_), .B(new_n3638_), .ZN(new_n3679_));
  INV_X1     g02675(.I(new_n3679_), .ZN(new_n3680_));
  INV_X1     g02676(.I(new_n3284_), .ZN(new_n3681_));
  NOR2_X1    g02677(.A1(new_n3681_), .A2(new_n3300_), .ZN(new_n3682_));
  INV_X1     g02678(.I(new_n3297_), .ZN(new_n3683_));
  AOI21_X1   g02679(.A1(new_n3285_), .A2(new_n3291_), .B(new_n3292_), .ZN(new_n3684_));
  NOR2_X1    g02680(.A1(new_n3683_), .A2(new_n3684_), .ZN(new_n3685_));
  NOR2_X1    g02681(.A1(new_n3685_), .A2(new_n3284_), .ZN(new_n3686_));
  OAI21_X1   g02682(.A1(new_n3682_), .A2(new_n3686_), .B(new_n3295_), .ZN(new_n3687_));
  OR2_X2     g02683(.A1(new_n3294_), .A2(new_n3290_), .Z(new_n3688_));
  NAND2_X1   g02684(.A1(new_n3685_), .A2(new_n3284_), .ZN(new_n3689_));
  NAND2_X1   g02685(.A1(new_n3681_), .A2(new_n3300_), .ZN(new_n3690_));
  NAND3_X1   g02686(.A1(new_n3690_), .A2(new_n3689_), .A3(new_n3688_), .ZN(new_n3691_));
  NAND2_X1   g02687(.A1(new_n3687_), .A2(new_n3691_), .ZN(new_n3692_));
  NOR4_X1    g02688(.A1(new_n3274_), .A2(new_n3284_), .A3(new_n3295_), .A4(new_n3300_), .ZN(new_n3693_));
  INV_X1     g02689(.I(new_n3693_), .ZN(new_n3694_));
  INV_X1     g02690(.I(new_n3270_), .ZN(new_n3695_));
  NAND2_X1   g02691(.A1(new_n3251_), .A2(\A[627] ), .ZN(new_n3696_));
  NAND2_X1   g02692(.A1(new_n3249_), .A2(\A[626] ), .ZN(new_n3697_));
  AOI21_X1   g02693(.A1(new_n3696_), .A2(new_n3697_), .B(new_n3254_), .ZN(new_n3698_));
  INV_X1     g02694(.I(new_n3257_), .ZN(new_n3699_));
  AOI21_X1   g02695(.A1(new_n3699_), .A2(new_n3255_), .B(\A[625] ), .ZN(new_n3700_));
  NOR2_X1    g02696(.A1(new_n3700_), .A2(new_n3698_), .ZN(new_n3701_));
  NAND2_X1   g02697(.A1(new_n3701_), .A2(new_n3273_), .ZN(new_n3702_));
  INV_X1     g02698(.I(new_n3702_), .ZN(new_n3703_));
  NOR2_X1    g02699(.A1(new_n3701_), .A2(new_n3273_), .ZN(new_n3704_));
  OAI21_X1   g02700(.A1(new_n3703_), .A2(new_n3704_), .B(new_n3695_), .ZN(new_n3705_));
  INV_X1     g02701(.I(new_n3273_), .ZN(new_n3706_));
  NAND2_X1   g02702(.A1(new_n3706_), .A2(new_n3259_), .ZN(new_n3707_));
  NAND3_X1   g02703(.A1(new_n3707_), .A2(new_n3702_), .A3(new_n3270_), .ZN(new_n3708_));
  NAND2_X1   g02704(.A1(new_n3705_), .A2(new_n3708_), .ZN(new_n3709_));
  XOR2_X1    g02705(.A1(new_n3701_), .A2(new_n3270_), .Z(new_n3710_));
  NOR2_X1    g02706(.A1(new_n3710_), .A2(new_n3706_), .ZN(new_n3711_));
  NOR2_X1    g02707(.A1(new_n3709_), .A2(new_n3711_), .ZN(new_n3712_));
  NAND2_X1   g02708(.A1(new_n3712_), .A2(new_n3694_), .ZN(new_n3713_));
  XOR2_X1    g02709(.A1(new_n3259_), .A2(new_n3270_), .Z(new_n3714_));
  NAND2_X1   g02710(.A1(new_n3714_), .A2(new_n3273_), .ZN(new_n3715_));
  NAND3_X1   g02711(.A1(new_n3715_), .A2(new_n3705_), .A3(new_n3708_), .ZN(new_n3716_));
  NAND2_X1   g02712(.A1(new_n3716_), .A2(new_n3693_), .ZN(new_n3717_));
  AOI21_X1   g02713(.A1(new_n3713_), .A2(new_n3717_), .B(new_n3692_), .ZN(new_n3718_));
  INV_X1     g02714(.I(new_n3718_), .ZN(new_n3719_));
  NOR2_X1    g02715(.A1(new_n3284_), .A2(new_n3295_), .ZN(new_n3720_));
  NOR2_X1    g02716(.A1(new_n3681_), .A2(new_n3688_), .ZN(new_n3721_));
  NOR2_X1    g02717(.A1(new_n3721_), .A2(new_n3720_), .ZN(new_n3722_));
  NOR3_X1    g02718(.A1(new_n3284_), .A2(new_n3295_), .A3(new_n3300_), .ZN(new_n3723_));
  NOR3_X1    g02719(.A1(new_n3722_), .A2(new_n3274_), .A3(new_n3723_), .ZN(new_n3724_));
  NAND4_X1   g02720(.A1(new_n3692_), .A2(new_n3724_), .A3(new_n3709_), .A4(new_n3715_), .ZN(new_n3725_));
  AOI21_X1   g02721(.A1(new_n3725_), .A2(new_n3716_), .B(new_n3694_), .ZN(new_n3726_));
  NOR4_X1    g02722(.A1(new_n3328_), .A2(new_n3338_), .A3(new_n3348_), .A4(new_n3353_), .ZN(new_n3727_));
  INV_X1     g02723(.I(new_n3727_), .ZN(new_n3728_));
  INV_X1     g02724(.I(new_n3324_), .ZN(new_n3729_));
  INV_X1     g02725(.I(new_n3327_), .ZN(new_n3730_));
  NOR2_X1    g02726(.A1(new_n3730_), .A2(new_n3313_), .ZN(new_n3731_));
  AND2_X2    g02727(.A1(new_n3307_), .A2(new_n3312_), .Z(new_n3732_));
  NOR2_X1    g02728(.A1(new_n3732_), .A2(new_n3327_), .ZN(new_n3733_));
  OAI21_X1   g02729(.A1(new_n3733_), .A2(new_n3731_), .B(new_n3729_), .ZN(new_n3734_));
  NOR3_X1    g02730(.A1(new_n3733_), .A2(new_n3729_), .A3(new_n3731_), .ZN(new_n3735_));
  INV_X1     g02731(.I(new_n3735_), .ZN(new_n3736_));
  XOR2_X1    g02732(.A1(new_n3313_), .A2(new_n3324_), .Z(new_n3737_));
  NAND2_X1   g02733(.A1(new_n3737_), .A2(new_n3327_), .ZN(new_n3738_));
  NAND4_X1   g02734(.A1(new_n3738_), .A2(new_n3736_), .A3(new_n3728_), .A4(new_n3734_), .ZN(new_n3739_));
  INV_X1     g02735(.I(new_n3348_), .ZN(new_n3740_));
  NAND3_X1   g02736(.A1(new_n3338_), .A2(new_n3350_), .A3(new_n3352_), .ZN(new_n3741_));
  INV_X1     g02737(.I(new_n3338_), .ZN(new_n3742_));
  NAND2_X1   g02738(.A1(new_n3742_), .A2(new_n3353_), .ZN(new_n3743_));
  AOI21_X1   g02739(.A1(new_n3743_), .A2(new_n3741_), .B(new_n3740_), .ZN(new_n3744_));
  INV_X1     g02740(.I(new_n3744_), .ZN(new_n3745_));
  NAND3_X1   g02741(.A1(new_n3743_), .A2(new_n3740_), .A3(new_n3741_), .ZN(new_n3746_));
  NAND2_X1   g02742(.A1(new_n3745_), .A2(new_n3746_), .ZN(new_n3747_));
  XNOR2_X1   g02743(.A1(new_n3338_), .A2(new_n3348_), .ZN(new_n3748_));
  NOR3_X1    g02744(.A1(new_n3338_), .A2(new_n3348_), .A3(new_n3353_), .ZN(new_n3749_));
  NAND4_X1   g02745(.A1(new_n3748_), .A2(new_n3313_), .A3(new_n3324_), .A4(new_n3327_), .ZN(new_n3750_));
  NAND4_X1   g02746(.A1(new_n3357_), .A2(new_n3739_), .A3(new_n3747_), .A4(new_n3750_), .ZN(new_n3751_));
  NOR2_X1    g02747(.A1(new_n3751_), .A2(new_n3726_), .ZN(new_n3752_));
  AND2_X2    g02748(.A1(new_n3687_), .A2(new_n3691_), .Z(new_n3753_));
  NAND3_X1   g02749(.A1(new_n3724_), .A2(new_n3709_), .A3(new_n3715_), .ZN(new_n3754_));
  NOR2_X1    g02750(.A1(new_n3754_), .A2(new_n3753_), .ZN(new_n3755_));
  OAI21_X1   g02751(.A1(new_n3755_), .A2(new_n3712_), .B(new_n3693_), .ZN(new_n3756_));
  NAND2_X1   g02752(.A1(new_n3302_), .A2(new_n3355_), .ZN(new_n3757_));
  NAND3_X1   g02753(.A1(new_n3739_), .A2(new_n3747_), .A3(new_n3750_), .ZN(new_n3758_));
  NOR2_X1    g02754(.A1(new_n3758_), .A2(new_n3757_), .ZN(new_n3759_));
  NOR2_X1    g02755(.A1(new_n3756_), .A2(new_n3759_), .ZN(new_n3760_));
  OAI21_X1   g02756(.A1(new_n3760_), .A2(new_n3752_), .B(new_n3719_), .ZN(new_n3761_));
  NAND2_X1   g02757(.A1(new_n3756_), .A2(new_n3759_), .ZN(new_n3762_));
  NAND2_X1   g02758(.A1(new_n3751_), .A2(new_n3726_), .ZN(new_n3763_));
  NAND3_X1   g02759(.A1(new_n3762_), .A2(new_n3718_), .A3(new_n3763_), .ZN(new_n3764_));
  AOI21_X1   g02760(.A1(new_n3761_), .A2(new_n3764_), .B(new_n3360_), .ZN(new_n3765_));
  NOR2_X1    g02761(.A1(new_n3680_), .A2(new_n3765_), .ZN(new_n3766_));
  NOR4_X1    g02762(.A1(new_n3388_), .A2(new_n3398_), .A3(new_n3409_), .A4(new_n3414_), .ZN(new_n3767_));
  INV_X1     g02763(.I(new_n3767_), .ZN(new_n3768_));
  INV_X1     g02764(.I(new_n3384_), .ZN(new_n3769_));
  INV_X1     g02765(.I(new_n3387_), .ZN(new_n3770_));
  NOR2_X1    g02766(.A1(new_n3770_), .A2(new_n3373_), .ZN(new_n3771_));
  NAND2_X1   g02767(.A1(new_n3365_), .A2(\A[603] ), .ZN(new_n3772_));
  NAND2_X1   g02768(.A1(new_n3363_), .A2(\A[602] ), .ZN(new_n3773_));
  AOI21_X1   g02769(.A1(new_n3772_), .A2(new_n3773_), .B(new_n3368_), .ZN(new_n3774_));
  INV_X1     g02770(.I(new_n3371_), .ZN(new_n3775_));
  AOI21_X1   g02771(.A1(new_n3775_), .A2(new_n3369_), .B(\A[601] ), .ZN(new_n3776_));
  NOR2_X1    g02772(.A1(new_n3776_), .A2(new_n3774_), .ZN(new_n3777_));
  NOR2_X1    g02773(.A1(new_n3777_), .A2(new_n3387_), .ZN(new_n3778_));
  OAI21_X1   g02774(.A1(new_n3771_), .A2(new_n3778_), .B(new_n3769_), .ZN(new_n3779_));
  NAND2_X1   g02775(.A1(new_n3777_), .A2(new_n3387_), .ZN(new_n3780_));
  NAND2_X1   g02776(.A1(new_n3770_), .A2(new_n3373_), .ZN(new_n3781_));
  NAND3_X1   g02777(.A1(new_n3781_), .A2(new_n3780_), .A3(new_n3384_), .ZN(new_n3782_));
  XOR2_X1    g02778(.A1(new_n3373_), .A2(new_n3384_), .Z(new_n3783_));
  NAND2_X1   g02779(.A1(new_n3783_), .A2(new_n3387_), .ZN(new_n3784_));
  NAND3_X1   g02780(.A1(new_n3784_), .A2(new_n3779_), .A3(new_n3782_), .ZN(new_n3785_));
  NAND2_X1   g02781(.A1(new_n3779_), .A2(new_n3782_), .ZN(new_n3786_));
  NOR2_X1    g02782(.A1(new_n3398_), .A2(new_n3409_), .ZN(new_n3787_));
  OR2_X2     g02783(.A1(new_n3397_), .A2(new_n3394_), .Z(new_n3788_));
  OR2_X2     g02784(.A1(new_n3408_), .A2(new_n3404_), .Z(new_n3789_));
  NOR2_X1    g02785(.A1(new_n3788_), .A2(new_n3789_), .ZN(new_n3790_));
  NOR2_X1    g02786(.A1(new_n3790_), .A2(new_n3787_), .ZN(new_n3791_));
  NOR3_X1    g02787(.A1(new_n3398_), .A2(new_n3414_), .A3(new_n3409_), .ZN(new_n3792_));
  NOR3_X1    g02788(.A1(new_n3791_), .A2(new_n3388_), .A3(new_n3792_), .ZN(new_n3793_));
  NOR2_X1    g02789(.A1(new_n3788_), .A2(new_n3414_), .ZN(new_n3794_));
  AND2_X2    g02790(.A1(new_n3410_), .A2(new_n3396_), .Z(new_n3795_));
  NOR2_X1    g02791(.A1(new_n3795_), .A2(new_n3412_), .ZN(new_n3796_));
  NOR2_X1    g02792(.A1(new_n3796_), .A2(new_n3398_), .ZN(new_n3797_));
  OAI21_X1   g02793(.A1(new_n3794_), .A2(new_n3797_), .B(new_n3409_), .ZN(new_n3798_));
  NAND2_X1   g02794(.A1(new_n3796_), .A2(new_n3398_), .ZN(new_n3799_));
  NAND2_X1   g02795(.A1(new_n3788_), .A2(new_n3414_), .ZN(new_n3800_));
  NAND3_X1   g02796(.A1(new_n3800_), .A2(new_n3799_), .A3(new_n3789_), .ZN(new_n3801_));
  NAND2_X1   g02797(.A1(new_n3798_), .A2(new_n3801_), .ZN(new_n3802_));
  NAND4_X1   g02798(.A1(new_n3793_), .A2(new_n3802_), .A3(new_n3786_), .A4(new_n3784_), .ZN(new_n3803_));
  AOI21_X1   g02799(.A1(new_n3803_), .A2(new_n3785_), .B(new_n3768_), .ZN(new_n3804_));
  INV_X1     g02800(.I(new_n3804_), .ZN(new_n3805_));
  AND2_X2    g02801(.A1(new_n3798_), .A2(new_n3801_), .Z(new_n3806_));
  XOR2_X1    g02802(.A1(new_n3785_), .A2(new_n3768_), .Z(new_n3807_));
  NAND2_X1   g02803(.A1(new_n3807_), .A2(new_n3806_), .ZN(new_n3808_));
  NOR4_X1    g02804(.A1(new_n3442_), .A2(new_n3452_), .A3(new_n3462_), .A4(new_n3467_), .ZN(new_n3809_));
  INV_X1     g02805(.I(new_n3809_), .ZN(new_n3810_));
  INV_X1     g02806(.I(new_n3438_), .ZN(new_n3811_));
  INV_X1     g02807(.I(new_n3441_), .ZN(new_n3812_));
  NOR2_X1    g02808(.A1(new_n3812_), .A2(new_n3427_), .ZN(new_n3813_));
  INV_X1     g02809(.I(new_n3427_), .ZN(new_n3814_));
  NOR2_X1    g02810(.A1(new_n3814_), .A2(new_n3441_), .ZN(new_n3815_));
  OAI21_X1   g02811(.A1(new_n3815_), .A2(new_n3813_), .B(new_n3811_), .ZN(new_n3816_));
  NOR3_X1    g02812(.A1(new_n3815_), .A2(new_n3811_), .A3(new_n3813_), .ZN(new_n3817_));
  INV_X1     g02813(.I(new_n3817_), .ZN(new_n3818_));
  XOR2_X1    g02814(.A1(new_n3427_), .A2(new_n3438_), .Z(new_n3819_));
  NAND2_X1   g02815(.A1(new_n3819_), .A2(new_n3441_), .ZN(new_n3820_));
  NAND3_X1   g02816(.A1(new_n3818_), .A2(new_n3820_), .A3(new_n3816_), .ZN(new_n3821_));
  INV_X1     g02817(.I(new_n3462_), .ZN(new_n3822_));
  NAND3_X1   g02818(.A1(new_n3452_), .A2(new_n3464_), .A3(new_n3466_), .ZN(new_n3823_));
  OR2_X2     g02819(.A1(new_n3451_), .A2(new_n3448_), .Z(new_n3824_));
  NAND2_X1   g02820(.A1(new_n3824_), .A2(new_n3467_), .ZN(new_n3825_));
  AOI21_X1   g02821(.A1(new_n3825_), .A2(new_n3823_), .B(new_n3822_), .ZN(new_n3826_));
  INV_X1     g02822(.I(new_n3826_), .ZN(new_n3827_));
  NAND3_X1   g02823(.A1(new_n3825_), .A2(new_n3822_), .A3(new_n3823_), .ZN(new_n3828_));
  NAND2_X1   g02824(.A1(new_n3827_), .A2(new_n3828_), .ZN(new_n3829_));
  XOR2_X1    g02825(.A1(new_n3452_), .A2(new_n3462_), .Z(new_n3830_));
  NOR3_X1    g02826(.A1(new_n3452_), .A2(new_n3462_), .A3(new_n3467_), .ZN(new_n3831_));
  NOR2_X1    g02827(.A1(new_n3830_), .A2(new_n3831_), .ZN(new_n3832_));
  NAND4_X1   g02828(.A1(new_n3832_), .A2(new_n3427_), .A3(new_n3438_), .A4(new_n3441_), .ZN(new_n3833_));
  NAND4_X1   g02829(.A1(new_n3833_), .A2(new_n3821_), .A3(new_n3829_), .A4(new_n3810_), .ZN(new_n3834_));
  NOR2_X1    g02830(.A1(new_n3834_), .A2(new_n3471_), .ZN(new_n3835_));
  NAND2_X1   g02831(.A1(new_n3808_), .A2(new_n3835_), .ZN(new_n3836_));
  INV_X1     g02832(.I(new_n3816_), .ZN(new_n3837_));
  XNOR2_X1   g02833(.A1(new_n3427_), .A2(new_n3438_), .ZN(new_n3838_));
  NOR2_X1    g02834(.A1(new_n3838_), .A2(new_n3812_), .ZN(new_n3839_));
  NOR4_X1    g02835(.A1(new_n3839_), .A2(new_n3837_), .A3(new_n3809_), .A4(new_n3817_), .ZN(new_n3840_));
  INV_X1     g02836(.I(new_n3828_), .ZN(new_n3841_));
  NOR2_X1    g02837(.A1(new_n3841_), .A2(new_n3826_), .ZN(new_n3842_));
  NOR4_X1    g02838(.A1(new_n3830_), .A2(new_n3814_), .A3(new_n3811_), .A4(new_n3812_), .ZN(new_n3843_));
  NOR3_X1    g02839(.A1(new_n3840_), .A2(new_n3842_), .A3(new_n3843_), .ZN(new_n3844_));
  NAND2_X1   g02840(.A1(new_n3844_), .A2(new_n3472_), .ZN(new_n3845_));
  NAND3_X1   g02841(.A1(new_n3845_), .A2(new_n3807_), .A3(new_n3806_), .ZN(new_n3846_));
  AOI21_X1   g02842(.A1(new_n3836_), .A2(new_n3846_), .B(new_n3805_), .ZN(new_n3847_));
  INV_X1     g02843(.I(new_n3847_), .ZN(new_n3848_));
  NAND2_X1   g02844(.A1(new_n3510_), .A2(new_n3524_), .ZN(new_n3849_));
  INV_X1     g02845(.I(new_n3849_), .ZN(new_n3850_));
  NOR2_X1    g02846(.A1(new_n3510_), .A2(new_n3524_), .ZN(new_n3851_));
  OAI21_X1   g02847(.A1(new_n3850_), .A2(new_n3851_), .B(new_n3521_), .ZN(new_n3852_));
  INV_X1     g02848(.I(new_n3521_), .ZN(new_n3853_));
  INV_X1     g02849(.I(new_n3851_), .ZN(new_n3854_));
  NAND3_X1   g02850(.A1(new_n3854_), .A2(new_n3849_), .A3(new_n3853_), .ZN(new_n3855_));
  NAND2_X1   g02851(.A1(new_n3852_), .A2(new_n3855_), .ZN(new_n3856_));
  NOR4_X1    g02852(.A1(new_n3499_), .A2(new_n3510_), .A3(new_n3521_), .A4(new_n3525_), .ZN(new_n3857_));
  INV_X1     g02853(.I(new_n3857_), .ZN(new_n3858_));
  INV_X1     g02854(.I(new_n3495_), .ZN(new_n3859_));
  INV_X1     g02855(.I(new_n3498_), .ZN(new_n3860_));
  NOR2_X1    g02856(.A1(new_n3860_), .A2(new_n3484_), .ZN(new_n3861_));
  NAND2_X1   g02857(.A1(new_n3476_), .A2(\A[579] ), .ZN(new_n3862_));
  NAND2_X1   g02858(.A1(new_n3474_), .A2(\A[578] ), .ZN(new_n3863_));
  AOI21_X1   g02859(.A1(new_n3862_), .A2(new_n3863_), .B(new_n3479_), .ZN(new_n3864_));
  INV_X1     g02860(.I(new_n3482_), .ZN(new_n3865_));
  AOI21_X1   g02861(.A1(new_n3865_), .A2(new_n3480_), .B(\A[577] ), .ZN(new_n3866_));
  NOR2_X1    g02862(.A1(new_n3866_), .A2(new_n3864_), .ZN(new_n3867_));
  NOR2_X1    g02863(.A1(new_n3867_), .A2(new_n3498_), .ZN(new_n3868_));
  OAI21_X1   g02864(.A1(new_n3861_), .A2(new_n3868_), .B(new_n3859_), .ZN(new_n3869_));
  NAND2_X1   g02865(.A1(new_n3867_), .A2(new_n3498_), .ZN(new_n3870_));
  NAND2_X1   g02866(.A1(new_n3860_), .A2(new_n3484_), .ZN(new_n3871_));
  NAND3_X1   g02867(.A1(new_n3871_), .A2(new_n3870_), .A3(new_n3495_), .ZN(new_n3872_));
  NAND2_X1   g02868(.A1(new_n3869_), .A2(new_n3872_), .ZN(new_n3873_));
  XOR2_X1    g02869(.A1(new_n3484_), .A2(new_n3495_), .Z(new_n3874_));
  AOI21_X1   g02870(.A1(new_n3498_), .A2(new_n3874_), .B(new_n3873_), .ZN(new_n3875_));
  NAND2_X1   g02871(.A1(new_n3875_), .A2(new_n3858_), .ZN(new_n3876_));
  NAND2_X1   g02872(.A1(new_n3874_), .A2(new_n3498_), .ZN(new_n3877_));
  NAND3_X1   g02873(.A1(new_n3877_), .A2(new_n3869_), .A3(new_n3872_), .ZN(new_n3878_));
  NAND2_X1   g02874(.A1(new_n3878_), .A2(new_n3857_), .ZN(new_n3879_));
  AOI21_X1   g02875(.A1(new_n3876_), .A2(new_n3879_), .B(new_n3856_), .ZN(new_n3880_));
  INV_X1     g02876(.I(new_n3880_), .ZN(new_n3881_));
  XOR2_X1    g02877(.A1(new_n3510_), .A2(new_n3521_), .Z(new_n3882_));
  NOR3_X1    g02878(.A1(new_n3525_), .A2(new_n3510_), .A3(new_n3521_), .ZN(new_n3883_));
  NOR3_X1    g02879(.A1(new_n3882_), .A2(new_n3499_), .A3(new_n3883_), .ZN(new_n3884_));
  NAND4_X1   g02880(.A1(new_n3856_), .A2(new_n3884_), .A3(new_n3877_), .A4(new_n3873_), .ZN(new_n3885_));
  AOI21_X1   g02881(.A1(new_n3885_), .A2(new_n3878_), .B(new_n3858_), .ZN(new_n3886_));
  NOR4_X1    g02882(.A1(new_n3553_), .A2(new_n3563_), .A3(new_n3573_), .A4(new_n3578_), .ZN(new_n3887_));
  INV_X1     g02883(.I(new_n3887_), .ZN(new_n3888_));
  INV_X1     g02884(.I(new_n3549_), .ZN(new_n3889_));
  INV_X1     g02885(.I(new_n3552_), .ZN(new_n3890_));
  NOR2_X1    g02886(.A1(new_n3890_), .A2(new_n3538_), .ZN(new_n3891_));
  INV_X1     g02887(.I(new_n3538_), .ZN(new_n3892_));
  NOR2_X1    g02888(.A1(new_n3892_), .A2(new_n3552_), .ZN(new_n3893_));
  OAI21_X1   g02889(.A1(new_n3893_), .A2(new_n3891_), .B(new_n3889_), .ZN(new_n3894_));
  NOR3_X1    g02890(.A1(new_n3893_), .A2(new_n3889_), .A3(new_n3891_), .ZN(new_n3895_));
  INV_X1     g02891(.I(new_n3895_), .ZN(new_n3896_));
  XOR2_X1    g02892(.A1(new_n3538_), .A2(new_n3549_), .Z(new_n3897_));
  NAND2_X1   g02893(.A1(new_n3897_), .A2(new_n3552_), .ZN(new_n3898_));
  NAND4_X1   g02894(.A1(new_n3896_), .A2(new_n3898_), .A3(new_n3888_), .A4(new_n3894_), .ZN(new_n3899_));
  INV_X1     g02895(.I(new_n3573_), .ZN(new_n3900_));
  NAND3_X1   g02896(.A1(new_n3563_), .A2(new_n3575_), .A3(new_n3577_), .ZN(new_n3901_));
  INV_X1     g02897(.I(new_n3563_), .ZN(new_n3902_));
  NAND2_X1   g02898(.A1(new_n3902_), .A2(new_n3578_), .ZN(new_n3903_));
  AOI21_X1   g02899(.A1(new_n3903_), .A2(new_n3901_), .B(new_n3900_), .ZN(new_n3904_));
  INV_X1     g02900(.I(new_n3904_), .ZN(new_n3905_));
  NAND3_X1   g02901(.A1(new_n3903_), .A2(new_n3900_), .A3(new_n3901_), .ZN(new_n3906_));
  NAND2_X1   g02902(.A1(new_n3905_), .A2(new_n3906_), .ZN(new_n3907_));
  NOR2_X1    g02903(.A1(new_n3563_), .A2(new_n3573_), .ZN(new_n3908_));
  NOR2_X1    g02904(.A1(new_n3902_), .A2(new_n3900_), .ZN(new_n3909_));
  OR2_X2     g02905(.A1(new_n3909_), .A2(new_n3908_), .Z(new_n3910_));
  NOR3_X1    g02906(.A1(new_n3563_), .A2(new_n3573_), .A3(new_n3578_), .ZN(new_n3911_));
  NAND4_X1   g02907(.A1(new_n3910_), .A2(new_n3538_), .A3(new_n3549_), .A4(new_n3552_), .ZN(new_n3912_));
  NAND4_X1   g02908(.A1(new_n3584_), .A2(new_n3899_), .A3(new_n3912_), .A4(new_n3907_), .ZN(new_n3913_));
  NOR2_X1    g02909(.A1(new_n3913_), .A2(new_n3886_), .ZN(new_n3914_));
  AND2_X2    g02910(.A1(new_n3852_), .A2(new_n3855_), .Z(new_n3915_));
  NAND3_X1   g02911(.A1(new_n3884_), .A2(new_n3877_), .A3(new_n3873_), .ZN(new_n3916_));
  NOR2_X1    g02912(.A1(new_n3916_), .A2(new_n3915_), .ZN(new_n3917_));
  OAI21_X1   g02913(.A1(new_n3917_), .A2(new_n3875_), .B(new_n3857_), .ZN(new_n3918_));
  NAND2_X1   g02914(.A1(new_n3527_), .A2(new_n3580_), .ZN(new_n3919_));
  INV_X1     g02915(.I(new_n3894_), .ZN(new_n3920_));
  XNOR2_X1   g02916(.A1(new_n3538_), .A2(new_n3549_), .ZN(new_n3921_));
  NOR2_X1    g02917(.A1(new_n3921_), .A2(new_n3890_), .ZN(new_n3922_));
  NOR4_X1    g02918(.A1(new_n3922_), .A2(new_n3920_), .A3(new_n3887_), .A4(new_n3895_), .ZN(new_n3923_));
  INV_X1     g02919(.I(new_n3906_), .ZN(new_n3924_));
  NOR2_X1    g02920(.A1(new_n3924_), .A2(new_n3904_), .ZN(new_n3925_));
  NOR2_X1    g02921(.A1(new_n3909_), .A2(new_n3908_), .ZN(new_n3926_));
  NOR4_X1    g02922(.A1(new_n3926_), .A2(new_n3892_), .A3(new_n3889_), .A4(new_n3890_), .ZN(new_n3927_));
  NOR4_X1    g02923(.A1(new_n3923_), .A2(new_n3919_), .A3(new_n3925_), .A4(new_n3927_), .ZN(new_n3928_));
  NOR2_X1    g02924(.A1(new_n3918_), .A2(new_n3928_), .ZN(new_n3929_));
  OAI21_X1   g02925(.A1(new_n3929_), .A2(new_n3914_), .B(new_n3881_), .ZN(new_n3930_));
  NAND2_X1   g02926(.A1(new_n3918_), .A2(new_n3928_), .ZN(new_n3931_));
  NAND2_X1   g02927(.A1(new_n3913_), .A2(new_n3886_), .ZN(new_n3932_));
  NAND3_X1   g02928(.A1(new_n3931_), .A2(new_n3880_), .A3(new_n3932_), .ZN(new_n3933_));
  AOI21_X1   g02929(.A1(new_n3930_), .A2(new_n3933_), .B(new_n3587_), .ZN(new_n3934_));
  NAND2_X1   g02930(.A1(new_n3848_), .A2(new_n3934_), .ZN(new_n3935_));
  NAND2_X1   g02931(.A1(new_n3934_), .A2(new_n3847_), .ZN(new_n3936_));
  AOI21_X1   g02932(.A1(new_n3935_), .A2(new_n3936_), .B(new_n3591_), .ZN(new_n3937_));
  INV_X1     g02933(.I(new_n3937_), .ZN(new_n3938_));
  NAND2_X1   g02934(.A1(new_n3938_), .A2(new_n3766_), .ZN(new_n3939_));
  INV_X1     g02935(.I(new_n3939_), .ZN(new_n3940_));
  NAND4_X1   g02936(.A1(new_n2961_), .A2(new_n2920_), .A3(new_n2931_), .A4(new_n2934_), .ZN(new_n3941_));
  INV_X1     g02937(.I(new_n2931_), .ZN(new_n3942_));
  INV_X1     g02938(.I(new_n2934_), .ZN(new_n3943_));
  NOR2_X1    g02939(.A1(new_n3943_), .A2(new_n2920_), .ZN(new_n3944_));
  INV_X1     g02940(.I(new_n2920_), .ZN(new_n3945_));
  NOR2_X1    g02941(.A1(new_n3945_), .A2(new_n2934_), .ZN(new_n3946_));
  OAI21_X1   g02942(.A1(new_n3946_), .A2(new_n3944_), .B(new_n3942_), .ZN(new_n3947_));
  NAND2_X1   g02943(.A1(new_n3945_), .A2(new_n2934_), .ZN(new_n3948_));
  NAND2_X1   g02944(.A1(new_n3943_), .A2(new_n2920_), .ZN(new_n3949_));
  NAND3_X1   g02945(.A1(new_n3948_), .A2(new_n2931_), .A3(new_n3949_), .ZN(new_n3950_));
  XOR2_X1    g02946(.A1(new_n2920_), .A2(new_n2931_), .Z(new_n3951_));
  NAND2_X1   g02947(.A1(new_n3951_), .A2(new_n2934_), .ZN(new_n3952_));
  NAND3_X1   g02948(.A1(new_n3952_), .A2(new_n3947_), .A3(new_n3950_), .ZN(new_n3953_));
  NAND2_X1   g02949(.A1(new_n3947_), .A2(new_n3950_), .ZN(new_n3954_));
  NOR3_X1    g02950(.A1(new_n2945_), .A2(new_n2955_), .A3(new_n2960_), .ZN(new_n3955_));
  NOR2_X1    g02951(.A1(new_n2945_), .A2(new_n2955_), .ZN(new_n3956_));
  INV_X1     g02952(.I(new_n2945_), .ZN(new_n3957_));
  INV_X1     g02953(.I(new_n2955_), .ZN(new_n3958_));
  NOR2_X1    g02954(.A1(new_n3957_), .A2(new_n3958_), .ZN(new_n3959_));
  NOR2_X1    g02955(.A1(new_n3959_), .A2(new_n3956_), .ZN(new_n3960_));
  NOR3_X1    g02956(.A1(new_n3960_), .A2(new_n2935_), .A3(new_n3955_), .ZN(new_n3961_));
  NOR2_X1    g02957(.A1(new_n3957_), .A2(new_n2960_), .ZN(new_n3962_));
  INV_X1     g02958(.I(new_n2960_), .ZN(new_n3963_));
  NOR2_X1    g02959(.A1(new_n3963_), .A2(new_n2945_), .ZN(new_n3964_));
  OAI21_X1   g02960(.A1(new_n3962_), .A2(new_n3964_), .B(new_n2955_), .ZN(new_n3965_));
  NAND2_X1   g02961(.A1(new_n3963_), .A2(new_n2945_), .ZN(new_n3966_));
  NAND2_X1   g02962(.A1(new_n3957_), .A2(new_n2960_), .ZN(new_n3967_));
  NAND3_X1   g02963(.A1(new_n3967_), .A2(new_n3966_), .A3(new_n3958_), .ZN(new_n3968_));
  NAND2_X1   g02964(.A1(new_n3965_), .A2(new_n3968_), .ZN(new_n3969_));
  NAND4_X1   g02965(.A1(new_n3969_), .A2(new_n3961_), .A3(new_n3954_), .A4(new_n3952_), .ZN(new_n3970_));
  AOI21_X1   g02966(.A1(new_n3970_), .A2(new_n3953_), .B(new_n3941_), .ZN(new_n3971_));
  INV_X1     g02967(.I(new_n3971_), .ZN(new_n3972_));
  INV_X1     g02968(.I(new_n3969_), .ZN(new_n3973_));
  XOR2_X1    g02969(.A1(new_n3953_), .A2(new_n3941_), .Z(new_n3974_));
  NAND2_X1   g02970(.A1(new_n3974_), .A2(new_n3973_), .ZN(new_n3975_));
  NOR2_X1    g02971(.A1(new_n2997_), .A2(new_n3007_), .ZN(new_n3976_));
  INV_X1     g02972(.I(new_n2997_), .ZN(new_n3977_));
  OR2_X2     g02973(.A1(new_n3006_), .A2(new_n3003_), .Z(new_n3978_));
  NOR2_X1    g02974(.A1(new_n3977_), .A2(new_n3978_), .ZN(new_n3979_));
  NOR2_X1    g02975(.A1(new_n3979_), .A2(new_n3976_), .ZN(new_n3980_));
  NOR3_X1    g02976(.A1(new_n2997_), .A2(new_n3007_), .A3(new_n3012_), .ZN(new_n3981_));
  INV_X1     g02977(.I(new_n3981_), .ZN(new_n3982_));
  NOR3_X1    g02978(.A1(new_n3980_), .A2(new_n2987_), .A3(new_n3982_), .ZN(new_n3983_));
  INV_X1     g02979(.I(new_n3983_), .ZN(new_n3984_));
  INV_X1     g02980(.I(new_n2982_), .ZN(new_n3985_));
  XNOR2_X1   g02981(.A1(new_n2985_), .A2(new_n2972_), .ZN(new_n3986_));
  NAND2_X1   g02982(.A1(new_n3986_), .A2(new_n3985_), .ZN(new_n3987_));
  XOR2_X1    g02983(.A1(new_n2985_), .A2(new_n2972_), .Z(new_n3988_));
  NAND2_X1   g02984(.A1(new_n3988_), .A2(new_n2982_), .ZN(new_n3989_));
  XOR2_X1    g02985(.A1(new_n2972_), .A2(new_n2982_), .Z(new_n3990_));
  NAND2_X1   g02986(.A1(new_n3990_), .A2(new_n2986_), .ZN(new_n3991_));
  NAND3_X1   g02987(.A1(new_n3987_), .A2(new_n3989_), .A3(new_n3991_), .ZN(new_n3992_));
  XOR2_X1    g02988(.A1(new_n2997_), .A2(new_n3012_), .Z(new_n3993_));
  XOR2_X1    g02989(.A1(new_n3993_), .A2(new_n3978_), .Z(new_n3994_));
  NOR2_X1    g02990(.A1(new_n3980_), .A2(new_n3981_), .ZN(new_n3995_));
  NAND4_X1   g02991(.A1(new_n3995_), .A2(new_n2972_), .A3(new_n2982_), .A4(new_n2986_), .ZN(new_n3996_));
  NAND4_X1   g02992(.A1(new_n3994_), .A2(new_n3996_), .A3(new_n3992_), .A4(new_n3984_), .ZN(new_n3997_));
  NOR2_X1    g02993(.A1(new_n3997_), .A2(new_n3015_), .ZN(new_n3998_));
  NAND2_X1   g02994(.A1(new_n3975_), .A2(new_n3998_), .ZN(new_n3999_));
  NOR2_X1    g02995(.A1(new_n3988_), .A2(new_n2982_), .ZN(new_n4000_));
  NOR2_X1    g02996(.A1(new_n3986_), .A2(new_n3985_), .ZN(new_n4001_));
  XNOR2_X1   g02997(.A1(new_n2972_), .A2(new_n2982_), .ZN(new_n4002_));
  NOR2_X1    g02998(.A1(new_n4002_), .A2(new_n2985_), .ZN(new_n4003_));
  NOR3_X1    g02999(.A1(new_n4001_), .A2(new_n4000_), .A3(new_n4003_), .ZN(new_n4004_));
  XOR2_X1    g03000(.A1(new_n3993_), .A2(new_n3007_), .Z(new_n4005_));
  INV_X1     g03001(.I(new_n2972_), .ZN(new_n4006_));
  OAI21_X1   g03002(.A1(new_n3976_), .A2(new_n3979_), .B(new_n3982_), .ZN(new_n4007_));
  NOR4_X1    g03003(.A1(new_n4007_), .A2(new_n4006_), .A3(new_n3985_), .A4(new_n2985_), .ZN(new_n4008_));
  NOR4_X1    g03004(.A1(new_n4004_), .A2(new_n4005_), .A3(new_n4008_), .A4(new_n3983_), .ZN(new_n4009_));
  NAND2_X1   g03005(.A1(new_n4009_), .A2(new_n3016_), .ZN(new_n4010_));
  NAND3_X1   g03006(.A1(new_n4010_), .A2(new_n3973_), .A3(new_n3974_), .ZN(new_n4011_));
  AOI21_X1   g03007(.A1(new_n3999_), .A2(new_n4011_), .B(new_n3972_), .ZN(new_n4012_));
  INV_X1     g03008(.I(new_n4012_), .ZN(new_n4013_));
  INV_X1     g03009(.I(new_n3054_), .ZN(new_n4014_));
  NOR2_X1    g03010(.A1(new_n4014_), .A2(new_n3069_), .ZN(new_n4015_));
  INV_X1     g03011(.I(new_n3069_), .ZN(new_n4016_));
  NOR2_X1    g03012(.A1(new_n4016_), .A2(new_n3054_), .ZN(new_n4017_));
  OAI21_X1   g03013(.A1(new_n4015_), .A2(new_n4017_), .B(new_n3064_), .ZN(new_n4018_));
  INV_X1     g03014(.I(new_n3064_), .ZN(new_n4019_));
  NAND2_X1   g03015(.A1(new_n4016_), .A2(new_n3054_), .ZN(new_n4020_));
  NAND2_X1   g03016(.A1(new_n4014_), .A2(new_n3069_), .ZN(new_n4021_));
  NAND3_X1   g03017(.A1(new_n4021_), .A2(new_n4020_), .A3(new_n4019_), .ZN(new_n4022_));
  NAND2_X1   g03018(.A1(new_n4018_), .A2(new_n4022_), .ZN(new_n4023_));
  INV_X1     g03019(.I(new_n4023_), .ZN(new_n4024_));
  NOR4_X1    g03020(.A1(new_n3044_), .A2(new_n3054_), .A3(new_n3064_), .A4(new_n3069_), .ZN(new_n4025_));
  INV_X1     g03021(.I(new_n4025_), .ZN(new_n4026_));
  INV_X1     g03022(.I(new_n3040_), .ZN(new_n4027_));
  NAND2_X1   g03023(.A1(new_n3021_), .A2(\A[531] ), .ZN(new_n4028_));
  NAND2_X1   g03024(.A1(new_n3019_), .A2(\A[530] ), .ZN(new_n4029_));
  AOI21_X1   g03025(.A1(new_n4028_), .A2(new_n4029_), .B(new_n3024_), .ZN(new_n4030_));
  INV_X1     g03026(.I(new_n3025_), .ZN(new_n4031_));
  AOI21_X1   g03027(.A1(new_n4031_), .A2(new_n3026_), .B(\A[529] ), .ZN(new_n4032_));
  NOR2_X1    g03028(.A1(new_n4032_), .A2(new_n4030_), .ZN(new_n4033_));
  NAND2_X1   g03029(.A1(new_n4033_), .A2(new_n3043_), .ZN(new_n4034_));
  INV_X1     g03030(.I(new_n4034_), .ZN(new_n4035_));
  NOR2_X1    g03031(.A1(new_n4033_), .A2(new_n3043_), .ZN(new_n4036_));
  OAI21_X1   g03032(.A1(new_n4035_), .A2(new_n4036_), .B(new_n4027_), .ZN(new_n4037_));
  INV_X1     g03033(.I(new_n3043_), .ZN(new_n4038_));
  NAND2_X1   g03034(.A1(new_n4038_), .A2(new_n3029_), .ZN(new_n4039_));
  NAND3_X1   g03035(.A1(new_n4039_), .A2(new_n4034_), .A3(new_n3040_), .ZN(new_n4040_));
  NAND2_X1   g03036(.A1(new_n4037_), .A2(new_n4040_), .ZN(new_n4041_));
  XOR2_X1    g03037(.A1(new_n4033_), .A2(new_n3040_), .Z(new_n4042_));
  NOR2_X1    g03038(.A1(new_n4042_), .A2(new_n4038_), .ZN(new_n4043_));
  NOR2_X1    g03039(.A1(new_n4041_), .A2(new_n4043_), .ZN(new_n4044_));
  NAND2_X1   g03040(.A1(new_n4044_), .A2(new_n4026_), .ZN(new_n4045_));
  OR2_X2     g03041(.A1(new_n4042_), .A2(new_n4038_), .Z(new_n4046_));
  NAND3_X1   g03042(.A1(new_n4046_), .A2(new_n4037_), .A3(new_n4040_), .ZN(new_n4047_));
  NAND2_X1   g03043(.A1(new_n4047_), .A2(new_n4025_), .ZN(new_n4048_));
  NAND2_X1   g03044(.A1(new_n4048_), .A2(new_n4045_), .ZN(new_n4049_));
  NAND2_X1   g03045(.A1(new_n4049_), .A2(new_n4024_), .ZN(new_n4050_));
  NOR3_X1    g03046(.A1(new_n3054_), .A2(new_n3064_), .A3(new_n3069_), .ZN(new_n4051_));
  NOR2_X1    g03047(.A1(new_n3054_), .A2(new_n3064_), .ZN(new_n4052_));
  NAND2_X1   g03048(.A1(new_n3054_), .A2(new_n3064_), .ZN(new_n4053_));
  INV_X1     g03049(.I(new_n4053_), .ZN(new_n4054_));
  NOR2_X1    g03050(.A1(new_n4054_), .A2(new_n4052_), .ZN(new_n4055_));
  NOR3_X1    g03051(.A1(new_n4055_), .A2(new_n3044_), .A3(new_n4051_), .ZN(new_n4056_));
  NAND4_X1   g03052(.A1(new_n4046_), .A2(new_n4023_), .A3(new_n4056_), .A4(new_n4041_), .ZN(new_n4057_));
  AOI21_X1   g03053(.A1(new_n4057_), .A2(new_n4047_), .B(new_n4026_), .ZN(new_n4058_));
  NOR4_X1    g03054(.A1(new_n3098_), .A2(new_n3108_), .A3(new_n3118_), .A4(new_n3123_), .ZN(new_n4059_));
  INV_X1     g03055(.I(new_n4059_), .ZN(new_n4060_));
  INV_X1     g03056(.I(new_n3092_), .ZN(new_n4061_));
  OAI22_X1   g03057(.A1(new_n3078_), .A2(new_n3093_), .B1(new_n3095_), .B2(new_n3088_), .ZN(new_n4062_));
  XNOR2_X1   g03058(.A1(new_n4062_), .A2(new_n3081_), .ZN(new_n4063_));
  NAND2_X1   g03059(.A1(new_n4063_), .A2(new_n4061_), .ZN(new_n4064_));
  XOR2_X1    g03060(.A1(new_n4062_), .A2(new_n3081_), .Z(new_n4065_));
  NAND2_X1   g03061(.A1(new_n4065_), .A2(new_n3092_), .ZN(new_n4066_));
  XOR2_X1    g03062(.A1(new_n3081_), .A2(new_n3092_), .Z(new_n4067_));
  NAND2_X1   g03063(.A1(new_n4067_), .A2(new_n3097_), .ZN(new_n4068_));
  NAND4_X1   g03064(.A1(new_n4060_), .A2(new_n4064_), .A3(new_n4066_), .A4(new_n4068_), .ZN(new_n4069_));
  INV_X1     g03065(.I(new_n3118_), .ZN(new_n4070_));
  XOR2_X1    g03066(.A1(new_n3108_), .A2(new_n3123_), .Z(new_n4071_));
  XOR2_X1    g03067(.A1(new_n4071_), .A2(new_n4070_), .Z(new_n4072_));
  INV_X1     g03068(.I(new_n3081_), .ZN(new_n4073_));
  INV_X1     g03069(.I(new_n3123_), .ZN(new_n4074_));
  NAND2_X1   g03070(.A1(new_n4070_), .A2(new_n4074_), .ZN(new_n4075_));
  NOR2_X1    g03071(.A1(new_n3108_), .A2(new_n3118_), .ZN(new_n4076_));
  INV_X1     g03072(.I(new_n3108_), .ZN(new_n4077_));
  NOR2_X1    g03073(.A1(new_n4077_), .A2(new_n4070_), .ZN(new_n4078_));
  OAI22_X1   g03074(.A1(new_n4076_), .A2(new_n4078_), .B1(new_n4075_), .B2(new_n3108_), .ZN(new_n4079_));
  NOR4_X1    g03075(.A1(new_n4079_), .A2(new_n4073_), .A3(new_n4061_), .A4(new_n4062_), .ZN(new_n4080_));
  NOR2_X1    g03076(.A1(new_n4080_), .A2(new_n4059_), .ZN(new_n4081_));
  NAND4_X1   g03077(.A1(new_n3127_), .A2(new_n4081_), .A3(new_n4069_), .A4(new_n4072_), .ZN(new_n4082_));
  NOR2_X1    g03078(.A1(new_n4082_), .A2(new_n4058_), .ZN(new_n4083_));
  INV_X1     g03079(.I(new_n4052_), .ZN(new_n4084_));
  AOI21_X1   g03080(.A1(new_n4084_), .A2(new_n4053_), .B(new_n4051_), .ZN(new_n4085_));
  NAND4_X1   g03081(.A1(new_n4085_), .A2(new_n3029_), .A3(new_n3040_), .A4(new_n3043_), .ZN(new_n4086_));
  NOR2_X1    g03082(.A1(new_n4024_), .A2(new_n4086_), .ZN(new_n4087_));
  OAI21_X1   g03083(.A1(new_n4087_), .A2(new_n4044_), .B(new_n4025_), .ZN(new_n4088_));
  NAND3_X1   g03084(.A1(new_n4064_), .A2(new_n4066_), .A3(new_n4068_), .ZN(new_n4089_));
  NOR3_X1    g03085(.A1(new_n3108_), .A2(new_n3118_), .A3(new_n3123_), .ZN(new_n4090_));
  NOR2_X1    g03086(.A1(new_n4078_), .A2(new_n4076_), .ZN(new_n4091_));
  NOR2_X1    g03087(.A1(new_n4091_), .A2(new_n4090_), .ZN(new_n4092_));
  NAND4_X1   g03088(.A1(new_n4092_), .A2(new_n3081_), .A3(new_n3092_), .A4(new_n3097_), .ZN(new_n4093_));
  NAND4_X1   g03089(.A1(new_n4093_), .A2(new_n4072_), .A3(new_n4089_), .A4(new_n4060_), .ZN(new_n4094_));
  NOR2_X1    g03090(.A1(new_n4094_), .A2(new_n3126_), .ZN(new_n4095_));
  NOR2_X1    g03091(.A1(new_n4095_), .A2(new_n4088_), .ZN(new_n4096_));
  OAI21_X1   g03092(.A1(new_n4096_), .A2(new_n4083_), .B(new_n4050_), .ZN(new_n4097_));
  AOI21_X1   g03093(.A1(new_n4048_), .A2(new_n4045_), .B(new_n4023_), .ZN(new_n4098_));
  NOR2_X1    g03094(.A1(new_n4065_), .A2(new_n3092_), .ZN(new_n4099_));
  NOR2_X1    g03095(.A1(new_n4063_), .A2(new_n4061_), .ZN(new_n4100_));
  XNOR2_X1   g03096(.A1(new_n3081_), .A2(new_n3092_), .ZN(new_n4101_));
  NOR2_X1    g03097(.A1(new_n4101_), .A2(new_n4062_), .ZN(new_n4102_));
  NOR3_X1    g03098(.A1(new_n4100_), .A2(new_n4099_), .A3(new_n4102_), .ZN(new_n4103_));
  XOR2_X1    g03099(.A1(new_n4071_), .A2(new_n3118_), .Z(new_n4104_));
  NOR4_X1    g03100(.A1(new_n4103_), .A2(new_n4104_), .A3(new_n4080_), .A4(new_n4059_), .ZN(new_n4105_));
  NAND3_X1   g03101(.A1(new_n4088_), .A2(new_n4105_), .A3(new_n3127_), .ZN(new_n4106_));
  NAND2_X1   g03102(.A1(new_n4082_), .A2(new_n4058_), .ZN(new_n4107_));
  NAND3_X1   g03103(.A1(new_n4107_), .A2(new_n4106_), .A3(new_n4098_), .ZN(new_n4108_));
  AOI21_X1   g03104(.A1(new_n4097_), .A2(new_n4108_), .B(new_n3130_), .ZN(new_n4109_));
  NOR2_X1    g03105(.A1(new_n4013_), .A2(new_n4109_), .ZN(new_n4110_));
  INV_X1     g03106(.I(new_n4110_), .ZN(new_n4111_));
  NOR4_X1    g03107(.A1(new_n2823_), .A2(new_n2833_), .A3(new_n2843_), .A4(new_n2848_), .ZN(new_n4112_));
  INV_X1     g03108(.I(new_n4112_), .ZN(new_n4113_));
  INV_X1     g03109(.I(new_n2818_), .ZN(new_n4114_));
  XNOR2_X1   g03110(.A1(new_n2821_), .A2(new_n2808_), .ZN(new_n4115_));
  NAND2_X1   g03111(.A1(new_n4115_), .A2(new_n4114_), .ZN(new_n4116_));
  XOR2_X1    g03112(.A1(new_n2821_), .A2(new_n2808_), .Z(new_n4117_));
  NAND2_X1   g03113(.A1(new_n4117_), .A2(new_n2818_), .ZN(new_n4118_));
  XOR2_X1    g03114(.A1(new_n2808_), .A2(new_n2818_), .Z(new_n4119_));
  NAND2_X1   g03115(.A1(new_n4119_), .A2(new_n2822_), .ZN(new_n4120_));
  NAND3_X1   g03116(.A1(new_n4116_), .A2(new_n4118_), .A3(new_n4120_), .ZN(new_n4121_));
  NAND2_X1   g03117(.A1(new_n4116_), .A2(new_n4118_), .ZN(new_n4122_));
  NOR3_X1    g03118(.A1(new_n2833_), .A2(new_n2843_), .A3(new_n2848_), .ZN(new_n4123_));
  NOR2_X1    g03119(.A1(new_n2833_), .A2(new_n2843_), .ZN(new_n4124_));
  OR2_X2     g03120(.A1(new_n2832_), .A2(new_n2829_), .Z(new_n4125_));
  INV_X1     g03121(.I(new_n2843_), .ZN(new_n4126_));
  NOR2_X1    g03122(.A1(new_n4126_), .A2(new_n4125_), .ZN(new_n4127_));
  NOR2_X1    g03123(.A1(new_n4127_), .A2(new_n4124_), .ZN(new_n4128_));
  XNOR2_X1   g03124(.A1(new_n2808_), .A2(new_n2818_), .ZN(new_n4129_));
  NOR2_X1    g03125(.A1(new_n4129_), .A2(new_n2821_), .ZN(new_n4130_));
  NOR4_X1    g03126(.A1(new_n4130_), .A2(new_n2823_), .A3(new_n4123_), .A4(new_n4128_), .ZN(new_n4131_));
  XOR2_X1    g03127(.A1(new_n2833_), .A2(new_n2848_), .Z(new_n4132_));
  XOR2_X1    g03128(.A1(new_n4132_), .A2(new_n4126_), .Z(new_n4133_));
  NAND3_X1   g03129(.A1(new_n4131_), .A2(new_n4133_), .A3(new_n4122_), .ZN(new_n4134_));
  AOI21_X1   g03130(.A1(new_n4134_), .A2(new_n4121_), .B(new_n4113_), .ZN(new_n4135_));
  INV_X1     g03131(.I(new_n4135_), .ZN(new_n4136_));
  XOR2_X1    g03132(.A1(new_n4132_), .A2(new_n2843_), .Z(new_n4137_));
  XOR2_X1    g03133(.A1(new_n4121_), .A2(new_n4113_), .Z(new_n4138_));
  NAND2_X1   g03134(.A1(new_n4138_), .A2(new_n4137_), .ZN(new_n4139_));
  NAND2_X1   g03135(.A1(new_n2850_), .A2(new_n2902_), .ZN(new_n4140_));
  NOR4_X1    g03136(.A1(new_n2875_), .A2(new_n2885_), .A3(new_n2895_), .A4(new_n2900_), .ZN(new_n4141_));
  INV_X1     g03137(.I(new_n4141_), .ZN(new_n4142_));
  INV_X1     g03138(.I(new_n2870_), .ZN(new_n4143_));
  XNOR2_X1   g03139(.A1(new_n2873_), .A2(new_n2860_), .ZN(new_n4144_));
  NAND2_X1   g03140(.A1(new_n4144_), .A2(new_n4143_), .ZN(new_n4145_));
  XOR2_X1    g03141(.A1(new_n2873_), .A2(new_n2860_), .Z(new_n4146_));
  NAND2_X1   g03142(.A1(new_n4146_), .A2(new_n2870_), .ZN(new_n4147_));
  XOR2_X1    g03143(.A1(new_n2860_), .A2(new_n2870_), .Z(new_n4148_));
  NAND2_X1   g03144(.A1(new_n4148_), .A2(new_n2874_), .ZN(new_n4149_));
  NAND3_X1   g03145(.A1(new_n4145_), .A2(new_n4147_), .A3(new_n4149_), .ZN(new_n4150_));
  OR2_X2     g03146(.A1(new_n2894_), .A2(new_n2891_), .Z(new_n4151_));
  XOR2_X1    g03147(.A1(new_n2885_), .A2(new_n2900_), .Z(new_n4152_));
  XOR2_X1    g03148(.A1(new_n4152_), .A2(new_n4151_), .Z(new_n4153_));
  NAND3_X1   g03149(.A1(new_n4151_), .A2(new_n2897_), .A3(new_n2899_), .ZN(new_n4154_));
  NOR2_X1    g03150(.A1(new_n4154_), .A2(new_n2885_), .ZN(new_n4155_));
  NOR2_X1    g03151(.A1(new_n2885_), .A2(new_n2895_), .ZN(new_n4156_));
  NOR3_X1    g03152(.A1(new_n4151_), .A2(new_n2881_), .A3(new_n2884_), .ZN(new_n4157_));
  NOR2_X1    g03153(.A1(new_n4157_), .A2(new_n4156_), .ZN(new_n4158_));
  NOR2_X1    g03154(.A1(new_n4158_), .A2(new_n4155_), .ZN(new_n4159_));
  NAND4_X1   g03155(.A1(new_n4159_), .A2(new_n2860_), .A3(new_n2870_), .A4(new_n2874_), .ZN(new_n4160_));
  NAND4_X1   g03156(.A1(new_n4160_), .A2(new_n4153_), .A3(new_n4150_), .A4(new_n4142_), .ZN(new_n4161_));
  NOR2_X1    g03157(.A1(new_n4161_), .A2(new_n4140_), .ZN(new_n4162_));
  NAND2_X1   g03158(.A1(new_n4139_), .A2(new_n4162_), .ZN(new_n4163_));
  NOR2_X1    g03159(.A1(new_n4146_), .A2(new_n2870_), .ZN(new_n4164_));
  NOR2_X1    g03160(.A1(new_n4144_), .A2(new_n4143_), .ZN(new_n4165_));
  XNOR2_X1   g03161(.A1(new_n2860_), .A2(new_n2870_), .ZN(new_n4166_));
  NOR2_X1    g03162(.A1(new_n4166_), .A2(new_n2873_), .ZN(new_n4167_));
  NOR3_X1    g03163(.A1(new_n4165_), .A2(new_n4164_), .A3(new_n4167_), .ZN(new_n4168_));
  XOR2_X1    g03164(.A1(new_n4152_), .A2(new_n2895_), .Z(new_n4169_));
  INV_X1     g03165(.I(new_n2860_), .ZN(new_n4170_));
  OAI22_X1   g03166(.A1(new_n4156_), .A2(new_n4157_), .B1(new_n4154_), .B2(new_n2885_), .ZN(new_n4171_));
  NOR4_X1    g03167(.A1(new_n4171_), .A2(new_n4170_), .A3(new_n4143_), .A4(new_n2873_), .ZN(new_n4172_));
  NOR4_X1    g03168(.A1(new_n4168_), .A2(new_n4169_), .A3(new_n4141_), .A4(new_n4172_), .ZN(new_n4173_));
  NAND2_X1   g03169(.A1(new_n4173_), .A2(new_n2903_), .ZN(new_n4174_));
  NAND3_X1   g03170(.A1(new_n4174_), .A2(new_n4138_), .A3(new_n4137_), .ZN(new_n4175_));
  AOI21_X1   g03171(.A1(new_n4163_), .A2(new_n4175_), .B(new_n4136_), .ZN(new_n4176_));
  INV_X1     g03172(.I(new_n4176_), .ZN(new_n4177_));
  OR2_X2     g03173(.A1(new_n2787_), .A2(new_n2784_), .Z(new_n4178_));
  NAND3_X1   g03174(.A1(new_n2778_), .A2(new_n2790_), .A3(new_n2792_), .ZN(new_n4179_));
  INV_X1     g03175(.I(new_n2778_), .ZN(new_n4180_));
  NAND2_X1   g03176(.A1(new_n4180_), .A2(new_n2793_), .ZN(new_n4181_));
  AOI21_X1   g03177(.A1(new_n4181_), .A2(new_n4179_), .B(new_n4178_), .ZN(new_n4182_));
  INV_X1     g03178(.I(new_n4182_), .ZN(new_n4183_));
  NAND3_X1   g03179(.A1(new_n4181_), .A2(new_n4178_), .A3(new_n4179_), .ZN(new_n4184_));
  NAND2_X1   g03180(.A1(new_n4183_), .A2(new_n4184_), .ZN(new_n4185_));
  NOR4_X1    g03181(.A1(new_n2768_), .A2(new_n2778_), .A3(new_n2788_), .A4(new_n2793_), .ZN(new_n4186_));
  INV_X1     g03182(.I(new_n4186_), .ZN(new_n4187_));
  INV_X1     g03183(.I(new_n2764_), .ZN(new_n4188_));
  NAND2_X1   g03184(.A1(new_n2745_), .A2(\A[483] ), .ZN(new_n4189_));
  NAND2_X1   g03185(.A1(new_n2743_), .A2(\A[482] ), .ZN(new_n4190_));
  AOI21_X1   g03186(.A1(new_n4189_), .A2(new_n4190_), .B(new_n2748_), .ZN(new_n4191_));
  INV_X1     g03187(.I(new_n2749_), .ZN(new_n4192_));
  AOI21_X1   g03188(.A1(new_n4192_), .A2(new_n2750_), .B(\A[481] ), .ZN(new_n4193_));
  NOR2_X1    g03189(.A1(new_n4193_), .A2(new_n4191_), .ZN(new_n4194_));
  NAND2_X1   g03190(.A1(new_n4194_), .A2(new_n2767_), .ZN(new_n4195_));
  INV_X1     g03191(.I(new_n4195_), .ZN(new_n4196_));
  NOR2_X1    g03192(.A1(new_n4194_), .A2(new_n2767_), .ZN(new_n4197_));
  OAI21_X1   g03193(.A1(new_n4196_), .A2(new_n4197_), .B(new_n4188_), .ZN(new_n4198_));
  INV_X1     g03194(.I(new_n2767_), .ZN(new_n4199_));
  NAND2_X1   g03195(.A1(new_n4199_), .A2(new_n2753_), .ZN(new_n4200_));
  NAND3_X1   g03196(.A1(new_n4200_), .A2(new_n4195_), .A3(new_n2764_), .ZN(new_n4201_));
  NAND2_X1   g03197(.A1(new_n4198_), .A2(new_n4201_), .ZN(new_n4202_));
  XOR2_X1    g03198(.A1(new_n2753_), .A2(new_n2764_), .Z(new_n4203_));
  AOI21_X1   g03199(.A1(new_n2767_), .A2(new_n4203_), .B(new_n4202_), .ZN(new_n4204_));
  NAND2_X1   g03200(.A1(new_n4204_), .A2(new_n4187_), .ZN(new_n4205_));
  NAND2_X1   g03201(.A1(new_n4203_), .A2(new_n2767_), .ZN(new_n4206_));
  NAND3_X1   g03202(.A1(new_n4206_), .A2(new_n4198_), .A3(new_n4201_), .ZN(new_n4207_));
  NAND2_X1   g03203(.A1(new_n4207_), .A2(new_n4186_), .ZN(new_n4208_));
  AOI21_X1   g03204(.A1(new_n4205_), .A2(new_n4208_), .B(new_n4185_), .ZN(new_n4209_));
  INV_X1     g03205(.I(new_n4209_), .ZN(new_n4210_));
  NOR3_X1    g03206(.A1(new_n2778_), .A2(new_n2788_), .A3(new_n2793_), .ZN(new_n4211_));
  NOR2_X1    g03207(.A1(new_n2778_), .A2(new_n2788_), .ZN(new_n4212_));
  NOR2_X1    g03208(.A1(new_n4180_), .A2(new_n4178_), .ZN(new_n4213_));
  NOR2_X1    g03209(.A1(new_n4213_), .A2(new_n4212_), .ZN(new_n4214_));
  NOR3_X1    g03210(.A1(new_n4214_), .A2(new_n2768_), .A3(new_n4211_), .ZN(new_n4215_));
  NAND4_X1   g03211(.A1(new_n4185_), .A2(new_n4202_), .A3(new_n4206_), .A4(new_n4215_), .ZN(new_n4216_));
  AOI21_X1   g03212(.A1(new_n4216_), .A2(new_n4207_), .B(new_n4187_), .ZN(new_n4217_));
  NAND4_X1   g03213(.A1(new_n2741_), .A2(new_n2699_), .A3(new_n2709_), .A4(new_n2714_), .ZN(new_n4218_));
  INV_X1     g03214(.I(new_n4218_), .ZN(new_n4219_));
  OAI22_X1   g03215(.A1(new_n2696_), .A2(new_n2710_), .B1(new_n2712_), .B2(new_n2706_), .ZN(new_n4220_));
  XOR2_X1    g03216(.A1(new_n4220_), .A2(new_n2699_), .Z(new_n4221_));
  NOR2_X1    g03217(.A1(new_n4221_), .A2(new_n2709_), .ZN(new_n4222_));
  INV_X1     g03218(.I(new_n2709_), .ZN(new_n4223_));
  XNOR2_X1   g03219(.A1(new_n4220_), .A2(new_n2699_), .ZN(new_n4224_));
  NOR2_X1    g03220(.A1(new_n4224_), .A2(new_n4223_), .ZN(new_n4225_));
  XNOR2_X1   g03221(.A1(new_n2699_), .A2(new_n2709_), .ZN(new_n4226_));
  NOR2_X1    g03222(.A1(new_n4226_), .A2(new_n4220_), .ZN(new_n4227_));
  NOR3_X1    g03223(.A1(new_n4225_), .A2(new_n4222_), .A3(new_n4227_), .ZN(new_n4228_));
  XOR2_X1    g03224(.A1(new_n2725_), .A2(new_n2740_), .Z(new_n4229_));
  XOR2_X1    g03225(.A1(new_n4229_), .A2(new_n2735_), .Z(new_n4230_));
  INV_X1     g03226(.I(new_n2699_), .ZN(new_n4231_));
  NAND4_X1   g03227(.A1(new_n2739_), .A2(new_n2726_), .A3(new_n2727_), .A4(new_n2729_), .ZN(new_n4232_));
  NOR2_X1    g03228(.A1(new_n2725_), .A2(new_n2735_), .ZN(new_n4233_));
  OR2_X2     g03229(.A1(new_n2734_), .A2(new_n2731_), .Z(new_n4234_));
  NOR3_X1    g03230(.A1(new_n4234_), .A2(new_n2721_), .A3(new_n2724_), .ZN(new_n4235_));
  OAI22_X1   g03231(.A1(new_n4235_), .A2(new_n4233_), .B1(new_n2725_), .B2(new_n4232_), .ZN(new_n4236_));
  NOR4_X1    g03232(.A1(new_n4236_), .A2(new_n4231_), .A3(new_n4223_), .A4(new_n4220_), .ZN(new_n4237_));
  NOR4_X1    g03233(.A1(new_n4228_), .A2(new_n4230_), .A3(new_n4219_), .A4(new_n4237_), .ZN(new_n4238_));
  NAND2_X1   g03234(.A1(new_n4238_), .A2(new_n2797_), .ZN(new_n4239_));
  NOR2_X1    g03235(.A1(new_n4239_), .A2(new_n4217_), .ZN(new_n4240_));
  INV_X1     g03236(.I(new_n4184_), .ZN(new_n4241_));
  NOR2_X1    g03237(.A1(new_n4241_), .A2(new_n4182_), .ZN(new_n4242_));
  NAND3_X1   g03238(.A1(new_n4215_), .A2(new_n4202_), .A3(new_n4206_), .ZN(new_n4243_));
  NOR2_X1    g03239(.A1(new_n4243_), .A2(new_n4242_), .ZN(new_n4244_));
  OAI21_X1   g03240(.A1(new_n4244_), .A2(new_n4204_), .B(new_n4186_), .ZN(new_n4245_));
  NOR4_X1    g03241(.A1(new_n4225_), .A2(new_n4222_), .A3(new_n4227_), .A4(new_n4219_), .ZN(new_n4246_));
  NOR2_X1    g03242(.A1(new_n4232_), .A2(new_n2725_), .ZN(new_n4247_));
  NOR2_X1    g03243(.A1(new_n4235_), .A2(new_n4233_), .ZN(new_n4248_));
  NOR2_X1    g03244(.A1(new_n4248_), .A2(new_n4247_), .ZN(new_n4249_));
  NAND4_X1   g03245(.A1(new_n4249_), .A2(new_n2699_), .A3(new_n2709_), .A4(new_n2714_), .ZN(new_n4250_));
  NAND2_X1   g03246(.A1(new_n4250_), .A2(new_n4218_), .ZN(new_n4251_));
  NOR4_X1    g03247(.A1(new_n4251_), .A2(new_n2796_), .A3(new_n4246_), .A4(new_n4230_), .ZN(new_n4252_));
  NOR2_X1    g03248(.A1(new_n4252_), .A2(new_n4245_), .ZN(new_n4253_));
  OAI21_X1   g03249(.A1(new_n4240_), .A2(new_n4253_), .B(new_n4210_), .ZN(new_n4254_));
  NAND2_X1   g03250(.A1(new_n4252_), .A2(new_n4245_), .ZN(new_n4255_));
  NAND2_X1   g03251(.A1(new_n4239_), .A2(new_n4217_), .ZN(new_n4256_));
  NAND3_X1   g03252(.A1(new_n4256_), .A2(new_n4255_), .A3(new_n4209_), .ZN(new_n4257_));
  AOI21_X1   g03253(.A1(new_n4254_), .A2(new_n4257_), .B(new_n2906_), .ZN(new_n4258_));
  NAND2_X1   g03254(.A1(new_n4177_), .A2(new_n4258_), .ZN(new_n4259_));
  NAND2_X1   g03255(.A1(new_n4258_), .A2(new_n4176_), .ZN(new_n4260_));
  AOI21_X1   g03256(.A1(new_n4259_), .A2(new_n4260_), .B(new_n3134_), .ZN(new_n4261_));
  NAND2_X1   g03257(.A1(new_n4261_), .A2(new_n4111_), .ZN(new_n4262_));
  NAND2_X1   g03258(.A1(new_n4261_), .A2(new_n4110_), .ZN(new_n4263_));
  NAND2_X1   g03259(.A1(new_n4262_), .A2(new_n4263_), .ZN(new_n4264_));
  NAND2_X1   g03260(.A1(new_n4264_), .A2(new_n3595_), .ZN(new_n4265_));
  NOR2_X1    g03261(.A1(new_n4265_), .A2(new_n3940_), .ZN(new_n4266_));
  NOR2_X1    g03262(.A1(new_n4265_), .A2(new_n3939_), .ZN(new_n4267_));
  NOR2_X1    g03263(.A1(new_n4266_), .A2(new_n4267_), .ZN(new_n4268_));
  INV_X1     g03264(.I(new_n4268_), .ZN(new_n4269_));
  OAI21_X1   g03265(.A1(new_n4269_), .A2(new_n3599_), .B(new_n2686_), .ZN(new_n4270_));
  OAI21_X1   g03266(.A1(new_n3595_), .A2(new_n4264_), .B(new_n3940_), .ZN(new_n4271_));
  NAND2_X1   g03267(.A1(new_n4271_), .A2(new_n4265_), .ZN(new_n4272_));
  INV_X1     g03268(.I(new_n4272_), .ZN(new_n4273_));
  NAND3_X1   g03269(.A1(new_n4259_), .A2(new_n4260_), .A3(new_n3134_), .ZN(new_n4274_));
  AOI21_X1   g03270(.A1(new_n4110_), .A2(new_n4274_), .B(new_n4261_), .ZN(new_n4275_));
  INV_X1     g03271(.I(new_n4275_), .ZN(new_n4276_));
  AOI21_X1   g03272(.A1(new_n4256_), .A2(new_n4255_), .B(new_n4209_), .ZN(new_n4277_));
  NOR3_X1    g03273(.A1(new_n4240_), .A2(new_n4253_), .A3(new_n4210_), .ZN(new_n4278_));
  OAI21_X1   g03274(.A1(new_n4277_), .A2(new_n4278_), .B(new_n2907_), .ZN(new_n4279_));
  NOR3_X1    g03275(.A1(new_n4277_), .A2(new_n4278_), .A3(new_n2907_), .ZN(new_n4280_));
  OAI21_X1   g03276(.A1(new_n4177_), .A2(new_n4280_), .B(new_n4279_), .ZN(new_n4281_));
  NOR2_X1    g03277(.A1(new_n4238_), .A2(new_n2797_), .ZN(new_n4282_));
  NAND4_X1   g03278(.A1(new_n4244_), .A2(new_n4242_), .A3(new_n4186_), .A4(new_n4207_), .ZN(new_n4283_));
  OAI21_X1   g03279(.A1(new_n4282_), .A2(new_n4283_), .B(new_n4239_), .ZN(new_n4284_));
  NAND2_X1   g03280(.A1(new_n2711_), .A2(new_n2713_), .ZN(new_n4285_));
  NAND3_X1   g03281(.A1(new_n4285_), .A2(new_n2699_), .A3(new_n2709_), .ZN(new_n4286_));
  NAND2_X1   g03282(.A1(new_n4286_), .A2(new_n4220_), .ZN(new_n4287_));
  OAI21_X1   g03283(.A1(new_n2737_), .A2(new_n2739_), .B(new_n4233_), .ZN(new_n4288_));
  NAND2_X1   g03284(.A1(new_n4288_), .A2(new_n2740_), .ZN(new_n4289_));
  XNOR2_X1   g03285(.A1(new_n4289_), .A2(new_n4287_), .ZN(new_n4290_));
  XOR2_X1    g03286(.A1(new_n4229_), .A2(new_n4234_), .Z(new_n4291_));
  OAI21_X1   g03287(.A1(new_n4228_), .A2(new_n4219_), .B(new_n4291_), .ZN(new_n4292_));
  AOI21_X1   g03288(.A1(new_n4292_), .A2(new_n4250_), .B(new_n4290_), .ZN(new_n4293_));
  INV_X1     g03289(.I(new_n4243_), .ZN(new_n4294_));
  NAND2_X1   g03290(.A1(new_n2765_), .A2(new_n2766_), .ZN(new_n4295_));
  NAND3_X1   g03291(.A1(new_n2753_), .A2(new_n2764_), .A3(new_n4295_), .ZN(new_n4296_));
  NAND2_X1   g03292(.A1(new_n4296_), .A2(new_n4199_), .ZN(new_n4297_));
  OAI21_X1   g03293(.A1(new_n2790_), .A2(new_n2792_), .B(new_n4212_), .ZN(new_n4298_));
  NAND2_X1   g03294(.A1(new_n4298_), .A2(new_n2793_), .ZN(new_n4299_));
  XOR2_X1    g03295(.A1(new_n4299_), .A2(new_n4297_), .Z(new_n4300_));
  AOI21_X1   g03296(.A1(new_n4187_), .A2(new_n4207_), .B(new_n4242_), .ZN(new_n4301_));
  OAI21_X1   g03297(.A1(new_n4301_), .A2(new_n4294_), .B(new_n4300_), .ZN(new_n4302_));
  NAND2_X1   g03298(.A1(new_n4293_), .A2(new_n4302_), .ZN(new_n4303_));
  INV_X1     g03299(.I(new_n4303_), .ZN(new_n4304_));
  NOR2_X1    g03300(.A1(new_n4293_), .A2(new_n4302_), .ZN(new_n4305_));
  OAI21_X1   g03301(.A1(new_n4304_), .A2(new_n4305_), .B(new_n4284_), .ZN(new_n4306_));
  NAND2_X1   g03302(.A1(new_n4224_), .A2(new_n4223_), .ZN(new_n4307_));
  NAND2_X1   g03303(.A1(new_n4221_), .A2(new_n2709_), .ZN(new_n4308_));
  XOR2_X1    g03304(.A1(new_n2699_), .A2(new_n2709_), .Z(new_n4309_));
  NAND2_X1   g03305(.A1(new_n4309_), .A2(new_n2714_), .ZN(new_n4310_));
  NAND4_X1   g03306(.A1(new_n4307_), .A2(new_n4308_), .A3(new_n4310_), .A4(new_n4218_), .ZN(new_n4311_));
  NOR2_X1    g03307(.A1(new_n4237_), .A2(new_n4219_), .ZN(new_n4312_));
  NAND3_X1   g03308(.A1(new_n4312_), .A2(new_n4311_), .A3(new_n4291_), .ZN(new_n4313_));
  NAND2_X1   g03309(.A1(new_n4313_), .A2(new_n2796_), .ZN(new_n4314_));
  NOR4_X1    g03310(.A1(new_n4216_), .A2(new_n4185_), .A3(new_n4187_), .A4(new_n4204_), .ZN(new_n4315_));
  AOI21_X1   g03311(.A1(new_n4314_), .A2(new_n4315_), .B(new_n4252_), .ZN(new_n4316_));
  XNOR2_X1   g03312(.A1(new_n4299_), .A2(new_n4297_), .ZN(new_n4317_));
  OAI21_X1   g03313(.A1(new_n4204_), .A2(new_n4186_), .B(new_n4185_), .ZN(new_n4318_));
  AOI21_X1   g03314(.A1(new_n4318_), .A2(new_n4243_), .B(new_n4317_), .ZN(new_n4319_));
  NOR2_X1    g03315(.A1(new_n4319_), .A2(new_n4293_), .ZN(new_n4320_));
  XOR2_X1    g03316(.A1(new_n4289_), .A2(new_n4287_), .Z(new_n4321_));
  NAND3_X1   g03317(.A1(new_n4307_), .A2(new_n4308_), .A3(new_n4310_), .ZN(new_n4322_));
  AOI21_X1   g03318(.A1(new_n4322_), .A2(new_n4218_), .B(new_n4230_), .ZN(new_n4323_));
  OAI21_X1   g03319(.A1(new_n4323_), .A2(new_n4237_), .B(new_n4321_), .ZN(new_n4324_));
  NOR2_X1    g03320(.A1(new_n4324_), .A2(new_n4302_), .ZN(new_n4325_));
  OAI21_X1   g03321(.A1(new_n4320_), .A2(new_n4325_), .B(new_n4316_), .ZN(new_n4326_));
  NAND2_X1   g03322(.A1(new_n4306_), .A2(new_n4326_), .ZN(new_n4327_));
  NAND2_X1   g03323(.A1(new_n4161_), .A2(new_n4140_), .ZN(new_n4328_));
  NOR2_X1    g03324(.A1(new_n4117_), .A2(new_n2818_), .ZN(new_n4329_));
  NOR2_X1    g03325(.A1(new_n4115_), .A2(new_n4114_), .ZN(new_n4330_));
  NOR3_X1    g03326(.A1(new_n4330_), .A2(new_n4329_), .A3(new_n4130_), .ZN(new_n4331_));
  NOR4_X1    g03327(.A1(new_n4134_), .A2(new_n4113_), .A3(new_n4331_), .A4(new_n4133_), .ZN(new_n4332_));
  AOI21_X1   g03328(.A1(new_n4332_), .A2(new_n4328_), .B(new_n4162_), .ZN(new_n4333_));
  NAND2_X1   g03329(.A1(new_n2860_), .A2(new_n2870_), .ZN(new_n4334_));
  NOR4_X1    g03330(.A1(new_n2871_), .A2(new_n2872_), .A3(new_n2857_), .A4(new_n2867_), .ZN(new_n4335_));
  OAI21_X1   g03331(.A1(new_n4334_), .A2(new_n4335_), .B(new_n2873_), .ZN(new_n4336_));
  OAI21_X1   g03332(.A1(new_n2897_), .A2(new_n2899_), .B(new_n4156_), .ZN(new_n4337_));
  NAND2_X1   g03333(.A1(new_n4337_), .A2(new_n2900_), .ZN(new_n4338_));
  XNOR2_X1   g03334(.A1(new_n4338_), .A2(new_n4336_), .ZN(new_n4339_));
  OAI21_X1   g03335(.A1(new_n4168_), .A2(new_n4141_), .B(new_n4153_), .ZN(new_n4340_));
  AOI21_X1   g03336(.A1(new_n4340_), .A2(new_n4160_), .B(new_n4339_), .ZN(new_n4341_));
  NOR2_X1    g03337(.A1(new_n4128_), .A2(new_n4123_), .ZN(new_n4342_));
  NAND4_X1   g03338(.A1(new_n4342_), .A2(new_n2808_), .A3(new_n2818_), .A4(new_n2822_), .ZN(new_n4343_));
  INV_X1     g03339(.I(new_n4343_), .ZN(new_n4344_));
  NAND2_X1   g03340(.A1(new_n2808_), .A2(new_n2818_), .ZN(new_n4345_));
  NOR4_X1    g03341(.A1(new_n2819_), .A2(new_n2820_), .A3(new_n2805_), .A4(new_n2816_), .ZN(new_n4346_));
  OAI21_X1   g03342(.A1(new_n4345_), .A2(new_n4346_), .B(new_n2821_), .ZN(new_n4347_));
  OAI21_X1   g03343(.A1(new_n2845_), .A2(new_n2847_), .B(new_n4124_), .ZN(new_n4348_));
  NAND2_X1   g03344(.A1(new_n4348_), .A2(new_n2848_), .ZN(new_n4349_));
  XOR2_X1    g03345(.A1(new_n4349_), .A2(new_n4347_), .Z(new_n4350_));
  AOI21_X1   g03346(.A1(new_n4113_), .A2(new_n4121_), .B(new_n4137_), .ZN(new_n4351_));
  OAI21_X1   g03347(.A1(new_n4351_), .A2(new_n4344_), .B(new_n4350_), .ZN(new_n4352_));
  NAND2_X1   g03348(.A1(new_n4352_), .A2(new_n4341_), .ZN(new_n4353_));
  XOR2_X1    g03349(.A1(new_n4338_), .A2(new_n4336_), .Z(new_n4354_));
  AOI21_X1   g03350(.A1(new_n4142_), .A2(new_n4150_), .B(new_n4169_), .ZN(new_n4355_));
  OAI21_X1   g03351(.A1(new_n4355_), .A2(new_n4172_), .B(new_n4354_), .ZN(new_n4356_));
  XNOR2_X1   g03352(.A1(new_n4349_), .A2(new_n4347_), .ZN(new_n4357_));
  OAI21_X1   g03353(.A1(new_n4331_), .A2(new_n4112_), .B(new_n4133_), .ZN(new_n4358_));
  AOI21_X1   g03354(.A1(new_n4358_), .A2(new_n4343_), .B(new_n4357_), .ZN(new_n4359_));
  NAND2_X1   g03355(.A1(new_n4359_), .A2(new_n4356_), .ZN(new_n4360_));
  AOI21_X1   g03356(.A1(new_n4353_), .A2(new_n4360_), .B(new_n4333_), .ZN(new_n4361_));
  NOR2_X1    g03357(.A1(new_n4173_), .A2(new_n2903_), .ZN(new_n4362_));
  NOR2_X1    g03358(.A1(new_n4343_), .A2(new_n4137_), .ZN(new_n4363_));
  NAND4_X1   g03359(.A1(new_n4363_), .A2(new_n4112_), .A3(new_n4121_), .A4(new_n4137_), .ZN(new_n4364_));
  OAI21_X1   g03360(.A1(new_n4362_), .A2(new_n4364_), .B(new_n4174_), .ZN(new_n4365_));
  NAND2_X1   g03361(.A1(new_n4356_), .A2(new_n4352_), .ZN(new_n4366_));
  NAND2_X1   g03362(.A1(new_n4359_), .A2(new_n4341_), .ZN(new_n4367_));
  AOI21_X1   g03363(.A1(new_n4366_), .A2(new_n4367_), .B(new_n4365_), .ZN(new_n4368_));
  NOR2_X1    g03364(.A1(new_n4368_), .A2(new_n4361_), .ZN(new_n4369_));
  NOR2_X1    g03365(.A1(new_n4369_), .A2(new_n4327_), .ZN(new_n4370_));
  NAND2_X1   g03366(.A1(new_n4324_), .A2(new_n4319_), .ZN(new_n4371_));
  AOI21_X1   g03367(.A1(new_n4303_), .A2(new_n4371_), .B(new_n4316_), .ZN(new_n4372_));
  NAND2_X1   g03368(.A1(new_n4324_), .A2(new_n4302_), .ZN(new_n4373_));
  NAND2_X1   g03369(.A1(new_n4319_), .A2(new_n4293_), .ZN(new_n4374_));
  AOI21_X1   g03370(.A1(new_n4373_), .A2(new_n4374_), .B(new_n4284_), .ZN(new_n4375_));
  NOR2_X1    g03371(.A1(new_n4375_), .A2(new_n4372_), .ZN(new_n4376_));
  NOR2_X1    g03372(.A1(new_n4359_), .A2(new_n4356_), .ZN(new_n4377_));
  NOR2_X1    g03373(.A1(new_n4352_), .A2(new_n4341_), .ZN(new_n4378_));
  OAI21_X1   g03374(.A1(new_n4377_), .A2(new_n4378_), .B(new_n4365_), .ZN(new_n4379_));
  NOR2_X1    g03375(.A1(new_n4359_), .A2(new_n4341_), .ZN(new_n4380_));
  NOR2_X1    g03376(.A1(new_n4356_), .A2(new_n4352_), .ZN(new_n4381_));
  OAI21_X1   g03377(.A1(new_n4381_), .A2(new_n4380_), .B(new_n4333_), .ZN(new_n4382_));
  NAND2_X1   g03378(.A1(new_n4379_), .A2(new_n4382_), .ZN(new_n4383_));
  NOR2_X1    g03379(.A1(new_n4383_), .A2(new_n4376_), .ZN(new_n4384_));
  OAI21_X1   g03380(.A1(new_n4384_), .A2(new_n4370_), .B(new_n4281_), .ZN(new_n4385_));
  NAND3_X1   g03381(.A1(new_n4254_), .A2(new_n4257_), .A3(new_n2906_), .ZN(new_n4386_));
  AOI21_X1   g03382(.A1(new_n4176_), .A2(new_n4386_), .B(new_n4258_), .ZN(new_n4387_));
  NOR2_X1    g03383(.A1(new_n4369_), .A2(new_n4376_), .ZN(new_n4388_));
  NOR2_X1    g03384(.A1(new_n4383_), .A2(new_n4327_), .ZN(new_n4389_));
  OAI21_X1   g03385(.A1(new_n4389_), .A2(new_n4388_), .B(new_n4387_), .ZN(new_n4390_));
  NAND2_X1   g03386(.A1(new_n4385_), .A2(new_n4390_), .ZN(new_n4391_));
  NAND3_X1   g03387(.A1(new_n4097_), .A2(new_n4108_), .A3(new_n3130_), .ZN(new_n4392_));
  AOI21_X1   g03388(.A1(new_n4012_), .A2(new_n4392_), .B(new_n4109_), .ZN(new_n4393_));
  NAND2_X1   g03389(.A1(new_n4094_), .A2(new_n3126_), .ZN(new_n4394_));
  NOR4_X1    g03390(.A1(new_n4057_), .A2(new_n4023_), .A3(new_n4026_), .A4(new_n4044_), .ZN(new_n4395_));
  AOI21_X1   g03391(.A1(new_n4394_), .A2(new_n4395_), .B(new_n4095_), .ZN(new_n4396_));
  NAND2_X1   g03392(.A1(new_n3094_), .A2(new_n3096_), .ZN(new_n4397_));
  NAND3_X1   g03393(.A1(new_n4397_), .A2(new_n3081_), .A3(new_n3092_), .ZN(new_n4398_));
  NAND2_X1   g03394(.A1(new_n4398_), .A2(new_n4062_), .ZN(new_n4399_));
  OAI21_X1   g03395(.A1(new_n3120_), .A2(new_n3122_), .B(new_n4076_), .ZN(new_n4400_));
  NAND2_X1   g03396(.A1(new_n4400_), .A2(new_n3123_), .ZN(new_n4401_));
  XNOR2_X1   g03397(.A1(new_n4401_), .A2(new_n4399_), .ZN(new_n4402_));
  OAI21_X1   g03398(.A1(new_n4103_), .A2(new_n4059_), .B(new_n4072_), .ZN(new_n4403_));
  AOI21_X1   g03399(.A1(new_n4403_), .A2(new_n4093_), .B(new_n4402_), .ZN(new_n4404_));
  NAND2_X1   g03400(.A1(new_n3041_), .A2(new_n3042_), .ZN(new_n4405_));
  NAND3_X1   g03401(.A1(new_n3029_), .A2(new_n3040_), .A3(new_n4405_), .ZN(new_n4406_));
  NAND2_X1   g03402(.A1(new_n4406_), .A2(new_n4038_), .ZN(new_n4407_));
  NOR2_X1    g03403(.A1(new_n3066_), .A2(new_n3068_), .ZN(new_n4408_));
  OAI21_X1   g03404(.A1(new_n4084_), .A2(new_n4408_), .B(new_n3069_), .ZN(new_n4409_));
  XNOR2_X1   g03405(.A1(new_n4409_), .A2(new_n4407_), .ZN(new_n4410_));
  OAI21_X1   g03406(.A1(new_n4044_), .A2(new_n4025_), .B(new_n4023_), .ZN(new_n4411_));
  AOI21_X1   g03407(.A1(new_n4411_), .A2(new_n4086_), .B(new_n4410_), .ZN(new_n4412_));
  INV_X1     g03408(.I(new_n4412_), .ZN(new_n4413_));
  NAND2_X1   g03409(.A1(new_n4413_), .A2(new_n4404_), .ZN(new_n4414_));
  XOR2_X1    g03410(.A1(new_n4401_), .A2(new_n4399_), .Z(new_n4415_));
  AOI21_X1   g03411(.A1(new_n4089_), .A2(new_n4060_), .B(new_n4104_), .ZN(new_n4416_));
  OAI21_X1   g03412(.A1(new_n4416_), .A2(new_n4080_), .B(new_n4415_), .ZN(new_n4417_));
  NAND2_X1   g03413(.A1(new_n4417_), .A2(new_n4412_), .ZN(new_n4418_));
  AOI21_X1   g03414(.A1(new_n4414_), .A2(new_n4418_), .B(new_n4396_), .ZN(new_n4419_));
  NOR2_X1    g03415(.A1(new_n4105_), .A2(new_n3127_), .ZN(new_n4420_));
  NAND4_X1   g03416(.A1(new_n4087_), .A2(new_n4047_), .A3(new_n4024_), .A4(new_n4025_), .ZN(new_n4421_));
  OAI21_X1   g03417(.A1(new_n4420_), .A2(new_n4421_), .B(new_n4082_), .ZN(new_n4422_));
  NAND2_X1   g03418(.A1(new_n4413_), .A2(new_n4417_), .ZN(new_n4423_));
  NAND2_X1   g03419(.A1(new_n4404_), .A2(new_n4412_), .ZN(new_n4424_));
  AOI21_X1   g03420(.A1(new_n4424_), .A2(new_n4423_), .B(new_n4422_), .ZN(new_n4425_));
  NOR2_X1    g03421(.A1(new_n4419_), .A2(new_n4425_), .ZN(new_n4426_));
  NOR2_X1    g03422(.A1(new_n4009_), .A2(new_n3016_), .ZN(new_n4427_));
  INV_X1     g03423(.I(new_n3953_), .ZN(new_n4428_));
  NOR4_X1    g03424(.A1(new_n3970_), .A2(new_n4428_), .A3(new_n3941_), .A4(new_n3969_), .ZN(new_n4429_));
  INV_X1     g03425(.I(new_n4429_), .ZN(new_n4430_));
  OAI21_X1   g03426(.A1(new_n4430_), .A2(new_n4427_), .B(new_n4010_), .ZN(new_n4431_));
  NAND2_X1   g03427(.A1(new_n2972_), .A2(new_n2982_), .ZN(new_n4432_));
  NOR4_X1    g03428(.A1(new_n2983_), .A2(new_n2984_), .A3(new_n2970_), .A4(new_n2980_), .ZN(new_n4433_));
  OAI21_X1   g03429(.A1(new_n4432_), .A2(new_n4433_), .B(new_n2985_), .ZN(new_n4434_));
  OAI21_X1   g03430(.A1(new_n3009_), .A2(new_n3011_), .B(new_n3976_), .ZN(new_n4435_));
  NAND2_X1   g03431(.A1(new_n4435_), .A2(new_n3012_), .ZN(new_n4436_));
  XNOR2_X1   g03432(.A1(new_n4436_), .A2(new_n4434_), .ZN(new_n4437_));
  OAI21_X1   g03433(.A1(new_n4004_), .A2(new_n3983_), .B(new_n3994_), .ZN(new_n4438_));
  AOI21_X1   g03434(.A1(new_n4438_), .A2(new_n3996_), .B(new_n4437_), .ZN(new_n4439_));
  NAND3_X1   g03435(.A1(new_n3961_), .A2(new_n3954_), .A3(new_n3952_), .ZN(new_n4440_));
  INV_X1     g03436(.I(new_n4440_), .ZN(new_n4441_));
  NAND2_X1   g03437(.A1(new_n2932_), .A2(new_n2933_), .ZN(new_n4442_));
  NAND3_X1   g03438(.A1(new_n2920_), .A2(new_n2931_), .A3(new_n4442_), .ZN(new_n4443_));
  NAND2_X1   g03439(.A1(new_n4443_), .A2(new_n3943_), .ZN(new_n4444_));
  OAI21_X1   g03440(.A1(new_n2957_), .A2(new_n2959_), .B(new_n3956_), .ZN(new_n4445_));
  NAND2_X1   g03441(.A1(new_n4445_), .A2(new_n2960_), .ZN(new_n4446_));
  XOR2_X1    g03442(.A1(new_n4446_), .A2(new_n4444_), .Z(new_n4447_));
  AOI21_X1   g03443(.A1(new_n3941_), .A2(new_n3953_), .B(new_n3973_), .ZN(new_n4448_));
  OAI21_X1   g03444(.A1(new_n4448_), .A2(new_n4441_), .B(new_n4447_), .ZN(new_n4449_));
  NAND2_X1   g03445(.A1(new_n4439_), .A2(new_n4449_), .ZN(new_n4450_));
  INV_X1     g03446(.I(new_n4450_), .ZN(new_n4451_));
  NOR2_X1    g03447(.A1(new_n4439_), .A2(new_n4449_), .ZN(new_n4452_));
  OAI21_X1   g03448(.A1(new_n4451_), .A2(new_n4452_), .B(new_n4431_), .ZN(new_n4453_));
  NAND2_X1   g03449(.A1(new_n3997_), .A2(new_n3015_), .ZN(new_n4454_));
  AOI21_X1   g03450(.A1(new_n4454_), .A2(new_n4429_), .B(new_n3998_), .ZN(new_n4455_));
  INV_X1     g03451(.I(new_n4444_), .ZN(new_n4456_));
  XOR2_X1    g03452(.A1(new_n4446_), .A2(new_n4456_), .Z(new_n4457_));
  NAND2_X1   g03453(.A1(new_n3953_), .A2(new_n3941_), .ZN(new_n4458_));
  NAND2_X1   g03454(.A1(new_n4458_), .A2(new_n3969_), .ZN(new_n4459_));
  AOI21_X1   g03455(.A1(new_n4459_), .A2(new_n4440_), .B(new_n4457_), .ZN(new_n4460_));
  NOR2_X1    g03456(.A1(new_n4460_), .A2(new_n4439_), .ZN(new_n4461_));
  XOR2_X1    g03457(.A1(new_n4436_), .A2(new_n4434_), .Z(new_n4462_));
  AOI21_X1   g03458(.A1(new_n3992_), .A2(new_n3984_), .B(new_n4005_), .ZN(new_n4463_));
  OAI21_X1   g03459(.A1(new_n4463_), .A2(new_n4008_), .B(new_n4462_), .ZN(new_n4464_));
  NOR2_X1    g03460(.A1(new_n4464_), .A2(new_n4449_), .ZN(new_n4465_));
  OAI21_X1   g03461(.A1(new_n4461_), .A2(new_n4465_), .B(new_n4455_), .ZN(new_n4466_));
  NAND2_X1   g03462(.A1(new_n4453_), .A2(new_n4466_), .ZN(new_n4467_));
  NAND2_X1   g03463(.A1(new_n4467_), .A2(new_n4426_), .ZN(new_n4468_));
  NAND2_X1   g03464(.A1(new_n4414_), .A2(new_n4418_), .ZN(new_n4469_));
  NAND2_X1   g03465(.A1(new_n4423_), .A2(new_n4424_), .ZN(new_n4470_));
  MUX2_X1    g03466(.I0(new_n4470_), .I1(new_n4469_), .S(new_n4422_), .Z(new_n4471_));
  NAND2_X1   g03467(.A1(new_n4460_), .A2(new_n4464_), .ZN(new_n4472_));
  AOI21_X1   g03468(.A1(new_n4450_), .A2(new_n4472_), .B(new_n4455_), .ZN(new_n4473_));
  NAND2_X1   g03469(.A1(new_n4464_), .A2(new_n4449_), .ZN(new_n4474_));
  NAND2_X1   g03470(.A1(new_n4460_), .A2(new_n4439_), .ZN(new_n4475_));
  AOI21_X1   g03471(.A1(new_n4474_), .A2(new_n4475_), .B(new_n4431_), .ZN(new_n4476_));
  NOR2_X1    g03472(.A1(new_n4473_), .A2(new_n4476_), .ZN(new_n4477_));
  NAND2_X1   g03473(.A1(new_n4471_), .A2(new_n4477_), .ZN(new_n4478_));
  AOI21_X1   g03474(.A1(new_n4478_), .A2(new_n4468_), .B(new_n4393_), .ZN(new_n4479_));
  AOI21_X1   g03475(.A1(new_n4107_), .A2(new_n4106_), .B(new_n4098_), .ZN(new_n4480_));
  NOR3_X1    g03476(.A1(new_n4096_), .A2(new_n4083_), .A3(new_n4050_), .ZN(new_n4481_));
  OAI21_X1   g03477(.A1(new_n4481_), .A2(new_n4480_), .B(new_n3131_), .ZN(new_n4482_));
  NOR3_X1    g03478(.A1(new_n4481_), .A2(new_n4480_), .A3(new_n3131_), .ZN(new_n4483_));
  OAI21_X1   g03479(.A1(new_n4013_), .A2(new_n4483_), .B(new_n4482_), .ZN(new_n4484_));
  NAND2_X1   g03480(.A1(new_n4471_), .A2(new_n4467_), .ZN(new_n4485_));
  NAND2_X1   g03481(.A1(new_n4477_), .A2(new_n4426_), .ZN(new_n4486_));
  AOI21_X1   g03482(.A1(new_n4485_), .A2(new_n4486_), .B(new_n4484_), .ZN(new_n4487_));
  NOR2_X1    g03483(.A1(new_n4479_), .A2(new_n4487_), .ZN(new_n4488_));
  NOR2_X1    g03484(.A1(new_n4488_), .A2(new_n4391_), .ZN(new_n4489_));
  NAND2_X1   g03485(.A1(new_n4383_), .A2(new_n4376_), .ZN(new_n4490_));
  NAND2_X1   g03486(.A1(new_n4369_), .A2(new_n4327_), .ZN(new_n4491_));
  AOI21_X1   g03487(.A1(new_n4491_), .A2(new_n4490_), .B(new_n4387_), .ZN(new_n4492_));
  NAND2_X1   g03488(.A1(new_n4383_), .A2(new_n4327_), .ZN(new_n4493_));
  NAND2_X1   g03489(.A1(new_n4369_), .A2(new_n4376_), .ZN(new_n4494_));
  AOI21_X1   g03490(.A1(new_n4494_), .A2(new_n4493_), .B(new_n4281_), .ZN(new_n4495_));
  NOR2_X1    g03491(.A1(new_n4495_), .A2(new_n4492_), .ZN(new_n4496_));
  NOR2_X1    g03492(.A1(new_n4471_), .A2(new_n4477_), .ZN(new_n4497_));
  NOR2_X1    g03493(.A1(new_n4467_), .A2(new_n4426_), .ZN(new_n4498_));
  OAI21_X1   g03494(.A1(new_n4497_), .A2(new_n4498_), .B(new_n4484_), .ZN(new_n4499_));
  NOR2_X1    g03495(.A1(new_n4477_), .A2(new_n4426_), .ZN(new_n4500_));
  NOR4_X1    g03496(.A1(new_n4473_), .A2(new_n4476_), .A3(new_n4419_), .A4(new_n4425_), .ZN(new_n4501_));
  OAI21_X1   g03497(.A1(new_n4500_), .A2(new_n4501_), .B(new_n4393_), .ZN(new_n4502_));
  NAND2_X1   g03498(.A1(new_n4499_), .A2(new_n4502_), .ZN(new_n4503_));
  NOR2_X1    g03499(.A1(new_n4496_), .A2(new_n4503_), .ZN(new_n4504_));
  OAI21_X1   g03500(.A1(new_n4489_), .A2(new_n4504_), .B(new_n4276_), .ZN(new_n4505_));
  AOI22_X1   g03501(.A1(new_n4385_), .A2(new_n4390_), .B1(new_n4499_), .B2(new_n4502_), .ZN(new_n4506_));
  NOR2_X1    g03502(.A1(new_n4391_), .A2(new_n4503_), .ZN(new_n4507_));
  OAI21_X1   g03503(.A1(new_n4507_), .A2(new_n4506_), .B(new_n4275_), .ZN(new_n4508_));
  NAND3_X1   g03504(.A1(new_n3935_), .A2(new_n3936_), .A3(new_n3591_), .ZN(new_n4509_));
  NAND2_X1   g03505(.A1(new_n4509_), .A2(new_n3766_), .ZN(new_n4510_));
  NAND2_X1   g03506(.A1(new_n4510_), .A2(new_n3938_), .ZN(new_n4511_));
  AOI21_X1   g03507(.A1(new_n3931_), .A2(new_n3932_), .B(new_n3880_), .ZN(new_n4512_));
  NOR3_X1    g03508(.A1(new_n3929_), .A2(new_n3881_), .A3(new_n3914_), .ZN(new_n4513_));
  OAI21_X1   g03509(.A1(new_n4513_), .A2(new_n4512_), .B(new_n3588_), .ZN(new_n4514_));
  NOR3_X1    g03510(.A1(new_n4513_), .A2(new_n4512_), .A3(new_n3588_), .ZN(new_n4515_));
  OAI21_X1   g03511(.A1(new_n3848_), .A2(new_n4515_), .B(new_n4514_), .ZN(new_n4516_));
  NOR3_X1    g03512(.A1(new_n3923_), .A2(new_n3925_), .A3(new_n3927_), .ZN(new_n4517_));
  NOR2_X1    g03513(.A1(new_n4517_), .A2(new_n3584_), .ZN(new_n4518_));
  NAND4_X1   g03514(.A1(new_n3917_), .A2(new_n3915_), .A3(new_n3857_), .A4(new_n3878_), .ZN(new_n4519_));
  OAI21_X1   g03515(.A1(new_n4518_), .A2(new_n4519_), .B(new_n3913_), .ZN(new_n4520_));
  NOR2_X1    g03516(.A1(new_n3926_), .A2(new_n3911_), .ZN(new_n4521_));
  NAND4_X1   g03517(.A1(new_n4521_), .A2(new_n3538_), .A3(new_n3549_), .A4(new_n3552_), .ZN(new_n4522_));
  INV_X1     g03518(.I(new_n4522_), .ZN(new_n4523_));
  NAND2_X1   g03519(.A1(new_n3550_), .A2(new_n3551_), .ZN(new_n4524_));
  NAND3_X1   g03520(.A1(new_n3538_), .A2(new_n3549_), .A3(new_n4524_), .ZN(new_n4525_));
  NAND2_X1   g03521(.A1(new_n4525_), .A2(new_n3890_), .ZN(new_n4526_));
  OAI21_X1   g03522(.A1(new_n3575_), .A2(new_n3577_), .B(new_n3908_), .ZN(new_n4527_));
  NAND2_X1   g03523(.A1(new_n4527_), .A2(new_n3578_), .ZN(new_n4528_));
  XOR2_X1    g03524(.A1(new_n4528_), .A2(new_n4526_), .Z(new_n4529_));
  NAND3_X1   g03525(.A1(new_n3896_), .A2(new_n3898_), .A3(new_n3894_), .ZN(new_n4530_));
  AOI21_X1   g03526(.A1(new_n4530_), .A2(new_n3888_), .B(new_n3925_), .ZN(new_n4531_));
  OAI21_X1   g03527(.A1(new_n4531_), .A2(new_n4523_), .B(new_n4529_), .ZN(new_n4532_));
  NAND2_X1   g03528(.A1(new_n3496_), .A2(new_n3497_), .ZN(new_n4533_));
  NAND3_X1   g03529(.A1(new_n3484_), .A2(new_n3495_), .A3(new_n4533_), .ZN(new_n4534_));
  NAND2_X1   g03530(.A1(new_n4534_), .A2(new_n3860_), .ZN(new_n4535_));
  NOR2_X1    g03531(.A1(new_n3510_), .A2(new_n3521_), .ZN(new_n4536_));
  NAND2_X1   g03532(.A1(new_n3522_), .A2(new_n3523_), .ZN(new_n4537_));
  NAND2_X1   g03533(.A1(new_n4536_), .A2(new_n4537_), .ZN(new_n4538_));
  NAND2_X1   g03534(.A1(new_n4538_), .A2(new_n3525_), .ZN(new_n4539_));
  XNOR2_X1   g03535(.A1(new_n4539_), .A2(new_n4535_), .ZN(new_n4540_));
  OAI21_X1   g03536(.A1(new_n3875_), .A2(new_n3857_), .B(new_n3856_), .ZN(new_n4541_));
  AOI21_X1   g03537(.A1(new_n4541_), .A2(new_n3916_), .B(new_n4540_), .ZN(new_n4542_));
  NOR2_X1    g03538(.A1(new_n4532_), .A2(new_n4542_), .ZN(new_n4543_));
  XNOR2_X1   g03539(.A1(new_n4528_), .A2(new_n4526_), .ZN(new_n4544_));
  NOR3_X1    g03540(.A1(new_n3922_), .A2(new_n3920_), .A3(new_n3895_), .ZN(new_n4545_));
  OAI21_X1   g03541(.A1(new_n4545_), .A2(new_n3887_), .B(new_n3907_), .ZN(new_n4546_));
  AOI21_X1   g03542(.A1(new_n4522_), .A2(new_n4546_), .B(new_n4544_), .ZN(new_n4547_));
  INV_X1     g03543(.I(new_n3916_), .ZN(new_n4548_));
  XOR2_X1    g03544(.A1(new_n4539_), .A2(new_n4535_), .Z(new_n4549_));
  AOI21_X1   g03545(.A1(new_n3878_), .A2(new_n3858_), .B(new_n3915_), .ZN(new_n4550_));
  OAI21_X1   g03546(.A1(new_n4550_), .A2(new_n4548_), .B(new_n4549_), .ZN(new_n4551_));
  NOR2_X1    g03547(.A1(new_n4547_), .A2(new_n4551_), .ZN(new_n4552_));
  OAI21_X1   g03548(.A1(new_n4543_), .A2(new_n4552_), .B(new_n4520_), .ZN(new_n4553_));
  NAND3_X1   g03549(.A1(new_n3899_), .A2(new_n3912_), .A3(new_n3907_), .ZN(new_n4554_));
  NAND2_X1   g03550(.A1(new_n4554_), .A2(new_n3919_), .ZN(new_n4555_));
  NOR4_X1    g03551(.A1(new_n3885_), .A2(new_n3856_), .A3(new_n3875_), .A4(new_n3858_), .ZN(new_n4556_));
  AOI21_X1   g03552(.A1(new_n4555_), .A2(new_n4556_), .B(new_n3928_), .ZN(new_n4557_));
  NOR2_X1    g03553(.A1(new_n4547_), .A2(new_n4542_), .ZN(new_n4558_));
  NOR2_X1    g03554(.A1(new_n4532_), .A2(new_n4551_), .ZN(new_n4559_));
  OAI21_X1   g03555(.A1(new_n4558_), .A2(new_n4559_), .B(new_n4557_), .ZN(new_n4560_));
  NAND2_X1   g03556(.A1(new_n4553_), .A2(new_n4560_), .ZN(new_n4561_));
  NOR2_X1    g03557(.A1(new_n3844_), .A2(new_n3472_), .ZN(new_n4562_));
  AOI21_X1   g03558(.A1(new_n3387_), .A2(new_n3783_), .B(new_n3786_), .ZN(new_n4563_));
  NOR4_X1    g03559(.A1(new_n3803_), .A2(new_n3768_), .A3(new_n4563_), .A4(new_n3802_), .ZN(new_n4564_));
  INV_X1     g03560(.I(new_n4564_), .ZN(new_n4565_));
  OAI21_X1   g03561(.A1(new_n4565_), .A2(new_n4562_), .B(new_n3845_), .ZN(new_n4566_));
  INV_X1     g03562(.I(new_n3833_), .ZN(new_n4567_));
  NAND2_X1   g03563(.A1(new_n3439_), .A2(new_n3440_), .ZN(new_n4568_));
  NAND3_X1   g03564(.A1(new_n3427_), .A2(new_n3438_), .A3(new_n4568_), .ZN(new_n4569_));
  NAND2_X1   g03565(.A1(new_n4569_), .A2(new_n3812_), .ZN(new_n4570_));
  NAND2_X1   g03566(.A1(new_n3822_), .A2(new_n3824_), .ZN(new_n4571_));
  NOR2_X1    g03567(.A1(new_n3464_), .A2(new_n3466_), .ZN(new_n4572_));
  OAI21_X1   g03568(.A1(new_n4571_), .A2(new_n4572_), .B(new_n3467_), .ZN(new_n4573_));
  XOR2_X1    g03569(.A1(new_n4573_), .A2(new_n4570_), .Z(new_n4574_));
  AOI21_X1   g03570(.A1(new_n3821_), .A2(new_n3810_), .B(new_n3842_), .ZN(new_n4575_));
  OAI21_X1   g03571(.A1(new_n4575_), .A2(new_n4567_), .B(new_n4574_), .ZN(new_n4576_));
  NAND3_X1   g03572(.A1(new_n3793_), .A2(new_n3786_), .A3(new_n3784_), .ZN(new_n4577_));
  NOR2_X1    g03573(.A1(new_n3769_), .A2(new_n3777_), .ZN(new_n4578_));
  NAND2_X1   g03574(.A1(new_n3385_), .A2(new_n3386_), .ZN(new_n4579_));
  AOI21_X1   g03575(.A1(new_n4578_), .A2(new_n4579_), .B(new_n3387_), .ZN(new_n4580_));
  NAND2_X1   g03576(.A1(new_n3795_), .A2(new_n3412_), .ZN(new_n4581_));
  AOI21_X1   g03577(.A1(new_n3787_), .A2(new_n4581_), .B(new_n3796_), .ZN(new_n4582_));
  XNOR2_X1   g03578(.A1(new_n4580_), .A2(new_n4582_), .ZN(new_n4583_));
  OAI21_X1   g03579(.A1(new_n4563_), .A2(new_n3767_), .B(new_n3802_), .ZN(new_n4584_));
  AOI21_X1   g03580(.A1(new_n4584_), .A2(new_n4577_), .B(new_n4583_), .ZN(new_n4585_));
  NOR2_X1    g03581(.A1(new_n4585_), .A2(new_n4576_), .ZN(new_n4586_));
  XNOR2_X1   g03582(.A1(new_n4573_), .A2(new_n4570_), .ZN(new_n4587_));
  NOR3_X1    g03583(.A1(new_n3839_), .A2(new_n3837_), .A3(new_n3817_), .ZN(new_n4588_));
  OAI21_X1   g03584(.A1(new_n4588_), .A2(new_n3809_), .B(new_n3829_), .ZN(new_n4589_));
  AOI21_X1   g03585(.A1(new_n4589_), .A2(new_n3833_), .B(new_n4587_), .ZN(new_n4590_));
  INV_X1     g03586(.I(new_n4577_), .ZN(new_n4591_));
  XOR2_X1    g03587(.A1(new_n4580_), .A2(new_n4582_), .Z(new_n4592_));
  AOI21_X1   g03588(.A1(new_n3785_), .A2(new_n3768_), .B(new_n3806_), .ZN(new_n4593_));
  OAI21_X1   g03589(.A1(new_n4593_), .A2(new_n4591_), .B(new_n4592_), .ZN(new_n4594_));
  NOR2_X1    g03590(.A1(new_n4590_), .A2(new_n4594_), .ZN(new_n4595_));
  NOR2_X1    g03591(.A1(new_n4595_), .A2(new_n4586_), .ZN(new_n4596_));
  NOR2_X1    g03592(.A1(new_n4590_), .A2(new_n4585_), .ZN(new_n4597_));
  NOR2_X1    g03593(.A1(new_n4594_), .A2(new_n4576_), .ZN(new_n4598_));
  NOR2_X1    g03594(.A1(new_n4597_), .A2(new_n4598_), .ZN(new_n4599_));
  MUX2_X1    g03595(.I0(new_n4599_), .I1(new_n4596_), .S(new_n4566_), .Z(new_n4600_));
  NOR2_X1    g03596(.A1(new_n4600_), .A2(new_n4561_), .ZN(new_n4601_));
  NAND2_X1   g03597(.A1(new_n4547_), .A2(new_n4551_), .ZN(new_n4602_));
  NAND2_X1   g03598(.A1(new_n4532_), .A2(new_n4542_), .ZN(new_n4603_));
  AOI21_X1   g03599(.A1(new_n4602_), .A2(new_n4603_), .B(new_n4557_), .ZN(new_n4604_));
  NAND2_X1   g03600(.A1(new_n4532_), .A2(new_n4551_), .ZN(new_n4605_));
  NAND2_X1   g03601(.A1(new_n4547_), .A2(new_n4542_), .ZN(new_n4606_));
  AOI21_X1   g03602(.A1(new_n4605_), .A2(new_n4606_), .B(new_n4520_), .ZN(new_n4607_));
  NOR2_X1    g03603(.A1(new_n4607_), .A2(new_n4604_), .ZN(new_n4608_));
  OAI21_X1   g03604(.A1(new_n4586_), .A2(new_n4595_), .B(new_n4566_), .ZN(new_n4609_));
  NAND2_X1   g03605(.A1(new_n3834_), .A2(new_n3471_), .ZN(new_n4610_));
  AOI21_X1   g03606(.A1(new_n4610_), .A2(new_n4564_), .B(new_n3835_), .ZN(new_n4611_));
  OAI21_X1   g03607(.A1(new_n4597_), .A2(new_n4598_), .B(new_n4611_), .ZN(new_n4612_));
  NAND2_X1   g03608(.A1(new_n4609_), .A2(new_n4612_), .ZN(new_n4613_));
  NOR2_X1    g03609(.A1(new_n4613_), .A2(new_n4608_), .ZN(new_n4614_));
  OAI21_X1   g03610(.A1(new_n4601_), .A2(new_n4614_), .B(new_n4516_), .ZN(new_n4615_));
  NAND3_X1   g03611(.A1(new_n3930_), .A2(new_n3933_), .A3(new_n3587_), .ZN(new_n4616_));
  AOI21_X1   g03612(.A1(new_n3847_), .A2(new_n4616_), .B(new_n3934_), .ZN(new_n4617_));
  AOI22_X1   g03613(.A1(new_n4609_), .A2(new_n4612_), .B1(new_n4553_), .B2(new_n4560_), .ZN(new_n4618_));
  NOR2_X1    g03614(.A1(new_n4613_), .A2(new_n4561_), .ZN(new_n4619_));
  OAI21_X1   g03615(.A1(new_n4619_), .A2(new_n4618_), .B(new_n4617_), .ZN(new_n4620_));
  NAND2_X1   g03616(.A1(new_n4615_), .A2(new_n4620_), .ZN(new_n4621_));
  NAND3_X1   g03617(.A1(new_n3761_), .A2(new_n3764_), .A3(new_n3360_), .ZN(new_n4622_));
  AOI21_X1   g03618(.A1(new_n3679_), .A2(new_n4622_), .B(new_n3765_), .ZN(new_n4623_));
  NAND2_X1   g03619(.A1(new_n3758_), .A2(new_n3757_), .ZN(new_n4624_));
  NOR4_X1    g03620(.A1(new_n3725_), .A2(new_n3692_), .A3(new_n3694_), .A4(new_n3712_), .ZN(new_n4625_));
  AOI21_X1   g03621(.A1(new_n4624_), .A2(new_n4625_), .B(new_n3759_), .ZN(new_n4626_));
  NOR2_X1    g03622(.A1(new_n3338_), .A2(new_n3348_), .ZN(new_n4627_));
  NOR2_X1    g03623(.A1(new_n3742_), .A2(new_n3740_), .ZN(new_n4628_));
  NOR2_X1    g03624(.A1(new_n4628_), .A2(new_n4627_), .ZN(new_n4629_));
  NOR2_X1    g03625(.A1(new_n4629_), .A2(new_n3749_), .ZN(new_n4630_));
  NAND4_X1   g03626(.A1(new_n4630_), .A2(new_n3313_), .A3(new_n3324_), .A4(new_n3327_), .ZN(new_n4631_));
  NAND2_X1   g03627(.A1(new_n3325_), .A2(new_n3326_), .ZN(new_n4632_));
  NAND3_X1   g03628(.A1(new_n3313_), .A2(new_n3324_), .A3(new_n4632_), .ZN(new_n4633_));
  NAND2_X1   g03629(.A1(new_n4633_), .A2(new_n3730_), .ZN(new_n4634_));
  OAI21_X1   g03630(.A1(new_n3350_), .A2(new_n3352_), .B(new_n4627_), .ZN(new_n4635_));
  NAND2_X1   g03631(.A1(new_n4635_), .A2(new_n3353_), .ZN(new_n4636_));
  XNOR2_X1   g03632(.A1(new_n4636_), .A2(new_n4634_), .ZN(new_n4637_));
  INV_X1     g03633(.I(new_n3734_), .ZN(new_n4638_));
  XNOR2_X1   g03634(.A1(new_n3313_), .A2(new_n3324_), .ZN(new_n4639_));
  NOR2_X1    g03635(.A1(new_n4639_), .A2(new_n3730_), .ZN(new_n4640_));
  NOR3_X1    g03636(.A1(new_n4640_), .A2(new_n4638_), .A3(new_n3735_), .ZN(new_n4641_));
  OAI21_X1   g03637(.A1(new_n4641_), .A2(new_n3727_), .B(new_n3747_), .ZN(new_n4642_));
  AOI21_X1   g03638(.A1(new_n4631_), .A2(new_n4642_), .B(new_n4637_), .ZN(new_n4643_));
  INV_X1     g03639(.I(new_n3754_), .ZN(new_n4644_));
  NAND2_X1   g03640(.A1(new_n3271_), .A2(new_n3272_), .ZN(new_n4645_));
  NAND3_X1   g03641(.A1(new_n3259_), .A2(new_n3270_), .A3(new_n4645_), .ZN(new_n4646_));
  NAND2_X1   g03642(.A1(new_n4646_), .A2(new_n3706_), .ZN(new_n4647_));
  NAND2_X1   g03643(.A1(new_n3683_), .A2(new_n3684_), .ZN(new_n4648_));
  NAND2_X1   g03644(.A1(new_n3720_), .A2(new_n4648_), .ZN(new_n4649_));
  NAND2_X1   g03645(.A1(new_n4649_), .A2(new_n3300_), .ZN(new_n4650_));
  XOR2_X1    g03646(.A1(new_n4650_), .A2(new_n4647_), .Z(new_n4651_));
  AOI21_X1   g03647(.A1(new_n3716_), .A2(new_n3694_), .B(new_n3753_), .ZN(new_n4652_));
  OAI21_X1   g03648(.A1(new_n4652_), .A2(new_n4644_), .B(new_n4651_), .ZN(new_n4653_));
  NAND2_X1   g03649(.A1(new_n4643_), .A2(new_n4653_), .ZN(new_n4654_));
  INV_X1     g03650(.I(new_n4631_), .ZN(new_n4655_));
  XOR2_X1    g03651(.A1(new_n4636_), .A2(new_n4634_), .Z(new_n4656_));
  NAND3_X1   g03652(.A1(new_n3738_), .A2(new_n3736_), .A3(new_n3734_), .ZN(new_n4657_));
  INV_X1     g03653(.I(new_n3746_), .ZN(new_n4658_));
  NOR2_X1    g03654(.A1(new_n4658_), .A2(new_n3744_), .ZN(new_n4659_));
  AOI21_X1   g03655(.A1(new_n4657_), .A2(new_n3728_), .B(new_n4659_), .ZN(new_n4660_));
  OAI21_X1   g03656(.A1(new_n4660_), .A2(new_n4655_), .B(new_n4656_), .ZN(new_n4661_));
  XNOR2_X1   g03657(.A1(new_n4650_), .A2(new_n4647_), .ZN(new_n4662_));
  OAI21_X1   g03658(.A1(new_n3712_), .A2(new_n3693_), .B(new_n3692_), .ZN(new_n4663_));
  AOI21_X1   g03659(.A1(new_n4663_), .A2(new_n3754_), .B(new_n4662_), .ZN(new_n4664_));
  NAND2_X1   g03660(.A1(new_n4661_), .A2(new_n4664_), .ZN(new_n4665_));
  AOI21_X1   g03661(.A1(new_n4654_), .A2(new_n4665_), .B(new_n4626_), .ZN(new_n4666_));
  NOR4_X1    g03662(.A1(new_n4640_), .A2(new_n4638_), .A3(new_n3727_), .A4(new_n3735_), .ZN(new_n4667_));
  INV_X1     g03663(.I(new_n3750_), .ZN(new_n4668_));
  NOR3_X1    g03664(.A1(new_n4667_), .A2(new_n4668_), .A3(new_n4659_), .ZN(new_n4669_));
  NOR2_X1    g03665(.A1(new_n4669_), .A2(new_n3357_), .ZN(new_n4670_));
  NAND4_X1   g03666(.A1(new_n3755_), .A2(new_n3753_), .A3(new_n3693_), .A4(new_n3716_), .ZN(new_n4671_));
  OAI21_X1   g03667(.A1(new_n4671_), .A2(new_n4670_), .B(new_n3751_), .ZN(new_n4672_));
  NAND2_X1   g03668(.A1(new_n4661_), .A2(new_n4653_), .ZN(new_n4673_));
  NAND2_X1   g03669(.A1(new_n4643_), .A2(new_n4664_), .ZN(new_n4674_));
  AOI21_X1   g03670(.A1(new_n4673_), .A2(new_n4674_), .B(new_n4672_), .ZN(new_n4675_));
  NOR2_X1    g03671(.A1(new_n4675_), .A2(new_n4666_), .ZN(new_n4676_));
  NOR2_X1    g03672(.A1(new_n3676_), .A2(new_n3247_), .ZN(new_n4677_));
  INV_X1     g03673(.I(new_n3636_), .ZN(new_n4678_));
  NAND4_X1   g03674(.A1(new_n4678_), .A2(new_n3600_), .A3(new_n3618_), .A4(new_n3639_), .ZN(new_n4679_));
  OAI21_X1   g03675(.A1(new_n4679_), .A2(new_n4677_), .B(new_n3677_), .ZN(new_n4680_));
  NOR2_X1    g03676(.A1(new_n3661_), .A2(new_n3662_), .ZN(new_n4681_));
  NAND4_X1   g03677(.A1(new_n4681_), .A2(new_n3202_), .A3(new_n3213_), .A4(new_n3216_), .ZN(new_n4682_));
  NAND2_X1   g03678(.A1(new_n3214_), .A2(new_n3215_), .ZN(new_n4683_));
  NAND3_X1   g03679(.A1(new_n3202_), .A2(new_n3213_), .A3(new_n4683_), .ZN(new_n4684_));
  NAND2_X1   g03680(.A1(new_n4684_), .A2(new_n3660_), .ZN(new_n4685_));
  NAND2_X1   g03681(.A1(new_n3653_), .A2(new_n3651_), .ZN(new_n4686_));
  NOR2_X1    g03682(.A1(new_n3239_), .A2(new_n3241_), .ZN(new_n4687_));
  OAI21_X1   g03683(.A1(new_n4686_), .A2(new_n4687_), .B(new_n3242_), .ZN(new_n4688_));
  XNOR2_X1   g03684(.A1(new_n4688_), .A2(new_n4685_), .ZN(new_n4689_));
  NOR3_X1    g03685(.A1(new_n3672_), .A2(new_n3669_), .A3(new_n3670_), .ZN(new_n4690_));
  OAI21_X1   g03686(.A1(new_n4690_), .A2(new_n3668_), .B(new_n3658_), .ZN(new_n4691_));
  AOI21_X1   g03687(.A1(new_n4691_), .A2(new_n4682_), .B(new_n4689_), .ZN(new_n4692_));
  NAND3_X1   g03688(.A1(new_n3626_), .A2(new_n3619_), .A3(new_n3617_), .ZN(new_n4693_));
  INV_X1     g03689(.I(new_n4693_), .ZN(new_n4694_));
  NOR2_X1    g03690(.A1(new_n3602_), .A2(new_n3610_), .ZN(new_n4695_));
  NAND2_X1   g03691(.A1(new_n3160_), .A2(new_n3161_), .ZN(new_n4696_));
  AOI21_X1   g03692(.A1(new_n4695_), .A2(new_n4696_), .B(new_n3162_), .ZN(new_n4697_));
  NAND2_X1   g03693(.A1(new_n3628_), .A2(new_n3187_), .ZN(new_n4698_));
  AOI21_X1   g03694(.A1(new_n3620_), .A2(new_n4698_), .B(new_n3629_), .ZN(new_n4699_));
  XOR2_X1    g03695(.A1(new_n4697_), .A2(new_n4699_), .Z(new_n4700_));
  AOI21_X1   g03696(.A1(new_n3618_), .A2(new_n3601_), .B(new_n3639_), .ZN(new_n4701_));
  OAI21_X1   g03697(.A1(new_n4701_), .A2(new_n4694_), .B(new_n4700_), .ZN(new_n4702_));
  NAND2_X1   g03698(.A1(new_n4702_), .A2(new_n4692_), .ZN(new_n4703_));
  INV_X1     g03699(.I(new_n4703_), .ZN(new_n4704_));
  NOR2_X1    g03700(.A1(new_n4702_), .A2(new_n4692_), .ZN(new_n4705_));
  OAI21_X1   g03701(.A1(new_n4704_), .A2(new_n4705_), .B(new_n4680_), .ZN(new_n4706_));
  NAND2_X1   g03702(.A1(new_n3665_), .A2(new_n3246_), .ZN(new_n4707_));
  AOI21_X1   g03703(.A1(new_n3162_), .A2(new_n3616_), .B(new_n3619_), .ZN(new_n4708_));
  NOR4_X1    g03704(.A1(new_n3636_), .A2(new_n3601_), .A3(new_n4708_), .A4(new_n3635_), .ZN(new_n4709_));
  AOI21_X1   g03705(.A1(new_n4707_), .A2(new_n4709_), .B(new_n3666_), .ZN(new_n4710_));
  XNOR2_X1   g03706(.A1(new_n4697_), .A2(new_n4699_), .ZN(new_n4711_));
  OAI21_X1   g03707(.A1(new_n4708_), .A2(new_n3600_), .B(new_n3635_), .ZN(new_n4712_));
  AOI21_X1   g03708(.A1(new_n4712_), .A2(new_n4693_), .B(new_n4711_), .ZN(new_n4713_));
  NOR2_X1    g03709(.A1(new_n4713_), .A2(new_n4692_), .ZN(new_n4714_));
  INV_X1     g03710(.I(new_n4682_), .ZN(new_n4715_));
  XOR2_X1    g03711(.A1(new_n4688_), .A2(new_n4685_), .Z(new_n4716_));
  NAND3_X1   g03712(.A1(new_n3649_), .A2(new_n3647_), .A3(new_n3645_), .ZN(new_n4717_));
  AOI21_X1   g03713(.A1(new_n4717_), .A2(new_n3642_), .B(new_n3675_), .ZN(new_n4718_));
  OAI21_X1   g03714(.A1(new_n4718_), .A2(new_n4715_), .B(new_n4716_), .ZN(new_n4719_));
  NOR2_X1    g03715(.A1(new_n4702_), .A2(new_n4719_), .ZN(new_n4720_));
  OAI21_X1   g03716(.A1(new_n4714_), .A2(new_n4720_), .B(new_n4710_), .ZN(new_n4721_));
  NAND2_X1   g03717(.A1(new_n4706_), .A2(new_n4721_), .ZN(new_n4722_));
  NAND2_X1   g03718(.A1(new_n4722_), .A2(new_n4676_), .ZN(new_n4723_));
  NOR2_X1    g03719(.A1(new_n4661_), .A2(new_n4664_), .ZN(new_n4724_));
  NOR2_X1    g03720(.A1(new_n4643_), .A2(new_n4653_), .ZN(new_n4725_));
  OAI21_X1   g03721(.A1(new_n4724_), .A2(new_n4725_), .B(new_n4672_), .ZN(new_n4726_));
  NOR2_X1    g03722(.A1(new_n4643_), .A2(new_n4664_), .ZN(new_n4727_));
  NOR2_X1    g03723(.A1(new_n4661_), .A2(new_n4653_), .ZN(new_n4728_));
  OAI21_X1   g03724(.A1(new_n4727_), .A2(new_n4728_), .B(new_n4626_), .ZN(new_n4729_));
  NAND2_X1   g03725(.A1(new_n4726_), .A2(new_n4729_), .ZN(new_n4730_));
  NAND2_X1   g03726(.A1(new_n4713_), .A2(new_n4719_), .ZN(new_n4731_));
  AOI21_X1   g03727(.A1(new_n4703_), .A2(new_n4731_), .B(new_n4710_), .ZN(new_n4732_));
  NAND2_X1   g03728(.A1(new_n4702_), .A2(new_n4719_), .ZN(new_n4733_));
  NAND2_X1   g03729(.A1(new_n4713_), .A2(new_n4692_), .ZN(new_n4734_));
  AOI21_X1   g03730(.A1(new_n4733_), .A2(new_n4734_), .B(new_n4680_), .ZN(new_n4735_));
  NOR2_X1    g03731(.A1(new_n4735_), .A2(new_n4732_), .ZN(new_n4736_));
  NAND2_X1   g03732(.A1(new_n4736_), .A2(new_n4730_), .ZN(new_n4737_));
  AOI21_X1   g03733(.A1(new_n4723_), .A2(new_n4737_), .B(new_n4623_), .ZN(new_n4738_));
  AOI21_X1   g03734(.A1(new_n3762_), .A2(new_n3763_), .B(new_n3718_), .ZN(new_n4739_));
  NOR3_X1    g03735(.A1(new_n3760_), .A2(new_n3719_), .A3(new_n3752_), .ZN(new_n4740_));
  OAI21_X1   g03736(.A1(new_n4740_), .A2(new_n4739_), .B(new_n3361_), .ZN(new_n4741_));
  NOR3_X1    g03737(.A1(new_n4740_), .A2(new_n4739_), .A3(new_n3361_), .ZN(new_n4742_));
  OAI21_X1   g03738(.A1(new_n3680_), .A2(new_n4742_), .B(new_n4741_), .ZN(new_n4743_));
  NAND2_X1   g03739(.A1(new_n4722_), .A2(new_n4730_), .ZN(new_n4744_));
  NAND2_X1   g03740(.A1(new_n4736_), .A2(new_n4676_), .ZN(new_n4745_));
  AOI21_X1   g03741(.A1(new_n4745_), .A2(new_n4744_), .B(new_n4743_), .ZN(new_n4746_));
  NOR2_X1    g03742(.A1(new_n4746_), .A2(new_n4738_), .ZN(new_n4747_));
  NOR2_X1    g03743(.A1(new_n4747_), .A2(new_n4621_), .ZN(new_n4748_));
  NAND2_X1   g03744(.A1(new_n4613_), .A2(new_n4608_), .ZN(new_n4749_));
  NAND2_X1   g03745(.A1(new_n4600_), .A2(new_n4561_), .ZN(new_n4750_));
  AOI21_X1   g03746(.A1(new_n4750_), .A2(new_n4749_), .B(new_n4617_), .ZN(new_n4751_));
  NAND2_X1   g03747(.A1(new_n4613_), .A2(new_n4561_), .ZN(new_n4752_));
  NAND2_X1   g03748(.A1(new_n4600_), .A2(new_n4608_), .ZN(new_n4753_));
  AOI21_X1   g03749(.A1(new_n4753_), .A2(new_n4752_), .B(new_n4516_), .ZN(new_n4754_));
  NOR2_X1    g03750(.A1(new_n4754_), .A2(new_n4751_), .ZN(new_n4755_));
  NOR2_X1    g03751(.A1(new_n4736_), .A2(new_n4730_), .ZN(new_n4756_));
  NOR2_X1    g03752(.A1(new_n4722_), .A2(new_n4676_), .ZN(new_n4757_));
  OAI21_X1   g03753(.A1(new_n4757_), .A2(new_n4756_), .B(new_n4743_), .ZN(new_n4758_));
  NOR2_X1    g03754(.A1(new_n4736_), .A2(new_n4676_), .ZN(new_n4759_));
  NOR2_X1    g03755(.A1(new_n4722_), .A2(new_n4730_), .ZN(new_n4760_));
  OAI21_X1   g03756(.A1(new_n4759_), .A2(new_n4760_), .B(new_n4623_), .ZN(new_n4761_));
  NAND2_X1   g03757(.A1(new_n4758_), .A2(new_n4761_), .ZN(new_n4762_));
  NOR2_X1    g03758(.A1(new_n4762_), .A2(new_n4755_), .ZN(new_n4763_));
  OAI21_X1   g03759(.A1(new_n4763_), .A2(new_n4748_), .B(new_n4511_), .ZN(new_n4764_));
  AOI21_X1   g03760(.A1(new_n3766_), .A2(new_n4509_), .B(new_n3937_), .ZN(new_n4765_));
  AOI22_X1   g03761(.A1(new_n4758_), .A2(new_n4761_), .B1(new_n4615_), .B2(new_n4620_), .ZN(new_n4766_));
  NOR2_X1    g03762(.A1(new_n4762_), .A2(new_n4621_), .ZN(new_n4767_));
  OAI21_X1   g03763(.A1(new_n4767_), .A2(new_n4766_), .B(new_n4765_), .ZN(new_n4768_));
  NAND2_X1   g03764(.A1(new_n4764_), .A2(new_n4768_), .ZN(new_n4769_));
  NAND3_X1   g03765(.A1(new_n4769_), .A2(new_n4505_), .A3(new_n4508_), .ZN(new_n4770_));
  NAND2_X1   g03766(.A1(new_n4505_), .A2(new_n4508_), .ZN(new_n4771_));
  NAND2_X1   g03767(.A1(new_n4762_), .A2(new_n4755_), .ZN(new_n4772_));
  NAND2_X1   g03768(.A1(new_n4747_), .A2(new_n4621_), .ZN(new_n4773_));
  AOI21_X1   g03769(.A1(new_n4772_), .A2(new_n4773_), .B(new_n4765_), .ZN(new_n4774_));
  OAI22_X1   g03770(.A1(new_n4738_), .A2(new_n4746_), .B1(new_n4754_), .B2(new_n4751_), .ZN(new_n4775_));
  NAND4_X1   g03771(.A1(new_n4615_), .A2(new_n4758_), .A3(new_n4761_), .A4(new_n4620_), .ZN(new_n4776_));
  AOI21_X1   g03772(.A1(new_n4775_), .A2(new_n4776_), .B(new_n4511_), .ZN(new_n4777_));
  NOR2_X1    g03773(.A1(new_n4774_), .A2(new_n4777_), .ZN(new_n4778_));
  NAND2_X1   g03774(.A1(new_n4771_), .A2(new_n4778_), .ZN(new_n4779_));
  AOI21_X1   g03775(.A1(new_n4779_), .A2(new_n4770_), .B(new_n4273_), .ZN(new_n4780_));
  NAND4_X1   g03776(.A1(new_n4505_), .A2(new_n4508_), .A3(new_n4764_), .A4(new_n4768_), .ZN(new_n4781_));
  NAND2_X1   g03777(.A1(new_n4496_), .A2(new_n4503_), .ZN(new_n4782_));
  NAND2_X1   g03778(.A1(new_n4488_), .A2(new_n4391_), .ZN(new_n4783_));
  AOI21_X1   g03779(.A1(new_n4783_), .A2(new_n4782_), .B(new_n4275_), .ZN(new_n4784_));
  INV_X1     g03780(.I(new_n4506_), .ZN(new_n4785_));
  NAND4_X1   g03781(.A1(new_n4385_), .A2(new_n4499_), .A3(new_n4390_), .A4(new_n4502_), .ZN(new_n4786_));
  AOI21_X1   g03782(.A1(new_n4785_), .A2(new_n4786_), .B(new_n4276_), .ZN(new_n4787_));
  OAI22_X1   g03783(.A1(new_n4787_), .A2(new_n4784_), .B1(new_n4774_), .B2(new_n4777_), .ZN(new_n4788_));
  AOI21_X1   g03784(.A1(new_n4788_), .A2(new_n4781_), .B(new_n4272_), .ZN(new_n4789_));
  NOR2_X1    g03785(.A1(new_n4780_), .A2(new_n4789_), .ZN(new_n4790_));
  NAND3_X1   g03786(.A1(new_n2677_), .A2(new_n2678_), .A3(new_n2684_), .ZN(new_n4791_));
  NAND2_X1   g03787(.A1(new_n4791_), .A2(new_n1824_), .ZN(new_n4792_));
  OAI21_X1   g03788(.A1(new_n2679_), .A2(new_n2684_), .B(new_n4792_), .ZN(new_n4793_));
  INV_X1     g03789(.I(new_n2676_), .ZN(new_n4794_));
  NAND3_X1   g03790(.A1(new_n2663_), .A2(new_n2668_), .A3(new_n2675_), .ZN(new_n4795_));
  NAND2_X1   g03791(.A1(new_n4795_), .A2(new_n2230_), .ZN(new_n4796_));
  NAND2_X1   g03792(.A1(new_n4796_), .A2(new_n4794_), .ZN(new_n4797_));
  NAND3_X1   g03793(.A1(new_n2653_), .A2(new_n2656_), .A3(new_n2661_), .ZN(new_n4798_));
  AOI21_X1   g03794(.A1(new_n2667_), .A2(new_n4798_), .B(new_n2662_), .ZN(new_n4799_));
  NAND2_X1   g03795(.A1(new_n2649_), .A2(new_n2650_), .ZN(new_n4800_));
  NOR4_X1    g03796(.A1(new_n2523_), .A2(new_n2453_), .A3(new_n2502_), .A4(new_n2510_), .ZN(new_n4801_));
  AOI21_X1   g03797(.A1(new_n4801_), .A2(new_n4800_), .B(new_n2651_), .ZN(new_n4802_));
  NAND2_X1   g03798(.A1(new_n2595_), .A2(new_n2596_), .ZN(new_n4803_));
  NAND2_X1   g03799(.A1(new_n2584_), .A2(new_n4803_), .ZN(new_n4804_));
  NAND2_X1   g03800(.A1(new_n4804_), .A2(new_n2605_), .ZN(new_n4805_));
  NAND2_X1   g03801(.A1(new_n2599_), .A2(new_n2600_), .ZN(new_n4806_));
  NAND2_X1   g03802(.A1(new_n2547_), .A2(new_n4806_), .ZN(new_n4807_));
  NAND2_X1   g03803(.A1(new_n4807_), .A2(new_n2618_), .ZN(new_n4808_));
  XNOR2_X1   g03804(.A1(new_n4805_), .A2(new_n4808_), .ZN(new_n4809_));
  NOR4_X1    g03805(.A1(new_n2593_), .A2(new_n2561_), .A3(new_n2598_), .A4(new_n2602_), .ZN(new_n4810_));
  OAI21_X1   g03806(.A1(new_n4810_), .A2(new_n2615_), .B(new_n2623_), .ZN(new_n4811_));
  AOI21_X1   g03807(.A1(new_n4811_), .A2(new_n2648_), .B(new_n4809_), .ZN(new_n4812_));
  NAND2_X1   g03808(.A1(new_n2484_), .A2(new_n2485_), .ZN(new_n4813_));
  NAND2_X1   g03809(.A1(new_n2490_), .A2(new_n4813_), .ZN(new_n4814_));
  NAND2_X1   g03810(.A1(new_n4814_), .A2(new_n2507_), .ZN(new_n4815_));
  NAND2_X1   g03811(.A1(new_n2449_), .A2(new_n2450_), .ZN(new_n4816_));
  NAND2_X1   g03812(.A1(new_n2499_), .A2(new_n4816_), .ZN(new_n4817_));
  NAND2_X1   g03813(.A1(new_n4817_), .A2(new_n2628_), .ZN(new_n4818_));
  XOR2_X1    g03814(.A1(new_n4815_), .A2(new_n4818_), .Z(new_n4819_));
  AOI21_X1   g03815(.A1(new_n2502_), .A2(new_n2517_), .B(new_n2640_), .ZN(new_n4820_));
  OAI21_X1   g03816(.A1(new_n4820_), .A2(new_n2522_), .B(new_n4819_), .ZN(new_n4821_));
  NAND2_X1   g03817(.A1(new_n4821_), .A2(new_n4812_), .ZN(new_n4822_));
  NAND2_X1   g03818(.A1(new_n2624_), .A2(new_n2602_), .ZN(new_n4823_));
  NOR4_X1    g03819(.A1(new_n4823_), .A2(new_n2572_), .A3(new_n2583_), .A4(new_n2605_), .ZN(new_n4824_));
  XOR2_X1    g03820(.A1(new_n4805_), .A2(new_n4808_), .Z(new_n4825_));
  AOI21_X1   g03821(.A1(new_n2646_), .A2(new_n2604_), .B(new_n2622_), .ZN(new_n4826_));
  OAI21_X1   g03822(.A1(new_n4826_), .A2(new_n4824_), .B(new_n4825_), .ZN(new_n4827_));
  XNOR2_X1   g03823(.A1(new_n4815_), .A2(new_n4818_), .ZN(new_n4828_));
  OAI21_X1   g03824(.A1(new_n2510_), .A2(new_n2512_), .B(new_n2453_), .ZN(new_n4829_));
  AOI21_X1   g03825(.A1(new_n4829_), .A2(new_n2641_), .B(new_n4828_), .ZN(new_n4830_));
  NAND2_X1   g03826(.A1(new_n4830_), .A2(new_n4827_), .ZN(new_n4831_));
  AOI21_X1   g03827(.A1(new_n4822_), .A2(new_n4831_), .B(new_n4802_), .ZN(new_n4832_));
  NOR4_X1    g03828(.A1(new_n4824_), .A2(new_n2615_), .A3(new_n4810_), .A4(new_n2622_), .ZN(new_n4833_));
  NOR2_X1    g03829(.A1(new_n4833_), .A2(new_n2634_), .ZN(new_n4834_));
  NAND4_X1   g03830(.A1(new_n2642_), .A2(new_n2640_), .A3(new_n2512_), .A4(new_n2517_), .ZN(new_n4835_));
  OAI21_X1   g03831(.A1(new_n4834_), .A2(new_n4835_), .B(new_n2635_), .ZN(new_n4836_));
  NAND2_X1   g03832(.A1(new_n4821_), .A2(new_n4827_), .ZN(new_n4837_));
  NAND2_X1   g03833(.A1(new_n4830_), .A2(new_n4812_), .ZN(new_n4838_));
  AOI21_X1   g03834(.A1(new_n4838_), .A2(new_n4837_), .B(new_n4836_), .ZN(new_n4839_));
  NOR2_X1    g03835(.A1(new_n4832_), .A2(new_n4839_), .ZN(new_n4840_));
  NOR2_X1    g03836(.A1(new_n2399_), .A2(new_n2407_), .ZN(new_n4841_));
  INV_X1     g03837(.I(new_n2299_), .ZN(new_n4842_));
  NAND4_X1   g03838(.A1(new_n4842_), .A2(new_n2258_), .A3(new_n2268_), .A4(new_n2272_), .ZN(new_n4843_));
  NOR2_X1    g03839(.A1(new_n4843_), .A2(new_n2410_), .ZN(new_n4844_));
  NAND4_X1   g03840(.A1(new_n4844_), .A2(new_n2290_), .A3(new_n2298_), .A4(new_n2410_), .ZN(new_n4845_));
  OAI21_X1   g03841(.A1(new_n4845_), .A2(new_n4841_), .B(new_n2408_), .ZN(new_n4846_));
  NAND2_X1   g03842(.A1(new_n2373_), .A2(new_n2374_), .ZN(new_n4847_));
  NAND2_X1   g03843(.A1(new_n2369_), .A2(new_n4847_), .ZN(new_n4848_));
  NAND2_X1   g03844(.A1(new_n4848_), .A2(new_n2387_), .ZN(new_n4849_));
  NAND2_X1   g03845(.A1(new_n2376_), .A2(new_n2377_), .ZN(new_n4850_));
  NAND2_X1   g03846(.A1(new_n2331_), .A2(new_n4850_), .ZN(new_n4851_));
  NAND2_X1   g03847(.A1(new_n4851_), .A2(new_n2379_), .ZN(new_n4852_));
  XOR2_X1    g03848(.A1(new_n4849_), .A2(new_n4852_), .Z(new_n4853_));
  AOI21_X1   g03849(.A1(new_n2413_), .A2(new_n2418_), .B(new_n2395_), .ZN(new_n4854_));
  OAI21_X1   g03850(.A1(new_n4854_), .A2(new_n2398_), .B(new_n4853_), .ZN(new_n4855_));
  NAND2_X1   g03851(.A1(new_n2258_), .A2(new_n2268_), .ZN(new_n4856_));
  NOR4_X1    g03852(.A1(new_n2269_), .A2(new_n2270_), .A3(new_n2255_), .A4(new_n2266_), .ZN(new_n4857_));
  OAI21_X1   g03853(.A1(new_n4856_), .A2(new_n4857_), .B(new_n2271_), .ZN(new_n4858_));
  INV_X1     g03854(.I(new_n2287_), .ZN(new_n4859_));
  NOR3_X1    g03855(.A1(new_n2246_), .A2(new_n2301_), .A3(new_n2283_), .ZN(new_n4860_));
  OAI21_X1   g03856(.A1(new_n4859_), .A2(new_n4860_), .B(new_n2302_), .ZN(new_n4861_));
  XNOR2_X1   g03857(.A1(new_n4861_), .A2(new_n4858_), .ZN(new_n4862_));
  NOR2_X1    g03858(.A1(new_n2294_), .A2(new_n2268_), .ZN(new_n4863_));
  NOR2_X1    g03859(.A1(new_n2292_), .A2(new_n2275_), .ZN(new_n4864_));
  XNOR2_X1   g03860(.A1(new_n2258_), .A2(new_n2268_), .ZN(new_n4865_));
  NOR2_X1    g03861(.A1(new_n4865_), .A2(new_n2271_), .ZN(new_n4866_));
  NOR3_X1    g03862(.A1(new_n4864_), .A2(new_n4863_), .A3(new_n4866_), .ZN(new_n4867_));
  OAI21_X1   g03863(.A1(new_n4867_), .A2(new_n2290_), .B(new_n2304_), .ZN(new_n4868_));
  AOI21_X1   g03864(.A1(new_n4868_), .A2(new_n4843_), .B(new_n4862_), .ZN(new_n4869_));
  NOR2_X1    g03865(.A1(new_n4869_), .A2(new_n4855_), .ZN(new_n4870_));
  XNOR2_X1   g03866(.A1(new_n4849_), .A2(new_n4852_), .ZN(new_n4871_));
  OAI21_X1   g03867(.A1(new_n2390_), .A2(new_n2382_), .B(new_n2419_), .ZN(new_n4872_));
  AOI21_X1   g03868(.A1(new_n4872_), .A2(new_n2420_), .B(new_n4871_), .ZN(new_n4873_));
  XOR2_X1    g03869(.A1(new_n4861_), .A2(new_n4858_), .Z(new_n4874_));
  AOI21_X1   g03870(.A1(new_n2298_), .A2(new_n2291_), .B(new_n2410_), .ZN(new_n4875_));
  OAI21_X1   g03871(.A1(new_n4875_), .A2(new_n2300_), .B(new_n4874_), .ZN(new_n4876_));
  NOR2_X1    g03872(.A1(new_n4876_), .A2(new_n4873_), .ZN(new_n4877_));
  OAI21_X1   g03873(.A1(new_n4877_), .A2(new_n4870_), .B(new_n4846_), .ZN(new_n4878_));
  NAND2_X1   g03874(.A1(new_n2421_), .A2(new_n2423_), .ZN(new_n4879_));
  NOR4_X1    g03875(.A1(new_n2305_), .A2(new_n2291_), .A3(new_n4867_), .A4(new_n2304_), .ZN(new_n4880_));
  AOI21_X1   g03876(.A1(new_n4879_), .A2(new_n4880_), .B(new_n2424_), .ZN(new_n4881_));
  NOR2_X1    g03877(.A1(new_n4869_), .A2(new_n4873_), .ZN(new_n4882_));
  NOR2_X1    g03878(.A1(new_n4876_), .A2(new_n4855_), .ZN(new_n4883_));
  OAI21_X1   g03879(.A1(new_n4882_), .A2(new_n4883_), .B(new_n4881_), .ZN(new_n4884_));
  NAND2_X1   g03880(.A1(new_n4884_), .A2(new_n4878_), .ZN(new_n4885_));
  NAND2_X1   g03881(.A1(new_n4885_), .A2(new_n4840_), .ZN(new_n4886_));
  NOR2_X1    g03882(.A1(new_n4830_), .A2(new_n4827_), .ZN(new_n4887_));
  NOR2_X1    g03883(.A1(new_n4821_), .A2(new_n4812_), .ZN(new_n4888_));
  OAI21_X1   g03884(.A1(new_n4888_), .A2(new_n4887_), .B(new_n4836_), .ZN(new_n4889_));
  NOR2_X1    g03885(.A1(new_n4830_), .A2(new_n4812_), .ZN(new_n4890_));
  NOR2_X1    g03886(.A1(new_n4821_), .A2(new_n4827_), .ZN(new_n4891_));
  OAI21_X1   g03887(.A1(new_n4890_), .A2(new_n4891_), .B(new_n4802_), .ZN(new_n4892_));
  NAND2_X1   g03888(.A1(new_n4892_), .A2(new_n4889_), .ZN(new_n4893_));
  NAND2_X1   g03889(.A1(new_n4876_), .A2(new_n4873_), .ZN(new_n4894_));
  NAND2_X1   g03890(.A1(new_n4869_), .A2(new_n4855_), .ZN(new_n4895_));
  AOI21_X1   g03891(.A1(new_n4895_), .A2(new_n4894_), .B(new_n4881_), .ZN(new_n4896_));
  NAND2_X1   g03892(.A1(new_n4876_), .A2(new_n4855_), .ZN(new_n4897_));
  NAND2_X1   g03893(.A1(new_n4869_), .A2(new_n4873_), .ZN(new_n4898_));
  AOI21_X1   g03894(.A1(new_n4898_), .A2(new_n4897_), .B(new_n4846_), .ZN(new_n4899_));
  NOR2_X1    g03895(.A1(new_n4896_), .A2(new_n4899_), .ZN(new_n4900_));
  NAND2_X1   g03896(.A1(new_n4900_), .A2(new_n4893_), .ZN(new_n4901_));
  AOI21_X1   g03897(.A1(new_n4901_), .A2(new_n4886_), .B(new_n4799_), .ZN(new_n4902_));
  AOI21_X1   g03898(.A1(new_n2654_), .A2(new_n2655_), .B(new_n2519_), .ZN(new_n4903_));
  NOR3_X1    g03899(.A1(new_n2652_), .A2(new_n2636_), .A3(new_n2520_), .ZN(new_n4904_));
  OAI21_X1   g03900(.A1(new_n4904_), .A2(new_n4903_), .B(new_n2672_), .ZN(new_n4905_));
  NOR3_X1    g03901(.A1(new_n4904_), .A2(new_n4903_), .A3(new_n2672_), .ZN(new_n4906_));
  OAI21_X1   g03902(.A1(new_n2426_), .A2(new_n4906_), .B(new_n4905_), .ZN(new_n4907_));
  NAND2_X1   g03903(.A1(new_n4885_), .A2(new_n4893_), .ZN(new_n4908_));
  NAND2_X1   g03904(.A1(new_n4900_), .A2(new_n4840_), .ZN(new_n4909_));
  AOI21_X1   g03905(.A1(new_n4909_), .A2(new_n4908_), .B(new_n4907_), .ZN(new_n4910_));
  NAND3_X1   g03906(.A1(new_n2215_), .A2(new_n2220_), .A3(new_n2228_), .ZN(new_n4911_));
  AOI21_X1   g03907(.A1(new_n2004_), .A2(new_n4911_), .B(new_n2229_), .ZN(new_n4912_));
  NAND2_X1   g03908(.A1(new_n2212_), .A2(new_n2213_), .ZN(new_n4913_));
  NOR2_X1    g03909(.A1(new_n2212_), .A2(new_n2213_), .ZN(new_n4914_));
  NAND3_X1   g03910(.A1(new_n2086_), .A2(new_n2041_), .A3(new_n2095_), .ZN(new_n4915_));
  OAI21_X1   g03911(.A1(new_n4914_), .A2(new_n4915_), .B(new_n4913_), .ZN(new_n4916_));
  NAND2_X1   g03912(.A1(new_n2170_), .A2(new_n2171_), .ZN(new_n4917_));
  NAND2_X1   g03913(.A1(new_n2155_), .A2(new_n4917_), .ZN(new_n4918_));
  NAND2_X1   g03914(.A1(new_n4918_), .A2(new_n2173_), .ZN(new_n4919_));
  NAND2_X1   g03915(.A1(new_n2175_), .A2(new_n2176_), .ZN(new_n4920_));
  NAND2_X1   g03916(.A1(new_n2118_), .A2(new_n4920_), .ZN(new_n4921_));
  NAND2_X1   g03917(.A1(new_n4921_), .A2(new_n2177_), .ZN(new_n4922_));
  XOR2_X1    g03918(.A1(new_n4919_), .A2(new_n4922_), .Z(new_n4923_));
  AOI21_X1   g03919(.A1(new_n2190_), .A2(new_n2181_), .B(new_n2211_), .ZN(new_n4924_));
  OAI21_X1   g03920(.A1(new_n4924_), .A2(new_n2198_), .B(new_n4923_), .ZN(new_n4925_));
  INV_X1     g03921(.I(new_n2089_), .ZN(new_n4926_));
  NOR3_X1    g03922(.A1(new_n4926_), .A2(new_n2053_), .A3(new_n2064_), .ZN(new_n4927_));
  NOR2_X1    g03923(.A1(new_n4927_), .A2(new_n2067_), .ZN(new_n4928_));
  NAND2_X1   g03924(.A1(new_n2036_), .A2(new_n2026_), .ZN(new_n4929_));
  NOR2_X1    g03925(.A1(new_n2028_), .A2(new_n2030_), .ZN(new_n4930_));
  OAI21_X1   g03926(.A1(new_n4929_), .A2(new_n4930_), .B(new_n2031_), .ZN(new_n4931_));
  XOR2_X1    g03927(.A1(new_n4931_), .A2(new_n4928_), .Z(new_n4932_));
  OAI21_X1   g03928(.A1(new_n2071_), .A2(new_n2085_), .B(new_n2040_), .ZN(new_n4933_));
  AOI21_X1   g03929(.A1(new_n2092_), .A2(new_n4933_), .B(new_n4932_), .ZN(new_n4934_));
  NOR2_X1    g03930(.A1(new_n4934_), .A2(new_n4925_), .ZN(new_n4935_));
  XNOR2_X1   g03931(.A1(new_n4919_), .A2(new_n4922_), .ZN(new_n4936_));
  OAI21_X1   g03932(.A1(new_n2210_), .A2(new_n2180_), .B(new_n2195_), .ZN(new_n4937_));
  AOI21_X1   g03933(.A1(new_n4937_), .A2(new_n2199_), .B(new_n4936_), .ZN(new_n4938_));
  XNOR2_X1   g03934(.A1(new_n4931_), .A2(new_n4928_), .ZN(new_n4939_));
  INV_X1     g03935(.I(new_n4933_), .ZN(new_n4940_));
  OAI21_X1   g03936(.A1(new_n4940_), .A2(new_n2091_), .B(new_n4939_), .ZN(new_n4941_));
  NOR2_X1    g03937(.A1(new_n4941_), .A2(new_n4938_), .ZN(new_n4942_));
  OAI21_X1   g03938(.A1(new_n4935_), .A2(new_n4942_), .B(new_n4916_), .ZN(new_n4943_));
  NOR2_X1    g03939(.A1(new_n2200_), .A2(new_n2205_), .ZN(new_n4944_));
  NAND2_X1   g03940(.A1(new_n2200_), .A2(new_n2205_), .ZN(new_n4945_));
  NOR3_X1    g03941(.A1(new_n2216_), .A2(new_n2040_), .A3(new_n2094_), .ZN(new_n4946_));
  AOI21_X1   g03942(.A1(new_n4945_), .A2(new_n4946_), .B(new_n4944_), .ZN(new_n4947_));
  NOR2_X1    g03943(.A1(new_n4938_), .A2(new_n4934_), .ZN(new_n4948_));
  NOR2_X1    g03944(.A1(new_n4941_), .A2(new_n4925_), .ZN(new_n4949_));
  OAI21_X1   g03945(.A1(new_n4948_), .A2(new_n4949_), .B(new_n4947_), .ZN(new_n4950_));
  NAND2_X1   g03946(.A1(new_n1980_), .A2(new_n1983_), .ZN(new_n4951_));
  AOI21_X1   g03947(.A1(new_n1995_), .A2(new_n1994_), .B(new_n1993_), .ZN(new_n4952_));
  NOR3_X1    g03948(.A1(new_n1989_), .A2(new_n1991_), .A3(new_n1930_), .ZN(new_n4953_));
  NOR2_X1    g03949(.A1(new_n4952_), .A2(new_n4953_), .ZN(new_n4954_));
  NOR3_X1    g03950(.A1(new_n4954_), .A2(new_n4951_), .A3(new_n1986_), .ZN(new_n4955_));
  NAND2_X1   g03951(.A1(new_n4955_), .A2(new_n2223_), .ZN(new_n4956_));
  NOR2_X1    g03952(.A1(new_n4955_), .A2(new_n2223_), .ZN(new_n4957_));
  NOR4_X1    g03953(.A1(new_n1906_), .A2(new_n1901_), .A3(new_n1878_), .A4(new_n1907_), .ZN(new_n4958_));
  INV_X1     g03954(.I(new_n4958_), .ZN(new_n4959_));
  OAI21_X1   g03955(.A1(new_n4959_), .A2(new_n4957_), .B(new_n4956_), .ZN(new_n4960_));
  NAND2_X1   g03956(.A1(new_n1999_), .A2(new_n4951_), .ZN(new_n4961_));
  INV_X1     g03957(.I(new_n4961_), .ZN(new_n4962_));
  NOR3_X1    g03958(.A1(new_n1998_), .A2(new_n1978_), .A3(new_n1970_), .ZN(new_n4963_));
  NOR2_X1    g03959(.A1(new_n4963_), .A2(new_n1961_), .ZN(new_n4964_));
  NOR2_X1    g03960(.A1(new_n1934_), .A2(new_n1932_), .ZN(new_n4965_));
  OR3_X2     g03961(.A1(new_n1919_), .A2(new_n1930_), .A3(new_n4965_), .Z(new_n4966_));
  NAND2_X1   g03962(.A1(new_n4966_), .A2(new_n1935_), .ZN(new_n4967_));
  XNOR2_X1   g03963(.A1(new_n4967_), .A2(new_n4964_), .ZN(new_n4968_));
  AOI21_X1   g03964(.A1(new_n1984_), .A2(new_n1987_), .B(new_n4954_), .ZN(new_n4969_));
  OAI21_X1   g03965(.A1(new_n4969_), .A2(new_n4962_), .B(new_n4968_), .ZN(new_n4970_));
  NAND2_X1   g03966(.A1(new_n1894_), .A2(new_n1907_), .ZN(new_n4971_));
  NAND3_X1   g03967(.A1(new_n1889_), .A2(new_n1884_), .A3(new_n1893_), .ZN(new_n4972_));
  NAND2_X1   g03968(.A1(new_n4972_), .A2(new_n1876_), .ZN(new_n4973_));
  NOR2_X1    g03969(.A1(new_n1835_), .A2(new_n1845_), .ZN(new_n4974_));
  INV_X1     g03970(.I(new_n1850_), .ZN(new_n4975_));
  NAND4_X1   g03971(.A1(new_n1846_), .A2(new_n1848_), .A3(new_n1833_), .A4(new_n1843_), .ZN(new_n4976_));
  AOI21_X1   g03972(.A1(new_n4974_), .A2(new_n4976_), .B(new_n4975_), .ZN(new_n4977_));
  XOR2_X1    g03973(.A1(new_n4973_), .A2(new_n4977_), .Z(new_n4978_));
  INV_X1     g03974(.I(new_n1878_), .ZN(new_n4979_));
  OAI22_X1   g03975(.A1(new_n1897_), .A2(new_n1899_), .B1(new_n1907_), .B2(new_n4979_), .ZN(new_n4980_));
  AOI21_X1   g03976(.A1(new_n4971_), .A2(new_n4980_), .B(new_n4978_), .ZN(new_n4981_));
  NOR2_X1    g03977(.A1(new_n4970_), .A2(new_n4981_), .ZN(new_n4982_));
  XOR2_X1    g03978(.A1(new_n4967_), .A2(new_n4964_), .Z(new_n4983_));
  OAI21_X1   g03979(.A1(new_n4951_), .A2(new_n1986_), .B(new_n1997_), .ZN(new_n4984_));
  AOI21_X1   g03980(.A1(new_n4984_), .A2(new_n4961_), .B(new_n4983_), .ZN(new_n4985_));
  INV_X1     g03981(.I(new_n4971_), .ZN(new_n4986_));
  XNOR2_X1   g03982(.A1(new_n4973_), .A2(new_n4977_), .ZN(new_n4987_));
  NOR2_X1    g03983(.A1(new_n1907_), .A2(new_n4979_), .ZN(new_n4988_));
  NOR2_X1    g03984(.A1(new_n1900_), .A2(new_n4988_), .ZN(new_n4989_));
  OAI21_X1   g03985(.A1(new_n4989_), .A2(new_n4986_), .B(new_n4987_), .ZN(new_n4990_));
  NOR2_X1    g03986(.A1(new_n4990_), .A2(new_n4985_), .ZN(new_n4991_));
  OAI21_X1   g03987(.A1(new_n4991_), .A2(new_n4982_), .B(new_n4960_), .ZN(new_n4992_));
  NAND2_X1   g03988(.A1(new_n2000_), .A2(new_n1964_), .ZN(new_n4993_));
  AOI21_X1   g03989(.A1(new_n4958_), .A2(new_n4993_), .B(new_n2001_), .ZN(new_n4994_));
  NOR2_X1    g03990(.A1(new_n4985_), .A2(new_n4981_), .ZN(new_n4995_));
  NOR2_X1    g03991(.A1(new_n4970_), .A2(new_n4990_), .ZN(new_n4996_));
  OAI21_X1   g03992(.A1(new_n4996_), .A2(new_n4995_), .B(new_n4994_), .ZN(new_n4997_));
  NAND2_X1   g03993(.A1(new_n4992_), .A2(new_n4997_), .ZN(new_n4998_));
  NAND3_X1   g03994(.A1(new_n4998_), .A2(new_n4943_), .A3(new_n4950_), .ZN(new_n4999_));
  NAND2_X1   g03995(.A1(new_n4941_), .A2(new_n4938_), .ZN(new_n5000_));
  NAND2_X1   g03996(.A1(new_n4934_), .A2(new_n4925_), .ZN(new_n5001_));
  AOI21_X1   g03997(.A1(new_n5000_), .A2(new_n5001_), .B(new_n4947_), .ZN(new_n5002_));
  NAND2_X1   g03998(.A1(new_n4941_), .A2(new_n4925_), .ZN(new_n5003_));
  NAND2_X1   g03999(.A1(new_n4938_), .A2(new_n4934_), .ZN(new_n5004_));
  AOI21_X1   g04000(.A1(new_n5003_), .A2(new_n5004_), .B(new_n4916_), .ZN(new_n5005_));
  NAND2_X1   g04001(.A1(new_n4990_), .A2(new_n4985_), .ZN(new_n5006_));
  NAND2_X1   g04002(.A1(new_n4970_), .A2(new_n4981_), .ZN(new_n5007_));
  AOI21_X1   g04003(.A1(new_n5006_), .A2(new_n5007_), .B(new_n4994_), .ZN(new_n5008_));
  NAND2_X1   g04004(.A1(new_n4970_), .A2(new_n4990_), .ZN(new_n5009_));
  NAND2_X1   g04005(.A1(new_n4985_), .A2(new_n4981_), .ZN(new_n5010_));
  AOI21_X1   g04006(.A1(new_n5009_), .A2(new_n5010_), .B(new_n4960_), .ZN(new_n5011_));
  NOR2_X1    g04007(.A1(new_n5011_), .A2(new_n5008_), .ZN(new_n5012_));
  OAI21_X1   g04008(.A1(new_n5002_), .A2(new_n5005_), .B(new_n5012_), .ZN(new_n5013_));
  AOI21_X1   g04009(.A1(new_n5013_), .A2(new_n4999_), .B(new_n4912_), .ZN(new_n5014_));
  AOI21_X1   g04010(.A1(new_n2219_), .A2(new_n2218_), .B(new_n2217_), .ZN(new_n5015_));
  NOR3_X1    g04011(.A1(new_n2206_), .A2(new_n2214_), .A3(new_n2087_), .ZN(new_n5016_));
  OAI21_X1   g04012(.A1(new_n5015_), .A2(new_n5016_), .B(new_n2669_), .ZN(new_n5017_));
  NOR3_X1    g04013(.A1(new_n5015_), .A2(new_n5016_), .A3(new_n2669_), .ZN(new_n5018_));
  OAI21_X1   g04014(.A1(new_n2005_), .A2(new_n5018_), .B(new_n5017_), .ZN(new_n5019_));
  OAI21_X1   g04015(.A1(new_n5002_), .A2(new_n5005_), .B(new_n4998_), .ZN(new_n5020_));
  NAND3_X1   g04016(.A1(new_n5012_), .A2(new_n4943_), .A3(new_n4950_), .ZN(new_n5021_));
  AOI21_X1   g04017(.A1(new_n5020_), .A2(new_n5021_), .B(new_n5019_), .ZN(new_n5022_));
  NOR2_X1    g04018(.A1(new_n5014_), .A2(new_n5022_), .ZN(new_n5023_));
  NOR3_X1    g04019(.A1(new_n5023_), .A2(new_n4902_), .A3(new_n4910_), .ZN(new_n5024_));
  NOR2_X1    g04020(.A1(new_n4900_), .A2(new_n4893_), .ZN(new_n5025_));
  NOR2_X1    g04021(.A1(new_n4885_), .A2(new_n4840_), .ZN(new_n5026_));
  OAI21_X1   g04022(.A1(new_n5025_), .A2(new_n5026_), .B(new_n4907_), .ZN(new_n5027_));
  NOR2_X1    g04023(.A1(new_n4900_), .A2(new_n4840_), .ZN(new_n5028_));
  NOR2_X1    g04024(.A1(new_n4885_), .A2(new_n4893_), .ZN(new_n5029_));
  OAI21_X1   g04025(.A1(new_n5028_), .A2(new_n5029_), .B(new_n4799_), .ZN(new_n5030_));
  NOR3_X1    g04026(.A1(new_n5012_), .A2(new_n5002_), .A3(new_n5005_), .ZN(new_n5031_));
  AOI21_X1   g04027(.A1(new_n4943_), .A2(new_n4950_), .B(new_n4998_), .ZN(new_n5032_));
  OAI21_X1   g04028(.A1(new_n5032_), .A2(new_n5031_), .B(new_n5019_), .ZN(new_n5033_));
  AOI22_X1   g04029(.A1(new_n4950_), .A2(new_n4943_), .B1(new_n4992_), .B2(new_n4997_), .ZN(new_n5034_));
  NOR3_X1    g04030(.A1(new_n4998_), .A2(new_n5002_), .A3(new_n5005_), .ZN(new_n5035_));
  OAI21_X1   g04031(.A1(new_n5035_), .A2(new_n5034_), .B(new_n4912_), .ZN(new_n5036_));
  NAND2_X1   g04032(.A1(new_n5033_), .A2(new_n5036_), .ZN(new_n5037_));
  AOI21_X1   g04033(.A1(new_n5027_), .A2(new_n5030_), .B(new_n5037_), .ZN(new_n5038_));
  OAI21_X1   g04034(.A1(new_n5038_), .A2(new_n5024_), .B(new_n4797_), .ZN(new_n5039_));
  AOI21_X1   g04035(.A1(new_n2230_), .A2(new_n4795_), .B(new_n2676_), .ZN(new_n5040_));
  AOI22_X1   g04036(.A1(new_n5030_), .A2(new_n5027_), .B1(new_n5033_), .B2(new_n5036_), .ZN(new_n5041_));
  NOR3_X1    g04037(.A1(new_n5037_), .A2(new_n4902_), .A3(new_n4910_), .ZN(new_n5042_));
  OAI21_X1   g04038(.A1(new_n5041_), .A2(new_n5042_), .B(new_n5040_), .ZN(new_n5043_));
  NAND2_X1   g04039(.A1(new_n5039_), .A2(new_n5043_), .ZN(new_n5044_));
  NOR2_X1    g04040(.A1(new_n1175_), .A2(new_n1365_), .ZN(new_n5045_));
  NAND3_X1   g04041(.A1(new_n1812_), .A2(new_n1815_), .A3(new_n1822_), .ZN(new_n5046_));
  AOI21_X1   g04042(.A1(new_n5045_), .A2(new_n5046_), .B(new_n1823_), .ZN(new_n5047_));
  INV_X1     g04043(.I(new_n1724_), .ZN(new_n5048_));
  AOI21_X1   g04044(.A1(new_n1808_), .A2(new_n1809_), .B(new_n1807_), .ZN(new_n5049_));
  NOR3_X1    g04045(.A1(new_n1784_), .A2(new_n1754_), .A3(new_n1805_), .ZN(new_n5050_));
  NOR2_X1    g04046(.A1(new_n5049_), .A2(new_n5050_), .ZN(new_n5051_));
  AOI21_X1   g04047(.A1(new_n5051_), .A2(new_n5048_), .B(new_n1604_), .ZN(new_n5052_));
  NOR2_X1    g04048(.A1(new_n1782_), .A2(new_n1723_), .ZN(new_n5053_));
  NAND4_X1   g04049(.A1(new_n1787_), .A2(new_n1733_), .A3(new_n1734_), .A4(new_n1755_), .ZN(new_n5054_));
  OAI21_X1   g04050(.A1(new_n5053_), .A2(new_n5054_), .B(new_n1783_), .ZN(new_n5055_));
  NAND2_X1   g04051(.A1(new_n1676_), .A2(new_n1686_), .ZN(new_n5056_));
  NOR2_X1    g04052(.A1(new_n1688_), .A2(new_n1690_), .ZN(new_n5057_));
  OAI21_X1   g04053(.A1(new_n5056_), .A2(new_n5057_), .B(new_n1691_), .ZN(new_n5058_));
  OAI21_X1   g04054(.A1(new_n1715_), .A2(new_n1717_), .B(new_n1775_), .ZN(new_n5059_));
  NAND2_X1   g04055(.A1(new_n5059_), .A2(new_n1718_), .ZN(new_n5060_));
  XOR2_X1    g04056(.A1(new_n5060_), .A2(new_n5058_), .Z(new_n5061_));
  AOI21_X1   g04057(.A1(new_n1789_), .A2(new_n1794_), .B(new_n1773_), .ZN(new_n5062_));
  OAI21_X1   g04058(.A1(new_n5062_), .A2(new_n1781_), .B(new_n5061_), .ZN(new_n5063_));
  NAND2_X1   g04059(.A1(new_n1636_), .A2(new_n1637_), .ZN(new_n5064_));
  NAND3_X1   g04060(.A1(new_n1624_), .A2(new_n1635_), .A3(new_n5064_), .ZN(new_n5065_));
  NAND2_X1   g04061(.A1(new_n5065_), .A2(new_n1736_), .ZN(new_n5066_));
  OAI21_X1   g04062(.A1(new_n1661_), .A2(new_n1663_), .B(new_n1756_), .ZN(new_n5067_));
  NAND2_X1   g04063(.A1(new_n5067_), .A2(new_n1664_), .ZN(new_n5068_));
  XNOR2_X1   g04064(.A1(new_n5068_), .A2(new_n5066_), .ZN(new_n5069_));
  OAI21_X1   g04065(.A1(new_n1752_), .A2(new_n1734_), .B(new_n1732_), .ZN(new_n5070_));
  AOI21_X1   g04066(.A1(new_n1786_), .A2(new_n5070_), .B(new_n5069_), .ZN(new_n5071_));
  NOR2_X1    g04067(.A1(new_n5063_), .A2(new_n5071_), .ZN(new_n5072_));
  XNOR2_X1   g04068(.A1(new_n5060_), .A2(new_n5058_), .ZN(new_n5073_));
  OAI21_X1   g04069(.A1(new_n1771_), .A2(new_n1763_), .B(new_n1798_), .ZN(new_n5074_));
  AOI21_X1   g04070(.A1(new_n5074_), .A2(new_n1802_), .B(new_n5073_), .ZN(new_n5075_));
  INV_X1     g04071(.I(new_n1786_), .ZN(new_n5076_));
  XOR2_X1    g04072(.A1(new_n5068_), .A2(new_n5066_), .Z(new_n5077_));
  INV_X1     g04073(.I(new_n5070_), .ZN(new_n5078_));
  OAI21_X1   g04074(.A1(new_n5078_), .A2(new_n5076_), .B(new_n5077_), .ZN(new_n5079_));
  NOR2_X1    g04075(.A1(new_n5079_), .A2(new_n5075_), .ZN(new_n5080_));
  OAI21_X1   g04076(.A1(new_n5072_), .A2(new_n5080_), .B(new_n5055_), .ZN(new_n5081_));
  NAND2_X1   g04077(.A1(new_n1803_), .A2(new_n1722_), .ZN(new_n5082_));
  INV_X1     g04078(.I(new_n1734_), .ZN(new_n5083_));
  NOR4_X1    g04079(.A1(new_n1761_), .A2(new_n1732_), .A3(new_n5083_), .A4(new_n1752_), .ZN(new_n5084_));
  AOI21_X1   g04080(.A1(new_n5082_), .A2(new_n5084_), .B(new_n1804_), .ZN(new_n5085_));
  NOR2_X1    g04081(.A1(new_n5075_), .A2(new_n5071_), .ZN(new_n5086_));
  NOR2_X1    g04082(.A1(new_n5079_), .A2(new_n5063_), .ZN(new_n5087_));
  OAI21_X1   g04083(.A1(new_n5086_), .A2(new_n5087_), .B(new_n5085_), .ZN(new_n5088_));
  NAND2_X1   g04084(.A1(new_n5081_), .A2(new_n5088_), .ZN(new_n5089_));
  INV_X1     g04085(.I(new_n1577_), .ZN(new_n5090_));
  XNOR2_X1   g04086(.A1(new_n1579_), .A2(new_n1581_), .ZN(new_n5091_));
  NOR2_X1    g04087(.A1(new_n5091_), .A2(new_n1585_), .ZN(new_n5092_));
  NAND2_X1   g04088(.A1(new_n5090_), .A2(new_n5092_), .ZN(new_n5093_));
  NAND2_X1   g04089(.A1(new_n1587_), .A2(new_n1577_), .ZN(new_n5094_));
  NAND4_X1   g04090(.A1(new_n1599_), .A2(new_n1410_), .A3(new_n1455_), .A4(new_n1591_), .ZN(new_n5095_));
  INV_X1     g04091(.I(new_n5095_), .ZN(new_n5096_));
  NAND2_X1   g04092(.A1(new_n5096_), .A2(new_n5094_), .ZN(new_n5097_));
  NAND2_X1   g04093(.A1(new_n5097_), .A2(new_n5093_), .ZN(new_n5098_));
  INV_X1     g04094(.I(new_n1598_), .ZN(new_n5099_));
  NAND2_X1   g04095(.A1(new_n1596_), .A2(new_n1437_), .ZN(new_n5100_));
  NAND2_X1   g04096(.A1(new_n1377_), .A2(new_n1381_), .ZN(new_n5101_));
  NAND2_X1   g04097(.A1(new_n1456_), .A2(new_n5101_), .ZN(new_n5102_));
  NAND2_X1   g04098(.A1(new_n5102_), .A2(new_n1392_), .ZN(new_n5103_));
  NAND2_X1   g04099(.A1(new_n5100_), .A2(new_n5103_), .ZN(new_n5104_));
  INV_X1     g04100(.I(new_n5104_), .ZN(new_n5105_));
  OAI21_X1   g04101(.A1(new_n1591_), .A2(new_n1589_), .B(new_n1409_), .ZN(new_n5106_));
  NAND2_X1   g04102(.A1(new_n5106_), .A2(new_n5105_), .ZN(new_n5107_));
  NAND2_X1   g04103(.A1(new_n1465_), .A2(new_n1455_), .ZN(new_n5108_));
  NAND3_X1   g04104(.A1(new_n5108_), .A2(new_n1409_), .A3(new_n5104_), .ZN(new_n5109_));
  AOI21_X1   g04105(.A1(new_n5107_), .A2(new_n5109_), .B(new_n5099_), .ZN(new_n5110_));
  AOI21_X1   g04106(.A1(new_n5108_), .A2(new_n1409_), .B(new_n5104_), .ZN(new_n5111_));
  NOR2_X1    g04107(.A1(new_n5106_), .A2(new_n5105_), .ZN(new_n5112_));
  NOR3_X1    g04108(.A1(new_n5112_), .A2(new_n5111_), .A3(new_n1598_), .ZN(new_n5113_));
  NOR2_X1    g04109(.A1(new_n5113_), .A2(new_n5110_), .ZN(new_n5114_));
  OAI21_X1   g04110(.A1(new_n1541_), .A2(new_n1547_), .B(new_n1557_), .ZN(new_n5115_));
  NAND2_X1   g04111(.A1(new_n1548_), .A2(new_n1549_), .ZN(new_n5116_));
  NAND2_X1   g04112(.A1(new_n1491_), .A2(new_n5116_), .ZN(new_n5117_));
  NAND2_X1   g04113(.A1(new_n5117_), .A2(new_n1551_), .ZN(new_n5118_));
  NAND2_X1   g04114(.A1(new_n5118_), .A2(new_n5115_), .ZN(new_n5119_));
  NAND2_X1   g04115(.A1(new_n1554_), .A2(new_n1562_), .ZN(new_n5120_));
  AOI21_X1   g04116(.A1(new_n5120_), .A2(new_n1568_), .B(new_n5119_), .ZN(new_n5121_));
  INV_X1     g04117(.I(new_n5119_), .ZN(new_n5122_));
  OAI21_X1   g04118(.A1(new_n1528_), .A2(new_n1573_), .B(new_n1578_), .ZN(new_n5123_));
  NOR2_X1    g04119(.A1(new_n1572_), .A2(new_n5123_), .ZN(new_n5124_));
  INV_X1     g04120(.I(new_n1559_), .ZN(new_n5125_));
  NAND2_X1   g04121(.A1(new_n5125_), .A2(new_n1560_), .ZN(new_n5126_));
  OAI21_X1   g04122(.A1(new_n5124_), .A2(new_n5126_), .B(new_n1568_), .ZN(new_n5127_));
  NOR2_X1    g04123(.A1(new_n5127_), .A2(new_n5122_), .ZN(new_n5128_));
  OAI21_X1   g04124(.A1(new_n5128_), .A2(new_n5121_), .B(new_n1576_), .ZN(new_n5129_));
  INV_X1     g04125(.I(new_n1576_), .ZN(new_n5130_));
  NAND2_X1   g04126(.A1(new_n5127_), .A2(new_n5122_), .ZN(new_n5131_));
  NAND3_X1   g04127(.A1(new_n5120_), .A2(new_n1568_), .A3(new_n5119_), .ZN(new_n5132_));
  NAND3_X1   g04128(.A1(new_n5131_), .A2(new_n5132_), .A3(new_n5130_), .ZN(new_n5133_));
  NAND2_X1   g04129(.A1(new_n5129_), .A2(new_n5133_), .ZN(new_n5134_));
  NOR2_X1    g04130(.A1(new_n5134_), .A2(new_n5114_), .ZN(new_n5135_));
  OAI21_X1   g04131(.A1(new_n5112_), .A2(new_n5111_), .B(new_n1598_), .ZN(new_n5136_));
  NAND3_X1   g04132(.A1(new_n5107_), .A2(new_n5109_), .A3(new_n5099_), .ZN(new_n5137_));
  NAND2_X1   g04133(.A1(new_n5136_), .A2(new_n5137_), .ZN(new_n5138_));
  AOI21_X1   g04134(.A1(new_n5131_), .A2(new_n5132_), .B(new_n5130_), .ZN(new_n5139_));
  NOR3_X1    g04135(.A1(new_n5128_), .A2(new_n5121_), .A3(new_n1576_), .ZN(new_n5140_));
  NOR2_X1    g04136(.A1(new_n5140_), .A2(new_n5139_), .ZN(new_n5141_));
  NOR2_X1    g04137(.A1(new_n5141_), .A2(new_n5138_), .ZN(new_n5142_));
  OAI21_X1   g04138(.A1(new_n5135_), .A2(new_n5142_), .B(new_n5098_), .ZN(new_n5143_));
  AOI21_X1   g04139(.A1(new_n5096_), .A2(new_n5094_), .B(new_n1588_), .ZN(new_n5144_));
  NOR2_X1    g04140(.A1(new_n5134_), .A2(new_n5138_), .ZN(new_n5145_));
  AOI22_X1   g04141(.A1(new_n5129_), .A2(new_n5133_), .B1(new_n5136_), .B2(new_n5137_), .ZN(new_n5146_));
  OAI21_X1   g04142(.A1(new_n5145_), .A2(new_n5146_), .B(new_n5144_), .ZN(new_n5147_));
  AOI21_X1   g04143(.A1(new_n5143_), .A2(new_n5147_), .B(new_n5089_), .ZN(new_n5148_));
  NAND2_X1   g04144(.A1(new_n5079_), .A2(new_n5075_), .ZN(new_n5149_));
  NAND2_X1   g04145(.A1(new_n5063_), .A2(new_n5071_), .ZN(new_n5150_));
  AOI21_X1   g04146(.A1(new_n5149_), .A2(new_n5150_), .B(new_n5085_), .ZN(new_n5151_));
  NAND2_X1   g04147(.A1(new_n5079_), .A2(new_n5063_), .ZN(new_n5152_));
  NAND2_X1   g04148(.A1(new_n5075_), .A2(new_n5071_), .ZN(new_n5153_));
  AOI21_X1   g04149(.A1(new_n5152_), .A2(new_n5153_), .B(new_n5055_), .ZN(new_n5154_));
  NOR2_X1    g04150(.A1(new_n5154_), .A2(new_n5151_), .ZN(new_n5155_));
  NAND2_X1   g04151(.A1(new_n5141_), .A2(new_n5138_), .ZN(new_n5156_));
  NAND2_X1   g04152(.A1(new_n5134_), .A2(new_n5114_), .ZN(new_n5157_));
  AOI21_X1   g04153(.A1(new_n5157_), .A2(new_n5156_), .B(new_n5144_), .ZN(new_n5158_));
  NAND2_X1   g04154(.A1(new_n5141_), .A2(new_n5114_), .ZN(new_n5159_));
  NAND2_X1   g04155(.A1(new_n5134_), .A2(new_n5138_), .ZN(new_n5160_));
  AOI21_X1   g04156(.A1(new_n5159_), .A2(new_n5160_), .B(new_n5098_), .ZN(new_n5161_));
  NOR3_X1    g04157(.A1(new_n5155_), .A2(new_n5161_), .A3(new_n5158_), .ZN(new_n5162_));
  OAI21_X1   g04158(.A1(new_n5148_), .A2(new_n5162_), .B(new_n5052_), .ZN(new_n5163_));
  OAI21_X1   g04159(.A1(new_n1811_), .A2(new_n1724_), .B(new_n1814_), .ZN(new_n5164_));
  NOR3_X1    g04160(.A1(new_n5089_), .A2(new_n5161_), .A3(new_n5158_), .ZN(new_n5165_));
  AOI21_X1   g04161(.A1(new_n5143_), .A2(new_n5147_), .B(new_n5155_), .ZN(new_n5166_));
  OAI21_X1   g04162(.A1(new_n5166_), .A2(new_n5165_), .B(new_n5164_), .ZN(new_n5167_));
  AOI21_X1   g04163(.A1(new_n1362_), .A2(new_n1363_), .B(new_n1361_), .ZN(new_n5168_));
  NOR3_X1    g04164(.A1(new_n1359_), .A2(new_n1349_), .A3(new_n1316_), .ZN(new_n5169_));
  OAI21_X1   g04165(.A1(new_n5168_), .A2(new_n5169_), .B(new_n1290_), .ZN(new_n5170_));
  NOR3_X1    g04166(.A1(new_n5168_), .A2(new_n5169_), .A3(new_n1290_), .ZN(new_n5171_));
  OAI21_X1   g04167(.A1(new_n1175_), .A2(new_n5171_), .B(new_n5170_), .ZN(new_n5172_));
  NOR3_X1    g04168(.A1(new_n1354_), .A2(new_n1357_), .A3(new_n1356_), .ZN(new_n5173_));
  NOR2_X1    g04169(.A1(new_n5173_), .A2(new_n1325_), .ZN(new_n5174_));
  NAND3_X1   g04170(.A1(new_n1315_), .A2(new_n1298_), .A3(new_n1324_), .ZN(new_n5175_));
  OAI21_X1   g04171(.A1(new_n5174_), .A2(new_n5175_), .B(new_n1348_), .ZN(new_n5176_));
  INV_X1     g04172(.I(new_n1346_), .ZN(new_n5177_));
  NAND2_X1   g04173(.A1(new_n1345_), .A2(new_n5177_), .ZN(new_n5178_));
  NOR4_X1    g04174(.A1(new_n5178_), .A2(new_n1331_), .A3(new_n1328_), .A4(new_n1329_), .ZN(new_n5179_));
  NAND2_X1   g04175(.A1(new_n1254_), .A2(new_n1255_), .ZN(new_n5180_));
  NAND3_X1   g04176(.A1(new_n1242_), .A2(new_n1253_), .A3(new_n5180_), .ZN(new_n5181_));
  NAND2_X1   g04177(.A1(new_n5181_), .A2(new_n1329_), .ZN(new_n5182_));
  NOR2_X1    g04178(.A1(new_n1267_), .A2(new_n1277_), .ZN(new_n5183_));
  OAI21_X1   g04179(.A1(new_n1279_), .A2(new_n1281_), .B(new_n5183_), .ZN(new_n5184_));
  NAND2_X1   g04180(.A1(new_n5184_), .A2(new_n1282_), .ZN(new_n5185_));
  XOR2_X1    g04181(.A1(new_n5185_), .A2(new_n5182_), .Z(new_n5186_));
  NAND3_X1   g04182(.A1(new_n1336_), .A2(new_n1334_), .A3(new_n1333_), .ZN(new_n5187_));
  AOI21_X1   g04183(.A1(new_n5187_), .A2(new_n1327_), .B(new_n1356_), .ZN(new_n5188_));
  OAI21_X1   g04184(.A1(new_n5188_), .A2(new_n5179_), .B(new_n5186_), .ZN(new_n5189_));
  NAND3_X1   g04185(.A1(new_n1310_), .A2(new_n1305_), .A3(new_n1318_), .ZN(new_n5190_));
  NAND2_X1   g04186(.A1(new_n5190_), .A2(new_n1229_), .ZN(new_n5191_));
  NAND2_X1   g04187(.A1(new_n1294_), .A2(new_n1292_), .ZN(new_n5192_));
  NOR2_X1    g04188(.A1(new_n1200_), .A2(new_n1202_), .ZN(new_n5193_));
  OAI21_X1   g04189(.A1(new_n5192_), .A2(new_n5193_), .B(new_n1203_), .ZN(new_n5194_));
  XNOR2_X1   g04190(.A1(new_n5194_), .A2(new_n5191_), .ZN(new_n5195_));
  OAI22_X1   g04191(.A1(new_n1297_), .A2(new_n1296_), .B1(new_n1314_), .B2(new_n1299_), .ZN(new_n5196_));
  AOI21_X1   g04192(.A1(new_n1321_), .A2(new_n5196_), .B(new_n5195_), .ZN(new_n5197_));
  NOR2_X1    g04193(.A1(new_n5189_), .A2(new_n5197_), .ZN(new_n5198_));
  INV_X1     g04194(.I(new_n5179_), .ZN(new_n5199_));
  XNOR2_X1   g04195(.A1(new_n5185_), .A2(new_n5182_), .ZN(new_n5200_));
  NOR3_X1    g04196(.A1(new_n1353_), .A2(new_n1350_), .A3(new_n1351_), .ZN(new_n5201_));
  OAI21_X1   g04197(.A1(new_n5201_), .A2(new_n1326_), .B(new_n1344_), .ZN(new_n5202_));
  AOI21_X1   g04198(.A1(new_n5199_), .A2(new_n5202_), .B(new_n5200_), .ZN(new_n5203_));
  XOR2_X1    g04199(.A1(new_n5194_), .A2(new_n5191_), .Z(new_n5204_));
  INV_X1     g04200(.I(new_n5196_), .ZN(new_n5205_));
  OAI21_X1   g04201(.A1(new_n5205_), .A2(new_n1320_), .B(new_n5204_), .ZN(new_n5206_));
  NOR2_X1    g04202(.A1(new_n5203_), .A2(new_n5206_), .ZN(new_n5207_));
  OAI21_X1   g04203(.A1(new_n5207_), .A2(new_n5198_), .B(new_n5176_), .ZN(new_n5208_));
  NAND3_X1   g04204(.A1(new_n1337_), .A2(new_n1344_), .A3(new_n1347_), .ZN(new_n5209_));
  NAND2_X1   g04205(.A1(new_n5209_), .A2(new_n1288_), .ZN(new_n5210_));
  INV_X1     g04206(.I(new_n1298_), .ZN(new_n5211_));
  XNOR2_X1   g04207(.A1(new_n1314_), .A2(new_n1299_), .ZN(new_n5212_));
  NOR3_X1    g04208(.A1(new_n5212_), .A2(new_n5211_), .A3(new_n1323_), .ZN(new_n5213_));
  AOI21_X1   g04209(.A1(new_n5213_), .A2(new_n5210_), .B(new_n1358_), .ZN(new_n5214_));
  NOR2_X1    g04210(.A1(new_n5203_), .A2(new_n5197_), .ZN(new_n5215_));
  NOR2_X1    g04211(.A1(new_n5189_), .A2(new_n5206_), .ZN(new_n5216_));
  OAI21_X1   g04212(.A1(new_n5215_), .A2(new_n5216_), .B(new_n5214_), .ZN(new_n5217_));
  NAND2_X1   g04213(.A1(new_n5217_), .A2(new_n5208_), .ZN(new_n5218_));
  AND2_X2    g04214(.A1(new_n1149_), .A2(new_n1153_), .Z(new_n5219_));
  OAI21_X1   g04215(.A1(new_n1165_), .A2(new_n1166_), .B(new_n1106_), .ZN(new_n5220_));
  NAND3_X1   g04216(.A1(new_n1163_), .A2(new_n1161_), .A3(new_n1157_), .ZN(new_n5221_));
  NAND2_X1   g04217(.A1(new_n5220_), .A2(new_n5221_), .ZN(new_n5222_));
  NAND3_X1   g04218(.A1(new_n5219_), .A2(new_n5222_), .A3(new_n1155_), .ZN(new_n5223_));
  NOR2_X1    g04219(.A1(new_n5223_), .A2(new_n1176_), .ZN(new_n5224_));
  NAND2_X1   g04220(.A1(new_n5223_), .A2(new_n1176_), .ZN(new_n5225_));
  NAND2_X1   g04221(.A1(new_n1074_), .A2(new_n1022_), .ZN(new_n5226_));
  NAND2_X1   g04222(.A1(new_n1072_), .A2(new_n1071_), .ZN(new_n5227_));
  NAND2_X1   g04223(.A1(new_n5227_), .A2(new_n5226_), .ZN(new_n5228_));
  NOR4_X1    g04224(.A1(new_n5228_), .A2(new_n1077_), .A3(new_n1056_), .A4(new_n1080_), .ZN(new_n5229_));
  AOI21_X1   g04225(.A1(new_n5225_), .A2(new_n5229_), .B(new_n5224_), .ZN(new_n5230_));
  NAND2_X1   g04226(.A1(new_n1154_), .A2(new_n1171_), .ZN(new_n5231_));
  NAND2_X1   g04227(.A1(new_n1150_), .A2(new_n1146_), .ZN(new_n5232_));
  OAI21_X1   g04228(.A1(new_n5232_), .A2(new_n1169_), .B(new_n1138_), .ZN(new_n5233_));
  NAND2_X1   g04229(.A1(new_n1158_), .A2(new_n1159_), .ZN(new_n5234_));
  NAND3_X1   g04230(.A1(new_n1162_), .A2(new_n1157_), .A3(new_n5234_), .ZN(new_n5235_));
  NAND2_X1   g04231(.A1(new_n5235_), .A2(new_n1111_), .ZN(new_n5236_));
  XNOR2_X1   g04232(.A1(new_n5236_), .A2(new_n5233_), .ZN(new_n5237_));
  OAI21_X1   g04233(.A1(new_n1154_), .A2(new_n1156_), .B(new_n5222_), .ZN(new_n5238_));
  AOI21_X1   g04234(.A1(new_n5231_), .A2(new_n5238_), .B(new_n5237_), .ZN(new_n5239_));
  NAND2_X1   g04235(.A1(new_n1080_), .A2(new_n1070_), .ZN(new_n5240_));
  INV_X1     g04236(.I(new_n5240_), .ZN(new_n5241_));
  NAND3_X1   g04237(.A1(new_n1063_), .A2(new_n1057_), .A3(new_n1068_), .ZN(new_n5242_));
  NAND2_X1   g04238(.A1(new_n5242_), .A2(new_n1054_), .ZN(new_n5243_));
  NOR2_X1    g04239(.A1(new_n1012_), .A2(new_n1022_), .ZN(new_n5244_));
  INV_X1     g04240(.I(new_n1027_), .ZN(new_n5245_));
  NAND4_X1   g04241(.A1(new_n1023_), .A2(new_n1025_), .A3(new_n1010_), .A4(new_n1020_), .ZN(new_n5246_));
  AOI21_X1   g04242(.A1(new_n5244_), .A2(new_n5246_), .B(new_n5245_), .ZN(new_n5247_));
  XNOR2_X1   g04243(.A1(new_n5243_), .A2(new_n5247_), .ZN(new_n5248_));
  OAI22_X1   g04244(.A1(new_n1080_), .A2(new_n1079_), .B1(new_n1073_), .B2(new_n1075_), .ZN(new_n5249_));
  INV_X1     g04245(.I(new_n5249_), .ZN(new_n5250_));
  OAI21_X1   g04246(.A1(new_n5250_), .A2(new_n5241_), .B(new_n5248_), .ZN(new_n5251_));
  NAND2_X1   g04247(.A1(new_n5251_), .A2(new_n5239_), .ZN(new_n5252_));
  INV_X1     g04248(.I(new_n5231_), .ZN(new_n5253_));
  XOR2_X1    g04249(.A1(new_n5236_), .A2(new_n5233_), .Z(new_n5254_));
  AOI21_X1   g04250(.A1(new_n5219_), .A2(new_n1155_), .B(new_n1168_), .ZN(new_n5255_));
  OAI21_X1   g04251(.A1(new_n5255_), .A2(new_n5253_), .B(new_n5254_), .ZN(new_n5256_));
  XOR2_X1    g04252(.A1(new_n5243_), .A2(new_n5247_), .Z(new_n5257_));
  AOI21_X1   g04253(.A1(new_n5240_), .A2(new_n5249_), .B(new_n5257_), .ZN(new_n5258_));
  NAND2_X1   g04254(.A1(new_n5256_), .A2(new_n5258_), .ZN(new_n5259_));
  AOI21_X1   g04255(.A1(new_n5252_), .A2(new_n5259_), .B(new_n5230_), .ZN(new_n5260_));
  NAND2_X1   g04256(.A1(new_n5225_), .A2(new_n5229_), .ZN(new_n5261_));
  NAND2_X1   g04257(.A1(new_n5261_), .A2(new_n1173_), .ZN(new_n5262_));
  NAND2_X1   g04258(.A1(new_n5251_), .A2(new_n5256_), .ZN(new_n5263_));
  NAND2_X1   g04259(.A1(new_n5239_), .A2(new_n5258_), .ZN(new_n5264_));
  AOI21_X1   g04260(.A1(new_n5263_), .A2(new_n5264_), .B(new_n5262_), .ZN(new_n5265_));
  NOR2_X1    g04261(.A1(new_n5265_), .A2(new_n5260_), .ZN(new_n5266_));
  NOR2_X1    g04262(.A1(new_n5218_), .A2(new_n5266_), .ZN(new_n5267_));
  NAND2_X1   g04263(.A1(new_n5203_), .A2(new_n5206_), .ZN(new_n5268_));
  NAND2_X1   g04264(.A1(new_n5189_), .A2(new_n5197_), .ZN(new_n5269_));
  AOI21_X1   g04265(.A1(new_n5268_), .A2(new_n5269_), .B(new_n5214_), .ZN(new_n5270_));
  NAND2_X1   g04266(.A1(new_n5189_), .A2(new_n5206_), .ZN(new_n5271_));
  NAND2_X1   g04267(.A1(new_n5203_), .A2(new_n5197_), .ZN(new_n5272_));
  AOI21_X1   g04268(.A1(new_n5272_), .A2(new_n5271_), .B(new_n5176_), .ZN(new_n5273_));
  NOR2_X1    g04269(.A1(new_n5270_), .A2(new_n5273_), .ZN(new_n5274_));
  NOR2_X1    g04270(.A1(new_n5256_), .A2(new_n5258_), .ZN(new_n5275_));
  NOR2_X1    g04271(.A1(new_n5251_), .A2(new_n5239_), .ZN(new_n5276_));
  OAI21_X1   g04272(.A1(new_n5276_), .A2(new_n5275_), .B(new_n5262_), .ZN(new_n5277_));
  NOR2_X1    g04273(.A1(new_n5239_), .A2(new_n5258_), .ZN(new_n5278_));
  NOR2_X1    g04274(.A1(new_n5251_), .A2(new_n5256_), .ZN(new_n5279_));
  OAI21_X1   g04275(.A1(new_n5279_), .A2(new_n5278_), .B(new_n5230_), .ZN(new_n5280_));
  NAND2_X1   g04276(.A1(new_n5277_), .A2(new_n5280_), .ZN(new_n5281_));
  NOR2_X1    g04277(.A1(new_n5274_), .A2(new_n5281_), .ZN(new_n5282_));
  OAI21_X1   g04278(.A1(new_n5282_), .A2(new_n5267_), .B(new_n5172_), .ZN(new_n5283_));
  XOR2_X1    g04279(.A1(new_n1084_), .A2(new_n5224_), .Z(new_n5284_));
  NOR3_X1    g04280(.A1(new_n5284_), .A2(new_n1056_), .A3(new_n1077_), .ZN(new_n5285_));
  NAND3_X1   g04281(.A1(new_n1364_), .A2(new_n1360_), .A3(new_n1291_), .ZN(new_n5286_));
  AOI21_X1   g04282(.A1(new_n5285_), .A2(new_n5286_), .B(new_n1365_), .ZN(new_n5287_));
  NOR2_X1    g04283(.A1(new_n5274_), .A2(new_n5266_), .ZN(new_n5288_));
  NOR3_X1    g04284(.A1(new_n5281_), .A2(new_n5270_), .A3(new_n5273_), .ZN(new_n5289_));
  OAI21_X1   g04285(.A1(new_n5288_), .A2(new_n5289_), .B(new_n5287_), .ZN(new_n5290_));
  NAND2_X1   g04286(.A1(new_n5283_), .A2(new_n5290_), .ZN(new_n5291_));
  NAND3_X1   g04287(.A1(new_n5291_), .A2(new_n5163_), .A3(new_n5167_), .ZN(new_n5292_));
  OAI21_X1   g04288(.A1(new_n5158_), .A2(new_n5161_), .B(new_n5155_), .ZN(new_n5293_));
  NAND3_X1   g04289(.A1(new_n5089_), .A2(new_n5143_), .A3(new_n5147_), .ZN(new_n5294_));
  AOI21_X1   g04290(.A1(new_n5293_), .A2(new_n5294_), .B(new_n5164_), .ZN(new_n5295_));
  NAND3_X1   g04291(.A1(new_n5155_), .A2(new_n5143_), .A3(new_n5147_), .ZN(new_n5296_));
  OAI21_X1   g04292(.A1(new_n5158_), .A2(new_n5161_), .B(new_n5089_), .ZN(new_n5297_));
  AOI21_X1   g04293(.A1(new_n5297_), .A2(new_n5296_), .B(new_n5052_), .ZN(new_n5298_));
  NAND2_X1   g04294(.A1(new_n5274_), .A2(new_n5281_), .ZN(new_n5299_));
  NAND2_X1   g04295(.A1(new_n5218_), .A2(new_n5266_), .ZN(new_n5300_));
  AOI21_X1   g04296(.A1(new_n5299_), .A2(new_n5300_), .B(new_n5287_), .ZN(new_n5301_));
  OAI22_X1   g04297(.A1(new_n5270_), .A2(new_n5273_), .B1(new_n5265_), .B2(new_n5260_), .ZN(new_n5302_));
  NAND2_X1   g04298(.A1(new_n5274_), .A2(new_n5266_), .ZN(new_n5303_));
  AOI21_X1   g04299(.A1(new_n5303_), .A2(new_n5302_), .B(new_n5172_), .ZN(new_n5304_));
  NOR2_X1    g04300(.A1(new_n5301_), .A2(new_n5304_), .ZN(new_n5305_));
  OAI21_X1   g04301(.A1(new_n5295_), .A2(new_n5298_), .B(new_n5305_), .ZN(new_n5306_));
  AOI21_X1   g04302(.A1(new_n5306_), .A2(new_n5292_), .B(new_n5047_), .ZN(new_n5307_));
  INV_X1     g04303(.I(new_n1823_), .ZN(new_n5308_));
  NAND2_X1   g04304(.A1(new_n5046_), .A2(new_n5045_), .ZN(new_n5309_));
  NAND2_X1   g04305(.A1(new_n5309_), .A2(new_n5308_), .ZN(new_n5310_));
  NAND3_X1   g04306(.A1(new_n5305_), .A2(new_n5163_), .A3(new_n5167_), .ZN(new_n5311_));
  OAI21_X1   g04307(.A1(new_n5295_), .A2(new_n5298_), .B(new_n5291_), .ZN(new_n5312_));
  AOI21_X1   g04308(.A1(new_n5312_), .A2(new_n5311_), .B(new_n5310_), .ZN(new_n5313_));
  NOR2_X1    g04309(.A1(new_n5313_), .A2(new_n5307_), .ZN(new_n5314_));
  NOR2_X1    g04310(.A1(new_n5314_), .A2(new_n5044_), .ZN(new_n5315_));
  NAND3_X1   g04311(.A1(new_n5037_), .A2(new_n5030_), .A3(new_n5027_), .ZN(new_n5316_));
  OAI21_X1   g04312(.A1(new_n4902_), .A2(new_n4910_), .B(new_n5023_), .ZN(new_n5317_));
  AOI21_X1   g04313(.A1(new_n5317_), .A2(new_n5316_), .B(new_n5040_), .ZN(new_n5318_));
  OAI22_X1   g04314(.A1(new_n4910_), .A2(new_n4902_), .B1(new_n5014_), .B2(new_n5022_), .ZN(new_n5319_));
  NAND3_X1   g04315(.A1(new_n5023_), .A2(new_n5027_), .A3(new_n5030_), .ZN(new_n5320_));
  AOI21_X1   g04316(.A1(new_n5320_), .A2(new_n5319_), .B(new_n4797_), .ZN(new_n5321_));
  NOR2_X1    g04317(.A1(new_n5318_), .A2(new_n5321_), .ZN(new_n5322_));
  NOR3_X1    g04318(.A1(new_n5305_), .A2(new_n5295_), .A3(new_n5298_), .ZN(new_n5323_));
  AOI21_X1   g04319(.A1(new_n5163_), .A2(new_n5167_), .B(new_n5291_), .ZN(new_n5324_));
  OAI21_X1   g04320(.A1(new_n5324_), .A2(new_n5323_), .B(new_n5310_), .ZN(new_n5325_));
  NOR3_X1    g04321(.A1(new_n5291_), .A2(new_n5295_), .A3(new_n5298_), .ZN(new_n5326_));
  AOI21_X1   g04322(.A1(new_n5163_), .A2(new_n5167_), .B(new_n5305_), .ZN(new_n5327_));
  OAI21_X1   g04323(.A1(new_n5327_), .A2(new_n5326_), .B(new_n5047_), .ZN(new_n5328_));
  NAND2_X1   g04324(.A1(new_n5325_), .A2(new_n5328_), .ZN(new_n5329_));
  NOR2_X1    g04325(.A1(new_n5329_), .A2(new_n5322_), .ZN(new_n5330_));
  OAI21_X1   g04326(.A1(new_n5315_), .A2(new_n5330_), .B(new_n4793_), .ZN(new_n5331_));
  INV_X1     g04327(.I(new_n4793_), .ZN(new_n5332_));
  NOR3_X1    g04328(.A1(new_n5044_), .A2(new_n5307_), .A3(new_n5313_), .ZN(new_n5333_));
  NOR2_X1    g04329(.A1(new_n5314_), .A2(new_n5322_), .ZN(new_n5334_));
  OAI21_X1   g04330(.A1(new_n5334_), .A2(new_n5333_), .B(new_n5332_), .ZN(new_n5335_));
  NAND2_X1   g04331(.A1(new_n5331_), .A2(new_n5335_), .ZN(new_n5336_));
  NAND2_X1   g04332(.A1(new_n4790_), .A2(new_n5336_), .ZN(new_n5337_));
  NAND2_X1   g04333(.A1(new_n5329_), .A2(new_n5322_), .ZN(new_n5338_));
  NAND3_X1   g04334(.A1(new_n5044_), .A2(new_n5325_), .A3(new_n5328_), .ZN(new_n5339_));
  AOI21_X1   g04335(.A1(new_n5338_), .A2(new_n5339_), .B(new_n5332_), .ZN(new_n5340_));
  NAND4_X1   g04336(.A1(new_n5325_), .A2(new_n5328_), .A3(new_n5039_), .A4(new_n5043_), .ZN(new_n5341_));
  OAI22_X1   g04337(.A1(new_n5313_), .A2(new_n5307_), .B1(new_n5318_), .B2(new_n5321_), .ZN(new_n5342_));
  AOI21_X1   g04338(.A1(new_n5342_), .A2(new_n5341_), .B(new_n4793_), .ZN(new_n5343_));
  NOR2_X1    g04339(.A1(new_n5340_), .A2(new_n5343_), .ZN(new_n5344_));
  OAI21_X1   g04340(.A1(new_n4780_), .A2(new_n4789_), .B(new_n5344_), .ZN(new_n5345_));
  AOI21_X1   g04341(.A1(new_n5345_), .A2(new_n5337_), .B(new_n4270_), .ZN(new_n5346_));
  INV_X1     g04342(.I(new_n4270_), .ZN(new_n5347_));
  NOR4_X1    g04343(.A1(new_n4780_), .A2(new_n4789_), .A3(new_n5340_), .A4(new_n5343_), .ZN(new_n5348_));
  INV_X1     g04344(.I(new_n5348_), .ZN(new_n5349_));
  OAI22_X1   g04345(.A1(new_n4780_), .A2(new_n4789_), .B1(new_n5340_), .B2(new_n5343_), .ZN(new_n5350_));
  AOI21_X1   g04346(.A1(new_n5349_), .A2(new_n5350_), .B(new_n5347_), .ZN(new_n5351_));
  NOR2_X1    g04347(.A1(new_n5351_), .A2(new_n5346_), .ZN(new_n5352_));
  INV_X1     g04348(.I(\A[939] ), .ZN(new_n5353_));
  NOR2_X1    g04349(.A1(new_n5353_), .A2(\A[938] ), .ZN(new_n5354_));
  INV_X1     g04350(.I(\A[938] ), .ZN(new_n5355_));
  NOR2_X1    g04351(.A1(new_n5355_), .A2(\A[939] ), .ZN(new_n5356_));
  OAI21_X1   g04352(.A1(new_n5354_), .A2(new_n5356_), .B(\A[937] ), .ZN(new_n5357_));
  INV_X1     g04353(.I(\A[937] ), .ZN(new_n5358_));
  NOR2_X1    g04354(.A1(\A[938] ), .A2(\A[939] ), .ZN(new_n5359_));
  NOR2_X1    g04355(.A1(new_n5355_), .A2(new_n5353_), .ZN(new_n5360_));
  OAI21_X1   g04356(.A1(new_n5360_), .A2(new_n5359_), .B(new_n5358_), .ZN(new_n5361_));
  NAND2_X1   g04357(.A1(new_n5361_), .A2(new_n5357_), .ZN(new_n5362_));
  INV_X1     g04358(.I(\A[942] ), .ZN(new_n5363_));
  NOR2_X1    g04359(.A1(new_n5363_), .A2(\A[941] ), .ZN(new_n5364_));
  INV_X1     g04360(.I(\A[941] ), .ZN(new_n5365_));
  NOR2_X1    g04361(.A1(new_n5365_), .A2(\A[942] ), .ZN(new_n5366_));
  OAI21_X1   g04362(.A1(new_n5364_), .A2(new_n5366_), .B(\A[940] ), .ZN(new_n5367_));
  INV_X1     g04363(.I(\A[940] ), .ZN(new_n5368_));
  NOR2_X1    g04364(.A1(new_n5365_), .A2(new_n5363_), .ZN(new_n5369_));
  NOR2_X1    g04365(.A1(\A[941] ), .A2(\A[942] ), .ZN(new_n5370_));
  OAI21_X1   g04366(.A1(new_n5369_), .A2(new_n5370_), .B(new_n5368_), .ZN(new_n5371_));
  NAND2_X1   g04367(.A1(new_n5371_), .A2(new_n5367_), .ZN(new_n5372_));
  INV_X1     g04368(.I(new_n5359_), .ZN(new_n5373_));
  OAI21_X1   g04369(.A1(\A[937] ), .A2(new_n5360_), .B(new_n5373_), .ZN(new_n5374_));
  INV_X1     g04370(.I(new_n5370_), .ZN(new_n5375_));
  OAI21_X1   g04371(.A1(\A[940] ), .A2(new_n5369_), .B(new_n5375_), .ZN(new_n5376_));
  NAND2_X1   g04372(.A1(new_n5374_), .A2(new_n5376_), .ZN(new_n5377_));
  INV_X1     g04373(.I(new_n5377_), .ZN(new_n5378_));
  NAND3_X1   g04374(.A1(new_n5378_), .A2(new_n5362_), .A3(new_n5372_), .ZN(new_n5379_));
  INV_X1     g04375(.I(\A[931] ), .ZN(new_n5380_));
  INV_X1     g04376(.I(\A[932] ), .ZN(new_n5381_));
  NAND2_X1   g04377(.A1(new_n5381_), .A2(\A[933] ), .ZN(new_n5382_));
  INV_X1     g04378(.I(\A[933] ), .ZN(new_n5383_));
  NAND2_X1   g04379(.A1(new_n5383_), .A2(\A[932] ), .ZN(new_n5384_));
  AOI21_X1   g04380(.A1(new_n5382_), .A2(new_n5384_), .B(new_n5380_), .ZN(new_n5385_));
  NAND2_X1   g04381(.A1(new_n5381_), .A2(new_n5383_), .ZN(new_n5386_));
  NAND2_X1   g04382(.A1(\A[932] ), .A2(\A[933] ), .ZN(new_n5387_));
  AOI21_X1   g04383(.A1(new_n5386_), .A2(new_n5387_), .B(\A[931] ), .ZN(new_n5388_));
  NOR2_X1    g04384(.A1(new_n5388_), .A2(new_n5385_), .ZN(new_n5389_));
  INV_X1     g04385(.I(\A[934] ), .ZN(new_n5390_));
  INV_X1     g04386(.I(\A[935] ), .ZN(new_n5391_));
  NAND2_X1   g04387(.A1(new_n5391_), .A2(\A[936] ), .ZN(new_n5392_));
  INV_X1     g04388(.I(\A[936] ), .ZN(new_n5393_));
  NAND2_X1   g04389(.A1(new_n5393_), .A2(\A[935] ), .ZN(new_n5394_));
  AOI21_X1   g04390(.A1(new_n5392_), .A2(new_n5394_), .B(new_n5390_), .ZN(new_n5395_));
  NAND2_X1   g04391(.A1(\A[935] ), .A2(\A[936] ), .ZN(new_n5396_));
  NAND2_X1   g04392(.A1(new_n5391_), .A2(new_n5393_), .ZN(new_n5397_));
  AOI21_X1   g04393(.A1(new_n5397_), .A2(new_n5396_), .B(\A[934] ), .ZN(new_n5398_));
  NOR2_X1    g04394(.A1(new_n5398_), .A2(new_n5395_), .ZN(new_n5399_));
  NAND2_X1   g04395(.A1(new_n5387_), .A2(new_n5380_), .ZN(new_n5400_));
  NAND2_X1   g04396(.A1(new_n5400_), .A2(new_n5386_), .ZN(new_n5401_));
  NAND2_X1   g04397(.A1(new_n5396_), .A2(new_n5390_), .ZN(new_n5402_));
  NAND2_X1   g04398(.A1(new_n5402_), .A2(new_n5397_), .ZN(new_n5403_));
  NAND2_X1   g04399(.A1(new_n5401_), .A2(new_n5403_), .ZN(new_n5404_));
  NOR3_X1    g04400(.A1(new_n5389_), .A2(new_n5399_), .A3(new_n5404_), .ZN(new_n5405_));
  XOR2_X1    g04401(.A1(new_n5379_), .A2(new_n5405_), .Z(new_n5406_));
  INV_X1     g04402(.I(\A[927] ), .ZN(new_n5407_));
  NOR2_X1    g04403(.A1(new_n5407_), .A2(\A[926] ), .ZN(new_n5408_));
  INV_X1     g04404(.I(\A[926] ), .ZN(new_n5409_));
  NOR2_X1    g04405(.A1(new_n5409_), .A2(\A[927] ), .ZN(new_n5410_));
  OAI21_X1   g04406(.A1(new_n5408_), .A2(new_n5410_), .B(\A[925] ), .ZN(new_n5411_));
  INV_X1     g04407(.I(\A[925] ), .ZN(new_n5412_));
  NOR2_X1    g04408(.A1(new_n5409_), .A2(new_n5407_), .ZN(new_n5413_));
  NOR2_X1    g04409(.A1(\A[926] ), .A2(\A[927] ), .ZN(new_n5414_));
  OAI21_X1   g04410(.A1(new_n5413_), .A2(new_n5414_), .B(new_n5412_), .ZN(new_n5415_));
  NAND2_X1   g04411(.A1(new_n5415_), .A2(new_n5411_), .ZN(new_n5416_));
  INV_X1     g04412(.I(\A[930] ), .ZN(new_n5417_));
  NOR2_X1    g04413(.A1(new_n5417_), .A2(\A[929] ), .ZN(new_n5418_));
  INV_X1     g04414(.I(\A[929] ), .ZN(new_n5419_));
  NOR2_X1    g04415(.A1(new_n5419_), .A2(\A[930] ), .ZN(new_n5420_));
  OAI21_X1   g04416(.A1(new_n5418_), .A2(new_n5420_), .B(\A[928] ), .ZN(new_n5421_));
  INV_X1     g04417(.I(\A[928] ), .ZN(new_n5422_));
  NOR2_X1    g04418(.A1(new_n5419_), .A2(new_n5417_), .ZN(new_n5423_));
  NOR2_X1    g04419(.A1(\A[929] ), .A2(\A[930] ), .ZN(new_n5424_));
  OAI21_X1   g04420(.A1(new_n5423_), .A2(new_n5424_), .B(new_n5422_), .ZN(new_n5425_));
  NAND2_X1   g04421(.A1(new_n5425_), .A2(new_n5421_), .ZN(new_n5426_));
  INV_X1     g04422(.I(new_n5414_), .ZN(new_n5427_));
  OAI21_X1   g04423(.A1(\A[925] ), .A2(new_n5413_), .B(new_n5427_), .ZN(new_n5428_));
  INV_X1     g04424(.I(new_n5424_), .ZN(new_n5429_));
  OAI21_X1   g04425(.A1(\A[928] ), .A2(new_n5423_), .B(new_n5429_), .ZN(new_n5430_));
  NAND2_X1   g04426(.A1(new_n5428_), .A2(new_n5430_), .ZN(new_n5431_));
  INV_X1     g04427(.I(new_n5431_), .ZN(new_n5432_));
  NAND3_X1   g04428(.A1(new_n5432_), .A2(new_n5416_), .A3(new_n5426_), .ZN(new_n5433_));
  INV_X1     g04429(.I(\A[919] ), .ZN(new_n5434_));
  INV_X1     g04430(.I(\A[920] ), .ZN(new_n5435_));
  NAND2_X1   g04431(.A1(new_n5435_), .A2(\A[921] ), .ZN(new_n5436_));
  INV_X1     g04432(.I(\A[921] ), .ZN(new_n5437_));
  NAND2_X1   g04433(.A1(new_n5437_), .A2(\A[920] ), .ZN(new_n5438_));
  AOI21_X1   g04434(.A1(new_n5436_), .A2(new_n5438_), .B(new_n5434_), .ZN(new_n5439_));
  NAND2_X1   g04435(.A1(\A[920] ), .A2(\A[921] ), .ZN(new_n5440_));
  NAND2_X1   g04436(.A1(new_n5435_), .A2(new_n5437_), .ZN(new_n5441_));
  AOI21_X1   g04437(.A1(new_n5441_), .A2(new_n5440_), .B(\A[919] ), .ZN(new_n5442_));
  NOR2_X1    g04438(.A1(new_n5442_), .A2(new_n5439_), .ZN(new_n5443_));
  INV_X1     g04439(.I(\A[922] ), .ZN(new_n5444_));
  INV_X1     g04440(.I(\A[923] ), .ZN(new_n5445_));
  NAND2_X1   g04441(.A1(new_n5445_), .A2(\A[924] ), .ZN(new_n5446_));
  INV_X1     g04442(.I(\A[924] ), .ZN(new_n5447_));
  NAND2_X1   g04443(.A1(new_n5447_), .A2(\A[923] ), .ZN(new_n5448_));
  AOI21_X1   g04444(.A1(new_n5446_), .A2(new_n5448_), .B(new_n5444_), .ZN(new_n5449_));
  NAND2_X1   g04445(.A1(\A[923] ), .A2(\A[924] ), .ZN(new_n5450_));
  NAND2_X1   g04446(.A1(new_n5445_), .A2(new_n5447_), .ZN(new_n5451_));
  AOI21_X1   g04447(.A1(new_n5451_), .A2(new_n5450_), .B(\A[922] ), .ZN(new_n5452_));
  NOR2_X1    g04448(.A1(new_n5452_), .A2(new_n5449_), .ZN(new_n5453_));
  NAND2_X1   g04449(.A1(new_n5440_), .A2(new_n5434_), .ZN(new_n5454_));
  NAND2_X1   g04450(.A1(new_n5454_), .A2(new_n5441_), .ZN(new_n5455_));
  NAND2_X1   g04451(.A1(new_n5450_), .A2(new_n5444_), .ZN(new_n5456_));
  NAND2_X1   g04452(.A1(new_n5456_), .A2(new_n5451_), .ZN(new_n5457_));
  NAND2_X1   g04453(.A1(new_n5455_), .A2(new_n5457_), .ZN(new_n5458_));
  NOR3_X1    g04454(.A1(new_n5443_), .A2(new_n5453_), .A3(new_n5458_), .ZN(new_n5459_));
  XOR2_X1    g04455(.A1(new_n5433_), .A2(new_n5459_), .Z(new_n5460_));
  XNOR2_X1   g04456(.A1(new_n5406_), .A2(new_n5460_), .ZN(new_n5461_));
  INV_X1     g04457(.I(\A[915] ), .ZN(new_n5462_));
  NOR2_X1    g04458(.A1(new_n5462_), .A2(\A[914] ), .ZN(new_n5463_));
  INV_X1     g04459(.I(\A[914] ), .ZN(new_n5464_));
  NOR2_X1    g04460(.A1(new_n5464_), .A2(\A[915] ), .ZN(new_n5465_));
  OAI21_X1   g04461(.A1(new_n5463_), .A2(new_n5465_), .B(\A[913] ), .ZN(new_n5466_));
  INV_X1     g04462(.I(\A[913] ), .ZN(new_n5467_));
  NOR2_X1    g04463(.A1(\A[914] ), .A2(\A[915] ), .ZN(new_n5468_));
  NOR2_X1    g04464(.A1(new_n5464_), .A2(new_n5462_), .ZN(new_n5469_));
  OAI21_X1   g04465(.A1(new_n5469_), .A2(new_n5468_), .B(new_n5467_), .ZN(new_n5470_));
  NAND2_X1   g04466(.A1(new_n5470_), .A2(new_n5466_), .ZN(new_n5471_));
  INV_X1     g04467(.I(\A[918] ), .ZN(new_n5472_));
  NOR2_X1    g04468(.A1(new_n5472_), .A2(\A[917] ), .ZN(new_n5473_));
  INV_X1     g04469(.I(\A[917] ), .ZN(new_n5474_));
  NOR2_X1    g04470(.A1(new_n5474_), .A2(\A[918] ), .ZN(new_n5475_));
  OAI21_X1   g04471(.A1(new_n5473_), .A2(new_n5475_), .B(\A[916] ), .ZN(new_n5476_));
  INV_X1     g04472(.I(\A[916] ), .ZN(new_n5477_));
  NOR2_X1    g04473(.A1(new_n5474_), .A2(new_n5472_), .ZN(new_n5478_));
  NOR2_X1    g04474(.A1(\A[917] ), .A2(\A[918] ), .ZN(new_n5479_));
  OAI21_X1   g04475(.A1(new_n5478_), .A2(new_n5479_), .B(new_n5477_), .ZN(new_n5480_));
  NAND2_X1   g04476(.A1(new_n5480_), .A2(new_n5476_), .ZN(new_n5481_));
  INV_X1     g04477(.I(new_n5468_), .ZN(new_n5482_));
  OAI21_X1   g04478(.A1(\A[913] ), .A2(new_n5469_), .B(new_n5482_), .ZN(new_n5483_));
  INV_X1     g04479(.I(new_n5479_), .ZN(new_n5484_));
  OAI21_X1   g04480(.A1(\A[916] ), .A2(new_n5478_), .B(new_n5484_), .ZN(new_n5485_));
  NAND2_X1   g04481(.A1(new_n5483_), .A2(new_n5485_), .ZN(new_n5486_));
  INV_X1     g04482(.I(new_n5486_), .ZN(new_n5487_));
  NAND3_X1   g04483(.A1(new_n5487_), .A2(new_n5471_), .A3(new_n5481_), .ZN(new_n5488_));
  INV_X1     g04484(.I(\A[907] ), .ZN(new_n5489_));
  INV_X1     g04485(.I(\A[908] ), .ZN(new_n5490_));
  NAND2_X1   g04486(.A1(new_n5490_), .A2(\A[909] ), .ZN(new_n5491_));
  INV_X1     g04487(.I(\A[909] ), .ZN(new_n5492_));
  NAND2_X1   g04488(.A1(new_n5492_), .A2(\A[908] ), .ZN(new_n5493_));
  AOI21_X1   g04489(.A1(new_n5491_), .A2(new_n5493_), .B(new_n5489_), .ZN(new_n5494_));
  NAND2_X1   g04490(.A1(new_n5490_), .A2(new_n5492_), .ZN(new_n5495_));
  NAND2_X1   g04491(.A1(\A[908] ), .A2(\A[909] ), .ZN(new_n5496_));
  AOI21_X1   g04492(.A1(new_n5495_), .A2(new_n5496_), .B(\A[907] ), .ZN(new_n5497_));
  NOR2_X1    g04493(.A1(new_n5497_), .A2(new_n5494_), .ZN(new_n5498_));
  INV_X1     g04494(.I(\A[910] ), .ZN(new_n5499_));
  INV_X1     g04495(.I(\A[911] ), .ZN(new_n5500_));
  NAND2_X1   g04496(.A1(new_n5500_), .A2(\A[912] ), .ZN(new_n5501_));
  INV_X1     g04497(.I(\A[912] ), .ZN(new_n5502_));
  NAND2_X1   g04498(.A1(new_n5502_), .A2(\A[911] ), .ZN(new_n5503_));
  AOI21_X1   g04499(.A1(new_n5501_), .A2(new_n5503_), .B(new_n5499_), .ZN(new_n5504_));
  NAND2_X1   g04500(.A1(\A[911] ), .A2(\A[912] ), .ZN(new_n5505_));
  NAND2_X1   g04501(.A1(new_n5500_), .A2(new_n5502_), .ZN(new_n5506_));
  AOI21_X1   g04502(.A1(new_n5506_), .A2(new_n5505_), .B(\A[910] ), .ZN(new_n5507_));
  NOR2_X1    g04503(.A1(new_n5507_), .A2(new_n5504_), .ZN(new_n5508_));
  NAND2_X1   g04504(.A1(new_n5496_), .A2(new_n5489_), .ZN(new_n5509_));
  NAND2_X1   g04505(.A1(new_n5509_), .A2(new_n5495_), .ZN(new_n5510_));
  NAND2_X1   g04506(.A1(new_n5505_), .A2(new_n5499_), .ZN(new_n5511_));
  NAND2_X1   g04507(.A1(new_n5511_), .A2(new_n5506_), .ZN(new_n5512_));
  NAND2_X1   g04508(.A1(new_n5510_), .A2(new_n5512_), .ZN(new_n5513_));
  NOR3_X1    g04509(.A1(new_n5498_), .A2(new_n5508_), .A3(new_n5513_), .ZN(new_n5514_));
  XOR2_X1    g04510(.A1(new_n5488_), .A2(new_n5514_), .Z(new_n5515_));
  INV_X1     g04511(.I(\A[903] ), .ZN(new_n5516_));
  NOR2_X1    g04512(.A1(new_n5516_), .A2(\A[902] ), .ZN(new_n5517_));
  INV_X1     g04513(.I(\A[902] ), .ZN(new_n5518_));
  NOR2_X1    g04514(.A1(new_n5518_), .A2(\A[903] ), .ZN(new_n5519_));
  OAI21_X1   g04515(.A1(new_n5517_), .A2(new_n5519_), .B(\A[901] ), .ZN(new_n5520_));
  INV_X1     g04516(.I(\A[901] ), .ZN(new_n5521_));
  NOR2_X1    g04517(.A1(\A[902] ), .A2(\A[903] ), .ZN(new_n5522_));
  NOR2_X1    g04518(.A1(new_n5518_), .A2(new_n5516_), .ZN(new_n5523_));
  OAI21_X1   g04519(.A1(new_n5523_), .A2(new_n5522_), .B(new_n5521_), .ZN(new_n5524_));
  NAND2_X1   g04520(.A1(new_n5524_), .A2(new_n5520_), .ZN(new_n5525_));
  INV_X1     g04521(.I(\A[906] ), .ZN(new_n5526_));
  NOR2_X1    g04522(.A1(new_n5526_), .A2(\A[905] ), .ZN(new_n5527_));
  INV_X1     g04523(.I(\A[905] ), .ZN(new_n5528_));
  NOR2_X1    g04524(.A1(new_n5528_), .A2(\A[906] ), .ZN(new_n5529_));
  OAI21_X1   g04525(.A1(new_n5527_), .A2(new_n5529_), .B(\A[904] ), .ZN(new_n5530_));
  INV_X1     g04526(.I(\A[904] ), .ZN(new_n5531_));
  NOR2_X1    g04527(.A1(\A[905] ), .A2(\A[906] ), .ZN(new_n5532_));
  NOR2_X1    g04528(.A1(new_n5528_), .A2(new_n5526_), .ZN(new_n5533_));
  OAI21_X1   g04529(.A1(new_n5533_), .A2(new_n5532_), .B(new_n5531_), .ZN(new_n5534_));
  NAND2_X1   g04530(.A1(new_n5534_), .A2(new_n5530_), .ZN(new_n5535_));
  INV_X1     g04531(.I(new_n5522_), .ZN(new_n5536_));
  OAI21_X1   g04532(.A1(\A[901] ), .A2(new_n5523_), .B(new_n5536_), .ZN(new_n5537_));
  INV_X1     g04533(.I(new_n5532_), .ZN(new_n5538_));
  OAI21_X1   g04534(.A1(\A[904] ), .A2(new_n5533_), .B(new_n5538_), .ZN(new_n5539_));
  NAND2_X1   g04535(.A1(new_n5537_), .A2(new_n5539_), .ZN(new_n5540_));
  INV_X1     g04536(.I(new_n5540_), .ZN(new_n5541_));
  NAND3_X1   g04537(.A1(new_n5541_), .A2(new_n5525_), .A3(new_n5535_), .ZN(new_n5542_));
  INV_X1     g04538(.I(\A[895] ), .ZN(new_n5543_));
  INV_X1     g04539(.I(\A[896] ), .ZN(new_n5544_));
  NAND2_X1   g04540(.A1(new_n5544_), .A2(\A[897] ), .ZN(new_n5545_));
  INV_X1     g04541(.I(\A[897] ), .ZN(new_n5546_));
  NAND2_X1   g04542(.A1(new_n5546_), .A2(\A[896] ), .ZN(new_n5547_));
  AOI21_X1   g04543(.A1(new_n5545_), .A2(new_n5547_), .B(new_n5543_), .ZN(new_n5548_));
  NAND2_X1   g04544(.A1(new_n5544_), .A2(new_n5546_), .ZN(new_n5549_));
  NAND2_X1   g04545(.A1(\A[896] ), .A2(\A[897] ), .ZN(new_n5550_));
  AOI21_X1   g04546(.A1(new_n5549_), .A2(new_n5550_), .B(\A[895] ), .ZN(new_n5551_));
  NOR2_X1    g04547(.A1(new_n5551_), .A2(new_n5548_), .ZN(new_n5552_));
  INV_X1     g04548(.I(\A[898] ), .ZN(new_n5553_));
  INV_X1     g04549(.I(\A[899] ), .ZN(new_n5554_));
  NAND2_X1   g04550(.A1(new_n5554_), .A2(\A[900] ), .ZN(new_n5555_));
  INV_X1     g04551(.I(\A[900] ), .ZN(new_n5556_));
  NAND2_X1   g04552(.A1(new_n5556_), .A2(\A[899] ), .ZN(new_n5557_));
  AOI21_X1   g04553(.A1(new_n5555_), .A2(new_n5557_), .B(new_n5553_), .ZN(new_n5558_));
  NAND2_X1   g04554(.A1(\A[899] ), .A2(\A[900] ), .ZN(new_n5559_));
  NAND2_X1   g04555(.A1(new_n5554_), .A2(new_n5556_), .ZN(new_n5560_));
  AOI21_X1   g04556(.A1(new_n5560_), .A2(new_n5559_), .B(\A[898] ), .ZN(new_n5561_));
  NOR2_X1    g04557(.A1(new_n5561_), .A2(new_n5558_), .ZN(new_n5562_));
  NAND2_X1   g04558(.A1(new_n5550_), .A2(new_n5543_), .ZN(new_n5563_));
  NAND2_X1   g04559(.A1(new_n5563_), .A2(new_n5549_), .ZN(new_n5564_));
  NAND2_X1   g04560(.A1(new_n5559_), .A2(new_n5553_), .ZN(new_n5565_));
  NAND2_X1   g04561(.A1(new_n5565_), .A2(new_n5560_), .ZN(new_n5566_));
  NAND2_X1   g04562(.A1(new_n5564_), .A2(new_n5566_), .ZN(new_n5567_));
  NOR3_X1    g04563(.A1(new_n5552_), .A2(new_n5562_), .A3(new_n5567_), .ZN(new_n5568_));
  XOR2_X1    g04564(.A1(new_n5542_), .A2(new_n5568_), .Z(new_n5569_));
  NAND2_X1   g04565(.A1(new_n5515_), .A2(new_n5569_), .ZN(new_n5570_));
  INV_X1     g04566(.I(new_n5570_), .ZN(new_n5571_));
  NOR2_X1    g04567(.A1(new_n5515_), .A2(new_n5569_), .ZN(new_n5572_));
  NOR3_X1    g04568(.A1(new_n5461_), .A2(new_n5571_), .A3(new_n5572_), .ZN(new_n5573_));
  INV_X1     g04569(.I(new_n5461_), .ZN(new_n5574_));
  NOR2_X1    g04570(.A1(new_n5571_), .A2(new_n5572_), .ZN(new_n5575_));
  NOR2_X1    g04571(.A1(new_n5574_), .A2(new_n5575_), .ZN(new_n5576_));
  NOR2_X1    g04572(.A1(new_n5576_), .A2(new_n5573_), .ZN(new_n5577_));
  INV_X1     g04573(.I(\A[891] ), .ZN(new_n5578_));
  NOR2_X1    g04574(.A1(new_n5578_), .A2(\A[890] ), .ZN(new_n5579_));
  INV_X1     g04575(.I(\A[890] ), .ZN(new_n5580_));
  NOR2_X1    g04576(.A1(new_n5580_), .A2(\A[891] ), .ZN(new_n5581_));
  OAI21_X1   g04577(.A1(new_n5579_), .A2(new_n5581_), .B(\A[889] ), .ZN(new_n5582_));
  NOR2_X1    g04578(.A1(\A[890] ), .A2(\A[891] ), .ZN(new_n5583_));
  NOR2_X1    g04579(.A1(new_n5580_), .A2(new_n5578_), .ZN(new_n5584_));
  NOR2_X1    g04580(.A1(new_n5584_), .A2(new_n5583_), .ZN(new_n5585_));
  OAI21_X1   g04581(.A1(\A[889] ), .A2(new_n5585_), .B(new_n5582_), .ZN(new_n5586_));
  INV_X1     g04582(.I(\A[894] ), .ZN(new_n5587_));
  NOR2_X1    g04583(.A1(new_n5587_), .A2(\A[893] ), .ZN(new_n5588_));
  INV_X1     g04584(.I(\A[893] ), .ZN(new_n5589_));
  NOR2_X1    g04585(.A1(new_n5589_), .A2(\A[894] ), .ZN(new_n5590_));
  OAI21_X1   g04586(.A1(new_n5588_), .A2(new_n5590_), .B(\A[892] ), .ZN(new_n5591_));
  INV_X1     g04587(.I(\A[892] ), .ZN(new_n5592_));
  NOR2_X1    g04588(.A1(new_n5589_), .A2(new_n5587_), .ZN(new_n5593_));
  NOR2_X1    g04589(.A1(\A[893] ), .A2(\A[894] ), .ZN(new_n5594_));
  OAI21_X1   g04590(.A1(new_n5593_), .A2(new_n5594_), .B(new_n5592_), .ZN(new_n5595_));
  NAND2_X1   g04591(.A1(new_n5595_), .A2(new_n5591_), .ZN(new_n5596_));
  NOR2_X1    g04592(.A1(new_n5584_), .A2(\A[889] ), .ZN(new_n5597_));
  NOR2_X1    g04593(.A1(new_n5593_), .A2(\A[892] ), .ZN(new_n5598_));
  OAI22_X1   g04594(.A1(new_n5583_), .A2(new_n5597_), .B1(new_n5598_), .B2(new_n5594_), .ZN(new_n5599_));
  INV_X1     g04595(.I(new_n5599_), .ZN(new_n5600_));
  NAND3_X1   g04596(.A1(new_n5600_), .A2(new_n5586_), .A3(new_n5596_), .ZN(new_n5601_));
  INV_X1     g04597(.I(\A[883] ), .ZN(new_n5602_));
  INV_X1     g04598(.I(\A[884] ), .ZN(new_n5603_));
  NAND2_X1   g04599(.A1(new_n5603_), .A2(\A[885] ), .ZN(new_n5604_));
  INV_X1     g04600(.I(\A[885] ), .ZN(new_n5605_));
  NAND2_X1   g04601(.A1(new_n5605_), .A2(\A[884] ), .ZN(new_n5606_));
  AOI21_X1   g04602(.A1(new_n5604_), .A2(new_n5606_), .B(new_n5602_), .ZN(new_n5607_));
  NAND2_X1   g04603(.A1(new_n5603_), .A2(new_n5605_), .ZN(new_n5608_));
  NAND2_X1   g04604(.A1(\A[884] ), .A2(\A[885] ), .ZN(new_n5609_));
  AOI21_X1   g04605(.A1(new_n5608_), .A2(new_n5609_), .B(\A[883] ), .ZN(new_n5610_));
  NOR2_X1    g04606(.A1(new_n5610_), .A2(new_n5607_), .ZN(new_n5611_));
  INV_X1     g04607(.I(\A[886] ), .ZN(new_n5612_));
  INV_X1     g04608(.I(\A[887] ), .ZN(new_n5613_));
  NAND2_X1   g04609(.A1(new_n5613_), .A2(\A[888] ), .ZN(new_n5614_));
  INV_X1     g04610(.I(\A[888] ), .ZN(new_n5615_));
  NAND2_X1   g04611(.A1(new_n5615_), .A2(\A[887] ), .ZN(new_n5616_));
  AOI21_X1   g04612(.A1(new_n5614_), .A2(new_n5616_), .B(new_n5612_), .ZN(new_n5617_));
  NAND2_X1   g04613(.A1(\A[887] ), .A2(\A[888] ), .ZN(new_n5618_));
  NAND2_X1   g04614(.A1(new_n5613_), .A2(new_n5615_), .ZN(new_n5619_));
  AOI21_X1   g04615(.A1(new_n5619_), .A2(new_n5618_), .B(\A[886] ), .ZN(new_n5620_));
  NOR2_X1    g04616(.A1(new_n5620_), .A2(new_n5617_), .ZN(new_n5621_));
  NAND2_X1   g04617(.A1(new_n5609_), .A2(new_n5602_), .ZN(new_n5622_));
  NAND2_X1   g04618(.A1(new_n5622_), .A2(new_n5608_), .ZN(new_n5623_));
  NAND2_X1   g04619(.A1(new_n5618_), .A2(new_n5612_), .ZN(new_n5624_));
  NAND2_X1   g04620(.A1(new_n5624_), .A2(new_n5619_), .ZN(new_n5625_));
  NAND2_X1   g04621(.A1(new_n5623_), .A2(new_n5625_), .ZN(new_n5626_));
  NOR3_X1    g04622(.A1(new_n5611_), .A2(new_n5621_), .A3(new_n5626_), .ZN(new_n5627_));
  XOR2_X1    g04623(.A1(new_n5601_), .A2(new_n5627_), .Z(new_n5628_));
  INV_X1     g04624(.I(\A[879] ), .ZN(new_n5629_));
  NOR2_X1    g04625(.A1(new_n5629_), .A2(\A[878] ), .ZN(new_n5630_));
  INV_X1     g04626(.I(\A[878] ), .ZN(new_n5631_));
  NOR2_X1    g04627(.A1(new_n5631_), .A2(\A[879] ), .ZN(new_n5632_));
  OAI21_X1   g04628(.A1(new_n5630_), .A2(new_n5632_), .B(\A[877] ), .ZN(new_n5633_));
  NOR2_X1    g04629(.A1(\A[878] ), .A2(\A[879] ), .ZN(new_n5634_));
  NOR2_X1    g04630(.A1(new_n5631_), .A2(new_n5629_), .ZN(new_n5635_));
  NOR2_X1    g04631(.A1(new_n5635_), .A2(new_n5634_), .ZN(new_n5636_));
  OAI21_X1   g04632(.A1(\A[877] ), .A2(new_n5636_), .B(new_n5633_), .ZN(new_n5637_));
  INV_X1     g04633(.I(\A[882] ), .ZN(new_n5638_));
  NOR2_X1    g04634(.A1(new_n5638_), .A2(\A[881] ), .ZN(new_n5639_));
  INV_X1     g04635(.I(\A[881] ), .ZN(new_n5640_));
  NOR2_X1    g04636(.A1(new_n5640_), .A2(\A[882] ), .ZN(new_n5641_));
  OAI21_X1   g04637(.A1(new_n5639_), .A2(new_n5641_), .B(\A[880] ), .ZN(new_n5642_));
  INV_X1     g04638(.I(\A[880] ), .ZN(new_n5643_));
  NOR2_X1    g04639(.A1(\A[881] ), .A2(\A[882] ), .ZN(new_n5644_));
  NOR2_X1    g04640(.A1(new_n5640_), .A2(new_n5638_), .ZN(new_n5645_));
  OAI21_X1   g04641(.A1(new_n5645_), .A2(new_n5644_), .B(new_n5643_), .ZN(new_n5646_));
  NAND2_X1   g04642(.A1(new_n5646_), .A2(new_n5642_), .ZN(new_n5647_));
  NOR2_X1    g04643(.A1(new_n5635_), .A2(\A[877] ), .ZN(new_n5648_));
  NOR2_X1    g04644(.A1(new_n5645_), .A2(\A[880] ), .ZN(new_n5649_));
  OAI22_X1   g04645(.A1(new_n5634_), .A2(new_n5648_), .B1(new_n5649_), .B2(new_n5644_), .ZN(new_n5650_));
  INV_X1     g04646(.I(new_n5650_), .ZN(new_n5651_));
  NAND3_X1   g04647(.A1(new_n5651_), .A2(new_n5637_), .A3(new_n5647_), .ZN(new_n5652_));
  INV_X1     g04648(.I(\A[871] ), .ZN(new_n5653_));
  INV_X1     g04649(.I(\A[872] ), .ZN(new_n5654_));
  NAND2_X1   g04650(.A1(new_n5654_), .A2(\A[873] ), .ZN(new_n5655_));
  INV_X1     g04651(.I(\A[873] ), .ZN(new_n5656_));
  NAND2_X1   g04652(.A1(new_n5656_), .A2(\A[872] ), .ZN(new_n5657_));
  AOI21_X1   g04653(.A1(new_n5655_), .A2(new_n5657_), .B(new_n5653_), .ZN(new_n5658_));
  NAND2_X1   g04654(.A1(new_n5654_), .A2(new_n5656_), .ZN(new_n5659_));
  NAND2_X1   g04655(.A1(\A[872] ), .A2(\A[873] ), .ZN(new_n5660_));
  AOI21_X1   g04656(.A1(new_n5659_), .A2(new_n5660_), .B(\A[871] ), .ZN(new_n5661_));
  NOR2_X1    g04657(.A1(new_n5661_), .A2(new_n5658_), .ZN(new_n5662_));
  INV_X1     g04658(.I(\A[874] ), .ZN(new_n5663_));
  INV_X1     g04659(.I(\A[875] ), .ZN(new_n5664_));
  NAND2_X1   g04660(.A1(new_n5664_), .A2(\A[876] ), .ZN(new_n5665_));
  INV_X1     g04661(.I(\A[876] ), .ZN(new_n5666_));
  NAND2_X1   g04662(.A1(new_n5666_), .A2(\A[875] ), .ZN(new_n5667_));
  AOI21_X1   g04663(.A1(new_n5665_), .A2(new_n5667_), .B(new_n5663_), .ZN(new_n5668_));
  NAND2_X1   g04664(.A1(\A[875] ), .A2(\A[876] ), .ZN(new_n5669_));
  NAND2_X1   g04665(.A1(new_n5664_), .A2(new_n5666_), .ZN(new_n5670_));
  AOI21_X1   g04666(.A1(new_n5670_), .A2(new_n5669_), .B(\A[874] ), .ZN(new_n5671_));
  NOR2_X1    g04667(.A1(new_n5671_), .A2(new_n5668_), .ZN(new_n5672_));
  NAND2_X1   g04668(.A1(new_n5660_), .A2(new_n5653_), .ZN(new_n5673_));
  NAND2_X1   g04669(.A1(new_n5673_), .A2(new_n5659_), .ZN(new_n5674_));
  NAND2_X1   g04670(.A1(new_n5669_), .A2(new_n5663_), .ZN(new_n5675_));
  NAND2_X1   g04671(.A1(new_n5675_), .A2(new_n5670_), .ZN(new_n5676_));
  NAND2_X1   g04672(.A1(new_n5674_), .A2(new_n5676_), .ZN(new_n5677_));
  NOR3_X1    g04673(.A1(new_n5662_), .A2(new_n5672_), .A3(new_n5677_), .ZN(new_n5678_));
  XOR2_X1    g04674(.A1(new_n5652_), .A2(new_n5678_), .Z(new_n5679_));
  XNOR2_X1   g04675(.A1(new_n5628_), .A2(new_n5679_), .ZN(new_n5680_));
  INV_X1     g04676(.I(\A[867] ), .ZN(new_n5681_));
  NOR2_X1    g04677(.A1(new_n5681_), .A2(\A[866] ), .ZN(new_n5682_));
  INV_X1     g04678(.I(\A[866] ), .ZN(new_n5683_));
  NOR2_X1    g04679(.A1(new_n5683_), .A2(\A[867] ), .ZN(new_n5684_));
  OAI21_X1   g04680(.A1(new_n5682_), .A2(new_n5684_), .B(\A[865] ), .ZN(new_n5685_));
  INV_X1     g04681(.I(\A[865] ), .ZN(new_n5686_));
  NOR2_X1    g04682(.A1(\A[866] ), .A2(\A[867] ), .ZN(new_n5687_));
  NOR2_X1    g04683(.A1(new_n5683_), .A2(new_n5681_), .ZN(new_n5688_));
  OAI21_X1   g04684(.A1(new_n5688_), .A2(new_n5687_), .B(new_n5686_), .ZN(new_n5689_));
  NAND2_X1   g04685(.A1(new_n5689_), .A2(new_n5685_), .ZN(new_n5690_));
  INV_X1     g04686(.I(\A[870] ), .ZN(new_n5691_));
  NOR2_X1    g04687(.A1(new_n5691_), .A2(\A[869] ), .ZN(new_n5692_));
  INV_X1     g04688(.I(\A[869] ), .ZN(new_n5693_));
  NOR2_X1    g04689(.A1(new_n5693_), .A2(\A[870] ), .ZN(new_n5694_));
  OAI21_X1   g04690(.A1(new_n5692_), .A2(new_n5694_), .B(\A[868] ), .ZN(new_n5695_));
  INV_X1     g04691(.I(\A[868] ), .ZN(new_n5696_));
  NOR2_X1    g04692(.A1(new_n5693_), .A2(new_n5691_), .ZN(new_n5697_));
  NOR2_X1    g04693(.A1(\A[869] ), .A2(\A[870] ), .ZN(new_n5698_));
  OAI21_X1   g04694(.A1(new_n5697_), .A2(new_n5698_), .B(new_n5696_), .ZN(new_n5699_));
  NAND2_X1   g04695(.A1(new_n5699_), .A2(new_n5695_), .ZN(new_n5700_));
  INV_X1     g04696(.I(new_n5687_), .ZN(new_n5701_));
  OAI21_X1   g04697(.A1(\A[865] ), .A2(new_n5688_), .B(new_n5701_), .ZN(new_n5702_));
  INV_X1     g04698(.I(new_n5698_), .ZN(new_n5703_));
  OAI21_X1   g04699(.A1(\A[868] ), .A2(new_n5697_), .B(new_n5703_), .ZN(new_n5704_));
  NAND2_X1   g04700(.A1(new_n5702_), .A2(new_n5704_), .ZN(new_n5705_));
  INV_X1     g04701(.I(new_n5705_), .ZN(new_n5706_));
  NAND3_X1   g04702(.A1(new_n5706_), .A2(new_n5690_), .A3(new_n5700_), .ZN(new_n5707_));
  INV_X1     g04703(.I(\A[859] ), .ZN(new_n5708_));
  INV_X1     g04704(.I(\A[860] ), .ZN(new_n5709_));
  NAND2_X1   g04705(.A1(new_n5709_), .A2(\A[861] ), .ZN(new_n5710_));
  INV_X1     g04706(.I(\A[861] ), .ZN(new_n5711_));
  NAND2_X1   g04707(.A1(new_n5711_), .A2(\A[860] ), .ZN(new_n5712_));
  AOI21_X1   g04708(.A1(new_n5710_), .A2(new_n5712_), .B(new_n5708_), .ZN(new_n5713_));
  NAND2_X1   g04709(.A1(new_n5709_), .A2(new_n5711_), .ZN(new_n5714_));
  NAND2_X1   g04710(.A1(\A[860] ), .A2(\A[861] ), .ZN(new_n5715_));
  AOI21_X1   g04711(.A1(new_n5714_), .A2(new_n5715_), .B(\A[859] ), .ZN(new_n5716_));
  NOR2_X1    g04712(.A1(new_n5716_), .A2(new_n5713_), .ZN(new_n5717_));
  INV_X1     g04713(.I(\A[862] ), .ZN(new_n5718_));
  INV_X1     g04714(.I(\A[863] ), .ZN(new_n5719_));
  NAND2_X1   g04715(.A1(new_n5719_), .A2(\A[864] ), .ZN(new_n5720_));
  INV_X1     g04716(.I(\A[864] ), .ZN(new_n5721_));
  NAND2_X1   g04717(.A1(new_n5721_), .A2(\A[863] ), .ZN(new_n5722_));
  AOI21_X1   g04718(.A1(new_n5720_), .A2(new_n5722_), .B(new_n5718_), .ZN(new_n5723_));
  NAND2_X1   g04719(.A1(\A[863] ), .A2(\A[864] ), .ZN(new_n5724_));
  NAND2_X1   g04720(.A1(new_n5719_), .A2(new_n5721_), .ZN(new_n5725_));
  AOI21_X1   g04721(.A1(new_n5725_), .A2(new_n5724_), .B(\A[862] ), .ZN(new_n5726_));
  NOR2_X1    g04722(.A1(new_n5726_), .A2(new_n5723_), .ZN(new_n5727_));
  NAND2_X1   g04723(.A1(new_n5715_), .A2(new_n5708_), .ZN(new_n5728_));
  NAND2_X1   g04724(.A1(new_n5728_), .A2(new_n5714_), .ZN(new_n5729_));
  NAND2_X1   g04725(.A1(new_n5724_), .A2(new_n5718_), .ZN(new_n5730_));
  NAND2_X1   g04726(.A1(new_n5730_), .A2(new_n5725_), .ZN(new_n5731_));
  NAND2_X1   g04727(.A1(new_n5729_), .A2(new_n5731_), .ZN(new_n5732_));
  NOR3_X1    g04728(.A1(new_n5717_), .A2(new_n5727_), .A3(new_n5732_), .ZN(new_n5733_));
  XOR2_X1    g04729(.A1(new_n5707_), .A2(new_n5733_), .Z(new_n5734_));
  INV_X1     g04730(.I(\A[855] ), .ZN(new_n5735_));
  NOR2_X1    g04731(.A1(new_n5735_), .A2(\A[854] ), .ZN(new_n5736_));
  INV_X1     g04732(.I(\A[854] ), .ZN(new_n5737_));
  NOR2_X1    g04733(.A1(new_n5737_), .A2(\A[855] ), .ZN(new_n5738_));
  OAI21_X1   g04734(.A1(new_n5736_), .A2(new_n5738_), .B(\A[853] ), .ZN(new_n5739_));
  NOR2_X1    g04735(.A1(\A[854] ), .A2(\A[855] ), .ZN(new_n5740_));
  NOR2_X1    g04736(.A1(new_n5737_), .A2(new_n5735_), .ZN(new_n5741_));
  NOR2_X1    g04737(.A1(new_n5741_), .A2(new_n5740_), .ZN(new_n5742_));
  OAI21_X1   g04738(.A1(\A[853] ), .A2(new_n5742_), .B(new_n5739_), .ZN(new_n5743_));
  INV_X1     g04739(.I(\A[858] ), .ZN(new_n5744_));
  NOR2_X1    g04740(.A1(new_n5744_), .A2(\A[857] ), .ZN(new_n5745_));
  INV_X1     g04741(.I(\A[857] ), .ZN(new_n5746_));
  NOR2_X1    g04742(.A1(new_n5746_), .A2(\A[858] ), .ZN(new_n5747_));
  OAI21_X1   g04743(.A1(new_n5745_), .A2(new_n5747_), .B(\A[856] ), .ZN(new_n5748_));
  INV_X1     g04744(.I(\A[856] ), .ZN(new_n5749_));
  NOR2_X1    g04745(.A1(\A[857] ), .A2(\A[858] ), .ZN(new_n5750_));
  NOR2_X1    g04746(.A1(new_n5746_), .A2(new_n5744_), .ZN(new_n5751_));
  OAI21_X1   g04747(.A1(new_n5751_), .A2(new_n5750_), .B(new_n5749_), .ZN(new_n5752_));
  NAND2_X1   g04748(.A1(new_n5752_), .A2(new_n5748_), .ZN(new_n5753_));
  INV_X1     g04749(.I(new_n5740_), .ZN(new_n5754_));
  OAI21_X1   g04750(.A1(\A[853] ), .A2(new_n5741_), .B(new_n5754_), .ZN(new_n5755_));
  INV_X1     g04751(.I(new_n5750_), .ZN(new_n5756_));
  OAI21_X1   g04752(.A1(\A[856] ), .A2(new_n5751_), .B(new_n5756_), .ZN(new_n5757_));
  NAND2_X1   g04753(.A1(new_n5755_), .A2(new_n5757_), .ZN(new_n5758_));
  INV_X1     g04754(.I(new_n5758_), .ZN(new_n5759_));
  NAND3_X1   g04755(.A1(new_n5759_), .A2(new_n5743_), .A3(new_n5753_), .ZN(new_n5760_));
  INV_X1     g04756(.I(\A[847] ), .ZN(new_n5761_));
  INV_X1     g04757(.I(\A[848] ), .ZN(new_n5762_));
  NAND2_X1   g04758(.A1(new_n5762_), .A2(\A[849] ), .ZN(new_n5763_));
  INV_X1     g04759(.I(\A[849] ), .ZN(new_n5764_));
  NAND2_X1   g04760(.A1(new_n5764_), .A2(\A[848] ), .ZN(new_n5765_));
  AOI21_X1   g04761(.A1(new_n5763_), .A2(new_n5765_), .B(new_n5761_), .ZN(new_n5766_));
  NAND2_X1   g04762(.A1(new_n5762_), .A2(new_n5764_), .ZN(new_n5767_));
  NAND2_X1   g04763(.A1(\A[848] ), .A2(\A[849] ), .ZN(new_n5768_));
  AOI21_X1   g04764(.A1(new_n5767_), .A2(new_n5768_), .B(\A[847] ), .ZN(new_n5769_));
  NOR2_X1    g04765(.A1(new_n5769_), .A2(new_n5766_), .ZN(new_n5770_));
  INV_X1     g04766(.I(\A[850] ), .ZN(new_n5771_));
  INV_X1     g04767(.I(\A[851] ), .ZN(new_n5772_));
  NAND2_X1   g04768(.A1(new_n5772_), .A2(\A[852] ), .ZN(new_n5773_));
  INV_X1     g04769(.I(\A[852] ), .ZN(new_n5774_));
  NAND2_X1   g04770(.A1(new_n5774_), .A2(\A[851] ), .ZN(new_n5775_));
  AOI21_X1   g04771(.A1(new_n5773_), .A2(new_n5775_), .B(new_n5771_), .ZN(new_n5776_));
  NAND2_X1   g04772(.A1(\A[851] ), .A2(\A[852] ), .ZN(new_n5777_));
  NAND2_X1   g04773(.A1(new_n5772_), .A2(new_n5774_), .ZN(new_n5778_));
  AOI21_X1   g04774(.A1(new_n5778_), .A2(new_n5777_), .B(\A[850] ), .ZN(new_n5779_));
  NOR2_X1    g04775(.A1(new_n5779_), .A2(new_n5776_), .ZN(new_n5780_));
  NAND2_X1   g04776(.A1(new_n5768_), .A2(new_n5761_), .ZN(new_n5781_));
  NAND2_X1   g04777(.A1(new_n5781_), .A2(new_n5767_), .ZN(new_n5782_));
  NAND2_X1   g04778(.A1(new_n5777_), .A2(new_n5771_), .ZN(new_n5783_));
  NAND2_X1   g04779(.A1(new_n5783_), .A2(new_n5778_), .ZN(new_n5784_));
  NAND2_X1   g04780(.A1(new_n5782_), .A2(new_n5784_), .ZN(new_n5785_));
  NOR3_X1    g04781(.A1(new_n5770_), .A2(new_n5780_), .A3(new_n5785_), .ZN(new_n5786_));
  XOR2_X1    g04782(.A1(new_n5760_), .A2(new_n5786_), .Z(new_n5787_));
  NAND2_X1   g04783(.A1(new_n5734_), .A2(new_n5787_), .ZN(new_n5788_));
  INV_X1     g04784(.I(new_n5788_), .ZN(new_n5789_));
  NOR2_X1    g04785(.A1(new_n5734_), .A2(new_n5787_), .ZN(new_n5790_));
  NOR3_X1    g04786(.A1(new_n5680_), .A2(new_n5789_), .A3(new_n5790_), .ZN(new_n5791_));
  INV_X1     g04787(.I(new_n5680_), .ZN(new_n5792_));
  NOR2_X1    g04788(.A1(new_n5789_), .A2(new_n5790_), .ZN(new_n5793_));
  NOR2_X1    g04789(.A1(new_n5792_), .A2(new_n5793_), .ZN(new_n5794_));
  NOR2_X1    g04790(.A1(new_n5794_), .A2(new_n5791_), .ZN(new_n5795_));
  NAND2_X1   g04791(.A1(new_n5795_), .A2(new_n5577_), .ZN(new_n5796_));
  INV_X1     g04792(.I(new_n5796_), .ZN(new_n5797_));
  NOR4_X1    g04793(.A1(new_n5601_), .A2(new_n5611_), .A3(new_n5621_), .A4(new_n5626_), .ZN(new_n5798_));
  INV_X1     g04794(.I(new_n5798_), .ZN(new_n5799_));
  INV_X1     g04795(.I(new_n5596_), .ZN(new_n5800_));
  XNOR2_X1   g04796(.A1(new_n5599_), .A2(new_n5586_), .ZN(new_n5801_));
  NAND2_X1   g04797(.A1(new_n5801_), .A2(new_n5800_), .ZN(new_n5802_));
  XOR2_X1    g04798(.A1(new_n5599_), .A2(new_n5586_), .Z(new_n5803_));
  NAND2_X1   g04799(.A1(new_n5803_), .A2(new_n5596_), .ZN(new_n5804_));
  XOR2_X1    g04800(.A1(new_n5586_), .A2(new_n5596_), .Z(new_n5805_));
  NAND2_X1   g04801(.A1(new_n5805_), .A2(new_n5600_), .ZN(new_n5806_));
  NAND3_X1   g04802(.A1(new_n5802_), .A2(new_n5804_), .A3(new_n5806_), .ZN(new_n5807_));
  NOR3_X1    g04803(.A1(new_n5611_), .A2(new_n5621_), .A3(new_n5626_), .ZN(new_n5808_));
  XOR2_X1    g04804(.A1(new_n5611_), .A2(new_n5621_), .Z(new_n5809_));
  NOR2_X1    g04805(.A1(new_n5809_), .A2(new_n5808_), .ZN(new_n5810_));
  NAND4_X1   g04806(.A1(new_n5810_), .A2(new_n5586_), .A3(new_n5596_), .A4(new_n5600_), .ZN(new_n5811_));
  XOR2_X1    g04807(.A1(new_n5611_), .A2(new_n5626_), .Z(new_n5812_));
  XOR2_X1    g04808(.A1(new_n5812_), .A2(new_n5621_), .Z(new_n5813_));
  NOR2_X1    g04809(.A1(new_n5813_), .A2(new_n5811_), .ZN(new_n5814_));
  INV_X1     g04810(.I(new_n5814_), .ZN(new_n5815_));
  AOI21_X1   g04811(.A1(new_n5815_), .A2(new_n5807_), .B(new_n5799_), .ZN(new_n5816_));
  INV_X1     g04812(.I(new_n5816_), .ZN(new_n5817_));
  OR2_X2     g04813(.A1(new_n5620_), .A2(new_n5617_), .Z(new_n5818_));
  XOR2_X1    g04814(.A1(new_n5812_), .A2(new_n5818_), .Z(new_n5819_));
  NOR2_X1    g04815(.A1(new_n5803_), .A2(new_n5596_), .ZN(new_n5820_));
  NOR2_X1    g04816(.A1(new_n5801_), .A2(new_n5800_), .ZN(new_n5821_));
  XNOR2_X1   g04817(.A1(new_n5586_), .A2(new_n5596_), .ZN(new_n5822_));
  NOR2_X1    g04818(.A1(new_n5822_), .A2(new_n5599_), .ZN(new_n5823_));
  NOR3_X1    g04819(.A1(new_n5821_), .A2(new_n5820_), .A3(new_n5823_), .ZN(new_n5824_));
  NAND2_X1   g04820(.A1(new_n5824_), .A2(new_n5799_), .ZN(new_n5825_));
  NAND2_X1   g04821(.A1(new_n5807_), .A2(new_n5798_), .ZN(new_n5826_));
  AOI21_X1   g04822(.A1(new_n5825_), .A2(new_n5826_), .B(new_n5819_), .ZN(new_n5827_));
  INV_X1     g04823(.I(new_n5827_), .ZN(new_n5828_));
  NAND2_X1   g04824(.A1(new_n5628_), .A2(new_n5679_), .ZN(new_n5829_));
  NOR4_X1    g04825(.A1(new_n5652_), .A2(new_n5662_), .A3(new_n5672_), .A4(new_n5677_), .ZN(new_n5830_));
  INV_X1     g04826(.I(new_n5830_), .ZN(new_n5831_));
  INV_X1     g04827(.I(new_n5647_), .ZN(new_n5832_));
  XNOR2_X1   g04828(.A1(new_n5650_), .A2(new_n5637_), .ZN(new_n5833_));
  NAND2_X1   g04829(.A1(new_n5833_), .A2(new_n5832_), .ZN(new_n5834_));
  XOR2_X1    g04830(.A1(new_n5650_), .A2(new_n5637_), .Z(new_n5835_));
  NAND2_X1   g04831(.A1(new_n5835_), .A2(new_n5647_), .ZN(new_n5836_));
  XOR2_X1    g04832(.A1(new_n5637_), .A2(new_n5647_), .Z(new_n5837_));
  NAND2_X1   g04833(.A1(new_n5837_), .A2(new_n5651_), .ZN(new_n5838_));
  NAND3_X1   g04834(.A1(new_n5834_), .A2(new_n5836_), .A3(new_n5838_), .ZN(new_n5839_));
  XOR2_X1    g04835(.A1(new_n5662_), .A2(new_n5677_), .Z(new_n5840_));
  XNOR2_X1   g04836(.A1(new_n5840_), .A2(new_n5672_), .ZN(new_n5841_));
  NOR3_X1    g04837(.A1(new_n5662_), .A2(new_n5672_), .A3(new_n5677_), .ZN(new_n5842_));
  XOR2_X1    g04838(.A1(new_n5662_), .A2(new_n5672_), .Z(new_n5843_));
  NOR2_X1    g04839(.A1(new_n5843_), .A2(new_n5842_), .ZN(new_n5844_));
  NAND4_X1   g04840(.A1(new_n5844_), .A2(new_n5637_), .A3(new_n5647_), .A4(new_n5651_), .ZN(new_n5845_));
  NAND4_X1   g04841(.A1(new_n5841_), .A2(new_n5839_), .A3(new_n5845_), .A4(new_n5831_), .ZN(new_n5846_));
  NOR2_X1    g04842(.A1(new_n5846_), .A2(new_n5829_), .ZN(new_n5847_));
  NAND2_X1   g04843(.A1(new_n5828_), .A2(new_n5847_), .ZN(new_n5848_));
  INV_X1     g04844(.I(new_n5847_), .ZN(new_n5849_));
  NAND2_X1   g04845(.A1(new_n5849_), .A2(new_n5827_), .ZN(new_n5850_));
  AOI21_X1   g04846(.A1(new_n5850_), .A2(new_n5848_), .B(new_n5817_), .ZN(new_n5851_));
  INV_X1     g04847(.I(new_n5727_), .ZN(new_n5852_));
  XOR2_X1    g04848(.A1(new_n5717_), .A2(new_n5732_), .Z(new_n5853_));
  XOR2_X1    g04849(.A1(new_n5853_), .A2(new_n5852_), .Z(new_n5854_));
  NAND4_X1   g04850(.A1(new_n5733_), .A2(new_n5690_), .A3(new_n5706_), .A4(new_n5700_), .ZN(new_n5855_));
  INV_X1     g04851(.I(new_n5700_), .ZN(new_n5856_));
  XNOR2_X1   g04852(.A1(new_n5705_), .A2(new_n5690_), .ZN(new_n5857_));
  NAND2_X1   g04853(.A1(new_n5857_), .A2(new_n5856_), .ZN(new_n5858_));
  XOR2_X1    g04854(.A1(new_n5705_), .A2(new_n5690_), .Z(new_n5859_));
  NAND2_X1   g04855(.A1(new_n5859_), .A2(new_n5700_), .ZN(new_n5860_));
  NAND2_X1   g04856(.A1(new_n5858_), .A2(new_n5860_), .ZN(new_n5861_));
  XNOR2_X1   g04857(.A1(new_n5690_), .A2(new_n5700_), .ZN(new_n5862_));
  NOR2_X1    g04858(.A1(new_n5862_), .A2(new_n5705_), .ZN(new_n5863_));
  NOR2_X1    g04859(.A1(new_n5861_), .A2(new_n5863_), .ZN(new_n5864_));
  NAND2_X1   g04860(.A1(new_n5864_), .A2(new_n5855_), .ZN(new_n5865_));
  INV_X1     g04861(.I(new_n5855_), .ZN(new_n5866_));
  INV_X1     g04862(.I(new_n5863_), .ZN(new_n5867_));
  NAND3_X1   g04863(.A1(new_n5867_), .A2(new_n5858_), .A3(new_n5860_), .ZN(new_n5868_));
  NAND2_X1   g04864(.A1(new_n5868_), .A2(new_n5866_), .ZN(new_n5869_));
  AOI21_X1   g04865(.A1(new_n5865_), .A2(new_n5869_), .B(new_n5854_), .ZN(new_n5870_));
  XOR2_X1    g04866(.A1(new_n5853_), .A2(new_n5727_), .Z(new_n5871_));
  NOR3_X1    g04867(.A1(new_n5717_), .A2(new_n5727_), .A3(new_n5732_), .ZN(new_n5872_));
  XOR2_X1    g04868(.A1(new_n5717_), .A2(new_n5727_), .Z(new_n5873_));
  NOR2_X1    g04869(.A1(new_n5873_), .A2(new_n5872_), .ZN(new_n5874_));
  NAND4_X1   g04870(.A1(new_n5874_), .A2(new_n5690_), .A3(new_n5700_), .A4(new_n5706_), .ZN(new_n5875_));
  NOR2_X1    g04871(.A1(new_n5871_), .A2(new_n5875_), .ZN(new_n5876_));
  OAI21_X1   g04872(.A1(new_n5876_), .A2(new_n5864_), .B(new_n5866_), .ZN(new_n5877_));
  NOR4_X1    g04873(.A1(new_n5760_), .A2(new_n5770_), .A3(new_n5780_), .A4(new_n5785_), .ZN(new_n5878_));
  XOR2_X1    g04874(.A1(new_n5743_), .A2(new_n5758_), .Z(new_n5879_));
  NOR2_X1    g04875(.A1(new_n5879_), .A2(new_n5753_), .ZN(new_n5880_));
  INV_X1     g04876(.I(new_n5753_), .ZN(new_n5881_));
  XNOR2_X1   g04877(.A1(new_n5743_), .A2(new_n5758_), .ZN(new_n5882_));
  NOR2_X1    g04878(.A1(new_n5882_), .A2(new_n5881_), .ZN(new_n5883_));
  XNOR2_X1   g04879(.A1(new_n5743_), .A2(new_n5753_), .ZN(new_n5884_));
  NOR2_X1    g04880(.A1(new_n5884_), .A2(new_n5758_), .ZN(new_n5885_));
  NOR4_X1    g04881(.A1(new_n5883_), .A2(new_n5885_), .A3(new_n5880_), .A4(new_n5878_), .ZN(new_n5886_));
  XOR2_X1    g04882(.A1(new_n5770_), .A2(new_n5785_), .Z(new_n5887_));
  XOR2_X1    g04883(.A1(new_n5887_), .A2(new_n5780_), .Z(new_n5888_));
  INV_X1     g04884(.I(new_n5878_), .ZN(new_n5889_));
  NOR3_X1    g04885(.A1(new_n5770_), .A2(new_n5780_), .A3(new_n5785_), .ZN(new_n5890_));
  XOR2_X1    g04886(.A1(new_n5770_), .A2(new_n5780_), .Z(new_n5891_));
  NOR2_X1    g04887(.A1(new_n5891_), .A2(new_n5890_), .ZN(new_n5892_));
  NAND4_X1   g04888(.A1(new_n5892_), .A2(new_n5743_), .A3(new_n5753_), .A4(new_n5759_), .ZN(new_n5893_));
  NAND2_X1   g04889(.A1(new_n5893_), .A2(new_n5889_), .ZN(new_n5894_));
  NOR4_X1    g04890(.A1(new_n5894_), .A2(new_n5788_), .A3(new_n5886_), .A4(new_n5888_), .ZN(new_n5895_));
  NAND2_X1   g04891(.A1(new_n5895_), .A2(new_n5877_), .ZN(new_n5896_));
  NOR2_X1    g04892(.A1(new_n5895_), .A2(new_n5877_), .ZN(new_n5897_));
  INV_X1     g04893(.I(new_n5897_), .ZN(new_n5898_));
  AOI21_X1   g04894(.A1(new_n5898_), .A2(new_n5896_), .B(new_n5870_), .ZN(new_n5899_));
  INV_X1     g04895(.I(new_n5870_), .ZN(new_n5900_));
  NOR4_X1    g04896(.A1(new_n5863_), .A2(new_n5707_), .A3(new_n5872_), .A4(new_n5873_), .ZN(new_n5901_));
  NAND3_X1   g04897(.A1(new_n5901_), .A2(new_n5854_), .A3(new_n5861_), .ZN(new_n5902_));
  AOI21_X1   g04898(.A1(new_n5902_), .A2(new_n5868_), .B(new_n5855_), .ZN(new_n5903_));
  OR3_X2     g04899(.A1(new_n5883_), .A2(new_n5880_), .A3(new_n5885_), .Z(new_n5904_));
  XNOR2_X1   g04900(.A1(new_n5887_), .A2(new_n5780_), .ZN(new_n5905_));
  NAND4_X1   g04901(.A1(new_n5904_), .A2(new_n5889_), .A3(new_n5905_), .A4(new_n5893_), .ZN(new_n5906_));
  NOR3_X1    g04902(.A1(new_n5903_), .A2(new_n5906_), .A3(new_n5788_), .ZN(new_n5907_));
  NOR3_X1    g04903(.A1(new_n5900_), .A2(new_n5907_), .A3(new_n5897_), .ZN(new_n5908_));
  OAI21_X1   g04904(.A1(new_n5899_), .A2(new_n5908_), .B(new_n5791_), .ZN(new_n5909_));
  NOR2_X1    g04905(.A1(new_n5909_), .A2(new_n5851_), .ZN(new_n5910_));
  INV_X1     g04906(.I(new_n5851_), .ZN(new_n5911_));
  NOR2_X1    g04907(.A1(new_n5909_), .A2(new_n5911_), .ZN(new_n5912_));
  OAI21_X1   g04908(.A1(new_n5910_), .A2(new_n5912_), .B(new_n5797_), .ZN(new_n5913_));
  NAND4_X1   g04909(.A1(new_n5405_), .A2(new_n5362_), .A3(new_n5378_), .A4(new_n5372_), .ZN(new_n5914_));
  INV_X1     g04910(.I(new_n5914_), .ZN(new_n5915_));
  XOR2_X1    g04911(.A1(new_n5377_), .A2(new_n5362_), .Z(new_n5916_));
  XNOR2_X1   g04912(.A1(new_n5916_), .A2(new_n5372_), .ZN(new_n5917_));
  XNOR2_X1   g04913(.A1(new_n5362_), .A2(new_n5372_), .ZN(new_n5918_));
  NOR2_X1    g04914(.A1(new_n5918_), .A2(new_n5377_), .ZN(new_n5919_));
  NOR2_X1    g04915(.A1(new_n5917_), .A2(new_n5919_), .ZN(new_n5920_));
  NOR3_X1    g04916(.A1(new_n5389_), .A2(new_n5399_), .A3(new_n5404_), .ZN(new_n5921_));
  XOR2_X1    g04917(.A1(new_n5389_), .A2(new_n5399_), .Z(new_n5922_));
  NOR2_X1    g04918(.A1(new_n5922_), .A2(new_n5921_), .ZN(new_n5923_));
  NAND4_X1   g04919(.A1(new_n5923_), .A2(new_n5362_), .A3(new_n5372_), .A4(new_n5378_), .ZN(new_n5924_));
  XOR2_X1    g04920(.A1(new_n5389_), .A2(new_n5404_), .Z(new_n5925_));
  XOR2_X1    g04921(.A1(new_n5925_), .A2(new_n5399_), .Z(new_n5926_));
  NOR2_X1    g04922(.A1(new_n5926_), .A2(new_n5924_), .ZN(new_n5927_));
  OAI21_X1   g04923(.A1(new_n5920_), .A2(new_n5927_), .B(new_n5915_), .ZN(new_n5928_));
  INV_X1     g04924(.I(new_n5928_), .ZN(new_n5929_));
  INV_X1     g04925(.I(new_n5926_), .ZN(new_n5930_));
  NAND2_X1   g04926(.A1(new_n5920_), .A2(new_n5914_), .ZN(new_n5931_));
  XOR2_X1    g04927(.A1(new_n5916_), .A2(new_n5372_), .Z(new_n5932_));
  INV_X1     g04928(.I(new_n5919_), .ZN(new_n5933_));
  NAND2_X1   g04929(.A1(new_n5932_), .A2(new_n5933_), .ZN(new_n5934_));
  NAND2_X1   g04930(.A1(new_n5934_), .A2(new_n5915_), .ZN(new_n5935_));
  AOI21_X1   g04931(.A1(new_n5931_), .A2(new_n5935_), .B(new_n5930_), .ZN(new_n5936_));
  NAND2_X1   g04932(.A1(new_n5406_), .A2(new_n5460_), .ZN(new_n5937_));
  NOR4_X1    g04933(.A1(new_n5433_), .A2(new_n5443_), .A3(new_n5453_), .A4(new_n5458_), .ZN(new_n5938_));
  INV_X1     g04934(.I(new_n5426_), .ZN(new_n5939_));
  XOR2_X1    g04935(.A1(new_n5431_), .A2(new_n5416_), .Z(new_n5940_));
  XOR2_X1    g04936(.A1(new_n5940_), .A2(new_n5939_), .Z(new_n5941_));
  XNOR2_X1   g04937(.A1(new_n5416_), .A2(new_n5426_), .ZN(new_n5942_));
  NOR2_X1    g04938(.A1(new_n5942_), .A2(new_n5431_), .ZN(new_n5943_));
  NOR3_X1    g04939(.A1(new_n5941_), .A2(new_n5938_), .A3(new_n5943_), .ZN(new_n5944_));
  XOR2_X1    g04940(.A1(new_n5443_), .A2(new_n5458_), .Z(new_n5945_));
  XOR2_X1    g04941(.A1(new_n5945_), .A2(new_n5453_), .Z(new_n5946_));
  INV_X1     g04942(.I(new_n5938_), .ZN(new_n5947_));
  XOR2_X1    g04943(.A1(new_n5443_), .A2(new_n5453_), .Z(new_n5948_));
  NOR3_X1    g04944(.A1(new_n5443_), .A2(new_n5453_), .A3(new_n5458_), .ZN(new_n5949_));
  NOR2_X1    g04945(.A1(new_n5948_), .A2(new_n5949_), .ZN(new_n5950_));
  NAND4_X1   g04946(.A1(new_n5950_), .A2(new_n5416_), .A3(new_n5426_), .A4(new_n5432_), .ZN(new_n5951_));
  NAND2_X1   g04947(.A1(new_n5951_), .A2(new_n5947_), .ZN(new_n5952_));
  NOR4_X1    g04948(.A1(new_n5944_), .A2(new_n5937_), .A3(new_n5952_), .A4(new_n5946_), .ZN(new_n5953_));
  XOR2_X1    g04949(.A1(new_n5936_), .A2(new_n5953_), .Z(new_n5954_));
  NAND2_X1   g04950(.A1(new_n5954_), .A2(new_n5929_), .ZN(new_n5955_));
  INV_X1     g04951(.I(new_n5573_), .ZN(new_n5956_));
  XOR2_X1    g04952(.A1(new_n5498_), .A2(new_n5513_), .Z(new_n5957_));
  XOR2_X1    g04953(.A1(new_n5957_), .A2(new_n5508_), .Z(new_n5958_));
  NAND4_X1   g04954(.A1(new_n5514_), .A2(new_n5471_), .A3(new_n5487_), .A4(new_n5481_), .ZN(new_n5959_));
  INV_X1     g04955(.I(new_n5959_), .ZN(new_n5960_));
  XOR2_X1    g04956(.A1(new_n5486_), .A2(new_n5471_), .Z(new_n5961_));
  NOR2_X1    g04957(.A1(new_n5961_), .A2(new_n5481_), .ZN(new_n5962_));
  AND2_X2    g04958(.A1(new_n5961_), .A2(new_n5481_), .Z(new_n5963_));
  XNOR2_X1   g04959(.A1(new_n5471_), .A2(new_n5481_), .ZN(new_n5964_));
  NOR2_X1    g04960(.A1(new_n5964_), .A2(new_n5486_), .ZN(new_n5965_));
  OR3_X2     g04961(.A1(new_n5963_), .A2(new_n5962_), .A3(new_n5965_), .Z(new_n5966_));
  NOR2_X1    g04962(.A1(new_n5966_), .A2(new_n5960_), .ZN(new_n5967_));
  INV_X1     g04963(.I(new_n5481_), .ZN(new_n5968_));
  XOR2_X1    g04964(.A1(new_n5961_), .A2(new_n5968_), .Z(new_n5969_));
  NOR2_X1    g04965(.A1(new_n5969_), .A2(new_n5965_), .ZN(new_n5970_));
  NOR2_X1    g04966(.A1(new_n5970_), .A2(new_n5959_), .ZN(new_n5971_));
  OAI21_X1   g04967(.A1(new_n5967_), .A2(new_n5971_), .B(new_n5958_), .ZN(new_n5972_));
  NOR3_X1    g04968(.A1(new_n5498_), .A2(new_n5508_), .A3(new_n5513_), .ZN(new_n5973_));
  XOR2_X1    g04969(.A1(new_n5498_), .A2(new_n5508_), .Z(new_n5974_));
  NOR2_X1    g04970(.A1(new_n5974_), .A2(new_n5973_), .ZN(new_n5975_));
  NAND4_X1   g04971(.A1(new_n5975_), .A2(new_n5471_), .A3(new_n5481_), .A4(new_n5487_), .ZN(new_n5976_));
  NOR2_X1    g04972(.A1(new_n5958_), .A2(new_n5976_), .ZN(new_n5977_));
  OAI21_X1   g04973(.A1(new_n5970_), .A2(new_n5977_), .B(new_n5960_), .ZN(new_n5978_));
  NOR4_X1    g04974(.A1(new_n5542_), .A2(new_n5552_), .A3(new_n5562_), .A4(new_n5567_), .ZN(new_n5979_));
  XOR2_X1    g04975(.A1(new_n5540_), .A2(new_n5525_), .Z(new_n5980_));
  NOR2_X1    g04976(.A1(new_n5980_), .A2(new_n5535_), .ZN(new_n5981_));
  INV_X1     g04977(.I(new_n5535_), .ZN(new_n5982_));
  XNOR2_X1   g04978(.A1(new_n5540_), .A2(new_n5525_), .ZN(new_n5983_));
  NOR2_X1    g04979(.A1(new_n5983_), .A2(new_n5982_), .ZN(new_n5984_));
  XNOR2_X1   g04980(.A1(new_n5525_), .A2(new_n5535_), .ZN(new_n5985_));
  NOR2_X1    g04981(.A1(new_n5985_), .A2(new_n5540_), .ZN(new_n5986_));
  NOR4_X1    g04982(.A1(new_n5984_), .A2(new_n5986_), .A3(new_n5981_), .A4(new_n5979_), .ZN(new_n5987_));
  XOR2_X1    g04983(.A1(new_n5552_), .A2(new_n5567_), .Z(new_n5988_));
  XOR2_X1    g04984(.A1(new_n5988_), .A2(new_n5562_), .Z(new_n5989_));
  INV_X1     g04985(.I(new_n5979_), .ZN(new_n5990_));
  NOR3_X1    g04986(.A1(new_n5552_), .A2(new_n5562_), .A3(new_n5567_), .ZN(new_n5991_));
  XOR2_X1    g04987(.A1(new_n5552_), .A2(new_n5562_), .Z(new_n5992_));
  NOR2_X1    g04988(.A1(new_n5992_), .A2(new_n5991_), .ZN(new_n5993_));
  NAND4_X1   g04989(.A1(new_n5993_), .A2(new_n5525_), .A3(new_n5535_), .A4(new_n5541_), .ZN(new_n5994_));
  NAND2_X1   g04990(.A1(new_n5994_), .A2(new_n5990_), .ZN(new_n5995_));
  NOR4_X1    g04991(.A1(new_n5995_), .A2(new_n5570_), .A3(new_n5987_), .A4(new_n5989_), .ZN(new_n5996_));
  NAND2_X1   g04992(.A1(new_n5978_), .A2(new_n5996_), .ZN(new_n5997_));
  INV_X1     g04993(.I(new_n5997_), .ZN(new_n5998_));
  NOR2_X1    g04994(.A1(new_n5978_), .A2(new_n5996_), .ZN(new_n5999_));
  OAI21_X1   g04995(.A1(new_n5998_), .A2(new_n5999_), .B(new_n5972_), .ZN(new_n6000_));
  XNOR2_X1   g04996(.A1(new_n5957_), .A2(new_n5508_), .ZN(new_n6001_));
  NAND2_X1   g04997(.A1(new_n5970_), .A2(new_n5959_), .ZN(new_n6002_));
  NAND2_X1   g04998(.A1(new_n5966_), .A2(new_n5960_), .ZN(new_n6003_));
  AOI21_X1   g04999(.A1(new_n6003_), .A2(new_n6002_), .B(new_n6001_), .ZN(new_n6004_));
  OR2_X2     g05000(.A1(new_n5978_), .A2(new_n5996_), .Z(new_n6005_));
  NAND3_X1   g05001(.A1(new_n6005_), .A2(new_n5997_), .A3(new_n6004_), .ZN(new_n6006_));
  AOI21_X1   g05002(.A1(new_n6000_), .A2(new_n6006_), .B(new_n5956_), .ZN(new_n6007_));
  NOR2_X1    g05003(.A1(new_n5955_), .A2(new_n6007_), .ZN(new_n6008_));
  INV_X1     g05004(.I(new_n5791_), .ZN(new_n6009_));
  OAI21_X1   g05005(.A1(new_n5897_), .A2(new_n5907_), .B(new_n5900_), .ZN(new_n6010_));
  NAND3_X1   g05006(.A1(new_n5898_), .A2(new_n5896_), .A3(new_n5870_), .ZN(new_n6011_));
  AOI21_X1   g05007(.A1(new_n6011_), .A2(new_n6010_), .B(new_n6009_), .ZN(new_n6012_));
  NAND2_X1   g05008(.A1(new_n6012_), .A2(new_n5911_), .ZN(new_n6013_));
  NAND2_X1   g05009(.A1(new_n6012_), .A2(new_n5851_), .ZN(new_n6014_));
  NAND3_X1   g05010(.A1(new_n6013_), .A2(new_n6014_), .A3(new_n5796_), .ZN(new_n6015_));
  NAND2_X1   g05011(.A1(new_n6015_), .A2(new_n6008_), .ZN(new_n6016_));
  NAND2_X1   g05012(.A1(new_n6016_), .A2(new_n5913_), .ZN(new_n6017_));
  INV_X1     g05013(.I(new_n6017_), .ZN(new_n6018_));
  NAND3_X1   g05014(.A1(new_n6011_), .A2(new_n6010_), .A3(new_n6009_), .ZN(new_n6019_));
  AOI21_X1   g05015(.A1(new_n5851_), .A2(new_n6019_), .B(new_n6012_), .ZN(new_n6020_));
  INV_X1     g05016(.I(new_n5895_), .ZN(new_n6021_));
  NOR3_X1    g05017(.A1(new_n5894_), .A2(new_n5886_), .A3(new_n5888_), .ZN(new_n6022_));
  NOR2_X1    g05018(.A1(new_n6022_), .A2(new_n5789_), .ZN(new_n6023_));
  NAND4_X1   g05019(.A1(new_n5876_), .A2(new_n5868_), .A3(new_n5871_), .A4(new_n5866_), .ZN(new_n6024_));
  OAI21_X1   g05020(.A1(new_n6023_), .A2(new_n6024_), .B(new_n6021_), .ZN(new_n6025_));
  INV_X1     g05021(.I(new_n5893_), .ZN(new_n6026_));
  NAND2_X1   g05022(.A1(new_n5743_), .A2(new_n5753_), .ZN(new_n6027_));
  NOR2_X1    g05023(.A1(new_n5755_), .A2(new_n5757_), .ZN(new_n6028_));
  OAI21_X1   g05024(.A1(new_n6027_), .A2(new_n6028_), .B(new_n5758_), .ZN(new_n6029_));
  NOR2_X1    g05025(.A1(new_n5770_), .A2(new_n5780_), .ZN(new_n6030_));
  OAI21_X1   g05026(.A1(new_n5782_), .A2(new_n5784_), .B(new_n6030_), .ZN(new_n6031_));
  NAND2_X1   g05027(.A1(new_n6031_), .A2(new_n5785_), .ZN(new_n6032_));
  XOR2_X1    g05028(.A1(new_n6032_), .A2(new_n6029_), .Z(new_n6033_));
  AOI21_X1   g05029(.A1(new_n5904_), .A2(new_n5889_), .B(new_n5888_), .ZN(new_n6034_));
  OAI21_X1   g05030(.A1(new_n6034_), .A2(new_n6026_), .B(new_n6033_), .ZN(new_n6035_));
  NAND2_X1   g05031(.A1(new_n5690_), .A2(new_n5700_), .ZN(new_n6036_));
  NOR2_X1    g05032(.A1(new_n5702_), .A2(new_n5704_), .ZN(new_n6037_));
  OAI21_X1   g05033(.A1(new_n6036_), .A2(new_n6037_), .B(new_n5705_), .ZN(new_n6038_));
  NOR2_X1    g05034(.A1(new_n5717_), .A2(new_n5727_), .ZN(new_n6039_));
  OAI21_X1   g05035(.A1(new_n5729_), .A2(new_n5731_), .B(new_n6039_), .ZN(new_n6040_));
  NAND2_X1   g05036(.A1(new_n6040_), .A2(new_n5732_), .ZN(new_n6041_));
  XOR2_X1    g05037(.A1(new_n6041_), .A2(new_n6038_), .Z(new_n6042_));
  INV_X1     g05038(.I(new_n6042_), .ZN(new_n6043_));
  OAI21_X1   g05039(.A1(new_n5864_), .A2(new_n5866_), .B(new_n5854_), .ZN(new_n6044_));
  AOI21_X1   g05040(.A1(new_n6044_), .A2(new_n5875_), .B(new_n6043_), .ZN(new_n6045_));
  NOR2_X1    g05041(.A1(new_n6045_), .A2(new_n6035_), .ZN(new_n6046_));
  XNOR2_X1   g05042(.A1(new_n6032_), .A2(new_n6029_), .ZN(new_n6047_));
  NOR3_X1    g05043(.A1(new_n5880_), .A2(new_n5883_), .A3(new_n5885_), .ZN(new_n6048_));
  OAI21_X1   g05044(.A1(new_n6048_), .A2(new_n5878_), .B(new_n5905_), .ZN(new_n6049_));
  AOI21_X1   g05045(.A1(new_n6049_), .A2(new_n5893_), .B(new_n6047_), .ZN(new_n6050_));
  INV_X1     g05046(.I(new_n5875_), .ZN(new_n6051_));
  AOI21_X1   g05047(.A1(new_n5868_), .A2(new_n5855_), .B(new_n5871_), .ZN(new_n6052_));
  OAI21_X1   g05048(.A1(new_n6052_), .A2(new_n6051_), .B(new_n6042_), .ZN(new_n6053_));
  NOR2_X1    g05049(.A1(new_n6053_), .A2(new_n6050_), .ZN(new_n6054_));
  NOR2_X1    g05050(.A1(new_n6046_), .A2(new_n6054_), .ZN(new_n6055_));
  NOR2_X1    g05051(.A1(new_n6045_), .A2(new_n6050_), .ZN(new_n6056_));
  NOR2_X1    g05052(.A1(new_n6035_), .A2(new_n6053_), .ZN(new_n6057_));
  NOR2_X1    g05053(.A1(new_n6056_), .A2(new_n6057_), .ZN(new_n6058_));
  MUX2_X1    g05054(.I0(new_n6058_), .I1(new_n6055_), .S(new_n6025_), .Z(new_n6059_));
  NAND2_X1   g05055(.A1(new_n5846_), .A2(new_n5829_), .ZN(new_n6060_));
  INV_X1     g05056(.I(new_n6060_), .ZN(new_n6061_));
  NAND4_X1   g05057(.A1(new_n5814_), .A2(new_n5798_), .A3(new_n5807_), .A4(new_n5813_), .ZN(new_n6062_));
  OAI21_X1   g05058(.A1(new_n6061_), .A2(new_n6062_), .B(new_n5849_), .ZN(new_n6063_));
  INV_X1     g05059(.I(new_n5845_), .ZN(new_n6064_));
  NAND2_X1   g05060(.A1(new_n5637_), .A2(new_n5647_), .ZN(new_n6065_));
  NOR4_X1    g05061(.A1(new_n5648_), .A2(new_n5649_), .A3(new_n5634_), .A4(new_n5644_), .ZN(new_n6066_));
  OAI21_X1   g05062(.A1(new_n6065_), .A2(new_n6066_), .B(new_n5650_), .ZN(new_n6067_));
  NOR2_X1    g05063(.A1(new_n5662_), .A2(new_n5672_), .ZN(new_n6068_));
  OAI21_X1   g05064(.A1(new_n5674_), .A2(new_n5676_), .B(new_n6068_), .ZN(new_n6069_));
  NAND2_X1   g05065(.A1(new_n6069_), .A2(new_n5677_), .ZN(new_n6070_));
  XOR2_X1    g05066(.A1(new_n6070_), .A2(new_n6067_), .Z(new_n6071_));
  XOR2_X1    g05067(.A1(new_n5840_), .A2(new_n5672_), .Z(new_n6072_));
  AOI21_X1   g05068(.A1(new_n5831_), .A2(new_n5839_), .B(new_n6072_), .ZN(new_n6073_));
  OAI21_X1   g05069(.A1(new_n6073_), .A2(new_n6064_), .B(new_n6071_), .ZN(new_n6074_));
  OR4_X2     g05070(.A1(new_n5583_), .A2(new_n5597_), .A3(new_n5598_), .A4(new_n5594_), .Z(new_n6075_));
  NAND3_X1   g05071(.A1(new_n6075_), .A2(new_n5586_), .A3(new_n5596_), .ZN(new_n6076_));
  NAND2_X1   g05072(.A1(new_n6076_), .A2(new_n5599_), .ZN(new_n6077_));
  NOR2_X1    g05073(.A1(new_n5611_), .A2(new_n5621_), .ZN(new_n6078_));
  OAI21_X1   g05074(.A1(new_n5623_), .A2(new_n5625_), .B(new_n6078_), .ZN(new_n6079_));
  NAND2_X1   g05075(.A1(new_n6079_), .A2(new_n5626_), .ZN(new_n6080_));
  XNOR2_X1   g05076(.A1(new_n6080_), .A2(new_n6077_), .ZN(new_n6081_));
  OAI21_X1   g05077(.A1(new_n5824_), .A2(new_n5798_), .B(new_n5819_), .ZN(new_n6082_));
  AOI21_X1   g05078(.A1(new_n6082_), .A2(new_n5811_), .B(new_n6081_), .ZN(new_n6083_));
  NOR2_X1    g05079(.A1(new_n6083_), .A2(new_n6074_), .ZN(new_n6084_));
  XNOR2_X1   g05080(.A1(new_n6070_), .A2(new_n6067_), .ZN(new_n6085_));
  NOR2_X1    g05081(.A1(new_n5835_), .A2(new_n5647_), .ZN(new_n6086_));
  NOR2_X1    g05082(.A1(new_n5833_), .A2(new_n5832_), .ZN(new_n6087_));
  XNOR2_X1   g05083(.A1(new_n5637_), .A2(new_n5647_), .ZN(new_n6088_));
  NOR2_X1    g05084(.A1(new_n6088_), .A2(new_n5650_), .ZN(new_n6089_));
  NOR3_X1    g05085(.A1(new_n6087_), .A2(new_n6086_), .A3(new_n6089_), .ZN(new_n6090_));
  OAI21_X1   g05086(.A1(new_n6090_), .A2(new_n5830_), .B(new_n5841_), .ZN(new_n6091_));
  AOI21_X1   g05087(.A1(new_n6091_), .A2(new_n5845_), .B(new_n6085_), .ZN(new_n6092_));
  INV_X1     g05088(.I(new_n5811_), .ZN(new_n6093_));
  XOR2_X1    g05089(.A1(new_n6080_), .A2(new_n6077_), .Z(new_n6094_));
  AOI21_X1   g05090(.A1(new_n5799_), .A2(new_n5807_), .B(new_n5813_), .ZN(new_n6095_));
  OAI21_X1   g05091(.A1(new_n6095_), .A2(new_n6093_), .B(new_n6094_), .ZN(new_n6096_));
  NOR2_X1    g05092(.A1(new_n6092_), .A2(new_n6096_), .ZN(new_n6097_));
  OAI21_X1   g05093(.A1(new_n6084_), .A2(new_n6097_), .B(new_n6063_), .ZN(new_n6098_));
  INV_X1     g05094(.I(new_n6062_), .ZN(new_n6099_));
  AOI21_X1   g05095(.A1(new_n6099_), .A2(new_n6060_), .B(new_n5847_), .ZN(new_n6100_));
  NOR2_X1    g05096(.A1(new_n6092_), .A2(new_n6083_), .ZN(new_n6101_));
  NOR2_X1    g05097(.A1(new_n6074_), .A2(new_n6096_), .ZN(new_n6102_));
  OAI21_X1   g05098(.A1(new_n6102_), .A2(new_n6101_), .B(new_n6100_), .ZN(new_n6103_));
  NAND2_X1   g05099(.A1(new_n6098_), .A2(new_n6103_), .ZN(new_n6104_));
  NAND2_X1   g05100(.A1(new_n6059_), .A2(new_n6104_), .ZN(new_n6105_));
  OAI21_X1   g05101(.A1(new_n6046_), .A2(new_n6054_), .B(new_n6025_), .ZN(new_n6106_));
  NAND2_X1   g05102(.A1(new_n5906_), .A2(new_n5788_), .ZN(new_n6107_));
  NOR4_X1    g05103(.A1(new_n5902_), .A2(new_n5854_), .A3(new_n5855_), .A4(new_n5864_), .ZN(new_n6108_));
  AOI21_X1   g05104(.A1(new_n6107_), .A2(new_n6108_), .B(new_n5895_), .ZN(new_n6109_));
  OAI21_X1   g05105(.A1(new_n6056_), .A2(new_n6057_), .B(new_n6109_), .ZN(new_n6110_));
  NAND2_X1   g05106(.A1(new_n6106_), .A2(new_n6110_), .ZN(new_n6111_));
  NOR2_X1    g05107(.A1(new_n6097_), .A2(new_n6084_), .ZN(new_n6112_));
  NOR2_X1    g05108(.A1(new_n6112_), .A2(new_n6100_), .ZN(new_n6113_));
  NOR2_X1    g05109(.A1(new_n6101_), .A2(new_n6102_), .ZN(new_n6114_));
  NOR2_X1    g05110(.A1(new_n6114_), .A2(new_n6063_), .ZN(new_n6115_));
  NOR2_X1    g05111(.A1(new_n6115_), .A2(new_n6113_), .ZN(new_n6116_));
  NAND2_X1   g05112(.A1(new_n6116_), .A2(new_n6111_), .ZN(new_n6117_));
  AOI21_X1   g05113(.A1(new_n6105_), .A2(new_n6117_), .B(new_n6020_), .ZN(new_n6118_));
  NOR3_X1    g05114(.A1(new_n5899_), .A2(new_n5908_), .A3(new_n5791_), .ZN(new_n6119_));
  OAI21_X1   g05115(.A1(new_n5911_), .A2(new_n6119_), .B(new_n5909_), .ZN(new_n6120_));
  AOI22_X1   g05116(.A1(new_n6098_), .A2(new_n6103_), .B1(new_n6106_), .B2(new_n6110_), .ZN(new_n6121_));
  INV_X1     g05117(.I(new_n6121_), .ZN(new_n6122_));
  NAND2_X1   g05118(.A1(new_n6059_), .A2(new_n6116_), .ZN(new_n6123_));
  AOI21_X1   g05119(.A1(new_n6122_), .A2(new_n6123_), .B(new_n6120_), .ZN(new_n6124_));
  NOR2_X1    g05120(.A1(new_n6124_), .A2(new_n6118_), .ZN(new_n6125_));
  AOI21_X1   g05121(.A1(new_n6005_), .A2(new_n5997_), .B(new_n6004_), .ZN(new_n6126_));
  NOR3_X1    g05122(.A1(new_n5998_), .A2(new_n5999_), .A3(new_n5972_), .ZN(new_n6127_));
  OAI21_X1   g05123(.A1(new_n6127_), .A2(new_n6126_), .B(new_n5573_), .ZN(new_n6128_));
  NOR3_X1    g05124(.A1(new_n6127_), .A2(new_n6126_), .A3(new_n5573_), .ZN(new_n6129_));
  OAI21_X1   g05125(.A1(new_n5955_), .A2(new_n6129_), .B(new_n6128_), .ZN(new_n6130_));
  INV_X1     g05126(.I(new_n5996_), .ZN(new_n6131_));
  NOR3_X1    g05127(.A1(new_n5995_), .A2(new_n5987_), .A3(new_n5989_), .ZN(new_n6132_));
  NOR2_X1    g05128(.A1(new_n6132_), .A2(new_n5571_), .ZN(new_n6133_));
  NAND4_X1   g05129(.A1(new_n5966_), .A2(new_n5977_), .A3(new_n5958_), .A4(new_n5960_), .ZN(new_n6134_));
  OAI21_X1   g05130(.A1(new_n6133_), .A2(new_n6134_), .B(new_n6131_), .ZN(new_n6135_));
  INV_X1     g05131(.I(new_n5994_), .ZN(new_n6136_));
  NAND2_X1   g05132(.A1(new_n5525_), .A2(new_n5535_), .ZN(new_n6137_));
  NOR2_X1    g05133(.A1(new_n5537_), .A2(new_n5539_), .ZN(new_n6138_));
  OAI21_X1   g05134(.A1(new_n6137_), .A2(new_n6138_), .B(new_n5540_), .ZN(new_n6139_));
  NOR2_X1    g05135(.A1(new_n5552_), .A2(new_n5562_), .ZN(new_n6140_));
  OAI21_X1   g05136(.A1(new_n5564_), .A2(new_n5566_), .B(new_n6140_), .ZN(new_n6141_));
  NAND2_X1   g05137(.A1(new_n6141_), .A2(new_n5567_), .ZN(new_n6142_));
  XNOR2_X1   g05138(.A1(new_n6142_), .A2(new_n6139_), .ZN(new_n6143_));
  INV_X1     g05139(.I(new_n6143_), .ZN(new_n6144_));
  NOR3_X1    g05140(.A1(new_n5984_), .A2(new_n5986_), .A3(new_n5981_), .ZN(new_n6145_));
  NOR2_X1    g05141(.A1(new_n6145_), .A2(new_n5979_), .ZN(new_n6146_));
  NOR2_X1    g05142(.A1(new_n6146_), .A2(new_n5989_), .ZN(new_n6147_));
  OAI21_X1   g05143(.A1(new_n6147_), .A2(new_n6136_), .B(new_n6144_), .ZN(new_n6148_));
  NAND2_X1   g05144(.A1(new_n5471_), .A2(new_n5481_), .ZN(new_n6149_));
  NOR2_X1    g05145(.A1(new_n5483_), .A2(new_n5485_), .ZN(new_n6150_));
  OAI21_X1   g05146(.A1(new_n6149_), .A2(new_n6150_), .B(new_n5486_), .ZN(new_n6151_));
  NOR2_X1    g05147(.A1(new_n5498_), .A2(new_n5508_), .ZN(new_n6152_));
  OAI21_X1   g05148(.A1(new_n5510_), .A2(new_n5512_), .B(new_n6152_), .ZN(new_n6153_));
  NAND2_X1   g05149(.A1(new_n6153_), .A2(new_n5513_), .ZN(new_n6154_));
  XNOR2_X1   g05150(.A1(new_n6154_), .A2(new_n6151_), .ZN(new_n6155_));
  OAI21_X1   g05151(.A1(new_n5969_), .A2(new_n5965_), .B(new_n5959_), .ZN(new_n6156_));
  NAND2_X1   g05152(.A1(new_n6156_), .A2(new_n6001_), .ZN(new_n6157_));
  AOI21_X1   g05153(.A1(new_n6157_), .A2(new_n5976_), .B(new_n6155_), .ZN(new_n6158_));
  NOR2_X1    g05154(.A1(new_n6158_), .A2(new_n6148_), .ZN(new_n6159_));
  XNOR2_X1   g05155(.A1(new_n5988_), .A2(new_n5562_), .ZN(new_n6160_));
  OR3_X2     g05156(.A1(new_n5984_), .A2(new_n5981_), .A3(new_n5986_), .Z(new_n6161_));
  NAND2_X1   g05157(.A1(new_n6161_), .A2(new_n5990_), .ZN(new_n6162_));
  NAND2_X1   g05158(.A1(new_n6162_), .A2(new_n6160_), .ZN(new_n6163_));
  AOI21_X1   g05159(.A1(new_n6163_), .A2(new_n5994_), .B(new_n6143_), .ZN(new_n6164_));
  INV_X1     g05160(.I(new_n5976_), .ZN(new_n6165_));
  INV_X1     g05161(.I(new_n6155_), .ZN(new_n6166_));
  AOI21_X1   g05162(.A1(new_n5966_), .A2(new_n5959_), .B(new_n5958_), .ZN(new_n6167_));
  OAI21_X1   g05163(.A1(new_n6167_), .A2(new_n6165_), .B(new_n6166_), .ZN(new_n6168_));
  NOR2_X1    g05164(.A1(new_n6164_), .A2(new_n6168_), .ZN(new_n6169_));
  OAI21_X1   g05165(.A1(new_n6169_), .A2(new_n6159_), .B(new_n6135_), .ZN(new_n6170_));
  NAND4_X1   g05166(.A1(new_n6161_), .A2(new_n5990_), .A3(new_n6160_), .A4(new_n5994_), .ZN(new_n6171_));
  NAND2_X1   g05167(.A1(new_n6171_), .A2(new_n5570_), .ZN(new_n6172_));
  INV_X1     g05168(.I(new_n6134_), .ZN(new_n6173_));
  AOI21_X1   g05169(.A1(new_n6173_), .A2(new_n6172_), .B(new_n5996_), .ZN(new_n6174_));
  NOR2_X1    g05170(.A1(new_n6164_), .A2(new_n6158_), .ZN(new_n6175_));
  NOR2_X1    g05171(.A1(new_n6168_), .A2(new_n6148_), .ZN(new_n6176_));
  OAI21_X1   g05172(.A1(new_n6175_), .A2(new_n6176_), .B(new_n6174_), .ZN(new_n6177_));
  NAND2_X1   g05173(.A1(new_n6177_), .A2(new_n6170_), .ZN(new_n6178_));
  XOR2_X1    g05174(.A1(new_n5940_), .A2(new_n5426_), .Z(new_n6179_));
  INV_X1     g05175(.I(new_n5943_), .ZN(new_n6180_));
  NAND2_X1   g05176(.A1(new_n6179_), .A2(new_n6180_), .ZN(new_n6181_));
  INV_X1     g05177(.I(new_n5946_), .ZN(new_n6182_));
  NAND4_X1   g05178(.A1(new_n6181_), .A2(new_n5947_), .A3(new_n6182_), .A4(new_n5951_), .ZN(new_n6183_));
  NAND2_X1   g05179(.A1(new_n6183_), .A2(new_n5937_), .ZN(new_n6184_));
  NAND4_X1   g05180(.A1(new_n5934_), .A2(new_n5927_), .A3(new_n5915_), .A4(new_n5926_), .ZN(new_n6185_));
  INV_X1     g05181(.I(new_n6185_), .ZN(new_n6186_));
  AOI21_X1   g05182(.A1(new_n6184_), .A2(new_n6186_), .B(new_n5953_), .ZN(new_n6187_));
  NAND2_X1   g05183(.A1(new_n5416_), .A2(new_n5426_), .ZN(new_n6188_));
  NOR2_X1    g05184(.A1(new_n5428_), .A2(new_n5430_), .ZN(new_n6189_));
  OAI21_X1   g05185(.A1(new_n6188_), .A2(new_n6189_), .B(new_n5431_), .ZN(new_n6190_));
  NOR2_X1    g05186(.A1(new_n5443_), .A2(new_n5453_), .ZN(new_n6191_));
  OAI21_X1   g05187(.A1(new_n5455_), .A2(new_n5457_), .B(new_n6191_), .ZN(new_n6192_));
  NAND2_X1   g05188(.A1(new_n6192_), .A2(new_n5458_), .ZN(new_n6193_));
  XNOR2_X1   g05189(.A1(new_n6193_), .A2(new_n6190_), .ZN(new_n6194_));
  OAI21_X1   g05190(.A1(new_n5941_), .A2(new_n5943_), .B(new_n5947_), .ZN(new_n6195_));
  NAND2_X1   g05191(.A1(new_n6195_), .A2(new_n6182_), .ZN(new_n6196_));
  AOI21_X1   g05192(.A1(new_n6196_), .A2(new_n5951_), .B(new_n6194_), .ZN(new_n6197_));
  INV_X1     g05193(.I(new_n5924_), .ZN(new_n6198_));
  NAND2_X1   g05194(.A1(new_n5362_), .A2(new_n5372_), .ZN(new_n6199_));
  NOR2_X1    g05195(.A1(new_n5374_), .A2(new_n5376_), .ZN(new_n6200_));
  OAI21_X1   g05196(.A1(new_n6199_), .A2(new_n6200_), .B(new_n5377_), .ZN(new_n6201_));
  NOR2_X1    g05197(.A1(new_n5389_), .A2(new_n5399_), .ZN(new_n6202_));
  OAI21_X1   g05198(.A1(new_n5401_), .A2(new_n5403_), .B(new_n6202_), .ZN(new_n6203_));
  NAND2_X1   g05199(.A1(new_n6203_), .A2(new_n5404_), .ZN(new_n6204_));
  XNOR2_X1   g05200(.A1(new_n6204_), .A2(new_n6201_), .ZN(new_n6205_));
  INV_X1     g05201(.I(new_n6205_), .ZN(new_n6206_));
  AOI21_X1   g05202(.A1(new_n5934_), .A2(new_n5914_), .B(new_n5926_), .ZN(new_n6207_));
  OAI21_X1   g05203(.A1(new_n6207_), .A2(new_n6198_), .B(new_n6206_), .ZN(new_n6208_));
  NAND2_X1   g05204(.A1(new_n6197_), .A2(new_n6208_), .ZN(new_n6209_));
  INV_X1     g05205(.I(new_n5951_), .ZN(new_n6210_));
  INV_X1     g05206(.I(new_n6194_), .ZN(new_n6211_));
  AOI21_X1   g05207(.A1(new_n6181_), .A2(new_n5947_), .B(new_n5946_), .ZN(new_n6212_));
  OAI21_X1   g05208(.A1(new_n6212_), .A2(new_n6210_), .B(new_n6211_), .ZN(new_n6213_));
  OAI21_X1   g05209(.A1(new_n5920_), .A2(new_n5915_), .B(new_n5930_), .ZN(new_n6214_));
  AOI21_X1   g05210(.A1(new_n6214_), .A2(new_n5924_), .B(new_n6205_), .ZN(new_n6215_));
  NAND2_X1   g05211(.A1(new_n6215_), .A2(new_n6213_), .ZN(new_n6216_));
  AOI21_X1   g05212(.A1(new_n6209_), .A2(new_n6216_), .B(new_n6187_), .ZN(new_n6217_));
  INV_X1     g05213(.I(new_n5937_), .ZN(new_n6218_));
  NAND3_X1   g05214(.A1(new_n6179_), .A2(new_n5947_), .A3(new_n6180_), .ZN(new_n6219_));
  INV_X1     g05215(.I(new_n5952_), .ZN(new_n6220_));
  NAND4_X1   g05216(.A1(new_n6220_), .A2(new_n6218_), .A3(new_n6219_), .A4(new_n6182_), .ZN(new_n6221_));
  NOR3_X1    g05217(.A1(new_n5944_), .A2(new_n5946_), .A3(new_n5952_), .ZN(new_n6222_));
  NOR2_X1    g05218(.A1(new_n6222_), .A2(new_n6218_), .ZN(new_n6223_));
  OAI21_X1   g05219(.A1(new_n6223_), .A2(new_n6185_), .B(new_n6221_), .ZN(new_n6224_));
  NAND2_X1   g05220(.A1(new_n6213_), .A2(new_n6208_), .ZN(new_n6225_));
  NAND2_X1   g05221(.A1(new_n6215_), .A2(new_n6197_), .ZN(new_n6226_));
  AOI21_X1   g05222(.A1(new_n6225_), .A2(new_n6226_), .B(new_n6224_), .ZN(new_n6227_));
  NOR2_X1    g05223(.A1(new_n6227_), .A2(new_n6217_), .ZN(new_n6228_));
  NOR2_X1    g05224(.A1(new_n6228_), .A2(new_n6178_), .ZN(new_n6229_));
  NAND2_X1   g05225(.A1(new_n6164_), .A2(new_n6168_), .ZN(new_n6230_));
  NAND2_X1   g05226(.A1(new_n6158_), .A2(new_n6148_), .ZN(new_n6231_));
  AOI21_X1   g05227(.A1(new_n6230_), .A2(new_n6231_), .B(new_n6174_), .ZN(new_n6232_));
  NAND2_X1   g05228(.A1(new_n6168_), .A2(new_n6148_), .ZN(new_n6233_));
  NAND2_X1   g05229(.A1(new_n6164_), .A2(new_n6158_), .ZN(new_n6234_));
  AOI21_X1   g05230(.A1(new_n6234_), .A2(new_n6233_), .B(new_n6135_), .ZN(new_n6235_));
  NOR2_X1    g05231(.A1(new_n6232_), .A2(new_n6235_), .ZN(new_n6236_));
  NOR2_X1    g05232(.A1(new_n6215_), .A2(new_n6213_), .ZN(new_n6237_));
  NOR2_X1    g05233(.A1(new_n6197_), .A2(new_n6208_), .ZN(new_n6238_));
  OAI21_X1   g05234(.A1(new_n6237_), .A2(new_n6238_), .B(new_n6224_), .ZN(new_n6239_));
  NOR2_X1    g05235(.A1(new_n6215_), .A2(new_n6197_), .ZN(new_n6240_));
  NOR2_X1    g05236(.A1(new_n6213_), .A2(new_n6208_), .ZN(new_n6241_));
  OAI21_X1   g05237(.A1(new_n6240_), .A2(new_n6241_), .B(new_n6187_), .ZN(new_n6242_));
  NAND2_X1   g05238(.A1(new_n6239_), .A2(new_n6242_), .ZN(new_n6243_));
  NOR2_X1    g05239(.A1(new_n6243_), .A2(new_n6236_), .ZN(new_n6244_));
  OAI21_X1   g05240(.A1(new_n6244_), .A2(new_n6229_), .B(new_n6130_), .ZN(new_n6245_));
  XOR2_X1    g05241(.A1(new_n5936_), .A2(new_n6221_), .Z(new_n6246_));
  NOR2_X1    g05242(.A1(new_n6246_), .A2(new_n5928_), .ZN(new_n6247_));
  NAND3_X1   g05243(.A1(new_n6000_), .A2(new_n6006_), .A3(new_n5956_), .ZN(new_n6248_));
  AOI21_X1   g05244(.A1(new_n6247_), .A2(new_n6248_), .B(new_n6007_), .ZN(new_n6249_));
  AOI22_X1   g05245(.A1(new_n6239_), .A2(new_n6242_), .B1(new_n6177_), .B2(new_n6170_), .ZN(new_n6250_));
  NOR4_X1    g05246(.A1(new_n6217_), .A2(new_n6227_), .A3(new_n6232_), .A4(new_n6235_), .ZN(new_n6251_));
  OAI21_X1   g05247(.A1(new_n6250_), .A2(new_n6251_), .B(new_n6249_), .ZN(new_n6252_));
  NAND2_X1   g05248(.A1(new_n6245_), .A2(new_n6252_), .ZN(new_n6253_));
  NAND2_X1   g05249(.A1(new_n6253_), .A2(new_n6125_), .ZN(new_n6254_));
  NOR2_X1    g05250(.A1(new_n6116_), .A2(new_n6111_), .ZN(new_n6255_));
  NOR2_X1    g05251(.A1(new_n6059_), .A2(new_n6104_), .ZN(new_n6256_));
  OAI21_X1   g05252(.A1(new_n6256_), .A2(new_n6255_), .B(new_n6120_), .ZN(new_n6257_));
  NOR2_X1    g05253(.A1(new_n6104_), .A2(new_n6111_), .ZN(new_n6258_));
  OAI21_X1   g05254(.A1(new_n6258_), .A2(new_n6121_), .B(new_n6020_), .ZN(new_n6259_));
  NAND2_X1   g05255(.A1(new_n6257_), .A2(new_n6259_), .ZN(new_n6260_));
  NAND2_X1   g05256(.A1(new_n6243_), .A2(new_n6236_), .ZN(new_n6261_));
  NAND2_X1   g05257(.A1(new_n6228_), .A2(new_n6178_), .ZN(new_n6262_));
  AOI21_X1   g05258(.A1(new_n6261_), .A2(new_n6262_), .B(new_n6249_), .ZN(new_n6263_));
  NAND2_X1   g05259(.A1(new_n6243_), .A2(new_n6178_), .ZN(new_n6264_));
  NAND4_X1   g05260(.A1(new_n6177_), .A2(new_n6239_), .A3(new_n6242_), .A4(new_n6170_), .ZN(new_n6265_));
  AOI21_X1   g05261(.A1(new_n6264_), .A2(new_n6265_), .B(new_n6130_), .ZN(new_n6266_));
  NOR2_X1    g05262(.A1(new_n6263_), .A2(new_n6266_), .ZN(new_n6267_));
  NAND2_X1   g05263(.A1(new_n6267_), .A2(new_n6260_), .ZN(new_n6268_));
  AOI21_X1   g05264(.A1(new_n6254_), .A2(new_n6268_), .B(new_n6018_), .ZN(new_n6269_));
  NAND2_X1   g05265(.A1(new_n6253_), .A2(new_n6260_), .ZN(new_n6270_));
  NAND4_X1   g05266(.A1(new_n6245_), .A2(new_n6252_), .A3(new_n6257_), .A4(new_n6259_), .ZN(new_n6271_));
  AOI21_X1   g05267(.A1(new_n6270_), .A2(new_n6271_), .B(new_n6017_), .ZN(new_n6272_));
  NOR2_X1    g05268(.A1(new_n6269_), .A2(new_n6272_), .ZN(new_n6273_));
  INV_X1     g05269(.I(\A[969] ), .ZN(new_n6274_));
  NOR2_X1    g05270(.A1(new_n6274_), .A2(\A[968] ), .ZN(new_n6275_));
  INV_X1     g05271(.I(\A[968] ), .ZN(new_n6276_));
  NOR2_X1    g05272(.A1(new_n6276_), .A2(\A[969] ), .ZN(new_n6277_));
  OAI21_X1   g05273(.A1(new_n6275_), .A2(new_n6277_), .B(\A[967] ), .ZN(new_n6278_));
  INV_X1     g05274(.I(\A[967] ), .ZN(new_n6279_));
  NAND2_X1   g05275(.A1(\A[968] ), .A2(\A[969] ), .ZN(new_n6280_));
  INV_X1     g05276(.I(new_n6280_), .ZN(new_n6281_));
  NOR2_X1    g05277(.A1(\A[968] ), .A2(\A[969] ), .ZN(new_n6282_));
  OAI21_X1   g05278(.A1(new_n6281_), .A2(new_n6282_), .B(new_n6279_), .ZN(new_n6283_));
  NAND2_X1   g05279(.A1(new_n6278_), .A2(new_n6283_), .ZN(new_n6284_));
  INV_X1     g05280(.I(\A[972] ), .ZN(new_n6285_));
  NOR2_X1    g05281(.A1(new_n6285_), .A2(\A[971] ), .ZN(new_n6286_));
  INV_X1     g05282(.I(\A[971] ), .ZN(new_n6287_));
  NOR2_X1    g05283(.A1(new_n6287_), .A2(\A[972] ), .ZN(new_n6288_));
  OAI21_X1   g05284(.A1(new_n6286_), .A2(new_n6288_), .B(\A[970] ), .ZN(new_n6289_));
  INV_X1     g05285(.I(\A[970] ), .ZN(new_n6290_));
  NAND2_X1   g05286(.A1(\A[971] ), .A2(\A[972] ), .ZN(new_n6291_));
  INV_X1     g05287(.I(new_n6291_), .ZN(new_n6292_));
  NOR2_X1    g05288(.A1(\A[971] ), .A2(\A[972] ), .ZN(new_n6293_));
  OAI21_X1   g05289(.A1(new_n6292_), .A2(new_n6293_), .B(new_n6290_), .ZN(new_n6294_));
  NAND2_X1   g05290(.A1(new_n6289_), .A2(new_n6294_), .ZN(new_n6295_));
  NAND2_X1   g05291(.A1(new_n6284_), .A2(new_n6295_), .ZN(new_n6296_));
  NAND2_X1   g05292(.A1(new_n6276_), .A2(\A[969] ), .ZN(new_n6297_));
  NAND2_X1   g05293(.A1(new_n6274_), .A2(\A[968] ), .ZN(new_n6298_));
  AOI21_X1   g05294(.A1(new_n6297_), .A2(new_n6298_), .B(new_n6279_), .ZN(new_n6299_));
  INV_X1     g05295(.I(new_n6282_), .ZN(new_n6300_));
  AOI21_X1   g05296(.A1(new_n6300_), .A2(new_n6280_), .B(\A[967] ), .ZN(new_n6301_));
  NOR2_X1    g05297(.A1(new_n6301_), .A2(new_n6299_), .ZN(new_n6302_));
  NAND2_X1   g05298(.A1(new_n6287_), .A2(\A[972] ), .ZN(new_n6303_));
  NAND2_X1   g05299(.A1(new_n6285_), .A2(\A[971] ), .ZN(new_n6304_));
  AOI21_X1   g05300(.A1(new_n6303_), .A2(new_n6304_), .B(new_n6290_), .ZN(new_n6305_));
  INV_X1     g05301(.I(new_n6293_), .ZN(new_n6306_));
  AOI21_X1   g05302(.A1(new_n6306_), .A2(new_n6291_), .B(\A[970] ), .ZN(new_n6307_));
  NOR2_X1    g05303(.A1(new_n6307_), .A2(new_n6305_), .ZN(new_n6308_));
  NAND2_X1   g05304(.A1(new_n6302_), .A2(new_n6308_), .ZN(new_n6309_));
  NAND2_X1   g05305(.A1(new_n6309_), .A2(new_n6296_), .ZN(new_n6310_));
  AOI21_X1   g05306(.A1(new_n6279_), .A2(new_n6280_), .B(new_n6282_), .ZN(new_n6311_));
  AOI21_X1   g05307(.A1(new_n6290_), .A2(new_n6291_), .B(new_n6293_), .ZN(new_n6312_));
  NOR2_X1    g05308(.A1(new_n6311_), .A2(new_n6312_), .ZN(new_n6313_));
  NAND3_X1   g05309(.A1(new_n6284_), .A2(new_n6295_), .A3(new_n6313_), .ZN(new_n6314_));
  INV_X1     g05310(.I(new_n6314_), .ZN(new_n6315_));
  NOR2_X1    g05311(.A1(new_n6310_), .A2(new_n6315_), .ZN(new_n6316_));
  INV_X1     g05312(.I(\A[973] ), .ZN(new_n6317_));
  INV_X1     g05313(.I(\A[974] ), .ZN(new_n6318_));
  NAND2_X1   g05314(.A1(new_n6318_), .A2(\A[975] ), .ZN(new_n6319_));
  INV_X1     g05315(.I(\A[975] ), .ZN(new_n6320_));
  NAND2_X1   g05316(.A1(new_n6320_), .A2(\A[974] ), .ZN(new_n6321_));
  AOI21_X1   g05317(.A1(new_n6319_), .A2(new_n6321_), .B(new_n6317_), .ZN(new_n6322_));
  NOR2_X1    g05318(.A1(\A[974] ), .A2(\A[975] ), .ZN(new_n6323_));
  INV_X1     g05319(.I(new_n6323_), .ZN(new_n6324_));
  NAND2_X1   g05320(.A1(\A[974] ), .A2(\A[975] ), .ZN(new_n6325_));
  AOI21_X1   g05321(.A1(new_n6324_), .A2(new_n6325_), .B(\A[973] ), .ZN(new_n6326_));
  NOR2_X1    g05322(.A1(new_n6326_), .A2(new_n6322_), .ZN(new_n6327_));
  INV_X1     g05323(.I(\A[976] ), .ZN(new_n6328_));
  INV_X1     g05324(.I(\A[977] ), .ZN(new_n6329_));
  NAND2_X1   g05325(.A1(new_n6329_), .A2(\A[978] ), .ZN(new_n6330_));
  INV_X1     g05326(.I(\A[978] ), .ZN(new_n6331_));
  NAND2_X1   g05327(.A1(new_n6331_), .A2(\A[977] ), .ZN(new_n6332_));
  AOI21_X1   g05328(.A1(new_n6330_), .A2(new_n6332_), .B(new_n6328_), .ZN(new_n6333_));
  NOR2_X1    g05329(.A1(\A[977] ), .A2(\A[978] ), .ZN(new_n6334_));
  INV_X1     g05330(.I(new_n6334_), .ZN(new_n6335_));
  NAND2_X1   g05331(.A1(\A[977] ), .A2(\A[978] ), .ZN(new_n6336_));
  AOI21_X1   g05332(.A1(new_n6335_), .A2(new_n6336_), .B(\A[976] ), .ZN(new_n6337_));
  NOR2_X1    g05333(.A1(new_n6337_), .A2(new_n6333_), .ZN(new_n6338_));
  NAND2_X1   g05334(.A1(new_n6327_), .A2(new_n6338_), .ZN(new_n6339_));
  AOI21_X1   g05335(.A1(new_n6328_), .A2(new_n6336_), .B(new_n6334_), .ZN(new_n6340_));
  INV_X1     g05336(.I(new_n6340_), .ZN(new_n6341_));
  AOI21_X1   g05337(.A1(new_n6317_), .A2(new_n6325_), .B(new_n6323_), .ZN(new_n6342_));
  INV_X1     g05338(.I(new_n6342_), .ZN(new_n6343_));
  NOR2_X1    g05339(.A1(new_n6341_), .A2(new_n6343_), .ZN(new_n6344_));
  INV_X1     g05340(.I(new_n6344_), .ZN(new_n6345_));
  NOR2_X1    g05341(.A1(new_n6339_), .A2(new_n6345_), .ZN(new_n6346_));
  NOR2_X1    g05342(.A1(new_n6320_), .A2(\A[974] ), .ZN(new_n6347_));
  NOR2_X1    g05343(.A1(new_n6318_), .A2(\A[975] ), .ZN(new_n6348_));
  OAI21_X1   g05344(.A1(new_n6347_), .A2(new_n6348_), .B(\A[973] ), .ZN(new_n6349_));
  INV_X1     g05345(.I(new_n6325_), .ZN(new_n6350_));
  OAI21_X1   g05346(.A1(new_n6350_), .A2(new_n6323_), .B(new_n6317_), .ZN(new_n6351_));
  NAND2_X1   g05347(.A1(new_n6349_), .A2(new_n6351_), .ZN(new_n6352_));
  NOR2_X1    g05348(.A1(new_n6331_), .A2(\A[977] ), .ZN(new_n6353_));
  NOR2_X1    g05349(.A1(new_n6329_), .A2(\A[978] ), .ZN(new_n6354_));
  OAI21_X1   g05350(.A1(new_n6353_), .A2(new_n6354_), .B(\A[976] ), .ZN(new_n6355_));
  INV_X1     g05351(.I(new_n6336_), .ZN(new_n6356_));
  OAI21_X1   g05352(.A1(new_n6356_), .A2(new_n6334_), .B(new_n6328_), .ZN(new_n6357_));
  NAND2_X1   g05353(.A1(new_n6355_), .A2(new_n6357_), .ZN(new_n6358_));
  NAND2_X1   g05354(.A1(new_n6352_), .A2(new_n6358_), .ZN(new_n6359_));
  NAND2_X1   g05355(.A1(new_n6339_), .A2(new_n6359_), .ZN(new_n6360_));
  NOR2_X1    g05356(.A1(new_n6360_), .A2(new_n6346_), .ZN(new_n6361_));
  INV_X1     g05357(.I(\A[987] ), .ZN(new_n6362_));
  NOR2_X1    g05358(.A1(new_n6362_), .A2(\A[986] ), .ZN(new_n6363_));
  INV_X1     g05359(.I(\A[986] ), .ZN(new_n6364_));
  NOR2_X1    g05360(.A1(new_n6364_), .A2(\A[987] ), .ZN(new_n6365_));
  OAI21_X1   g05361(.A1(new_n6363_), .A2(new_n6365_), .B(\A[985] ), .ZN(new_n6366_));
  INV_X1     g05362(.I(\A[985] ), .ZN(new_n6367_));
  NOR2_X1    g05363(.A1(\A[986] ), .A2(\A[987] ), .ZN(new_n6368_));
  NAND2_X1   g05364(.A1(\A[986] ), .A2(\A[987] ), .ZN(new_n6369_));
  INV_X1     g05365(.I(new_n6369_), .ZN(new_n6370_));
  OAI21_X1   g05366(.A1(new_n6370_), .A2(new_n6368_), .B(new_n6367_), .ZN(new_n6371_));
  NAND2_X1   g05367(.A1(new_n6366_), .A2(new_n6371_), .ZN(new_n6372_));
  INV_X1     g05368(.I(\A[990] ), .ZN(new_n6373_));
  NOR2_X1    g05369(.A1(new_n6373_), .A2(\A[989] ), .ZN(new_n6374_));
  INV_X1     g05370(.I(\A[989] ), .ZN(new_n6375_));
  NOR2_X1    g05371(.A1(new_n6375_), .A2(\A[990] ), .ZN(new_n6376_));
  OAI21_X1   g05372(.A1(new_n6374_), .A2(new_n6376_), .B(\A[988] ), .ZN(new_n6377_));
  INV_X1     g05373(.I(\A[988] ), .ZN(new_n6378_));
  NOR2_X1    g05374(.A1(\A[989] ), .A2(\A[990] ), .ZN(new_n6379_));
  NAND2_X1   g05375(.A1(\A[989] ), .A2(\A[990] ), .ZN(new_n6380_));
  INV_X1     g05376(.I(new_n6380_), .ZN(new_n6381_));
  OAI21_X1   g05377(.A1(new_n6381_), .A2(new_n6379_), .B(new_n6378_), .ZN(new_n6382_));
  NAND2_X1   g05378(.A1(new_n6377_), .A2(new_n6382_), .ZN(new_n6383_));
  NOR2_X1    g05379(.A1(new_n6372_), .A2(new_n6383_), .ZN(new_n6384_));
  AOI21_X1   g05380(.A1(new_n6378_), .A2(new_n6380_), .B(new_n6379_), .ZN(new_n6385_));
  INV_X1     g05381(.I(new_n6385_), .ZN(new_n6386_));
  AOI21_X1   g05382(.A1(new_n6367_), .A2(new_n6369_), .B(new_n6368_), .ZN(new_n6387_));
  INV_X1     g05383(.I(new_n6387_), .ZN(new_n6388_));
  NOR2_X1    g05384(.A1(new_n6386_), .A2(new_n6388_), .ZN(new_n6389_));
  NAND2_X1   g05385(.A1(new_n6384_), .A2(new_n6389_), .ZN(new_n6390_));
  NAND2_X1   g05386(.A1(new_n6364_), .A2(\A[987] ), .ZN(new_n6391_));
  NAND2_X1   g05387(.A1(new_n6362_), .A2(\A[986] ), .ZN(new_n6392_));
  AOI21_X1   g05388(.A1(new_n6391_), .A2(new_n6392_), .B(new_n6367_), .ZN(new_n6393_));
  INV_X1     g05389(.I(new_n6368_), .ZN(new_n6394_));
  AOI21_X1   g05390(.A1(new_n6394_), .A2(new_n6369_), .B(\A[985] ), .ZN(new_n6395_));
  NOR2_X1    g05391(.A1(new_n6395_), .A2(new_n6393_), .ZN(new_n6396_));
  NAND2_X1   g05392(.A1(new_n6375_), .A2(\A[990] ), .ZN(new_n6397_));
  NAND2_X1   g05393(.A1(new_n6373_), .A2(\A[989] ), .ZN(new_n6398_));
  AOI21_X1   g05394(.A1(new_n6397_), .A2(new_n6398_), .B(new_n6378_), .ZN(new_n6399_));
  INV_X1     g05395(.I(new_n6379_), .ZN(new_n6400_));
  AOI21_X1   g05396(.A1(new_n6400_), .A2(new_n6380_), .B(\A[988] ), .ZN(new_n6401_));
  NOR2_X1    g05397(.A1(new_n6401_), .A2(new_n6399_), .ZN(new_n6402_));
  NOR2_X1    g05398(.A1(new_n6396_), .A2(new_n6402_), .ZN(new_n6403_));
  NOR2_X1    g05399(.A1(new_n6403_), .A2(new_n6384_), .ZN(new_n6404_));
  NAND2_X1   g05400(.A1(new_n6404_), .A2(new_n6390_), .ZN(new_n6405_));
  INV_X1     g05401(.I(\A[981] ), .ZN(new_n6406_));
  NOR2_X1    g05402(.A1(new_n6406_), .A2(\A[980] ), .ZN(new_n6407_));
  INV_X1     g05403(.I(\A[980] ), .ZN(new_n6408_));
  NOR2_X1    g05404(.A1(new_n6408_), .A2(\A[981] ), .ZN(new_n6409_));
  OAI21_X1   g05405(.A1(new_n6407_), .A2(new_n6409_), .B(\A[979] ), .ZN(new_n6410_));
  INV_X1     g05406(.I(\A[979] ), .ZN(new_n6411_));
  NAND2_X1   g05407(.A1(\A[980] ), .A2(\A[981] ), .ZN(new_n6412_));
  INV_X1     g05408(.I(new_n6412_), .ZN(new_n6413_));
  NOR2_X1    g05409(.A1(\A[980] ), .A2(\A[981] ), .ZN(new_n6414_));
  OAI21_X1   g05410(.A1(new_n6413_), .A2(new_n6414_), .B(new_n6411_), .ZN(new_n6415_));
  NAND2_X1   g05411(.A1(new_n6410_), .A2(new_n6415_), .ZN(new_n6416_));
  INV_X1     g05412(.I(\A[984] ), .ZN(new_n6417_));
  NOR2_X1    g05413(.A1(new_n6417_), .A2(\A[983] ), .ZN(new_n6418_));
  INV_X1     g05414(.I(\A[983] ), .ZN(new_n6419_));
  NOR2_X1    g05415(.A1(new_n6419_), .A2(\A[984] ), .ZN(new_n6420_));
  OAI21_X1   g05416(.A1(new_n6418_), .A2(new_n6420_), .B(\A[982] ), .ZN(new_n6421_));
  INV_X1     g05417(.I(\A[982] ), .ZN(new_n6422_));
  NAND2_X1   g05418(.A1(\A[983] ), .A2(\A[984] ), .ZN(new_n6423_));
  INV_X1     g05419(.I(new_n6423_), .ZN(new_n6424_));
  NOR2_X1    g05420(.A1(\A[983] ), .A2(\A[984] ), .ZN(new_n6425_));
  OAI21_X1   g05421(.A1(new_n6424_), .A2(new_n6425_), .B(new_n6422_), .ZN(new_n6426_));
  NAND2_X1   g05422(.A1(new_n6421_), .A2(new_n6426_), .ZN(new_n6427_));
  NAND2_X1   g05423(.A1(new_n6416_), .A2(new_n6427_), .ZN(new_n6428_));
  NAND2_X1   g05424(.A1(new_n6408_), .A2(\A[981] ), .ZN(new_n6429_));
  NAND2_X1   g05425(.A1(new_n6406_), .A2(\A[980] ), .ZN(new_n6430_));
  AOI21_X1   g05426(.A1(new_n6429_), .A2(new_n6430_), .B(new_n6411_), .ZN(new_n6431_));
  INV_X1     g05427(.I(new_n6414_), .ZN(new_n6432_));
  AOI21_X1   g05428(.A1(new_n6432_), .A2(new_n6412_), .B(\A[979] ), .ZN(new_n6433_));
  NOR2_X1    g05429(.A1(new_n6433_), .A2(new_n6431_), .ZN(new_n6434_));
  NAND2_X1   g05430(.A1(new_n6419_), .A2(\A[984] ), .ZN(new_n6435_));
  NAND2_X1   g05431(.A1(new_n6417_), .A2(\A[983] ), .ZN(new_n6436_));
  AOI21_X1   g05432(.A1(new_n6435_), .A2(new_n6436_), .B(new_n6422_), .ZN(new_n6437_));
  INV_X1     g05433(.I(new_n6425_), .ZN(new_n6438_));
  AOI21_X1   g05434(.A1(new_n6438_), .A2(new_n6423_), .B(\A[982] ), .ZN(new_n6439_));
  NOR2_X1    g05435(.A1(new_n6439_), .A2(new_n6437_), .ZN(new_n6440_));
  NAND2_X1   g05436(.A1(new_n6434_), .A2(new_n6440_), .ZN(new_n6441_));
  AOI21_X1   g05437(.A1(new_n6422_), .A2(new_n6423_), .B(new_n6425_), .ZN(new_n6442_));
  NOR4_X1    g05438(.A1(new_n6442_), .A2(\A[979] ), .A3(\A[980] ), .A4(\A[981] ), .ZN(new_n6443_));
  NAND2_X1   g05439(.A1(new_n6427_), .A2(new_n6443_), .ZN(new_n6444_));
  AND3_X2    g05440(.A1(new_n6441_), .A2(new_n6428_), .A3(new_n6444_), .Z(new_n6445_));
  NAND2_X1   g05441(.A1(new_n6405_), .A2(new_n6445_), .ZN(new_n6446_));
  NAND2_X1   g05442(.A1(new_n6396_), .A2(new_n6402_), .ZN(new_n6447_));
  NAND2_X1   g05443(.A1(new_n6372_), .A2(new_n6383_), .ZN(new_n6448_));
  NAND2_X1   g05444(.A1(new_n6447_), .A2(new_n6448_), .ZN(new_n6449_));
  AOI21_X1   g05445(.A1(new_n6384_), .A2(new_n6389_), .B(new_n6449_), .ZN(new_n6450_));
  NOR2_X1    g05446(.A1(new_n6434_), .A2(new_n6440_), .ZN(new_n6451_));
  NOR2_X1    g05447(.A1(new_n6416_), .A2(new_n6427_), .ZN(new_n6452_));
  NOR2_X1    g05448(.A1(new_n6451_), .A2(new_n6452_), .ZN(new_n6453_));
  NAND2_X1   g05449(.A1(new_n6453_), .A2(new_n6444_), .ZN(new_n6454_));
  NAND2_X1   g05450(.A1(new_n6450_), .A2(new_n6454_), .ZN(new_n6455_));
  AOI21_X1   g05451(.A1(new_n6455_), .A2(new_n6446_), .B(new_n6361_), .ZN(new_n6456_));
  INV_X1     g05452(.I(new_n6456_), .ZN(new_n6457_));
  NAND3_X1   g05453(.A1(new_n6455_), .A2(new_n6446_), .A3(new_n6361_), .ZN(new_n6458_));
  AOI21_X1   g05454(.A1(new_n6457_), .A2(new_n6458_), .B(new_n6316_), .ZN(new_n6459_));
  NAND3_X1   g05455(.A1(new_n6457_), .A2(new_n6458_), .A3(new_n6316_), .ZN(new_n6460_));
  INV_X1     g05456(.I(new_n6460_), .ZN(new_n6461_));
  INV_X1     g05457(.I(\A[963] ), .ZN(new_n6462_));
  NOR2_X1    g05458(.A1(new_n6462_), .A2(\A[962] ), .ZN(new_n6463_));
  INV_X1     g05459(.I(\A[962] ), .ZN(new_n6464_));
  NOR2_X1    g05460(.A1(new_n6464_), .A2(\A[963] ), .ZN(new_n6465_));
  OAI21_X1   g05461(.A1(new_n6463_), .A2(new_n6465_), .B(\A[961] ), .ZN(new_n6466_));
  INV_X1     g05462(.I(\A[961] ), .ZN(new_n6467_));
  NAND2_X1   g05463(.A1(\A[962] ), .A2(\A[963] ), .ZN(new_n6468_));
  INV_X1     g05464(.I(new_n6468_), .ZN(new_n6469_));
  NOR2_X1    g05465(.A1(\A[962] ), .A2(\A[963] ), .ZN(new_n6470_));
  OAI21_X1   g05466(.A1(new_n6469_), .A2(new_n6470_), .B(new_n6467_), .ZN(new_n6471_));
  NAND2_X1   g05467(.A1(new_n6466_), .A2(new_n6471_), .ZN(new_n6472_));
  INV_X1     g05468(.I(\A[966] ), .ZN(new_n6473_));
  NOR2_X1    g05469(.A1(new_n6473_), .A2(\A[965] ), .ZN(new_n6474_));
  INV_X1     g05470(.I(\A[965] ), .ZN(new_n6475_));
  NOR2_X1    g05471(.A1(new_n6475_), .A2(\A[966] ), .ZN(new_n6476_));
  OAI21_X1   g05472(.A1(new_n6474_), .A2(new_n6476_), .B(\A[964] ), .ZN(new_n6477_));
  INV_X1     g05473(.I(\A[964] ), .ZN(new_n6478_));
  NAND2_X1   g05474(.A1(\A[965] ), .A2(\A[966] ), .ZN(new_n6479_));
  INV_X1     g05475(.I(new_n6479_), .ZN(new_n6480_));
  NOR2_X1    g05476(.A1(\A[965] ), .A2(\A[966] ), .ZN(new_n6481_));
  OAI21_X1   g05477(.A1(new_n6480_), .A2(new_n6481_), .B(new_n6478_), .ZN(new_n6482_));
  NAND2_X1   g05478(.A1(new_n6477_), .A2(new_n6482_), .ZN(new_n6483_));
  AOI21_X1   g05479(.A1(new_n6467_), .A2(new_n6468_), .B(new_n6470_), .ZN(new_n6484_));
  AOI21_X1   g05480(.A1(new_n6478_), .A2(new_n6479_), .B(new_n6481_), .ZN(new_n6485_));
  NOR2_X1    g05481(.A1(new_n6484_), .A2(new_n6485_), .ZN(new_n6486_));
  NAND3_X1   g05482(.A1(new_n6472_), .A2(new_n6483_), .A3(new_n6486_), .ZN(new_n6487_));
  INV_X1     g05483(.I(\A[957] ), .ZN(new_n6488_));
  NOR2_X1    g05484(.A1(new_n6488_), .A2(\A[956] ), .ZN(new_n6489_));
  INV_X1     g05485(.I(\A[956] ), .ZN(new_n6490_));
  NOR2_X1    g05486(.A1(new_n6490_), .A2(\A[957] ), .ZN(new_n6491_));
  OAI21_X1   g05487(.A1(new_n6489_), .A2(new_n6491_), .B(\A[955] ), .ZN(new_n6492_));
  INV_X1     g05488(.I(\A[955] ), .ZN(new_n6493_));
  NAND2_X1   g05489(.A1(\A[956] ), .A2(\A[957] ), .ZN(new_n6494_));
  INV_X1     g05490(.I(new_n6494_), .ZN(new_n6495_));
  NOR2_X1    g05491(.A1(\A[956] ), .A2(\A[957] ), .ZN(new_n6496_));
  OAI21_X1   g05492(.A1(new_n6495_), .A2(new_n6496_), .B(new_n6493_), .ZN(new_n6497_));
  NAND2_X1   g05493(.A1(new_n6492_), .A2(new_n6497_), .ZN(new_n6498_));
  INV_X1     g05494(.I(\A[960] ), .ZN(new_n6499_));
  NOR2_X1    g05495(.A1(new_n6499_), .A2(\A[959] ), .ZN(new_n6500_));
  INV_X1     g05496(.I(\A[959] ), .ZN(new_n6501_));
  NOR2_X1    g05497(.A1(new_n6501_), .A2(\A[960] ), .ZN(new_n6502_));
  OAI21_X1   g05498(.A1(new_n6500_), .A2(new_n6502_), .B(\A[958] ), .ZN(new_n6503_));
  INV_X1     g05499(.I(\A[958] ), .ZN(new_n6504_));
  NAND2_X1   g05500(.A1(\A[959] ), .A2(\A[960] ), .ZN(new_n6505_));
  INV_X1     g05501(.I(new_n6505_), .ZN(new_n6506_));
  NOR2_X1    g05502(.A1(\A[959] ), .A2(\A[960] ), .ZN(new_n6507_));
  OAI21_X1   g05503(.A1(new_n6506_), .A2(new_n6507_), .B(new_n6504_), .ZN(new_n6508_));
  NAND2_X1   g05504(.A1(new_n6503_), .A2(new_n6508_), .ZN(new_n6509_));
  AOI21_X1   g05505(.A1(new_n6493_), .A2(new_n6494_), .B(new_n6496_), .ZN(new_n6510_));
  AOI21_X1   g05506(.A1(new_n6504_), .A2(new_n6505_), .B(new_n6507_), .ZN(new_n6511_));
  NOR2_X1    g05507(.A1(new_n6510_), .A2(new_n6511_), .ZN(new_n6512_));
  NAND3_X1   g05508(.A1(new_n6498_), .A2(new_n6509_), .A3(new_n6512_), .ZN(new_n6513_));
  XOR2_X1    g05509(.A1(new_n6487_), .A2(new_n6513_), .Z(new_n6514_));
  INV_X1     g05510(.I(\A[951] ), .ZN(new_n6515_));
  NOR2_X1    g05511(.A1(new_n6515_), .A2(\A[950] ), .ZN(new_n6516_));
  INV_X1     g05512(.I(\A[950] ), .ZN(new_n6517_));
  NOR2_X1    g05513(.A1(new_n6517_), .A2(\A[951] ), .ZN(new_n6518_));
  OAI21_X1   g05514(.A1(new_n6516_), .A2(new_n6518_), .B(\A[949] ), .ZN(new_n6519_));
  INV_X1     g05515(.I(\A[949] ), .ZN(new_n6520_));
  NAND2_X1   g05516(.A1(\A[950] ), .A2(\A[951] ), .ZN(new_n6521_));
  INV_X1     g05517(.I(new_n6521_), .ZN(new_n6522_));
  NOR2_X1    g05518(.A1(\A[950] ), .A2(\A[951] ), .ZN(new_n6523_));
  OAI21_X1   g05519(.A1(new_n6522_), .A2(new_n6523_), .B(new_n6520_), .ZN(new_n6524_));
  NAND2_X1   g05520(.A1(new_n6519_), .A2(new_n6524_), .ZN(new_n6525_));
  INV_X1     g05521(.I(\A[954] ), .ZN(new_n6526_));
  NOR2_X1    g05522(.A1(new_n6526_), .A2(\A[953] ), .ZN(new_n6527_));
  INV_X1     g05523(.I(\A[953] ), .ZN(new_n6528_));
  NOR2_X1    g05524(.A1(new_n6528_), .A2(\A[954] ), .ZN(new_n6529_));
  OAI21_X1   g05525(.A1(new_n6527_), .A2(new_n6529_), .B(\A[952] ), .ZN(new_n6530_));
  INV_X1     g05526(.I(\A[952] ), .ZN(new_n6531_));
  NAND2_X1   g05527(.A1(\A[953] ), .A2(\A[954] ), .ZN(new_n6532_));
  INV_X1     g05528(.I(new_n6532_), .ZN(new_n6533_));
  NOR2_X1    g05529(.A1(\A[953] ), .A2(\A[954] ), .ZN(new_n6534_));
  OAI21_X1   g05530(.A1(new_n6533_), .A2(new_n6534_), .B(new_n6531_), .ZN(new_n6535_));
  NAND2_X1   g05531(.A1(new_n6530_), .A2(new_n6535_), .ZN(new_n6536_));
  AOI21_X1   g05532(.A1(new_n6520_), .A2(new_n6521_), .B(new_n6523_), .ZN(new_n6537_));
  AOI21_X1   g05533(.A1(new_n6531_), .A2(new_n6532_), .B(new_n6534_), .ZN(new_n6538_));
  NOR2_X1    g05534(.A1(new_n6537_), .A2(new_n6538_), .ZN(new_n6539_));
  NAND3_X1   g05535(.A1(new_n6525_), .A2(new_n6536_), .A3(new_n6539_), .ZN(new_n6540_));
  INV_X1     g05536(.I(\A[945] ), .ZN(new_n6541_));
  NOR2_X1    g05537(.A1(new_n6541_), .A2(\A[944] ), .ZN(new_n6542_));
  INV_X1     g05538(.I(\A[944] ), .ZN(new_n6543_));
  NOR2_X1    g05539(.A1(new_n6543_), .A2(\A[945] ), .ZN(new_n6544_));
  OAI21_X1   g05540(.A1(new_n6542_), .A2(new_n6544_), .B(\A[943] ), .ZN(new_n6545_));
  INV_X1     g05541(.I(\A[943] ), .ZN(new_n6546_));
  NAND2_X1   g05542(.A1(\A[944] ), .A2(\A[945] ), .ZN(new_n6547_));
  INV_X1     g05543(.I(new_n6547_), .ZN(new_n6548_));
  NOR2_X1    g05544(.A1(\A[944] ), .A2(\A[945] ), .ZN(new_n6549_));
  OAI21_X1   g05545(.A1(new_n6548_), .A2(new_n6549_), .B(new_n6546_), .ZN(new_n6550_));
  NAND2_X1   g05546(.A1(new_n6545_), .A2(new_n6550_), .ZN(new_n6551_));
  INV_X1     g05547(.I(\A[948] ), .ZN(new_n6552_));
  NOR2_X1    g05548(.A1(new_n6552_), .A2(\A[947] ), .ZN(new_n6553_));
  INV_X1     g05549(.I(\A[947] ), .ZN(new_n6554_));
  NOR2_X1    g05550(.A1(new_n6554_), .A2(\A[948] ), .ZN(new_n6555_));
  OAI21_X1   g05551(.A1(new_n6553_), .A2(new_n6555_), .B(\A[946] ), .ZN(new_n6556_));
  INV_X1     g05552(.I(\A[946] ), .ZN(new_n6557_));
  NAND2_X1   g05553(.A1(\A[947] ), .A2(\A[948] ), .ZN(new_n6558_));
  INV_X1     g05554(.I(new_n6558_), .ZN(new_n6559_));
  NOR2_X1    g05555(.A1(\A[947] ), .A2(\A[948] ), .ZN(new_n6560_));
  OAI21_X1   g05556(.A1(new_n6559_), .A2(new_n6560_), .B(new_n6557_), .ZN(new_n6561_));
  NAND2_X1   g05557(.A1(new_n6556_), .A2(new_n6561_), .ZN(new_n6562_));
  AOI21_X1   g05558(.A1(new_n6546_), .A2(new_n6547_), .B(new_n6549_), .ZN(new_n6563_));
  AOI21_X1   g05559(.A1(new_n6557_), .A2(new_n6558_), .B(new_n6560_), .ZN(new_n6564_));
  NOR2_X1    g05560(.A1(new_n6563_), .A2(new_n6564_), .ZN(new_n6565_));
  NAND3_X1   g05561(.A1(new_n6551_), .A2(new_n6562_), .A3(new_n6565_), .ZN(new_n6566_));
  XOR2_X1    g05562(.A1(new_n6540_), .A2(new_n6566_), .Z(new_n6567_));
  NAND2_X1   g05563(.A1(new_n6514_), .A2(new_n6567_), .ZN(new_n6568_));
  NAND2_X1   g05564(.A1(new_n6490_), .A2(\A[957] ), .ZN(new_n6569_));
  NAND2_X1   g05565(.A1(new_n6488_), .A2(\A[956] ), .ZN(new_n6570_));
  AOI21_X1   g05566(.A1(new_n6569_), .A2(new_n6570_), .B(new_n6493_), .ZN(new_n6571_));
  INV_X1     g05567(.I(new_n6496_), .ZN(new_n6572_));
  AOI21_X1   g05568(.A1(new_n6572_), .A2(new_n6494_), .B(\A[955] ), .ZN(new_n6573_));
  NOR2_X1    g05569(.A1(new_n6573_), .A2(new_n6571_), .ZN(new_n6574_));
  NAND2_X1   g05570(.A1(new_n6501_), .A2(\A[960] ), .ZN(new_n6575_));
  NAND2_X1   g05571(.A1(new_n6499_), .A2(\A[959] ), .ZN(new_n6576_));
  AOI21_X1   g05572(.A1(new_n6575_), .A2(new_n6576_), .B(new_n6504_), .ZN(new_n6577_));
  INV_X1     g05573(.I(new_n6507_), .ZN(new_n6578_));
  AOI21_X1   g05574(.A1(new_n6578_), .A2(new_n6505_), .B(\A[958] ), .ZN(new_n6579_));
  NOR2_X1    g05575(.A1(new_n6579_), .A2(new_n6577_), .ZN(new_n6580_));
  OR2_X2     g05576(.A1(new_n6510_), .A2(new_n6511_), .Z(new_n6581_));
  NOR3_X1    g05577(.A1(new_n6581_), .A2(new_n6574_), .A3(new_n6580_), .ZN(new_n6582_));
  XOR2_X1    g05578(.A1(new_n6582_), .A2(new_n6487_), .Z(new_n6583_));
  NAND2_X1   g05579(.A1(new_n6543_), .A2(\A[945] ), .ZN(new_n6584_));
  NAND2_X1   g05580(.A1(new_n6541_), .A2(\A[944] ), .ZN(new_n6585_));
  AOI21_X1   g05581(.A1(new_n6584_), .A2(new_n6585_), .B(new_n6546_), .ZN(new_n6586_));
  INV_X1     g05582(.I(new_n6549_), .ZN(new_n6587_));
  AOI21_X1   g05583(.A1(new_n6587_), .A2(new_n6547_), .B(\A[943] ), .ZN(new_n6588_));
  NOR2_X1    g05584(.A1(new_n6588_), .A2(new_n6586_), .ZN(new_n6589_));
  NAND2_X1   g05585(.A1(new_n6554_), .A2(\A[948] ), .ZN(new_n6590_));
  NAND2_X1   g05586(.A1(new_n6552_), .A2(\A[947] ), .ZN(new_n6591_));
  AOI21_X1   g05587(.A1(new_n6590_), .A2(new_n6591_), .B(new_n6557_), .ZN(new_n6592_));
  INV_X1     g05588(.I(new_n6560_), .ZN(new_n6593_));
  AOI21_X1   g05589(.A1(new_n6593_), .A2(new_n6558_), .B(\A[946] ), .ZN(new_n6594_));
  NOR2_X1    g05590(.A1(new_n6594_), .A2(new_n6592_), .ZN(new_n6595_));
  INV_X1     g05591(.I(new_n6565_), .ZN(new_n6596_));
  NOR3_X1    g05592(.A1(new_n6596_), .A2(new_n6589_), .A3(new_n6595_), .ZN(new_n6597_));
  XOR2_X1    g05593(.A1(new_n6597_), .A2(new_n6540_), .Z(new_n6598_));
  NAND2_X1   g05594(.A1(new_n6598_), .A2(new_n6583_), .ZN(new_n6599_));
  NAND2_X1   g05595(.A1(new_n6599_), .A2(new_n6568_), .ZN(new_n6600_));
  NOR3_X1    g05596(.A1(new_n6461_), .A2(new_n6459_), .A3(new_n6600_), .ZN(new_n6601_));
  AOI21_X1   g05597(.A1(new_n6411_), .A2(new_n6412_), .B(new_n6414_), .ZN(new_n6602_));
  NOR2_X1    g05598(.A1(new_n6602_), .A2(new_n6442_), .ZN(new_n6603_));
  INV_X1     g05599(.I(new_n6603_), .ZN(new_n6604_));
  NOR2_X1    g05600(.A1(new_n6604_), .A2(new_n6416_), .ZN(new_n6605_));
  NOR2_X1    g05601(.A1(new_n6434_), .A2(new_n6603_), .ZN(new_n6606_));
  OAI21_X1   g05602(.A1(new_n6605_), .A2(new_n6606_), .B(new_n6440_), .ZN(new_n6607_));
  NAND2_X1   g05603(.A1(new_n6434_), .A2(new_n6603_), .ZN(new_n6608_));
  NAND2_X1   g05604(.A1(new_n6604_), .A2(new_n6416_), .ZN(new_n6609_));
  NAND3_X1   g05605(.A1(new_n6609_), .A2(new_n6608_), .A3(new_n6427_), .ZN(new_n6610_));
  AND2_X2    g05606(.A1(new_n6607_), .A2(new_n6610_), .Z(new_n6611_));
  NAND2_X1   g05607(.A1(new_n6441_), .A2(new_n6428_), .ZN(new_n6612_));
  INV_X1     g05608(.I(new_n6389_), .ZN(new_n6613_));
  OAI21_X1   g05609(.A1(new_n6447_), .A2(new_n6613_), .B(new_n6444_), .ZN(new_n6614_));
  NOR3_X1    g05610(.A1(new_n6614_), .A2(new_n6449_), .A3(new_n6612_), .ZN(new_n6615_));
  NOR2_X1    g05611(.A1(new_n6385_), .A2(new_n6387_), .ZN(new_n6616_));
  INV_X1     g05612(.I(new_n6616_), .ZN(new_n6617_));
  NOR2_X1    g05613(.A1(new_n6617_), .A2(new_n6372_), .ZN(new_n6618_));
  NOR2_X1    g05614(.A1(new_n6396_), .A2(new_n6616_), .ZN(new_n6619_));
  OAI21_X1   g05615(.A1(new_n6618_), .A2(new_n6619_), .B(new_n6402_), .ZN(new_n6620_));
  NAND2_X1   g05616(.A1(new_n6396_), .A2(new_n6616_), .ZN(new_n6621_));
  NAND2_X1   g05617(.A1(new_n6617_), .A2(new_n6372_), .ZN(new_n6622_));
  NAND3_X1   g05618(.A1(new_n6622_), .A2(new_n6621_), .A3(new_n6383_), .ZN(new_n6623_));
  NAND2_X1   g05619(.A1(new_n6620_), .A2(new_n6623_), .ZN(new_n6624_));
  XOR2_X1    g05620(.A1(new_n6615_), .A2(new_n6624_), .Z(new_n6625_));
  NAND2_X1   g05621(.A1(new_n6625_), .A2(new_n6611_), .ZN(new_n6626_));
  AOI21_X1   g05622(.A1(new_n6622_), .A2(new_n6621_), .B(new_n6383_), .ZN(new_n6627_));
  NOR3_X1    g05623(.A1(new_n6618_), .A2(new_n6619_), .A3(new_n6402_), .ZN(new_n6628_));
  NOR2_X1    g05624(.A1(new_n6628_), .A2(new_n6627_), .ZN(new_n6629_));
  NAND2_X1   g05625(.A1(new_n6607_), .A2(new_n6610_), .ZN(new_n6630_));
  NOR2_X1    g05626(.A1(new_n6449_), .A2(new_n6612_), .ZN(new_n6631_));
  XOR2_X1    g05627(.A1(new_n6385_), .A2(new_n6387_), .Z(new_n6632_));
  NAND2_X1   g05628(.A1(new_n6384_), .A2(new_n6632_), .ZN(new_n6633_));
  OAI21_X1   g05629(.A1(new_n6389_), .A2(new_n6616_), .B(new_n6447_), .ZN(new_n6634_));
  NAND2_X1   g05630(.A1(new_n6634_), .A2(new_n6633_), .ZN(new_n6635_));
  NAND2_X1   g05631(.A1(new_n6403_), .A2(new_n6613_), .ZN(new_n6636_));
  NOR2_X1    g05632(.A1(new_n6636_), .A2(new_n6444_), .ZN(new_n6637_));
  NAND4_X1   g05633(.A1(new_n6630_), .A2(new_n6635_), .A3(new_n6631_), .A4(new_n6637_), .ZN(new_n6638_));
  NAND2_X1   g05634(.A1(new_n6638_), .A2(new_n6629_), .ZN(new_n6639_));
  NAND2_X1   g05635(.A1(new_n6639_), .A2(new_n6615_), .ZN(new_n6640_));
  NOR2_X1    g05636(.A1(new_n6302_), .A2(new_n6308_), .ZN(new_n6641_));
  NOR2_X1    g05637(.A1(new_n6284_), .A2(new_n6295_), .ZN(new_n6642_));
  NOR2_X1    g05638(.A1(new_n6641_), .A2(new_n6642_), .ZN(new_n6643_));
  NOR2_X1    g05639(.A1(new_n6352_), .A2(new_n6358_), .ZN(new_n6644_));
  NAND2_X1   g05640(.A1(new_n6644_), .A2(new_n6344_), .ZN(new_n6645_));
  NOR2_X1    g05641(.A1(new_n6327_), .A2(new_n6338_), .ZN(new_n6646_));
  NOR2_X1    g05642(.A1(new_n6646_), .A2(new_n6644_), .ZN(new_n6647_));
  NAND4_X1   g05643(.A1(new_n6643_), .A2(new_n6647_), .A3(new_n6645_), .A4(new_n6314_), .ZN(new_n6648_));
  NOR2_X1    g05644(.A1(new_n6340_), .A2(new_n6342_), .ZN(new_n6649_));
  NAND2_X1   g05645(.A1(new_n6327_), .A2(new_n6649_), .ZN(new_n6650_));
  INV_X1     g05646(.I(new_n6649_), .ZN(new_n6651_));
  NAND2_X1   g05647(.A1(new_n6651_), .A2(new_n6352_), .ZN(new_n6652_));
  AOI21_X1   g05648(.A1(new_n6652_), .A2(new_n6650_), .B(new_n6358_), .ZN(new_n6653_));
  NOR2_X1    g05649(.A1(new_n6651_), .A2(new_n6352_), .ZN(new_n6654_));
  NOR2_X1    g05650(.A1(new_n6327_), .A2(new_n6649_), .ZN(new_n6655_));
  NOR3_X1    g05651(.A1(new_n6654_), .A2(new_n6655_), .A3(new_n6338_), .ZN(new_n6656_));
  NOR2_X1    g05652(.A1(new_n6656_), .A2(new_n6653_), .ZN(new_n6657_));
  INV_X1     g05653(.I(new_n6313_), .ZN(new_n6658_));
  NOR2_X1    g05654(.A1(new_n6658_), .A2(new_n6284_), .ZN(new_n6659_));
  NOR2_X1    g05655(.A1(new_n6302_), .A2(new_n6313_), .ZN(new_n6660_));
  OAI21_X1   g05656(.A1(new_n6659_), .A2(new_n6660_), .B(new_n6308_), .ZN(new_n6661_));
  NAND2_X1   g05657(.A1(new_n6302_), .A2(new_n6313_), .ZN(new_n6662_));
  NAND2_X1   g05658(.A1(new_n6658_), .A2(new_n6284_), .ZN(new_n6663_));
  NAND3_X1   g05659(.A1(new_n6663_), .A2(new_n6662_), .A3(new_n6295_), .ZN(new_n6664_));
  NAND2_X1   g05660(.A1(new_n6661_), .A2(new_n6664_), .ZN(new_n6665_));
  NOR2_X1    g05661(.A1(new_n6310_), .A2(new_n6360_), .ZN(new_n6666_));
  XOR2_X1    g05662(.A1(new_n6340_), .A2(new_n6342_), .Z(new_n6667_));
  NAND2_X1   g05663(.A1(new_n6644_), .A2(new_n6667_), .ZN(new_n6668_));
  OAI21_X1   g05664(.A1(new_n6344_), .A2(new_n6649_), .B(new_n6339_), .ZN(new_n6669_));
  NAND2_X1   g05665(.A1(new_n6669_), .A2(new_n6668_), .ZN(new_n6670_));
  NAND2_X1   g05666(.A1(new_n6646_), .A2(new_n6345_), .ZN(new_n6671_));
  NOR2_X1    g05667(.A1(new_n6671_), .A2(new_n6314_), .ZN(new_n6672_));
  NAND3_X1   g05668(.A1(new_n6670_), .A2(new_n6666_), .A3(new_n6672_), .ZN(new_n6673_));
  NAND4_X1   g05669(.A1(new_n6673_), .A2(new_n6648_), .A3(new_n6657_), .A4(new_n6665_), .ZN(new_n6674_));
  NOR2_X1    g05670(.A1(new_n6454_), .A2(new_n6316_), .ZN(new_n6675_));
  NAND2_X1   g05671(.A1(new_n6643_), .A2(new_n6314_), .ZN(new_n6676_));
  NOR2_X1    g05672(.A1(new_n6676_), .A2(new_n6445_), .ZN(new_n6677_));
  NAND2_X1   g05673(.A1(new_n6647_), .A2(new_n6645_), .ZN(new_n6678_));
  NOR2_X1    g05674(.A1(new_n6450_), .A2(new_n6678_), .ZN(new_n6679_));
  NOR2_X1    g05675(.A1(new_n6361_), .A2(new_n6405_), .ZN(new_n6680_));
  OAI22_X1   g05676(.A1(new_n6679_), .A2(new_n6680_), .B1(new_n6675_), .B2(new_n6677_), .ZN(new_n6681_));
  NOR2_X1    g05677(.A1(new_n6681_), .A2(new_n6674_), .ZN(new_n6682_));
  NAND2_X1   g05678(.A1(new_n6682_), .A2(new_n6640_), .ZN(new_n6683_));
  INV_X1     g05679(.I(new_n6682_), .ZN(new_n6684_));
  NAND3_X1   g05680(.A1(new_n6684_), .A2(new_n6615_), .A3(new_n6639_), .ZN(new_n6685_));
  AOI21_X1   g05681(.A1(new_n6685_), .A2(new_n6683_), .B(new_n6626_), .ZN(new_n6686_));
  NAND2_X1   g05682(.A1(new_n6574_), .A2(new_n6512_), .ZN(new_n6687_));
  NAND2_X1   g05683(.A1(new_n6581_), .A2(new_n6498_), .ZN(new_n6688_));
  AOI21_X1   g05684(.A1(new_n6688_), .A2(new_n6687_), .B(new_n6509_), .ZN(new_n6689_));
  NOR2_X1    g05685(.A1(new_n6581_), .A2(new_n6498_), .ZN(new_n6690_));
  NOR2_X1    g05686(.A1(new_n6574_), .A2(new_n6512_), .ZN(new_n6691_));
  NOR3_X1    g05687(.A1(new_n6690_), .A2(new_n6691_), .A3(new_n6580_), .ZN(new_n6692_));
  OR2_X2     g05688(.A1(new_n6692_), .A2(new_n6689_), .Z(new_n6693_));
  NOR2_X1    g05689(.A1(new_n6487_), .A2(new_n6513_), .ZN(new_n6694_));
  INV_X1     g05690(.I(new_n6483_), .ZN(new_n6695_));
  INV_X1     g05691(.I(new_n6486_), .ZN(new_n6696_));
  NOR2_X1    g05692(.A1(new_n6696_), .A2(new_n6472_), .ZN(new_n6697_));
  NAND2_X1   g05693(.A1(new_n6464_), .A2(\A[963] ), .ZN(new_n6698_));
  NAND2_X1   g05694(.A1(new_n6462_), .A2(\A[962] ), .ZN(new_n6699_));
  AOI21_X1   g05695(.A1(new_n6698_), .A2(new_n6699_), .B(new_n6467_), .ZN(new_n6700_));
  INV_X1     g05696(.I(new_n6470_), .ZN(new_n6701_));
  AOI21_X1   g05697(.A1(new_n6701_), .A2(new_n6468_), .B(\A[961] ), .ZN(new_n6702_));
  NOR2_X1    g05698(.A1(new_n6702_), .A2(new_n6700_), .ZN(new_n6703_));
  NOR2_X1    g05699(.A1(new_n6703_), .A2(new_n6486_), .ZN(new_n6704_));
  OAI21_X1   g05700(.A1(new_n6697_), .A2(new_n6704_), .B(new_n6695_), .ZN(new_n6705_));
  NAND2_X1   g05701(.A1(new_n6703_), .A2(new_n6486_), .ZN(new_n6706_));
  NAND2_X1   g05702(.A1(new_n6696_), .A2(new_n6472_), .ZN(new_n6707_));
  NAND3_X1   g05703(.A1(new_n6707_), .A2(new_n6706_), .A3(new_n6483_), .ZN(new_n6708_));
  NOR2_X1    g05704(.A1(new_n6695_), .A2(new_n6472_), .ZN(new_n6709_));
  NOR2_X1    g05705(.A1(new_n6703_), .A2(new_n6483_), .ZN(new_n6710_));
  OAI21_X1   g05706(.A1(new_n6709_), .A2(new_n6710_), .B(new_n6486_), .ZN(new_n6711_));
  NAND3_X1   g05707(.A1(new_n6711_), .A2(new_n6705_), .A3(new_n6708_), .ZN(new_n6712_));
  XOR2_X1    g05708(.A1(new_n6712_), .A2(new_n6694_), .Z(new_n6713_));
  NOR2_X1    g05709(.A1(new_n6713_), .A2(new_n6693_), .ZN(new_n6714_));
  INV_X1     g05710(.I(new_n6714_), .ZN(new_n6715_));
  AOI21_X1   g05711(.A1(new_n6707_), .A2(new_n6706_), .B(new_n6483_), .ZN(new_n6716_));
  NOR3_X1    g05712(.A1(new_n6697_), .A2(new_n6704_), .A3(new_n6695_), .ZN(new_n6717_));
  NAND2_X1   g05713(.A1(new_n6703_), .A2(new_n6483_), .ZN(new_n6718_));
  NAND2_X1   g05714(.A1(new_n6695_), .A2(new_n6472_), .ZN(new_n6719_));
  AOI21_X1   g05715(.A1(new_n6719_), .A2(new_n6718_), .B(new_n6696_), .ZN(new_n6720_));
  NOR3_X1    g05716(.A1(new_n6720_), .A2(new_n6716_), .A3(new_n6717_), .ZN(new_n6721_));
  NOR2_X1    g05717(.A1(new_n6692_), .A2(new_n6689_), .ZN(new_n6722_));
  NAND2_X1   g05718(.A1(new_n6498_), .A2(new_n6509_), .ZN(new_n6723_));
  NAND2_X1   g05719(.A1(new_n6574_), .A2(new_n6580_), .ZN(new_n6724_));
  NOR2_X1    g05720(.A1(new_n6581_), .A2(new_n6574_), .ZN(new_n6725_));
  AOI22_X1   g05721(.A1(new_n6723_), .A2(new_n6724_), .B1(new_n6725_), .B2(new_n6509_), .ZN(new_n6726_));
  NAND4_X1   g05722(.A1(new_n6726_), .A2(new_n6472_), .A3(new_n6483_), .A4(new_n6486_), .ZN(new_n6727_));
  NOR2_X1    g05723(.A1(new_n6727_), .A2(new_n6722_), .ZN(new_n6728_));
  OAI21_X1   g05724(.A1(new_n6728_), .A2(new_n6721_), .B(new_n6694_), .ZN(new_n6729_));
  NOR2_X1    g05725(.A1(new_n6540_), .A2(new_n6566_), .ZN(new_n6730_));
  INV_X1     g05726(.I(new_n6536_), .ZN(new_n6731_));
  OR2_X2     g05727(.A1(new_n6537_), .A2(new_n6538_), .Z(new_n6732_));
  NOR2_X1    g05728(.A1(new_n6732_), .A2(new_n6525_), .ZN(new_n6733_));
  NAND2_X1   g05729(.A1(new_n6517_), .A2(\A[951] ), .ZN(new_n6734_));
  NAND2_X1   g05730(.A1(new_n6515_), .A2(\A[950] ), .ZN(new_n6735_));
  AOI21_X1   g05731(.A1(new_n6734_), .A2(new_n6735_), .B(new_n6520_), .ZN(new_n6736_));
  INV_X1     g05732(.I(new_n6523_), .ZN(new_n6737_));
  AOI21_X1   g05733(.A1(new_n6737_), .A2(new_n6521_), .B(\A[949] ), .ZN(new_n6738_));
  NOR2_X1    g05734(.A1(new_n6738_), .A2(new_n6736_), .ZN(new_n6739_));
  NOR2_X1    g05735(.A1(new_n6739_), .A2(new_n6539_), .ZN(new_n6740_));
  OAI21_X1   g05736(.A1(new_n6733_), .A2(new_n6740_), .B(new_n6731_), .ZN(new_n6741_));
  NAND2_X1   g05737(.A1(new_n6739_), .A2(new_n6539_), .ZN(new_n6742_));
  NAND2_X1   g05738(.A1(new_n6732_), .A2(new_n6525_), .ZN(new_n6743_));
  NAND3_X1   g05739(.A1(new_n6743_), .A2(new_n6742_), .A3(new_n6536_), .ZN(new_n6744_));
  NAND2_X1   g05740(.A1(new_n6741_), .A2(new_n6744_), .ZN(new_n6745_));
  NAND2_X1   g05741(.A1(new_n6739_), .A2(new_n6536_), .ZN(new_n6746_));
  NOR2_X1    g05742(.A1(new_n6739_), .A2(new_n6536_), .ZN(new_n6747_));
  INV_X1     g05743(.I(new_n6747_), .ZN(new_n6748_));
  AOI21_X1   g05744(.A1(new_n6748_), .A2(new_n6746_), .B(new_n6732_), .ZN(new_n6749_));
  NOR3_X1    g05745(.A1(new_n6745_), .A2(new_n6730_), .A3(new_n6749_), .ZN(new_n6750_));
  NAND2_X1   g05746(.A1(new_n6589_), .A2(new_n6565_), .ZN(new_n6751_));
  NAND2_X1   g05747(.A1(new_n6596_), .A2(new_n6551_), .ZN(new_n6752_));
  AOI21_X1   g05748(.A1(new_n6752_), .A2(new_n6751_), .B(new_n6562_), .ZN(new_n6753_));
  INV_X1     g05749(.I(new_n6751_), .ZN(new_n6754_));
  NOR2_X1    g05750(.A1(new_n6589_), .A2(new_n6565_), .ZN(new_n6755_));
  NOR3_X1    g05751(.A1(new_n6754_), .A2(new_n6755_), .A3(new_n6595_), .ZN(new_n6756_));
  NOR2_X1    g05752(.A1(new_n6756_), .A2(new_n6753_), .ZN(new_n6757_));
  NAND2_X1   g05753(.A1(new_n6551_), .A2(new_n6562_), .ZN(new_n6758_));
  NAND2_X1   g05754(.A1(new_n6589_), .A2(new_n6595_), .ZN(new_n6759_));
  NAND2_X1   g05755(.A1(new_n6759_), .A2(new_n6758_), .ZN(new_n6760_));
  NOR3_X1    g05756(.A1(new_n6596_), .A2(new_n6589_), .A3(new_n6595_), .ZN(new_n6761_));
  NAND4_X1   g05757(.A1(new_n6760_), .A2(new_n6525_), .A3(new_n6536_), .A4(new_n6539_), .ZN(new_n6762_));
  INV_X1     g05758(.I(new_n6762_), .ZN(new_n6763_));
  NOR4_X1    g05759(.A1(new_n6599_), .A2(new_n6750_), .A3(new_n6757_), .A4(new_n6763_), .ZN(new_n6764_));
  NAND2_X1   g05760(.A1(new_n6764_), .A2(new_n6729_), .ZN(new_n6765_));
  NOR2_X1    g05761(.A1(new_n6574_), .A2(new_n6580_), .ZN(new_n6766_));
  NOR2_X1    g05762(.A1(new_n6498_), .A2(new_n6509_), .ZN(new_n6767_));
  NAND2_X1   g05763(.A1(new_n6498_), .A2(new_n6512_), .ZN(new_n6768_));
  OAI22_X1   g05764(.A1(new_n6766_), .A2(new_n6767_), .B1(new_n6768_), .B2(new_n6580_), .ZN(new_n6769_));
  NOR4_X1    g05765(.A1(new_n6769_), .A2(new_n6703_), .A3(new_n6695_), .A4(new_n6696_), .ZN(new_n6770_));
  NAND2_X1   g05766(.A1(new_n6693_), .A2(new_n6770_), .ZN(new_n6771_));
  NAND2_X1   g05767(.A1(new_n6771_), .A2(new_n6712_), .ZN(new_n6772_));
  NOR2_X1    g05768(.A1(new_n6514_), .A2(new_n6567_), .ZN(new_n6773_));
  INV_X1     g05769(.I(new_n6730_), .ZN(new_n6774_));
  AOI21_X1   g05770(.A1(new_n6743_), .A2(new_n6742_), .B(new_n6536_), .ZN(new_n6775_));
  NOR3_X1    g05771(.A1(new_n6733_), .A2(new_n6740_), .A3(new_n6731_), .ZN(new_n6776_));
  NOR2_X1    g05772(.A1(new_n6776_), .A2(new_n6775_), .ZN(new_n6777_));
  INV_X1     g05773(.I(new_n6746_), .ZN(new_n6778_));
  OAI21_X1   g05774(.A1(new_n6778_), .A2(new_n6747_), .B(new_n6539_), .ZN(new_n6779_));
  NAND3_X1   g05775(.A1(new_n6777_), .A2(new_n6774_), .A3(new_n6779_), .ZN(new_n6780_));
  INV_X1     g05776(.I(new_n6757_), .ZN(new_n6781_));
  NAND4_X1   g05777(.A1(new_n6773_), .A2(new_n6780_), .A3(new_n6781_), .A4(new_n6762_), .ZN(new_n6782_));
  NAND3_X1   g05778(.A1(new_n6782_), .A2(new_n6772_), .A3(new_n6694_), .ZN(new_n6783_));
  NAND2_X1   g05779(.A1(new_n6783_), .A2(new_n6765_), .ZN(new_n6784_));
  NAND2_X1   g05780(.A1(new_n6784_), .A2(new_n6715_), .ZN(new_n6785_));
  NAND3_X1   g05781(.A1(new_n6714_), .A2(new_n6783_), .A3(new_n6765_), .ZN(new_n6786_));
  NAND2_X1   g05782(.A1(new_n6785_), .A2(new_n6786_), .ZN(new_n6787_));
  OAI21_X1   g05783(.A1(new_n6787_), .A2(new_n6601_), .B(new_n6686_), .ZN(new_n6788_));
  NOR3_X1    g05784(.A1(new_n6750_), .A2(new_n6763_), .A3(new_n6757_), .ZN(new_n6789_));
  NOR2_X1    g05785(.A1(new_n6789_), .A2(new_n6773_), .ZN(new_n6790_));
  NAND4_X1   g05786(.A1(new_n6728_), .A2(new_n6722_), .A3(new_n6694_), .A4(new_n6712_), .ZN(new_n6791_));
  OAI21_X1   g05787(.A1(new_n6790_), .A2(new_n6791_), .B(new_n6782_), .ZN(new_n6792_));
  NAND3_X1   g05788(.A1(new_n6551_), .A2(new_n6562_), .A3(new_n6565_), .ZN(new_n6793_));
  NAND2_X1   g05789(.A1(new_n6760_), .A2(new_n6793_), .ZN(new_n6794_));
  NOR4_X1    g05790(.A1(new_n6794_), .A2(new_n6739_), .A3(new_n6731_), .A4(new_n6732_), .ZN(new_n6795_));
  NAND2_X1   g05791(.A1(new_n6537_), .A2(new_n6538_), .ZN(new_n6796_));
  NAND3_X1   g05792(.A1(new_n6525_), .A2(new_n6536_), .A3(new_n6796_), .ZN(new_n6797_));
  NAND2_X1   g05793(.A1(new_n6797_), .A2(new_n6732_), .ZN(new_n6798_));
  NOR2_X1    g05794(.A1(new_n6589_), .A2(new_n6595_), .ZN(new_n6799_));
  NAND2_X1   g05795(.A1(new_n6563_), .A2(new_n6564_), .ZN(new_n6800_));
  AOI21_X1   g05796(.A1(new_n6799_), .A2(new_n6800_), .B(new_n6565_), .ZN(new_n6801_));
  XNOR2_X1   g05797(.A1(new_n6801_), .A2(new_n6798_), .ZN(new_n6802_));
  AOI21_X1   g05798(.A1(new_n6777_), .A2(new_n6779_), .B(new_n6730_), .ZN(new_n6803_));
  NOR2_X1    g05799(.A1(new_n6803_), .A2(new_n6757_), .ZN(new_n6804_));
  OAI21_X1   g05800(.A1(new_n6804_), .A2(new_n6795_), .B(new_n6802_), .ZN(new_n6805_));
  NAND2_X1   g05801(.A1(new_n6484_), .A2(new_n6485_), .ZN(new_n6806_));
  NAND3_X1   g05802(.A1(new_n6472_), .A2(new_n6483_), .A3(new_n6806_), .ZN(new_n6807_));
  NAND2_X1   g05803(.A1(new_n6807_), .A2(new_n6696_), .ZN(new_n6808_));
  NAND2_X1   g05804(.A1(new_n6510_), .A2(new_n6511_), .ZN(new_n6809_));
  AOI21_X1   g05805(.A1(new_n6766_), .A2(new_n6809_), .B(new_n6512_), .ZN(new_n6810_));
  XNOR2_X1   g05806(.A1(new_n6810_), .A2(new_n6808_), .ZN(new_n6811_));
  INV_X1     g05807(.I(new_n6694_), .ZN(new_n6812_));
  AOI21_X1   g05808(.A1(new_n6712_), .A2(new_n6812_), .B(new_n6722_), .ZN(new_n6813_));
  OAI21_X1   g05809(.A1(new_n6813_), .A2(new_n6770_), .B(new_n6811_), .ZN(new_n6814_));
  XOR2_X1    g05810(.A1(new_n6805_), .A2(new_n6814_), .Z(new_n6815_));
  NAND2_X1   g05811(.A1(new_n6815_), .A2(new_n6792_), .ZN(new_n6816_));
  NAND3_X1   g05812(.A1(new_n6781_), .A2(new_n6780_), .A3(new_n6762_), .ZN(new_n6817_));
  NAND2_X1   g05813(.A1(new_n6817_), .A2(new_n6599_), .ZN(new_n6818_));
  NOR4_X1    g05814(.A1(new_n6771_), .A2(new_n6693_), .A3(new_n6812_), .A4(new_n6721_), .ZN(new_n6819_));
  AOI21_X1   g05815(.A1(new_n6818_), .A2(new_n6819_), .B(new_n6764_), .ZN(new_n6820_));
  NAND2_X1   g05816(.A1(new_n6805_), .A2(new_n6814_), .ZN(new_n6821_));
  AOI21_X1   g05817(.A1(new_n6758_), .A2(new_n6759_), .B(new_n6761_), .ZN(new_n6822_));
  NAND4_X1   g05818(.A1(new_n6822_), .A2(new_n6525_), .A3(new_n6536_), .A4(new_n6539_), .ZN(new_n6823_));
  XOR2_X1    g05819(.A1(new_n6801_), .A2(new_n6798_), .Z(new_n6824_));
  OAI21_X1   g05820(.A1(new_n6745_), .A2(new_n6749_), .B(new_n6774_), .ZN(new_n6825_));
  NAND2_X1   g05821(.A1(new_n6781_), .A2(new_n6825_), .ZN(new_n6826_));
  AOI21_X1   g05822(.A1(new_n6826_), .A2(new_n6823_), .B(new_n6824_), .ZN(new_n6827_));
  XOR2_X1    g05823(.A1(new_n6810_), .A2(new_n6808_), .Z(new_n6828_));
  OAI21_X1   g05824(.A1(new_n6721_), .A2(new_n6694_), .B(new_n6693_), .ZN(new_n6829_));
  AOI21_X1   g05825(.A1(new_n6829_), .A2(new_n6727_), .B(new_n6828_), .ZN(new_n6830_));
  NAND2_X1   g05826(.A1(new_n6827_), .A2(new_n6830_), .ZN(new_n6831_));
  NAND2_X1   g05827(.A1(new_n6831_), .A2(new_n6821_), .ZN(new_n6832_));
  NAND2_X1   g05828(.A1(new_n6832_), .A2(new_n6820_), .ZN(new_n6833_));
  NAND2_X1   g05829(.A1(new_n6816_), .A2(new_n6833_), .ZN(new_n6834_));
  NAND2_X1   g05830(.A1(new_n6681_), .A2(new_n6674_), .ZN(new_n6835_));
  NAND4_X1   g05831(.A1(new_n6404_), .A2(new_n6453_), .A3(new_n6390_), .A4(new_n6444_), .ZN(new_n6836_));
  NOR4_X1    g05832(.A1(new_n6638_), .A2(new_n6630_), .A3(new_n6836_), .A4(new_n6624_), .ZN(new_n6837_));
  AOI21_X1   g05833(.A1(new_n6835_), .A2(new_n6837_), .B(new_n6682_), .ZN(new_n6838_));
  INV_X1     g05834(.I(new_n6673_), .ZN(new_n6839_));
  NOR4_X1    g05835(.A1(new_n6310_), .A2(new_n6360_), .A3(new_n6346_), .A4(new_n6315_), .ZN(new_n6840_));
  OAI21_X1   g05836(.A1(new_n6654_), .A2(new_n6655_), .B(new_n6338_), .ZN(new_n6841_));
  NAND3_X1   g05837(.A1(new_n6652_), .A2(new_n6650_), .A3(new_n6358_), .ZN(new_n6842_));
  NAND2_X1   g05838(.A1(new_n6841_), .A2(new_n6842_), .ZN(new_n6843_));
  OAI21_X1   g05839(.A1(new_n6840_), .A2(new_n6843_), .B(new_n6665_), .ZN(new_n6844_));
  AOI21_X1   g05840(.A1(new_n6646_), .A2(new_n6345_), .B(new_n6649_), .ZN(new_n6845_));
  NAND2_X1   g05841(.A1(new_n6311_), .A2(new_n6312_), .ZN(new_n6846_));
  AOI21_X1   g05842(.A1(new_n6641_), .A2(new_n6846_), .B(new_n6313_), .ZN(new_n6847_));
  NOR2_X1    g05843(.A1(new_n6845_), .A2(new_n6847_), .ZN(new_n6848_));
  NAND2_X1   g05844(.A1(new_n6844_), .A2(new_n6848_), .ZN(new_n6849_));
  NAND2_X1   g05845(.A1(new_n6648_), .A2(new_n6657_), .ZN(new_n6850_));
  INV_X1     g05846(.I(new_n6848_), .ZN(new_n6851_));
  NAND3_X1   g05847(.A1(new_n6850_), .A2(new_n6665_), .A3(new_n6851_), .ZN(new_n6852_));
  AOI21_X1   g05848(.A1(new_n6849_), .A2(new_n6852_), .B(new_n6839_), .ZN(new_n6853_));
  AOI21_X1   g05849(.A1(new_n6850_), .A2(new_n6665_), .B(new_n6851_), .ZN(new_n6854_));
  NOR2_X1    g05850(.A1(new_n6844_), .A2(new_n6848_), .ZN(new_n6855_));
  NOR3_X1    g05851(.A1(new_n6855_), .A2(new_n6854_), .A3(new_n6673_), .ZN(new_n6856_));
  NOR2_X1    g05852(.A1(new_n6856_), .A2(new_n6853_), .ZN(new_n6857_));
  NAND3_X1   g05853(.A1(new_n6635_), .A2(new_n6631_), .A3(new_n6637_), .ZN(new_n6858_));
  NAND2_X1   g05854(.A1(new_n6836_), .A2(new_n6629_), .ZN(new_n6859_));
  AOI21_X1   g05855(.A1(new_n6403_), .A2(new_n6613_), .B(new_n6616_), .ZN(new_n6860_));
  NAND2_X1   g05856(.A1(new_n6602_), .A2(new_n6442_), .ZN(new_n6861_));
  AOI21_X1   g05857(.A1(new_n6451_), .A2(new_n6861_), .B(new_n6603_), .ZN(new_n6862_));
  NOR2_X1    g05858(.A1(new_n6860_), .A2(new_n6862_), .ZN(new_n6863_));
  INV_X1     g05859(.I(new_n6863_), .ZN(new_n6864_));
  AOI21_X1   g05860(.A1(new_n6859_), .A2(new_n6630_), .B(new_n6864_), .ZN(new_n6865_));
  OAI21_X1   g05861(.A1(new_n6615_), .A2(new_n6624_), .B(new_n6630_), .ZN(new_n6866_));
  NOR2_X1    g05862(.A1(new_n6866_), .A2(new_n6863_), .ZN(new_n6867_));
  OAI21_X1   g05863(.A1(new_n6867_), .A2(new_n6865_), .B(new_n6858_), .ZN(new_n6868_));
  INV_X1     g05864(.I(new_n6858_), .ZN(new_n6869_));
  NAND2_X1   g05865(.A1(new_n6866_), .A2(new_n6863_), .ZN(new_n6870_));
  NAND3_X1   g05866(.A1(new_n6859_), .A2(new_n6630_), .A3(new_n6864_), .ZN(new_n6871_));
  NAND3_X1   g05867(.A1(new_n6870_), .A2(new_n6871_), .A3(new_n6869_), .ZN(new_n6872_));
  NAND2_X1   g05868(.A1(new_n6868_), .A2(new_n6872_), .ZN(new_n6873_));
  NAND2_X1   g05869(.A1(new_n6857_), .A2(new_n6873_), .ZN(new_n6874_));
  OAI21_X1   g05870(.A1(new_n6855_), .A2(new_n6854_), .B(new_n6673_), .ZN(new_n6875_));
  NAND3_X1   g05871(.A1(new_n6849_), .A2(new_n6852_), .A3(new_n6839_), .ZN(new_n6876_));
  NAND2_X1   g05872(.A1(new_n6875_), .A2(new_n6876_), .ZN(new_n6877_));
  AOI21_X1   g05873(.A1(new_n6870_), .A2(new_n6871_), .B(new_n6869_), .ZN(new_n6878_));
  NOR3_X1    g05874(.A1(new_n6867_), .A2(new_n6865_), .A3(new_n6858_), .ZN(new_n6879_));
  NOR2_X1    g05875(.A1(new_n6879_), .A2(new_n6878_), .ZN(new_n6880_));
  NAND2_X1   g05876(.A1(new_n6880_), .A2(new_n6877_), .ZN(new_n6881_));
  AOI21_X1   g05877(.A1(new_n6874_), .A2(new_n6881_), .B(new_n6838_), .ZN(new_n6882_));
  NAND2_X1   g05878(.A1(new_n6835_), .A2(new_n6837_), .ZN(new_n6883_));
  NAND2_X1   g05879(.A1(new_n6883_), .A2(new_n6684_), .ZN(new_n6884_));
  NAND2_X1   g05880(.A1(new_n6877_), .A2(new_n6873_), .ZN(new_n6885_));
  NAND4_X1   g05881(.A1(new_n6875_), .A2(new_n6876_), .A3(new_n6868_), .A4(new_n6872_), .ZN(new_n6886_));
  AOI21_X1   g05882(.A1(new_n6885_), .A2(new_n6886_), .B(new_n6884_), .ZN(new_n6887_));
  NOR2_X1    g05883(.A1(new_n6882_), .A2(new_n6887_), .ZN(new_n6888_));
  XOR2_X1    g05884(.A1(new_n6888_), .A2(new_n6834_), .Z(new_n6889_));
  OAI21_X1   g05885(.A1(new_n6882_), .A2(new_n6887_), .B(new_n6834_), .ZN(new_n6890_));
  AOI21_X1   g05886(.A1(new_n6821_), .A2(new_n6831_), .B(new_n6792_), .ZN(new_n6891_));
  AOI21_X1   g05887(.A1(new_n6792_), .A2(new_n6815_), .B(new_n6891_), .ZN(new_n6892_));
  NOR2_X1    g05888(.A1(new_n6880_), .A2(new_n6877_), .ZN(new_n6893_));
  NOR2_X1    g05889(.A1(new_n6857_), .A2(new_n6873_), .ZN(new_n6894_));
  OAI21_X1   g05890(.A1(new_n6893_), .A2(new_n6894_), .B(new_n6884_), .ZN(new_n6895_));
  NOR2_X1    g05891(.A1(new_n6857_), .A2(new_n6880_), .ZN(new_n6896_));
  NOR4_X1    g05892(.A1(new_n6853_), .A2(new_n6856_), .A3(new_n6879_), .A4(new_n6878_), .ZN(new_n6897_));
  OAI21_X1   g05893(.A1(new_n6896_), .A2(new_n6897_), .B(new_n6838_), .ZN(new_n6898_));
  NAND3_X1   g05894(.A1(new_n6895_), .A2(new_n6892_), .A3(new_n6898_), .ZN(new_n6899_));
  NAND2_X1   g05895(.A1(new_n6890_), .A2(new_n6899_), .ZN(new_n6900_));
  NAND2_X1   g05896(.A1(new_n6900_), .A2(new_n6788_), .ZN(new_n6901_));
  OAI21_X1   g05897(.A1(new_n6788_), .A2(new_n6889_), .B(new_n6901_), .ZN(new_n6902_));
  INV_X1     g05898(.I(new_n6902_), .ZN(new_n6903_));
  INV_X1     g05899(.I(\A[27] ), .ZN(new_n6904_));
  NOR2_X1    g05900(.A1(new_n6904_), .A2(\A[26] ), .ZN(new_n6905_));
  INV_X1     g05901(.I(\A[26] ), .ZN(new_n6906_));
  NOR2_X1    g05902(.A1(new_n6906_), .A2(\A[27] ), .ZN(new_n6907_));
  OAI21_X1   g05903(.A1(new_n6905_), .A2(new_n6907_), .B(\A[25] ), .ZN(new_n6908_));
  INV_X1     g05904(.I(\A[25] ), .ZN(new_n6909_));
  NOR2_X1    g05905(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n6910_));
  AND2_X2    g05906(.A1(\A[26] ), .A2(\A[27] ), .Z(new_n6911_));
  OAI21_X1   g05907(.A1(new_n6911_), .A2(new_n6910_), .B(new_n6909_), .ZN(new_n6912_));
  NAND2_X1   g05908(.A1(new_n6908_), .A2(new_n6912_), .ZN(new_n6913_));
  INV_X1     g05909(.I(\A[30] ), .ZN(new_n6914_));
  NOR2_X1    g05910(.A1(new_n6914_), .A2(\A[29] ), .ZN(new_n6915_));
  INV_X1     g05911(.I(\A[29] ), .ZN(new_n6916_));
  NOR2_X1    g05912(.A1(new_n6916_), .A2(\A[30] ), .ZN(new_n6917_));
  OAI21_X1   g05913(.A1(new_n6915_), .A2(new_n6917_), .B(\A[28] ), .ZN(new_n6918_));
  INV_X1     g05914(.I(\A[28] ), .ZN(new_n6919_));
  NAND2_X1   g05915(.A1(\A[29] ), .A2(\A[30] ), .ZN(new_n6920_));
  INV_X1     g05916(.I(new_n6920_), .ZN(new_n6921_));
  NOR2_X1    g05917(.A1(\A[29] ), .A2(\A[30] ), .ZN(new_n6922_));
  OAI21_X1   g05918(.A1(new_n6921_), .A2(new_n6922_), .B(new_n6919_), .ZN(new_n6923_));
  NAND2_X1   g05919(.A1(new_n6918_), .A2(new_n6923_), .ZN(new_n6924_));
  AOI21_X1   g05920(.A1(\A[26] ), .A2(\A[27] ), .B(\A[25] ), .ZN(new_n6925_));
  AOI21_X1   g05921(.A1(\A[29] ), .A2(\A[30] ), .B(\A[28] ), .ZN(new_n6926_));
  OAI22_X1   g05922(.A1(new_n6910_), .A2(new_n6925_), .B1(new_n6926_), .B2(new_n6922_), .ZN(new_n6927_));
  XOR2_X1    g05923(.A1(new_n6924_), .A2(new_n6913_), .Z(new_n6929_));
  INV_X1     g05924(.I(\A[19] ), .ZN(new_n6930_));
  INV_X1     g05925(.I(\A[20] ), .ZN(new_n6931_));
  NAND2_X1   g05926(.A1(new_n6931_), .A2(\A[21] ), .ZN(new_n6932_));
  INV_X1     g05927(.I(\A[21] ), .ZN(new_n6933_));
  NAND2_X1   g05928(.A1(new_n6933_), .A2(\A[20] ), .ZN(new_n6934_));
  AOI21_X1   g05929(.A1(new_n6932_), .A2(new_n6934_), .B(new_n6930_), .ZN(new_n6935_));
  NOR2_X1    g05930(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n6936_));
  INV_X1     g05931(.I(new_n6936_), .ZN(new_n6937_));
  NAND2_X1   g05932(.A1(\A[20] ), .A2(\A[21] ), .ZN(new_n6938_));
  AOI21_X1   g05933(.A1(new_n6937_), .A2(new_n6938_), .B(\A[19] ), .ZN(new_n6939_));
  NOR2_X1    g05934(.A1(new_n6939_), .A2(new_n6935_), .ZN(new_n6940_));
  INV_X1     g05935(.I(\A[24] ), .ZN(new_n6941_));
  NOR2_X1    g05936(.A1(new_n6941_), .A2(\A[23] ), .ZN(new_n6942_));
  INV_X1     g05937(.I(\A[23] ), .ZN(new_n6943_));
  NOR2_X1    g05938(.A1(new_n6943_), .A2(\A[24] ), .ZN(new_n6944_));
  OAI21_X1   g05939(.A1(new_n6942_), .A2(new_n6944_), .B(\A[22] ), .ZN(new_n6945_));
  INV_X1     g05940(.I(\A[22] ), .ZN(new_n6946_));
  NAND2_X1   g05941(.A1(\A[23] ), .A2(\A[24] ), .ZN(new_n6947_));
  INV_X1     g05942(.I(new_n6947_), .ZN(new_n6948_));
  NOR2_X1    g05943(.A1(\A[23] ), .A2(\A[24] ), .ZN(new_n6949_));
  OAI21_X1   g05944(.A1(new_n6948_), .A2(new_n6949_), .B(new_n6946_), .ZN(new_n6950_));
  NAND2_X1   g05945(.A1(new_n6945_), .A2(new_n6950_), .ZN(new_n6951_));
  AOI21_X1   g05946(.A1(\A[20] ), .A2(\A[21] ), .B(\A[19] ), .ZN(new_n6952_));
  AOI21_X1   g05947(.A1(\A[23] ), .A2(\A[24] ), .B(\A[22] ), .ZN(new_n6953_));
  OAI22_X1   g05948(.A1(new_n6936_), .A2(new_n6952_), .B1(new_n6953_), .B2(new_n6949_), .ZN(new_n6954_));
  INV_X1     g05949(.I(new_n6954_), .ZN(new_n6955_));
  XOR2_X1    g05950(.A1(new_n6940_), .A2(new_n6951_), .Z(new_n6956_));
  XOR2_X1    g05951(.A1(new_n6956_), .A2(new_n6929_), .Z(new_n6957_));
  INV_X1     g05952(.I(\A[15] ), .ZN(new_n6958_));
  NOR2_X1    g05953(.A1(new_n6958_), .A2(\A[14] ), .ZN(new_n6959_));
  INV_X1     g05954(.I(\A[14] ), .ZN(new_n6960_));
  NOR2_X1    g05955(.A1(new_n6960_), .A2(\A[15] ), .ZN(new_n6961_));
  OAI21_X1   g05956(.A1(new_n6959_), .A2(new_n6961_), .B(\A[13] ), .ZN(new_n6962_));
  INV_X1     g05957(.I(\A[13] ), .ZN(new_n6963_));
  NOR2_X1    g05958(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n6964_));
  NAND2_X1   g05959(.A1(\A[14] ), .A2(\A[15] ), .ZN(new_n6965_));
  INV_X1     g05960(.I(new_n6965_), .ZN(new_n6966_));
  OAI21_X1   g05961(.A1(new_n6966_), .A2(new_n6964_), .B(new_n6963_), .ZN(new_n6967_));
  NAND2_X1   g05962(.A1(new_n6962_), .A2(new_n6967_), .ZN(new_n6968_));
  INV_X1     g05963(.I(\A[18] ), .ZN(new_n6969_));
  NOR2_X1    g05964(.A1(new_n6969_), .A2(\A[17] ), .ZN(new_n6970_));
  INV_X1     g05965(.I(\A[17] ), .ZN(new_n6971_));
  NOR2_X1    g05966(.A1(new_n6971_), .A2(\A[18] ), .ZN(new_n6972_));
  OAI21_X1   g05967(.A1(new_n6970_), .A2(new_n6972_), .B(\A[16] ), .ZN(new_n6973_));
  INV_X1     g05968(.I(\A[16] ), .ZN(new_n6974_));
  NAND2_X1   g05969(.A1(\A[17] ), .A2(\A[18] ), .ZN(new_n6975_));
  INV_X1     g05970(.I(new_n6975_), .ZN(new_n6976_));
  NOR2_X1    g05971(.A1(\A[17] ), .A2(\A[18] ), .ZN(new_n6977_));
  OAI21_X1   g05972(.A1(new_n6976_), .A2(new_n6977_), .B(new_n6974_), .ZN(new_n6978_));
  NAND2_X1   g05973(.A1(new_n6973_), .A2(new_n6978_), .ZN(new_n6979_));
  AOI21_X1   g05974(.A1(\A[14] ), .A2(\A[15] ), .B(\A[13] ), .ZN(new_n6980_));
  NOR2_X1    g05975(.A1(new_n6980_), .A2(new_n6964_), .ZN(new_n6981_));
  AOI21_X1   g05976(.A1(\A[17] ), .A2(\A[18] ), .B(\A[16] ), .ZN(new_n6982_));
  NOR2_X1    g05977(.A1(new_n6982_), .A2(new_n6977_), .ZN(new_n6983_));
  NOR2_X1    g05978(.A1(new_n6981_), .A2(new_n6983_), .ZN(new_n6984_));
  XOR2_X1    g05979(.A1(new_n6968_), .A2(new_n6979_), .Z(new_n6985_));
  INV_X1     g05980(.I(\A[9] ), .ZN(new_n6986_));
  NOR2_X1    g05981(.A1(new_n6986_), .A2(\A[8] ), .ZN(new_n6987_));
  INV_X1     g05982(.I(\A[8] ), .ZN(new_n6988_));
  NOR2_X1    g05983(.A1(new_n6988_), .A2(\A[9] ), .ZN(new_n6989_));
  OAI21_X1   g05984(.A1(new_n6987_), .A2(new_n6989_), .B(\A[7] ), .ZN(new_n6990_));
  INV_X1     g05985(.I(\A[7] ), .ZN(new_n6991_));
  NOR2_X1    g05986(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n6992_));
  NAND2_X1   g05987(.A1(\A[8] ), .A2(\A[9] ), .ZN(new_n6993_));
  INV_X1     g05988(.I(new_n6993_), .ZN(new_n6994_));
  OAI21_X1   g05989(.A1(new_n6994_), .A2(new_n6992_), .B(new_n6991_), .ZN(new_n6995_));
  NAND2_X1   g05990(.A1(new_n6990_), .A2(new_n6995_), .ZN(new_n6996_));
  INV_X1     g05991(.I(\A[12] ), .ZN(new_n6997_));
  NOR2_X1    g05992(.A1(new_n6997_), .A2(\A[11] ), .ZN(new_n6998_));
  INV_X1     g05993(.I(\A[11] ), .ZN(new_n6999_));
  NOR2_X1    g05994(.A1(new_n6999_), .A2(\A[12] ), .ZN(new_n7000_));
  OAI21_X1   g05995(.A1(new_n6998_), .A2(new_n7000_), .B(\A[10] ), .ZN(new_n7001_));
  INV_X1     g05996(.I(\A[10] ), .ZN(new_n7002_));
  NAND2_X1   g05997(.A1(\A[11] ), .A2(\A[12] ), .ZN(new_n7003_));
  INV_X1     g05998(.I(new_n7003_), .ZN(new_n7004_));
  NOR2_X1    g05999(.A1(\A[11] ), .A2(\A[12] ), .ZN(new_n7005_));
  OAI21_X1   g06000(.A1(new_n7004_), .A2(new_n7005_), .B(new_n7002_), .ZN(new_n7006_));
  NAND2_X1   g06001(.A1(new_n7001_), .A2(new_n7006_), .ZN(new_n7007_));
  AOI21_X1   g06002(.A1(\A[8] ), .A2(\A[9] ), .B(\A[7] ), .ZN(new_n7008_));
  AOI21_X1   g06003(.A1(\A[11] ), .A2(\A[12] ), .B(\A[10] ), .ZN(new_n7009_));
  OAI22_X1   g06004(.A1(new_n6992_), .A2(new_n7008_), .B1(new_n7009_), .B2(new_n7005_), .ZN(new_n7010_));
  INV_X1     g06005(.I(new_n7010_), .ZN(new_n7011_));
  XOR2_X1    g06006(.A1(new_n6996_), .A2(new_n7007_), .Z(new_n7012_));
  XOR2_X1    g06007(.A1(new_n6985_), .A2(new_n7012_), .Z(new_n7013_));
  INV_X1     g06008(.I(\A[994] ), .ZN(new_n7014_));
  NOR2_X1    g06009(.A1(\A[995] ), .A2(\A[996] ), .ZN(new_n7015_));
  NAND2_X1   g06010(.A1(\A[995] ), .A2(\A[996] ), .ZN(new_n7016_));
  AOI21_X1   g06011(.A1(new_n7014_), .A2(new_n7016_), .B(new_n7015_), .ZN(new_n7017_));
  INV_X1     g06012(.I(\A[991] ), .ZN(new_n7018_));
  NOR2_X1    g06013(.A1(\A[992] ), .A2(\A[993] ), .ZN(new_n7019_));
  NAND2_X1   g06014(.A1(\A[992] ), .A2(\A[993] ), .ZN(new_n7020_));
  AOI21_X1   g06015(.A1(new_n7018_), .A2(new_n7020_), .B(new_n7019_), .ZN(new_n7021_));
  XNOR2_X1   g06016(.A1(new_n7017_), .A2(new_n7021_), .ZN(new_n7022_));
  INV_X1     g06017(.I(\A[0] ), .ZN(new_n7023_));
  INV_X1     g06018(.I(\A[6] ), .ZN(new_n7024_));
  XOR2_X1    g06019(.A1(\A[1] ), .A2(\A[2] ), .Z(new_n7025_));
  NAND2_X1   g06020(.A1(new_n7025_), .A2(new_n7024_), .ZN(new_n7026_));
  XNOR2_X1   g06021(.A1(\A[1] ), .A2(\A[2] ), .ZN(new_n7027_));
  NAND2_X1   g06022(.A1(new_n7027_), .A2(\A[6] ), .ZN(new_n7028_));
  AOI21_X1   g06023(.A1(new_n7028_), .A2(new_n7026_), .B(new_n7023_), .ZN(new_n7029_));
  NAND2_X1   g06024(.A1(new_n7023_), .A2(\A[1] ), .ZN(new_n7030_));
  INV_X1     g06025(.I(\A[1] ), .ZN(new_n7031_));
  NAND2_X1   g06026(.A1(new_n7031_), .A2(\A[0] ), .ZN(new_n7032_));
  AOI21_X1   g06027(.A1(new_n7030_), .A2(new_n7032_), .B(\A[2] ), .ZN(new_n7033_));
  INV_X1     g06028(.I(\A[2] ), .ZN(new_n7034_));
  NOR2_X1    g06029(.A1(new_n7031_), .A2(\A[0] ), .ZN(new_n7035_));
  NOR2_X1    g06030(.A1(new_n7023_), .A2(\A[1] ), .ZN(new_n7036_));
  NOR3_X1    g06031(.A1(new_n7035_), .A2(new_n7036_), .A3(new_n7034_), .ZN(new_n7037_));
  OAI21_X1   g06032(.A1(new_n7033_), .A2(new_n7037_), .B(\A[6] ), .ZN(new_n7038_));
  INV_X1     g06033(.I(\A[3] ), .ZN(new_n7039_));
  INV_X1     g06034(.I(\A[4] ), .ZN(new_n7040_));
  NAND2_X1   g06035(.A1(new_n7040_), .A2(\A[5] ), .ZN(new_n7041_));
  INV_X1     g06036(.I(\A[5] ), .ZN(new_n7042_));
  NAND2_X1   g06037(.A1(new_n7042_), .A2(\A[4] ), .ZN(new_n7043_));
  AOI21_X1   g06038(.A1(new_n7041_), .A2(new_n7043_), .B(new_n7039_), .ZN(new_n7044_));
  NAND2_X1   g06039(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n7045_));
  NOR2_X1    g06040(.A1(\A[4] ), .A2(\A[5] ), .ZN(new_n7046_));
  INV_X1     g06041(.I(new_n7046_), .ZN(new_n7047_));
  AOI21_X1   g06042(.A1(new_n7047_), .A2(new_n7045_), .B(\A[3] ), .ZN(new_n7048_));
  NOR2_X1    g06043(.A1(new_n7048_), .A2(new_n7044_), .ZN(new_n7049_));
  INV_X1     g06044(.I(\A[997] ), .ZN(new_n7050_));
  INV_X1     g06045(.I(\A[998] ), .ZN(new_n7051_));
  NAND2_X1   g06046(.A1(new_n7051_), .A2(\A[999] ), .ZN(new_n7052_));
  INV_X1     g06047(.I(\A[999] ), .ZN(new_n7053_));
  NAND2_X1   g06048(.A1(new_n7053_), .A2(\A[998] ), .ZN(new_n7054_));
  AOI21_X1   g06049(.A1(new_n7052_), .A2(new_n7054_), .B(new_n7050_), .ZN(new_n7055_));
  NAND2_X1   g06050(.A1(\A[998] ), .A2(\A[999] ), .ZN(new_n7056_));
  NAND2_X1   g06051(.A1(new_n7051_), .A2(new_n7053_), .ZN(new_n7057_));
  AOI21_X1   g06052(.A1(new_n7057_), .A2(new_n7056_), .B(\A[997] ), .ZN(new_n7058_));
  NOR2_X1    g06053(.A1(new_n7058_), .A2(new_n7055_), .ZN(new_n7059_));
  NOR2_X1    g06054(.A1(new_n7049_), .A2(new_n7059_), .ZN(new_n7060_));
  NAND2_X1   g06055(.A1(new_n7060_), .A2(new_n7038_), .ZN(new_n7061_));
  OAI21_X1   g06056(.A1(new_n7035_), .A2(new_n7036_), .B(new_n7034_), .ZN(new_n7062_));
  NAND3_X1   g06057(.A1(new_n7030_), .A2(new_n7032_), .A3(\A[2] ), .ZN(new_n7063_));
  AOI21_X1   g06058(.A1(new_n7062_), .A2(new_n7063_), .B(new_n7024_), .ZN(new_n7064_));
  OAI22_X1   g06059(.A1(new_n7044_), .A2(new_n7048_), .B1(new_n7058_), .B2(new_n7055_), .ZN(new_n7065_));
  NAND2_X1   g06060(.A1(new_n7065_), .A2(new_n7064_), .ZN(new_n7066_));
  AOI21_X1   g06061(.A1(new_n7061_), .A2(new_n7066_), .B(new_n7029_), .ZN(new_n7067_));
  NOR2_X1    g06062(.A1(new_n7027_), .A2(\A[6] ), .ZN(new_n7068_));
  NOR2_X1    g06063(.A1(new_n7025_), .A2(new_n7024_), .ZN(new_n7069_));
  OAI21_X1   g06064(.A1(new_n7068_), .A2(new_n7069_), .B(\A[0] ), .ZN(new_n7070_));
  NOR2_X1    g06065(.A1(new_n7065_), .A2(new_n7064_), .ZN(new_n7071_));
  INV_X1     g06066(.I(new_n7066_), .ZN(new_n7072_));
  NOR3_X1    g06067(.A1(new_n7072_), .A2(new_n7070_), .A3(new_n7071_), .ZN(new_n7073_));
  OAI21_X1   g06068(.A1(new_n7073_), .A2(new_n7067_), .B(new_n7022_), .ZN(new_n7074_));
  INV_X1     g06069(.I(new_n7022_), .ZN(new_n7075_));
  OAI21_X1   g06070(.A1(new_n7072_), .A2(new_n7071_), .B(new_n7070_), .ZN(new_n7076_));
  NAND3_X1   g06071(.A1(new_n7061_), .A2(new_n7029_), .A3(new_n7066_), .ZN(new_n7077_));
  NAND3_X1   g06072(.A1(new_n7076_), .A2(new_n7077_), .A3(new_n7075_), .ZN(new_n7078_));
  NAND2_X1   g06073(.A1(new_n7074_), .A2(new_n7078_), .ZN(new_n7079_));
  XOR2_X1    g06074(.A1(new_n7079_), .A2(new_n7013_), .Z(new_n7080_));
  NAND2_X1   g06075(.A1(new_n7080_), .A2(new_n6957_), .ZN(new_n7081_));
  XOR2_X1    g06076(.A1(new_n7079_), .A2(new_n7013_), .Z(new_n7082_));
  OAI21_X1   g06077(.A1(new_n6957_), .A2(new_n7082_), .B(new_n7081_), .ZN(new_n7083_));
  INV_X1     g06078(.I(\A[55] ), .ZN(new_n7084_));
  INV_X1     g06079(.I(\A[56] ), .ZN(new_n7085_));
  NAND2_X1   g06080(.A1(new_n7085_), .A2(\A[57] ), .ZN(new_n7086_));
  INV_X1     g06081(.I(\A[57] ), .ZN(new_n7087_));
  NAND2_X1   g06082(.A1(new_n7087_), .A2(\A[56] ), .ZN(new_n7088_));
  AOI21_X1   g06083(.A1(new_n7086_), .A2(new_n7088_), .B(new_n7084_), .ZN(new_n7089_));
  NOR2_X1    g06084(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n7090_));
  INV_X1     g06085(.I(new_n7090_), .ZN(new_n7091_));
  NAND2_X1   g06086(.A1(\A[56] ), .A2(\A[57] ), .ZN(new_n7092_));
  AOI21_X1   g06087(.A1(new_n7091_), .A2(new_n7092_), .B(\A[55] ), .ZN(new_n7093_));
  NOR2_X1    g06088(.A1(new_n7093_), .A2(new_n7089_), .ZN(new_n7094_));
  INV_X1     g06089(.I(\A[60] ), .ZN(new_n7095_));
  NOR2_X1    g06090(.A1(new_n7095_), .A2(\A[59] ), .ZN(new_n7096_));
  INV_X1     g06091(.I(\A[59] ), .ZN(new_n7097_));
  NOR2_X1    g06092(.A1(new_n7097_), .A2(\A[60] ), .ZN(new_n7098_));
  OAI21_X1   g06093(.A1(new_n7096_), .A2(new_n7098_), .B(\A[58] ), .ZN(new_n7099_));
  INV_X1     g06094(.I(\A[58] ), .ZN(new_n7100_));
  NAND2_X1   g06095(.A1(\A[59] ), .A2(\A[60] ), .ZN(new_n7101_));
  INV_X1     g06096(.I(new_n7101_), .ZN(new_n7102_));
  NOR2_X1    g06097(.A1(\A[59] ), .A2(\A[60] ), .ZN(new_n7103_));
  OAI21_X1   g06098(.A1(new_n7102_), .A2(new_n7103_), .B(new_n7100_), .ZN(new_n7104_));
  NAND2_X1   g06099(.A1(new_n7099_), .A2(new_n7104_), .ZN(new_n7105_));
  AOI21_X1   g06100(.A1(new_n7084_), .A2(new_n7092_), .B(new_n7090_), .ZN(new_n7106_));
  AOI21_X1   g06101(.A1(new_n7100_), .A2(new_n7101_), .B(new_n7103_), .ZN(new_n7107_));
  NOR2_X1    g06102(.A1(new_n7106_), .A2(new_n7107_), .ZN(new_n7108_));
  XOR2_X1    g06103(.A1(new_n7094_), .A2(new_n7105_), .Z(new_n7109_));
  INV_X1     g06104(.I(new_n7109_), .ZN(new_n7110_));
  INV_X1     g06105(.I(\A[67] ), .ZN(new_n7111_));
  INV_X1     g06106(.I(\A[68] ), .ZN(new_n7112_));
  NAND2_X1   g06107(.A1(new_n7112_), .A2(\A[69] ), .ZN(new_n7113_));
  INV_X1     g06108(.I(\A[69] ), .ZN(new_n7114_));
  NAND2_X1   g06109(.A1(new_n7114_), .A2(\A[68] ), .ZN(new_n7115_));
  AOI21_X1   g06110(.A1(new_n7113_), .A2(new_n7115_), .B(new_n7111_), .ZN(new_n7116_));
  NOR2_X1    g06111(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n7117_));
  INV_X1     g06112(.I(new_n7117_), .ZN(new_n7118_));
  NAND2_X1   g06113(.A1(\A[68] ), .A2(\A[69] ), .ZN(new_n7119_));
  AOI21_X1   g06114(.A1(new_n7118_), .A2(new_n7119_), .B(\A[67] ), .ZN(new_n7120_));
  NOR2_X1    g06115(.A1(new_n7120_), .A2(new_n7116_), .ZN(new_n7121_));
  INV_X1     g06116(.I(\A[72] ), .ZN(new_n7122_));
  NOR2_X1    g06117(.A1(new_n7122_), .A2(\A[71] ), .ZN(new_n7123_));
  INV_X1     g06118(.I(\A[71] ), .ZN(new_n7124_));
  NOR2_X1    g06119(.A1(new_n7124_), .A2(\A[72] ), .ZN(new_n7125_));
  OAI21_X1   g06120(.A1(new_n7123_), .A2(new_n7125_), .B(\A[70] ), .ZN(new_n7126_));
  INV_X1     g06121(.I(\A[70] ), .ZN(new_n7127_));
  NAND2_X1   g06122(.A1(\A[71] ), .A2(\A[72] ), .ZN(new_n7128_));
  INV_X1     g06123(.I(new_n7128_), .ZN(new_n7129_));
  NOR2_X1    g06124(.A1(\A[71] ), .A2(\A[72] ), .ZN(new_n7130_));
  OAI21_X1   g06125(.A1(new_n7129_), .A2(new_n7130_), .B(new_n7127_), .ZN(new_n7131_));
  NAND2_X1   g06126(.A1(new_n7126_), .A2(new_n7131_), .ZN(new_n7132_));
  AOI21_X1   g06127(.A1(new_n7111_), .A2(new_n7119_), .B(new_n7117_), .ZN(new_n7133_));
  AOI21_X1   g06128(.A1(new_n7127_), .A2(new_n7128_), .B(new_n7130_), .ZN(new_n7134_));
  NOR2_X1    g06129(.A1(new_n7133_), .A2(new_n7134_), .ZN(new_n7135_));
  XOR2_X1    g06130(.A1(new_n7121_), .A2(new_n7132_), .Z(new_n7136_));
  INV_X1     g06131(.I(\A[75] ), .ZN(new_n7137_));
  NOR2_X1    g06132(.A1(new_n7137_), .A2(\A[74] ), .ZN(new_n7138_));
  INV_X1     g06133(.I(\A[74] ), .ZN(new_n7139_));
  NOR2_X1    g06134(.A1(new_n7139_), .A2(\A[75] ), .ZN(new_n7140_));
  OAI21_X1   g06135(.A1(new_n7138_), .A2(new_n7140_), .B(\A[73] ), .ZN(new_n7141_));
  INV_X1     g06136(.I(\A[73] ), .ZN(new_n7142_));
  NOR2_X1    g06137(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n7143_));
  AND2_X2    g06138(.A1(\A[74] ), .A2(\A[75] ), .Z(new_n7144_));
  OAI21_X1   g06139(.A1(new_n7144_), .A2(new_n7143_), .B(new_n7142_), .ZN(new_n7145_));
  NAND2_X1   g06140(.A1(new_n7141_), .A2(new_n7145_), .ZN(new_n7146_));
  INV_X1     g06141(.I(\A[76] ), .ZN(new_n7147_));
  INV_X1     g06142(.I(\A[77] ), .ZN(new_n7148_));
  NAND2_X1   g06143(.A1(new_n7148_), .A2(\A[78] ), .ZN(new_n7149_));
  INV_X1     g06144(.I(\A[78] ), .ZN(new_n7150_));
  NAND2_X1   g06145(.A1(new_n7150_), .A2(\A[77] ), .ZN(new_n7151_));
  AOI21_X1   g06146(.A1(new_n7149_), .A2(new_n7151_), .B(new_n7147_), .ZN(new_n7152_));
  NAND2_X1   g06147(.A1(\A[77] ), .A2(\A[78] ), .ZN(new_n7153_));
  NOR2_X1    g06148(.A1(\A[77] ), .A2(\A[78] ), .ZN(new_n7154_));
  INV_X1     g06149(.I(new_n7154_), .ZN(new_n7155_));
  AOI21_X1   g06150(.A1(new_n7155_), .A2(new_n7153_), .B(\A[76] ), .ZN(new_n7156_));
  NOR2_X1    g06151(.A1(new_n7156_), .A2(new_n7152_), .ZN(new_n7157_));
  AOI21_X1   g06152(.A1(\A[74] ), .A2(\A[75] ), .B(\A[73] ), .ZN(new_n7158_));
  AOI21_X1   g06153(.A1(\A[77] ), .A2(\A[78] ), .B(\A[76] ), .ZN(new_n7159_));
  OAI22_X1   g06154(.A1(new_n7143_), .A2(new_n7158_), .B1(new_n7159_), .B2(new_n7154_), .ZN(new_n7160_));
  INV_X1     g06155(.I(new_n7160_), .ZN(new_n7161_));
  XOR2_X1    g06156(.A1(new_n7157_), .A2(new_n7146_), .Z(new_n7162_));
  INV_X1     g06157(.I(\A[63] ), .ZN(new_n7163_));
  NOR2_X1    g06158(.A1(new_n7163_), .A2(\A[62] ), .ZN(new_n7164_));
  INV_X1     g06159(.I(\A[62] ), .ZN(new_n7165_));
  NOR2_X1    g06160(.A1(new_n7165_), .A2(\A[63] ), .ZN(new_n7166_));
  OAI21_X1   g06161(.A1(new_n7164_), .A2(new_n7166_), .B(\A[61] ), .ZN(new_n7167_));
  INV_X1     g06162(.I(\A[61] ), .ZN(new_n7168_));
  NOR2_X1    g06163(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n7169_));
  AND2_X2    g06164(.A1(\A[62] ), .A2(\A[63] ), .Z(new_n7170_));
  OAI21_X1   g06165(.A1(new_n7170_), .A2(new_n7169_), .B(new_n7168_), .ZN(new_n7171_));
  NAND2_X1   g06166(.A1(new_n7167_), .A2(new_n7171_), .ZN(new_n7172_));
  INV_X1     g06167(.I(\A[64] ), .ZN(new_n7173_));
  INV_X1     g06168(.I(\A[65] ), .ZN(new_n7174_));
  NAND2_X1   g06169(.A1(new_n7174_), .A2(\A[66] ), .ZN(new_n7175_));
  INV_X1     g06170(.I(\A[66] ), .ZN(new_n7176_));
  NAND2_X1   g06171(.A1(new_n7176_), .A2(\A[65] ), .ZN(new_n7177_));
  AOI21_X1   g06172(.A1(new_n7175_), .A2(new_n7177_), .B(new_n7173_), .ZN(new_n7178_));
  NAND2_X1   g06173(.A1(\A[65] ), .A2(\A[66] ), .ZN(new_n7179_));
  NOR2_X1    g06174(.A1(\A[65] ), .A2(\A[66] ), .ZN(new_n7180_));
  INV_X1     g06175(.I(new_n7180_), .ZN(new_n7181_));
  AOI21_X1   g06176(.A1(new_n7181_), .A2(new_n7179_), .B(\A[64] ), .ZN(new_n7182_));
  NOR2_X1    g06177(.A1(new_n7182_), .A2(new_n7178_), .ZN(new_n7183_));
  AOI21_X1   g06178(.A1(\A[62] ), .A2(\A[63] ), .B(\A[61] ), .ZN(new_n7184_));
  AOI21_X1   g06179(.A1(\A[65] ), .A2(\A[66] ), .B(\A[64] ), .ZN(new_n7185_));
  OAI22_X1   g06180(.A1(new_n7169_), .A2(new_n7184_), .B1(new_n7185_), .B2(new_n7180_), .ZN(new_n7186_));
  INV_X1     g06181(.I(new_n7186_), .ZN(new_n7187_));
  XOR2_X1    g06182(.A1(new_n7183_), .A2(new_n7172_), .Z(new_n7188_));
  XOR2_X1    g06183(.A1(new_n7162_), .A2(new_n7188_), .Z(new_n7189_));
  NAND2_X1   g06184(.A1(new_n7189_), .A2(new_n7136_), .ZN(new_n7190_));
  NOR2_X1    g06185(.A1(new_n7114_), .A2(\A[68] ), .ZN(new_n7191_));
  NOR2_X1    g06186(.A1(new_n7112_), .A2(\A[69] ), .ZN(new_n7192_));
  OAI21_X1   g06187(.A1(new_n7191_), .A2(new_n7192_), .B(\A[67] ), .ZN(new_n7193_));
  INV_X1     g06188(.I(new_n7119_), .ZN(new_n7194_));
  OAI21_X1   g06189(.A1(new_n7194_), .A2(new_n7117_), .B(new_n7111_), .ZN(new_n7195_));
  NAND2_X1   g06190(.A1(new_n7193_), .A2(new_n7195_), .ZN(new_n7196_));
  XOR2_X1    g06191(.A1(new_n7196_), .A2(new_n7132_), .Z(new_n7197_));
  XNOR2_X1   g06192(.A1(new_n7162_), .A2(new_n7188_), .ZN(new_n7198_));
  NAND2_X1   g06193(.A1(new_n7198_), .A2(new_n7197_), .ZN(new_n7199_));
  AOI21_X1   g06194(.A1(new_n7199_), .A2(new_n7190_), .B(new_n7110_), .ZN(new_n7200_));
  NOR2_X1    g06195(.A1(new_n7198_), .A2(new_n7197_), .ZN(new_n7201_));
  NOR2_X1    g06196(.A1(new_n7189_), .A2(new_n7136_), .ZN(new_n7202_));
  NOR3_X1    g06197(.A1(new_n7201_), .A2(new_n7202_), .A3(new_n7109_), .ZN(new_n7203_));
  INV_X1     g06198(.I(\A[34] ), .ZN(new_n7204_));
  NOR2_X1    g06199(.A1(\A[35] ), .A2(\A[36] ), .ZN(new_n7205_));
  NAND2_X1   g06200(.A1(\A[35] ), .A2(\A[36] ), .ZN(new_n7206_));
  AOI21_X1   g06201(.A1(new_n7204_), .A2(new_n7206_), .B(new_n7205_), .ZN(new_n7207_));
  INV_X1     g06202(.I(\A[31] ), .ZN(new_n7208_));
  NOR2_X1    g06203(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n7209_));
  NAND2_X1   g06204(.A1(\A[32] ), .A2(\A[33] ), .ZN(new_n7210_));
  AOI21_X1   g06205(.A1(new_n7208_), .A2(new_n7210_), .B(new_n7209_), .ZN(new_n7211_));
  XOR2_X1    g06206(.A1(new_n7207_), .A2(new_n7211_), .Z(new_n7212_));
  NOR2_X1    g06207(.A1(\A[47] ), .A2(\A[48] ), .ZN(new_n7213_));
  AOI21_X1   g06208(.A1(\A[47] ), .A2(\A[48] ), .B(\A[46] ), .ZN(new_n7214_));
  NOR2_X1    g06209(.A1(new_n7214_), .A2(new_n7213_), .ZN(new_n7215_));
  NOR2_X1    g06210(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n7216_));
  AOI21_X1   g06211(.A1(\A[44] ), .A2(\A[45] ), .B(\A[43] ), .ZN(new_n7217_));
  NOR2_X1    g06212(.A1(new_n7217_), .A2(new_n7216_), .ZN(new_n7218_));
  XOR2_X1    g06213(.A1(new_n7215_), .A2(new_n7218_), .Z(new_n7219_));
  INV_X1     g06214(.I(new_n7219_), .ZN(new_n7220_));
  NOR2_X1    g06215(.A1(\A[53] ), .A2(\A[54] ), .ZN(new_n7221_));
  AOI21_X1   g06216(.A1(\A[53] ), .A2(\A[54] ), .B(\A[52] ), .ZN(new_n7222_));
  NOR2_X1    g06217(.A1(new_n7222_), .A2(new_n7221_), .ZN(new_n7223_));
  NOR2_X1    g06218(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n7224_));
  AOI21_X1   g06219(.A1(\A[50] ), .A2(\A[51] ), .B(\A[49] ), .ZN(new_n7225_));
  NOR2_X1    g06220(.A1(new_n7225_), .A2(new_n7224_), .ZN(new_n7226_));
  XNOR2_X1   g06221(.A1(new_n7223_), .A2(new_n7226_), .ZN(new_n7227_));
  NOR2_X1    g06222(.A1(\A[41] ), .A2(\A[42] ), .ZN(new_n7228_));
  AOI21_X1   g06223(.A1(\A[41] ), .A2(\A[42] ), .B(\A[40] ), .ZN(new_n7229_));
  NOR2_X1    g06224(.A1(new_n7229_), .A2(new_n7228_), .ZN(new_n7230_));
  NOR2_X1    g06225(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n7231_));
  AOI21_X1   g06226(.A1(\A[38] ), .A2(\A[39] ), .B(\A[37] ), .ZN(new_n7232_));
  NOR2_X1    g06227(.A1(new_n7232_), .A2(new_n7231_), .ZN(new_n7233_));
  XOR2_X1    g06228(.A1(new_n7230_), .A2(new_n7233_), .Z(new_n7234_));
  XNOR2_X1   g06229(.A1(new_n7227_), .A2(new_n7234_), .ZN(new_n7235_));
  NAND2_X1   g06230(.A1(new_n7235_), .A2(new_n7220_), .ZN(new_n7236_));
  XOR2_X1    g06231(.A1(new_n7227_), .A2(new_n7234_), .Z(new_n7237_));
  NAND2_X1   g06232(.A1(new_n7237_), .A2(new_n7219_), .ZN(new_n7238_));
  AOI21_X1   g06233(.A1(new_n7236_), .A2(new_n7238_), .B(new_n7212_), .ZN(new_n7239_));
  INV_X1     g06234(.I(new_n7212_), .ZN(new_n7240_));
  NOR2_X1    g06235(.A1(new_n7237_), .A2(new_n7219_), .ZN(new_n7241_));
  NOR2_X1    g06236(.A1(new_n7235_), .A2(new_n7220_), .ZN(new_n7242_));
  NOR3_X1    g06237(.A1(new_n7242_), .A2(new_n7241_), .A3(new_n7240_), .ZN(new_n7243_));
  NOR2_X1    g06238(.A1(new_n7239_), .A2(new_n7243_), .ZN(new_n7244_));
  INV_X1     g06239(.I(new_n7244_), .ZN(new_n7245_));
  OAI21_X1   g06240(.A1(new_n7200_), .A2(new_n7203_), .B(new_n7245_), .ZN(new_n7246_));
  OAI21_X1   g06241(.A1(new_n7201_), .A2(new_n7202_), .B(new_n7109_), .ZN(new_n7247_));
  NAND3_X1   g06242(.A1(new_n7199_), .A2(new_n7190_), .A3(new_n7110_), .ZN(new_n7248_));
  NAND3_X1   g06243(.A1(new_n7247_), .A2(new_n7248_), .A3(new_n7244_), .ZN(new_n7249_));
  NAND2_X1   g06244(.A1(new_n7246_), .A2(new_n7249_), .ZN(new_n7250_));
  NOR2_X1    g06245(.A1(new_n7083_), .A2(new_n7250_), .ZN(new_n7251_));
  NOR2_X1    g06246(.A1(new_n6933_), .A2(\A[20] ), .ZN(new_n7252_));
  NOR2_X1    g06247(.A1(new_n6931_), .A2(\A[21] ), .ZN(new_n7253_));
  OAI21_X1   g06248(.A1(new_n7252_), .A2(new_n7253_), .B(\A[19] ), .ZN(new_n7254_));
  INV_X1     g06249(.I(new_n6938_), .ZN(new_n7255_));
  OAI21_X1   g06250(.A1(new_n7255_), .A2(new_n6936_), .B(new_n6930_), .ZN(new_n7256_));
  NAND3_X1   g06251(.A1(new_n6955_), .A2(new_n7254_), .A3(new_n7256_), .ZN(new_n7257_));
  OAI21_X1   g06252(.A1(new_n6935_), .A2(new_n6939_), .B(new_n6954_), .ZN(new_n7258_));
  AOI21_X1   g06253(.A1(new_n7257_), .A2(new_n7258_), .B(new_n6951_), .ZN(new_n7259_));
  NAND2_X1   g06254(.A1(new_n6943_), .A2(\A[24] ), .ZN(new_n7260_));
  NAND2_X1   g06255(.A1(new_n6941_), .A2(\A[23] ), .ZN(new_n7261_));
  AOI21_X1   g06256(.A1(new_n7260_), .A2(new_n7261_), .B(new_n6946_), .ZN(new_n7262_));
  INV_X1     g06257(.I(new_n6949_), .ZN(new_n7263_));
  AOI21_X1   g06258(.A1(new_n7263_), .A2(new_n6947_), .B(\A[22] ), .ZN(new_n7264_));
  NOR2_X1    g06259(.A1(new_n7264_), .A2(new_n7262_), .ZN(new_n7265_));
  NOR3_X1    g06260(.A1(new_n6939_), .A2(new_n6954_), .A3(new_n6935_), .ZN(new_n7266_));
  NOR2_X1    g06261(.A1(new_n6940_), .A2(new_n6955_), .ZN(new_n7267_));
  NOR3_X1    g06262(.A1(new_n7267_), .A2(new_n7265_), .A3(new_n7266_), .ZN(new_n7268_));
  NOR2_X1    g06263(.A1(new_n7268_), .A2(new_n7259_), .ZN(new_n7269_));
  NOR2_X1    g06264(.A1(new_n7265_), .A2(new_n6924_), .ZN(new_n7270_));
  NAND2_X1   g06265(.A1(new_n6916_), .A2(\A[30] ), .ZN(new_n7271_));
  NAND2_X1   g06266(.A1(new_n6914_), .A2(\A[29] ), .ZN(new_n7272_));
  AOI21_X1   g06267(.A1(new_n7271_), .A2(new_n7272_), .B(new_n6919_), .ZN(new_n7273_));
  INV_X1     g06268(.I(new_n6922_), .ZN(new_n7274_));
  AOI21_X1   g06269(.A1(new_n7274_), .A2(new_n6920_), .B(\A[28] ), .ZN(new_n7275_));
  NOR2_X1    g06270(.A1(new_n7275_), .A2(new_n7273_), .ZN(new_n7276_));
  NOR2_X1    g06271(.A1(new_n7276_), .A2(new_n6951_), .ZN(new_n7277_));
  NAND2_X1   g06272(.A1(new_n6906_), .A2(\A[27] ), .ZN(new_n7278_));
  NAND2_X1   g06273(.A1(new_n6904_), .A2(\A[26] ), .ZN(new_n7279_));
  AOI21_X1   g06274(.A1(new_n7278_), .A2(new_n7279_), .B(new_n6909_), .ZN(new_n7280_));
  INV_X1     g06275(.I(new_n6910_), .ZN(new_n7281_));
  NAND2_X1   g06276(.A1(\A[26] ), .A2(\A[27] ), .ZN(new_n7282_));
  AOI21_X1   g06277(.A1(new_n7281_), .A2(new_n7282_), .B(\A[25] ), .ZN(new_n7283_));
  NOR2_X1    g06278(.A1(new_n7283_), .A2(new_n7280_), .ZN(new_n7284_));
  NAND2_X1   g06279(.A1(new_n7254_), .A2(new_n7256_), .ZN(new_n7285_));
  NOR2_X1    g06280(.A1(new_n7284_), .A2(new_n7285_), .ZN(new_n7286_));
  NOR2_X1    g06281(.A1(new_n6940_), .A2(new_n6913_), .ZN(new_n7287_));
  OAI22_X1   g06282(.A1(new_n7270_), .A2(new_n7277_), .B1(new_n7286_), .B2(new_n7287_), .ZN(new_n7288_));
  AOI21_X1   g06283(.A1(new_n6918_), .A2(new_n6923_), .B(new_n6927_), .ZN(new_n7289_));
  AOI21_X1   g06284(.A1(new_n6945_), .A2(new_n6950_), .B(new_n6954_), .ZN(new_n7290_));
  AOI22_X1   g06285(.A1(new_n6913_), .A2(new_n7289_), .B1(new_n7290_), .B2(new_n7285_), .ZN(new_n7291_));
  INV_X1     g06286(.I(new_n7291_), .ZN(new_n7292_));
  NOR2_X1    g06287(.A1(new_n7288_), .A2(new_n7292_), .ZN(new_n7293_));
  NOR2_X1    g06288(.A1(new_n6925_), .A2(new_n6910_), .ZN(new_n7294_));
  INV_X1     g06289(.I(new_n7294_), .ZN(new_n7295_));
  NAND2_X1   g06290(.A1(new_n6920_), .A2(new_n6919_), .ZN(new_n7296_));
  NAND2_X1   g06291(.A1(new_n7296_), .A2(new_n7274_), .ZN(new_n7297_));
  NAND4_X1   g06292(.A1(new_n6908_), .A2(new_n7295_), .A3(new_n7297_), .A4(new_n6912_), .ZN(new_n7298_));
  OAI21_X1   g06293(.A1(new_n7280_), .A2(new_n7283_), .B(new_n6927_), .ZN(new_n7299_));
  AOI21_X1   g06294(.A1(new_n7298_), .A2(new_n7299_), .B(new_n6924_), .ZN(new_n7300_));
  NOR3_X1    g06295(.A1(new_n7283_), .A2(new_n6927_), .A3(new_n7280_), .ZN(new_n7301_));
  AOI22_X1   g06296(.A1(new_n7295_), .A2(new_n7297_), .B1(new_n6908_), .B2(new_n6912_), .ZN(new_n7302_));
  NOR3_X1    g06297(.A1(new_n7302_), .A2(new_n7301_), .A3(new_n7276_), .ZN(new_n7303_));
  NOR2_X1    g06298(.A1(new_n7303_), .A2(new_n7300_), .ZN(new_n7304_));
  NOR2_X1    g06299(.A1(new_n7293_), .A2(new_n7304_), .ZN(new_n7305_));
  NAND2_X1   g06300(.A1(new_n7276_), .A2(new_n6951_), .ZN(new_n7306_));
  NAND2_X1   g06301(.A1(new_n7265_), .A2(new_n6924_), .ZN(new_n7307_));
  NAND2_X1   g06302(.A1(new_n6940_), .A2(new_n6913_), .ZN(new_n7308_));
  NAND2_X1   g06303(.A1(new_n7284_), .A2(new_n7285_), .ZN(new_n7309_));
  AOI22_X1   g06304(.A1(new_n7306_), .A2(new_n7307_), .B1(new_n7309_), .B2(new_n7308_), .ZN(new_n7310_));
  NAND2_X1   g06305(.A1(new_n7310_), .A2(new_n7291_), .ZN(new_n7311_));
  OAI21_X1   g06306(.A1(new_n7302_), .A2(new_n7301_), .B(new_n7276_), .ZN(new_n7312_));
  NAND3_X1   g06307(.A1(new_n7298_), .A2(new_n7299_), .A3(new_n6924_), .ZN(new_n7313_));
  NAND2_X1   g06308(.A1(new_n7312_), .A2(new_n7313_), .ZN(new_n7314_));
  NOR2_X1    g06309(.A1(new_n7311_), .A2(new_n7314_), .ZN(new_n7315_));
  OAI21_X1   g06310(.A1(new_n7305_), .A2(new_n7315_), .B(new_n7269_), .ZN(new_n7316_));
  NAND3_X1   g06311(.A1(new_n7294_), .A2(new_n7274_), .A3(new_n7296_), .ZN(new_n7317_));
  NOR2_X1    g06312(.A1(new_n7276_), .A2(new_n7284_), .ZN(new_n7318_));
  NAND4_X1   g06313(.A1(new_n7318_), .A2(new_n7285_), .A3(new_n7290_), .A4(new_n7317_), .ZN(new_n7319_));
  NOR4_X1    g06314(.A1(new_n7269_), .A2(new_n7288_), .A3(new_n7304_), .A4(new_n7319_), .ZN(new_n7320_));
  OAI21_X1   g06315(.A1(new_n7320_), .A2(new_n7314_), .B(new_n7293_), .ZN(new_n7321_));
  NAND3_X1   g06316(.A1(new_n6984_), .A2(new_n6962_), .A3(new_n6967_), .ZN(new_n7322_));
  NAND2_X1   g06317(.A1(new_n6960_), .A2(\A[15] ), .ZN(new_n7323_));
  NAND2_X1   g06318(.A1(new_n6958_), .A2(\A[14] ), .ZN(new_n7324_));
  AOI21_X1   g06319(.A1(new_n7323_), .A2(new_n7324_), .B(new_n6963_), .ZN(new_n7325_));
  INV_X1     g06320(.I(new_n6964_), .ZN(new_n7326_));
  AOI21_X1   g06321(.A1(new_n7326_), .A2(new_n6965_), .B(\A[13] ), .ZN(new_n7327_));
  OAI22_X1   g06322(.A1(new_n6964_), .A2(new_n6980_), .B1(new_n6982_), .B2(new_n6977_), .ZN(new_n7328_));
  OAI21_X1   g06323(.A1(new_n7325_), .A2(new_n7327_), .B(new_n7328_), .ZN(new_n7329_));
  AOI21_X1   g06324(.A1(new_n7322_), .A2(new_n7329_), .B(new_n6979_), .ZN(new_n7330_));
  NAND2_X1   g06325(.A1(new_n6971_), .A2(\A[18] ), .ZN(new_n7331_));
  NAND2_X1   g06326(.A1(new_n6969_), .A2(\A[17] ), .ZN(new_n7332_));
  AOI21_X1   g06327(.A1(new_n7331_), .A2(new_n7332_), .B(new_n6974_), .ZN(new_n7333_));
  INV_X1     g06328(.I(new_n6977_), .ZN(new_n7334_));
  AOI21_X1   g06329(.A1(new_n7334_), .A2(new_n6975_), .B(\A[16] ), .ZN(new_n7335_));
  NOR2_X1    g06330(.A1(new_n7335_), .A2(new_n7333_), .ZN(new_n7336_));
  NOR3_X1    g06331(.A1(new_n7327_), .A2(new_n7328_), .A3(new_n7325_), .ZN(new_n7337_));
  AOI21_X1   g06332(.A1(new_n6962_), .A2(new_n6967_), .B(new_n6984_), .ZN(new_n7338_));
  NOR3_X1    g06333(.A1(new_n7338_), .A2(new_n7336_), .A3(new_n7337_), .ZN(new_n7339_));
  NOR2_X1    g06334(.A1(new_n7339_), .A2(new_n7330_), .ZN(new_n7340_));
  NAND2_X1   g06335(.A1(new_n7336_), .A2(new_n7007_), .ZN(new_n7341_));
  NAND2_X1   g06336(.A1(new_n6999_), .A2(\A[12] ), .ZN(new_n7342_));
  NAND2_X1   g06337(.A1(new_n6997_), .A2(\A[11] ), .ZN(new_n7343_));
  AOI21_X1   g06338(.A1(new_n7342_), .A2(new_n7343_), .B(new_n7002_), .ZN(new_n7344_));
  INV_X1     g06339(.I(new_n7005_), .ZN(new_n7345_));
  AOI21_X1   g06340(.A1(new_n7345_), .A2(new_n7003_), .B(\A[10] ), .ZN(new_n7346_));
  NOR2_X1    g06341(.A1(new_n7346_), .A2(new_n7344_), .ZN(new_n7347_));
  NAND2_X1   g06342(.A1(new_n7347_), .A2(new_n6979_), .ZN(new_n7348_));
  NAND2_X1   g06343(.A1(new_n7341_), .A2(new_n7348_), .ZN(new_n7349_));
  NAND2_X1   g06344(.A1(new_n6988_), .A2(\A[9] ), .ZN(new_n7350_));
  NAND2_X1   g06345(.A1(new_n6986_), .A2(\A[8] ), .ZN(new_n7351_));
  AOI21_X1   g06346(.A1(new_n7350_), .A2(new_n7351_), .B(new_n6991_), .ZN(new_n7352_));
  INV_X1     g06347(.I(new_n6992_), .ZN(new_n7353_));
  AOI21_X1   g06348(.A1(new_n7353_), .A2(new_n6993_), .B(\A[7] ), .ZN(new_n7354_));
  NOR2_X1    g06349(.A1(new_n7354_), .A2(new_n7352_), .ZN(new_n7355_));
  NAND2_X1   g06350(.A1(new_n7355_), .A2(new_n6968_), .ZN(new_n7356_));
  NOR2_X1    g06351(.A1(new_n7327_), .A2(new_n7325_), .ZN(new_n7357_));
  NAND2_X1   g06352(.A1(new_n7357_), .A2(new_n6996_), .ZN(new_n7358_));
  NAND2_X1   g06353(.A1(new_n7356_), .A2(new_n7358_), .ZN(new_n7359_));
  AOI21_X1   g06354(.A1(new_n6973_), .A2(new_n6978_), .B(new_n7328_), .ZN(new_n7360_));
  AOI21_X1   g06355(.A1(new_n7001_), .A2(new_n7006_), .B(new_n7010_), .ZN(new_n7361_));
  AOI22_X1   g06356(.A1(new_n6968_), .A2(new_n7360_), .B1(new_n7361_), .B2(new_n6996_), .ZN(new_n7362_));
  NAND3_X1   g06357(.A1(new_n7349_), .A2(new_n7359_), .A3(new_n7362_), .ZN(new_n7363_));
  NOR2_X1    g06358(.A1(new_n6996_), .A2(new_n7010_), .ZN(new_n7364_));
  OAI21_X1   g06359(.A1(new_n7352_), .A2(new_n7354_), .B(new_n7010_), .ZN(new_n7365_));
  INV_X1     g06360(.I(new_n7365_), .ZN(new_n7366_));
  OAI21_X1   g06361(.A1(new_n7366_), .A2(new_n7364_), .B(new_n7347_), .ZN(new_n7367_));
  NAND2_X1   g06362(.A1(new_n7355_), .A2(new_n7011_), .ZN(new_n7368_));
  NAND3_X1   g06363(.A1(new_n7368_), .A2(new_n7007_), .A3(new_n7365_), .ZN(new_n7369_));
  NAND2_X1   g06364(.A1(new_n7367_), .A2(new_n7369_), .ZN(new_n7370_));
  NOR2_X1    g06365(.A1(new_n7347_), .A2(new_n6979_), .ZN(new_n7371_));
  NOR2_X1    g06366(.A1(new_n7336_), .A2(new_n7007_), .ZN(new_n7372_));
  NOR2_X1    g06367(.A1(new_n7357_), .A2(new_n6996_), .ZN(new_n7373_));
  NOR2_X1    g06368(.A1(new_n7355_), .A2(new_n6968_), .ZN(new_n7374_));
  OAI22_X1   g06369(.A1(new_n7371_), .A2(new_n7372_), .B1(new_n7373_), .B2(new_n7374_), .ZN(new_n7375_));
  NAND2_X1   g06370(.A1(new_n6981_), .A2(new_n6983_), .ZN(new_n7376_));
  NOR2_X1    g06371(.A1(new_n7357_), .A2(new_n7336_), .ZN(new_n7377_));
  NAND4_X1   g06372(.A1(new_n7377_), .A2(new_n6996_), .A3(new_n7361_), .A4(new_n7376_), .ZN(new_n7378_));
  NAND3_X1   g06373(.A1(new_n7363_), .A2(new_n7370_), .A3(new_n7340_), .ZN(new_n7380_));
  INV_X1     g06374(.I(new_n7380_), .ZN(new_n7381_));
  XOR2_X1    g06375(.A1(new_n7285_), .A2(new_n6951_), .Z(new_n7382_));
  XOR2_X1    g06376(.A1(new_n7355_), .A2(new_n7007_), .Z(new_n7383_));
  NAND2_X1   g06377(.A1(new_n7382_), .A2(new_n7383_), .ZN(new_n7384_));
  NAND2_X1   g06378(.A1(new_n6956_), .A2(new_n7012_), .ZN(new_n7385_));
  XOR2_X1    g06379(.A1(new_n7276_), .A2(new_n6913_), .Z(new_n7386_));
  NAND2_X1   g06380(.A1(new_n6985_), .A2(new_n7386_), .ZN(new_n7387_));
  XOR2_X1    g06381(.A1(new_n7357_), .A2(new_n6979_), .Z(new_n7388_));
  NAND2_X1   g06382(.A1(new_n7388_), .A2(new_n6929_), .ZN(new_n7389_));
  AOI22_X1   g06383(.A1(new_n7384_), .A2(new_n7385_), .B1(new_n7387_), .B2(new_n7389_), .ZN(new_n7390_));
  NAND3_X1   g06384(.A1(new_n7321_), .A2(new_n7381_), .A3(new_n7390_), .ZN(new_n7391_));
  OAI21_X1   g06385(.A1(new_n7267_), .A2(new_n7266_), .B(new_n7265_), .ZN(new_n7392_));
  NAND3_X1   g06386(.A1(new_n7257_), .A2(new_n7258_), .A3(new_n6951_), .ZN(new_n7393_));
  NAND2_X1   g06387(.A1(new_n7392_), .A2(new_n7393_), .ZN(new_n7394_));
  NAND3_X1   g06388(.A1(new_n6924_), .A2(new_n6913_), .A3(new_n7317_), .ZN(new_n7395_));
  NOR4_X1    g06389(.A1(new_n7395_), .A2(new_n6940_), .A3(new_n7265_), .A4(new_n6954_), .ZN(new_n7396_));
  NAND4_X1   g06390(.A1(new_n7394_), .A2(new_n7310_), .A3(new_n7314_), .A4(new_n7396_), .ZN(new_n7397_));
  AOI21_X1   g06391(.A1(new_n7397_), .A2(new_n7304_), .B(new_n7311_), .ZN(new_n7398_));
  NOR2_X1    g06392(.A1(new_n6956_), .A2(new_n7012_), .ZN(new_n7399_));
  NOR2_X1    g06393(.A1(new_n7382_), .A2(new_n7383_), .ZN(new_n7400_));
  NOR2_X1    g06394(.A1(new_n7388_), .A2(new_n6929_), .ZN(new_n7401_));
  NOR2_X1    g06395(.A1(new_n6985_), .A2(new_n7386_), .ZN(new_n7402_));
  OAI22_X1   g06396(.A1(new_n7399_), .A2(new_n7400_), .B1(new_n7402_), .B2(new_n7401_), .ZN(new_n7403_));
  OAI21_X1   g06397(.A1(new_n7380_), .A2(new_n7403_), .B(new_n7398_), .ZN(new_n7404_));
  AOI21_X1   g06398(.A1(new_n7404_), .A2(new_n7391_), .B(new_n7316_), .ZN(new_n7405_));
  XOR2_X1    g06399(.A1(new_n7382_), .A2(new_n6929_), .Z(new_n7406_));
  XOR2_X1    g06400(.A1(new_n6985_), .A2(new_n7383_), .Z(new_n7407_));
  NAND2_X1   g06401(.A1(new_n7407_), .A2(new_n7406_), .ZN(new_n7408_));
  NAND2_X1   g06402(.A1(new_n7013_), .A2(new_n6957_), .ZN(new_n7409_));
  AOI21_X1   g06403(.A1(new_n7409_), .A2(new_n7408_), .B(new_n7079_), .ZN(new_n7410_));
  INV_X1     g06404(.I(new_n7410_), .ZN(new_n7411_));
  OAI21_X1   g06405(.A1(new_n7029_), .A2(new_n7064_), .B(new_n7049_), .ZN(new_n7412_));
  AOI21_X1   g06406(.A1(\A[4] ), .A2(\A[5] ), .B(\A[3] ), .ZN(new_n7413_));
  NOR2_X1    g06407(.A1(new_n7413_), .A2(new_n7046_), .ZN(new_n7414_));
  NOR2_X1    g06408(.A1(\A[1] ), .A2(\A[2] ), .ZN(new_n7415_));
  AOI21_X1   g06409(.A1(\A[1] ), .A2(\A[2] ), .B(\A[0] ), .ZN(new_n7416_));
  NOR2_X1    g06410(.A1(new_n7416_), .A2(new_n7415_), .ZN(new_n7417_));
  NOR2_X1    g06411(.A1(new_n7414_), .A2(new_n7417_), .ZN(new_n7418_));
  NOR4_X1    g06412(.A1(new_n7413_), .A2(new_n7416_), .A3(new_n7046_), .A4(new_n7415_), .ZN(new_n7419_));
  NOR2_X1    g06413(.A1(new_n7418_), .A2(new_n7419_), .ZN(new_n7420_));
  NOR2_X1    g06414(.A1(new_n7420_), .A2(new_n7038_), .ZN(new_n7421_));
  NAND3_X1   g06415(.A1(new_n7421_), .A2(new_n7060_), .A3(new_n7070_), .ZN(new_n7422_));
  OAI22_X1   g06416(.A1(new_n7046_), .A2(new_n7413_), .B1(new_n7416_), .B2(new_n7415_), .ZN(new_n7423_));
  NAND2_X1   g06417(.A1(new_n7414_), .A2(new_n7417_), .ZN(new_n7424_));
  NAND2_X1   g06418(.A1(new_n7424_), .A2(new_n7423_), .ZN(new_n7425_));
  NAND2_X1   g06419(.A1(new_n7425_), .A2(new_n7064_), .ZN(new_n7426_));
  OAI21_X1   g06420(.A1(new_n7426_), .A2(new_n7060_), .B(new_n7029_), .ZN(new_n7427_));
  AOI21_X1   g06421(.A1(new_n7427_), .A2(new_n7422_), .B(new_n7412_), .ZN(new_n7428_));
  NAND2_X1   g06422(.A1(new_n7056_), .A2(new_n7050_), .ZN(new_n7429_));
  AND2_X2    g06423(.A1(new_n7429_), .A2(new_n7057_), .Z(new_n7430_));
  NOR2_X1    g06424(.A1(new_n7428_), .A2(new_n7430_), .ZN(new_n7431_));
  NAND2_X1   g06425(.A1(new_n7428_), .A2(new_n7430_), .ZN(new_n7432_));
  INV_X1     g06426(.I(\A[995] ), .ZN(new_n7433_));
  NAND2_X1   g06427(.A1(new_n7433_), .A2(\A[996] ), .ZN(new_n7434_));
  INV_X1     g06428(.I(\A[996] ), .ZN(new_n7435_));
  NAND2_X1   g06429(.A1(new_n7435_), .A2(\A[995] ), .ZN(new_n7436_));
  AOI21_X1   g06430(.A1(new_n7434_), .A2(new_n7436_), .B(new_n7014_), .ZN(new_n7437_));
  INV_X1     g06431(.I(new_n7015_), .ZN(new_n7438_));
  AOI21_X1   g06432(.A1(new_n7438_), .A2(new_n7016_), .B(\A[994] ), .ZN(new_n7439_));
  NOR2_X1    g06433(.A1(new_n7439_), .A2(new_n7437_), .ZN(new_n7440_));
  INV_X1     g06434(.I(new_n7440_), .ZN(new_n7441_));
  INV_X1     g06435(.I(\A[992] ), .ZN(new_n7442_));
  NAND2_X1   g06436(.A1(new_n7442_), .A2(\A[993] ), .ZN(new_n7443_));
  INV_X1     g06437(.I(\A[993] ), .ZN(new_n7444_));
  NAND2_X1   g06438(.A1(new_n7444_), .A2(\A[992] ), .ZN(new_n7445_));
  AOI21_X1   g06439(.A1(new_n7443_), .A2(new_n7445_), .B(new_n7018_), .ZN(new_n7446_));
  INV_X1     g06440(.I(new_n7019_), .ZN(new_n7447_));
  AOI21_X1   g06441(.A1(new_n7447_), .A2(new_n7020_), .B(\A[991] ), .ZN(new_n7448_));
  NOR2_X1    g06442(.A1(new_n7448_), .A2(new_n7446_), .ZN(new_n7449_));
  NOR2_X1    g06443(.A1(new_n7017_), .A2(new_n7021_), .ZN(new_n7450_));
  NAND2_X1   g06444(.A1(new_n7449_), .A2(new_n7450_), .ZN(new_n7451_));
  OAI22_X1   g06445(.A1(new_n7448_), .A2(new_n7446_), .B1(new_n7017_), .B2(new_n7021_), .ZN(new_n7452_));
  AOI21_X1   g06446(.A1(new_n7451_), .A2(new_n7452_), .B(new_n7441_), .ZN(new_n7453_));
  NOR4_X1    g06447(.A1(new_n7448_), .A2(new_n7446_), .A3(new_n7017_), .A4(new_n7021_), .ZN(new_n7454_));
  INV_X1     g06448(.I(new_n7452_), .ZN(new_n7455_));
  NOR3_X1    g06449(.A1(new_n7455_), .A2(new_n7440_), .A3(new_n7454_), .ZN(new_n7456_));
  NOR2_X1    g06450(.A1(new_n7456_), .A2(new_n7453_), .ZN(new_n7457_));
  NOR4_X1    g06451(.A1(new_n7073_), .A2(new_n7457_), .A3(new_n7067_), .A4(new_n7022_), .ZN(new_n7458_));
  NAND2_X1   g06452(.A1(new_n7458_), .A2(new_n7432_), .ZN(new_n7459_));
  INV_X1     g06453(.I(new_n7049_), .ZN(new_n7460_));
  AOI21_X1   g06454(.A1(new_n7070_), .A2(new_n7038_), .B(new_n7460_), .ZN(new_n7461_));
  NOR3_X1    g06455(.A1(new_n7426_), .A2(new_n7029_), .A3(new_n7065_), .ZN(new_n7462_));
  AOI21_X1   g06456(.A1(new_n7421_), .A2(new_n7065_), .B(new_n7070_), .ZN(new_n7463_));
  OAI21_X1   g06457(.A1(new_n7463_), .A2(new_n7462_), .B(new_n7461_), .ZN(new_n7464_));
  INV_X1     g06458(.I(new_n7430_), .ZN(new_n7465_));
  NOR2_X1    g06459(.A1(new_n7464_), .A2(new_n7465_), .ZN(new_n7466_));
  OAI21_X1   g06460(.A1(new_n7455_), .A2(new_n7454_), .B(new_n7440_), .ZN(new_n7467_));
  NAND3_X1   g06461(.A1(new_n7451_), .A2(new_n7441_), .A3(new_n7452_), .ZN(new_n7468_));
  NAND2_X1   g06462(.A1(new_n7467_), .A2(new_n7468_), .ZN(new_n7469_));
  NAND4_X1   g06463(.A1(new_n7076_), .A2(new_n7469_), .A3(new_n7077_), .A4(new_n7075_), .ZN(new_n7470_));
  NAND2_X1   g06464(.A1(new_n7470_), .A2(new_n7466_), .ZN(new_n7471_));
  AOI21_X1   g06465(.A1(new_n7459_), .A2(new_n7471_), .B(new_n7431_), .ZN(new_n7472_));
  NOR3_X1    g06466(.A1(new_n7458_), .A2(new_n7428_), .A3(new_n7430_), .ZN(new_n7473_));
  NOR2_X1    g06467(.A1(new_n7472_), .A2(new_n7473_), .ZN(new_n7474_));
  NOR2_X1    g06468(.A1(new_n7411_), .A2(new_n7474_), .ZN(new_n7475_));
  INV_X1     g06469(.I(new_n7475_), .ZN(new_n7476_));
  NOR2_X1    g06470(.A1(new_n7476_), .A2(new_n7405_), .ZN(new_n7477_));
  INV_X1     g06471(.I(new_n7316_), .ZN(new_n7478_));
  NOR3_X1    g06472(.A1(new_n7398_), .A2(new_n7403_), .A3(new_n7380_), .ZN(new_n7479_));
  NOR2_X1    g06473(.A1(new_n7399_), .A2(new_n7400_), .ZN(new_n7480_));
  NOR2_X1    g06474(.A1(new_n7402_), .A2(new_n7401_), .ZN(new_n7481_));
  NOR3_X1    g06475(.A1(new_n7480_), .A2(new_n7481_), .A3(new_n7380_), .ZN(new_n7482_));
  NOR2_X1    g06476(.A1(new_n7482_), .A2(new_n7321_), .ZN(new_n7483_));
  OAI21_X1   g06477(.A1(new_n7483_), .A2(new_n7479_), .B(new_n7478_), .ZN(new_n7484_));
  NOR2_X1    g06478(.A1(new_n7476_), .A2(new_n7484_), .ZN(new_n7485_));
  OAI21_X1   g06479(.A1(new_n7477_), .A2(new_n7485_), .B(new_n7251_), .ZN(new_n7486_));
  NAND2_X1   g06480(.A1(new_n7121_), .A2(new_n7135_), .ZN(new_n7487_));
  OR2_X2     g06481(.A1(new_n7133_), .A2(new_n7134_), .Z(new_n7488_));
  NAND2_X1   g06482(.A1(new_n7488_), .A2(new_n7196_), .ZN(new_n7489_));
  AOI21_X1   g06483(.A1(new_n7489_), .A2(new_n7487_), .B(new_n7132_), .ZN(new_n7490_));
  INV_X1     g06484(.I(new_n7132_), .ZN(new_n7491_));
  NOR2_X1    g06485(.A1(new_n7488_), .A2(new_n7196_), .ZN(new_n7492_));
  NOR2_X1    g06486(.A1(new_n7121_), .A2(new_n7135_), .ZN(new_n7493_));
  NOR3_X1    g06487(.A1(new_n7492_), .A2(new_n7493_), .A3(new_n7491_), .ZN(new_n7494_));
  NOR2_X1    g06488(.A1(new_n7494_), .A2(new_n7490_), .ZN(new_n7495_));
  NOR2_X1    g06489(.A1(new_n7150_), .A2(\A[77] ), .ZN(new_n7496_));
  NOR2_X1    g06490(.A1(new_n7148_), .A2(\A[78] ), .ZN(new_n7497_));
  OAI21_X1   g06491(.A1(new_n7496_), .A2(new_n7497_), .B(\A[76] ), .ZN(new_n7498_));
  INV_X1     g06492(.I(new_n7153_), .ZN(new_n7499_));
  OAI21_X1   g06493(.A1(new_n7499_), .A2(new_n7154_), .B(new_n7147_), .ZN(new_n7500_));
  NAND2_X1   g06494(.A1(new_n7498_), .A2(new_n7500_), .ZN(new_n7501_));
  NOR2_X1    g06495(.A1(new_n7491_), .A2(new_n7501_), .ZN(new_n7502_));
  NOR2_X1    g06496(.A1(new_n7157_), .A2(new_n7132_), .ZN(new_n7503_));
  AOI21_X1   g06497(.A1(new_n7141_), .A2(new_n7145_), .B(new_n7196_), .ZN(new_n7504_));
  NOR2_X1    g06498(.A1(new_n7121_), .A2(new_n7146_), .ZN(new_n7505_));
  OAI22_X1   g06499(.A1(new_n7502_), .A2(new_n7503_), .B1(new_n7504_), .B2(new_n7505_), .ZN(new_n7506_));
  NAND3_X1   g06500(.A1(new_n7196_), .A2(new_n7132_), .A3(new_n7135_), .ZN(new_n7507_));
  NAND3_X1   g06501(.A1(new_n7501_), .A2(new_n7146_), .A3(new_n7161_), .ZN(new_n7508_));
  NAND2_X1   g06502(.A1(new_n7507_), .A2(new_n7508_), .ZN(new_n7509_));
  NOR2_X1    g06503(.A1(new_n7506_), .A2(new_n7509_), .ZN(new_n7510_));
  NAND2_X1   g06504(.A1(new_n7139_), .A2(\A[75] ), .ZN(new_n7511_));
  NAND2_X1   g06505(.A1(new_n7137_), .A2(\A[74] ), .ZN(new_n7512_));
  AOI21_X1   g06506(.A1(new_n7511_), .A2(new_n7512_), .B(new_n7142_), .ZN(new_n7513_));
  INV_X1     g06507(.I(new_n7143_), .ZN(new_n7514_));
  NAND2_X1   g06508(.A1(\A[74] ), .A2(\A[75] ), .ZN(new_n7515_));
  AOI21_X1   g06509(.A1(new_n7514_), .A2(new_n7515_), .B(\A[73] ), .ZN(new_n7516_));
  NOR3_X1    g06510(.A1(new_n7516_), .A2(new_n7160_), .A3(new_n7513_), .ZN(new_n7517_));
  NOR2_X1    g06511(.A1(new_n7158_), .A2(new_n7143_), .ZN(new_n7518_));
  INV_X1     g06512(.I(new_n7518_), .ZN(new_n7519_));
  NOR2_X1    g06513(.A1(new_n7159_), .A2(new_n7154_), .ZN(new_n7520_));
  INV_X1     g06514(.I(new_n7520_), .ZN(new_n7521_));
  AOI22_X1   g06515(.A1(new_n7519_), .A2(new_n7521_), .B1(new_n7141_), .B2(new_n7145_), .ZN(new_n7522_));
  OAI21_X1   g06516(.A1(new_n7522_), .A2(new_n7517_), .B(new_n7157_), .ZN(new_n7523_));
  NAND4_X1   g06517(.A1(new_n7519_), .A2(new_n7521_), .A3(new_n7141_), .A4(new_n7145_), .ZN(new_n7524_));
  OAI21_X1   g06518(.A1(new_n7513_), .A2(new_n7516_), .B(new_n7160_), .ZN(new_n7525_));
  NAND3_X1   g06519(.A1(new_n7524_), .A2(new_n7525_), .A3(new_n7501_), .ZN(new_n7526_));
  NAND2_X1   g06520(.A1(new_n7523_), .A2(new_n7526_), .ZN(new_n7527_));
  XOR2_X1    g06521(.A1(new_n7510_), .A2(new_n7527_), .Z(new_n7528_));
  NAND2_X1   g06522(.A1(new_n7528_), .A2(new_n7495_), .ZN(new_n7529_));
  INV_X1     g06523(.I(new_n7510_), .ZN(new_n7530_));
  AOI21_X1   g06524(.A1(new_n7524_), .A2(new_n7525_), .B(new_n7501_), .ZN(new_n7531_));
  NOR3_X1    g06525(.A1(new_n7522_), .A2(new_n7517_), .A3(new_n7157_), .ZN(new_n7532_));
  NOR2_X1    g06526(.A1(new_n7532_), .A2(new_n7531_), .ZN(new_n7533_));
  OR2_X2     g06527(.A1(new_n7494_), .A2(new_n7490_), .Z(new_n7534_));
  NAND2_X1   g06528(.A1(new_n7518_), .A2(new_n7520_), .ZN(new_n7535_));
  NAND3_X1   g06529(.A1(new_n7501_), .A2(new_n7146_), .A3(new_n7535_), .ZN(new_n7536_));
  OR2_X2     g06530(.A1(new_n7507_), .A2(new_n7536_), .Z(new_n7537_));
  NOR3_X1    g06531(.A1(new_n7506_), .A2(new_n7537_), .A3(new_n7533_), .ZN(new_n7538_));
  NAND2_X1   g06532(.A1(new_n7538_), .A2(new_n7534_), .ZN(new_n7539_));
  AOI21_X1   g06533(.A1(new_n7539_), .A2(new_n7533_), .B(new_n7530_), .ZN(new_n7540_));
  XOR2_X1    g06534(.A1(new_n7109_), .A2(new_n7136_), .Z(new_n7541_));
  NAND2_X1   g06535(.A1(new_n7165_), .A2(\A[63] ), .ZN(new_n7542_));
  NAND2_X1   g06536(.A1(new_n7163_), .A2(\A[62] ), .ZN(new_n7543_));
  AOI21_X1   g06537(.A1(new_n7542_), .A2(new_n7543_), .B(new_n7168_), .ZN(new_n7544_));
  INV_X1     g06538(.I(new_n7169_), .ZN(new_n7545_));
  NAND2_X1   g06539(.A1(\A[62] ), .A2(\A[63] ), .ZN(new_n7546_));
  AOI21_X1   g06540(.A1(new_n7545_), .A2(new_n7546_), .B(\A[61] ), .ZN(new_n7547_));
  NOR3_X1    g06541(.A1(new_n7547_), .A2(new_n7186_), .A3(new_n7544_), .ZN(new_n7548_));
  NOR2_X1    g06542(.A1(new_n7184_), .A2(new_n7169_), .ZN(new_n7549_));
  INV_X1     g06543(.I(new_n7549_), .ZN(new_n7550_));
  NAND2_X1   g06544(.A1(new_n7179_), .A2(new_n7173_), .ZN(new_n7551_));
  NAND2_X1   g06545(.A1(new_n7551_), .A2(new_n7181_), .ZN(new_n7552_));
  AOI22_X1   g06546(.A1(new_n7550_), .A2(new_n7552_), .B1(new_n7167_), .B2(new_n7171_), .ZN(new_n7553_));
  OAI21_X1   g06547(.A1(new_n7553_), .A2(new_n7548_), .B(new_n7183_), .ZN(new_n7554_));
  NOR2_X1    g06548(.A1(new_n7176_), .A2(\A[65] ), .ZN(new_n7555_));
  NOR2_X1    g06549(.A1(new_n7174_), .A2(\A[66] ), .ZN(new_n7556_));
  OAI21_X1   g06550(.A1(new_n7555_), .A2(new_n7556_), .B(\A[64] ), .ZN(new_n7557_));
  INV_X1     g06551(.I(new_n7179_), .ZN(new_n7558_));
  OAI21_X1   g06552(.A1(new_n7558_), .A2(new_n7180_), .B(new_n7173_), .ZN(new_n7559_));
  NAND2_X1   g06553(.A1(new_n7557_), .A2(new_n7559_), .ZN(new_n7560_));
  NAND4_X1   g06554(.A1(new_n7167_), .A2(new_n7550_), .A3(new_n7552_), .A4(new_n7171_), .ZN(new_n7561_));
  OAI21_X1   g06555(.A1(new_n7544_), .A2(new_n7547_), .B(new_n7186_), .ZN(new_n7562_));
  NAND3_X1   g06556(.A1(new_n7561_), .A2(new_n7562_), .A3(new_n7560_), .ZN(new_n7563_));
  NAND2_X1   g06557(.A1(new_n7554_), .A2(new_n7563_), .ZN(new_n7564_));
  INV_X1     g06558(.I(new_n7105_), .ZN(new_n7565_));
  NOR2_X1    g06559(.A1(new_n7565_), .A2(new_n7560_), .ZN(new_n7566_));
  NOR2_X1    g06560(.A1(new_n7183_), .A2(new_n7105_), .ZN(new_n7567_));
  NOR2_X1    g06561(.A1(new_n7087_), .A2(\A[56] ), .ZN(new_n7568_));
  NOR2_X1    g06562(.A1(new_n7085_), .A2(\A[57] ), .ZN(new_n7569_));
  OAI21_X1   g06563(.A1(new_n7568_), .A2(new_n7569_), .B(\A[55] ), .ZN(new_n7570_));
  INV_X1     g06564(.I(new_n7092_), .ZN(new_n7571_));
  OAI21_X1   g06565(.A1(new_n7571_), .A2(new_n7090_), .B(new_n7084_), .ZN(new_n7572_));
  NAND2_X1   g06566(.A1(new_n7570_), .A2(new_n7572_), .ZN(new_n7573_));
  AOI21_X1   g06567(.A1(new_n7167_), .A2(new_n7171_), .B(new_n7573_), .ZN(new_n7574_));
  NOR2_X1    g06568(.A1(new_n7094_), .A2(new_n7172_), .ZN(new_n7575_));
  OAI22_X1   g06569(.A1(new_n7566_), .A2(new_n7567_), .B1(new_n7574_), .B2(new_n7575_), .ZN(new_n7576_));
  NOR4_X1    g06570(.A1(new_n7106_), .A2(\A[58] ), .A3(\A[59] ), .A4(\A[60] ), .ZN(new_n7577_));
  NAND2_X1   g06571(.A1(new_n7573_), .A2(new_n7577_), .ZN(new_n7578_));
  NAND3_X1   g06572(.A1(new_n7560_), .A2(new_n7172_), .A3(new_n7187_), .ZN(new_n7579_));
  NAND2_X1   g06573(.A1(new_n7579_), .A2(new_n7578_), .ZN(new_n7580_));
  NOR2_X1    g06574(.A1(new_n7576_), .A2(new_n7580_), .ZN(new_n7581_));
  NAND2_X1   g06575(.A1(new_n7094_), .A2(new_n7108_), .ZN(new_n7582_));
  INV_X1     g06576(.I(new_n7108_), .ZN(new_n7583_));
  NAND2_X1   g06577(.A1(new_n7583_), .A2(new_n7573_), .ZN(new_n7584_));
  AOI21_X1   g06578(.A1(new_n7584_), .A2(new_n7582_), .B(new_n7105_), .ZN(new_n7585_));
  INV_X1     g06579(.I(new_n7582_), .ZN(new_n7586_));
  NOR2_X1    g06580(.A1(new_n7094_), .A2(new_n7108_), .ZN(new_n7587_));
  NOR3_X1    g06581(.A1(new_n7586_), .A2(new_n7587_), .A3(new_n7565_), .ZN(new_n7588_));
  NOR2_X1    g06582(.A1(new_n7588_), .A2(new_n7585_), .ZN(new_n7589_));
  NAND3_X1   g06583(.A1(new_n7549_), .A2(new_n7181_), .A3(new_n7551_), .ZN(new_n7590_));
  NAND3_X1   g06584(.A1(new_n7560_), .A2(new_n7172_), .A3(new_n7590_), .ZN(new_n7591_));
  OR2_X2     g06585(.A1(new_n7591_), .A2(new_n7578_), .Z(new_n7592_));
  NOR2_X1    g06586(.A1(new_n7576_), .A2(new_n7592_), .ZN(new_n7593_));
  NOR3_X1    g06587(.A1(new_n7581_), .A2(new_n7589_), .A3(new_n7564_), .ZN(new_n7594_));
  NAND3_X1   g06588(.A1(new_n7594_), .A2(new_n7541_), .A3(new_n7189_), .ZN(new_n7595_));
  XOR2_X1    g06589(.A1(new_n7595_), .A2(new_n7540_), .Z(new_n7596_));
  NOR2_X1    g06590(.A1(new_n7596_), .A2(new_n7529_), .ZN(new_n7597_));
  INV_X1     g06591(.I(new_n7249_), .ZN(new_n7598_));
  INV_X1     g06592(.I(\A[46] ), .ZN(new_n7599_));
  INV_X1     g06593(.I(\A[47] ), .ZN(new_n7600_));
  NAND2_X1   g06594(.A1(new_n7600_), .A2(\A[48] ), .ZN(new_n7601_));
  INV_X1     g06595(.I(\A[48] ), .ZN(new_n7602_));
  NAND2_X1   g06596(.A1(new_n7602_), .A2(\A[47] ), .ZN(new_n7603_));
  AOI21_X1   g06597(.A1(new_n7601_), .A2(new_n7603_), .B(new_n7599_), .ZN(new_n7604_));
  INV_X1     g06598(.I(new_n7213_), .ZN(new_n7605_));
  NAND2_X1   g06599(.A1(\A[47] ), .A2(\A[48] ), .ZN(new_n7606_));
  AOI21_X1   g06600(.A1(new_n7605_), .A2(new_n7606_), .B(\A[46] ), .ZN(new_n7607_));
  NOR2_X1    g06601(.A1(new_n7607_), .A2(new_n7604_), .ZN(new_n7608_));
  INV_X1     g06602(.I(\A[45] ), .ZN(new_n7609_));
  NOR2_X1    g06603(.A1(new_n7609_), .A2(\A[44] ), .ZN(new_n7610_));
  INV_X1     g06604(.I(\A[44] ), .ZN(new_n7611_));
  NOR2_X1    g06605(.A1(new_n7611_), .A2(\A[45] ), .ZN(new_n7612_));
  OAI21_X1   g06606(.A1(new_n7610_), .A2(new_n7612_), .B(\A[43] ), .ZN(new_n7613_));
  INV_X1     g06607(.I(\A[43] ), .ZN(new_n7614_));
  NAND2_X1   g06608(.A1(\A[44] ), .A2(\A[45] ), .ZN(new_n7615_));
  INV_X1     g06609(.I(new_n7615_), .ZN(new_n7616_));
  OAI21_X1   g06610(.A1(new_n7616_), .A2(new_n7216_), .B(new_n7614_), .ZN(new_n7617_));
  NAND2_X1   g06611(.A1(new_n7613_), .A2(new_n7617_), .ZN(new_n7618_));
  NOR2_X1    g06612(.A1(new_n7215_), .A2(new_n7218_), .ZN(new_n7619_));
  INV_X1     g06613(.I(new_n7619_), .ZN(new_n7620_));
  NOR2_X1    g06614(.A1(new_n7620_), .A2(new_n7618_), .ZN(new_n7621_));
  NAND2_X1   g06615(.A1(new_n7611_), .A2(\A[45] ), .ZN(new_n7622_));
  NAND2_X1   g06616(.A1(new_n7609_), .A2(\A[44] ), .ZN(new_n7623_));
  AOI21_X1   g06617(.A1(new_n7622_), .A2(new_n7623_), .B(new_n7614_), .ZN(new_n7624_));
  INV_X1     g06618(.I(new_n7216_), .ZN(new_n7625_));
  AOI21_X1   g06619(.A1(new_n7625_), .A2(new_n7615_), .B(\A[43] ), .ZN(new_n7626_));
  NOR2_X1    g06620(.A1(new_n7626_), .A2(new_n7624_), .ZN(new_n7627_));
  NOR2_X1    g06621(.A1(new_n7627_), .A2(new_n7619_), .ZN(new_n7628_));
  OAI21_X1   g06622(.A1(new_n7621_), .A2(new_n7628_), .B(new_n7608_), .ZN(new_n7629_));
  NOR2_X1    g06623(.A1(new_n7602_), .A2(\A[47] ), .ZN(new_n7630_));
  NOR2_X1    g06624(.A1(new_n7600_), .A2(\A[48] ), .ZN(new_n7631_));
  OAI21_X1   g06625(.A1(new_n7630_), .A2(new_n7631_), .B(\A[46] ), .ZN(new_n7632_));
  INV_X1     g06626(.I(new_n7606_), .ZN(new_n7633_));
  OAI21_X1   g06627(.A1(new_n7633_), .A2(new_n7213_), .B(new_n7599_), .ZN(new_n7634_));
  NAND2_X1   g06628(.A1(new_n7632_), .A2(new_n7634_), .ZN(new_n7635_));
  NAND2_X1   g06629(.A1(new_n7627_), .A2(new_n7619_), .ZN(new_n7636_));
  NAND2_X1   g06630(.A1(new_n7620_), .A2(new_n7618_), .ZN(new_n7637_));
  NAND3_X1   g06631(.A1(new_n7637_), .A2(new_n7636_), .A3(new_n7635_), .ZN(new_n7638_));
  NAND2_X1   g06632(.A1(new_n7629_), .A2(new_n7638_), .ZN(new_n7639_));
  INV_X1     g06633(.I(new_n7639_), .ZN(new_n7640_));
  INV_X1     g06634(.I(\A[52] ), .ZN(new_n7641_));
  INV_X1     g06635(.I(\A[53] ), .ZN(new_n7642_));
  NAND2_X1   g06636(.A1(new_n7642_), .A2(\A[54] ), .ZN(new_n7643_));
  INV_X1     g06637(.I(\A[54] ), .ZN(new_n7644_));
  NAND2_X1   g06638(.A1(new_n7644_), .A2(\A[53] ), .ZN(new_n7645_));
  AOI21_X1   g06639(.A1(new_n7643_), .A2(new_n7645_), .B(new_n7641_), .ZN(new_n7646_));
  INV_X1     g06640(.I(new_n7221_), .ZN(new_n7647_));
  NAND2_X1   g06641(.A1(\A[53] ), .A2(\A[54] ), .ZN(new_n7648_));
  AOI21_X1   g06642(.A1(new_n7647_), .A2(new_n7648_), .B(\A[52] ), .ZN(new_n7649_));
  NOR2_X1    g06643(.A1(new_n7649_), .A2(new_n7646_), .ZN(new_n7650_));
  INV_X1     g06644(.I(\A[51] ), .ZN(new_n7651_));
  NOR2_X1    g06645(.A1(new_n7651_), .A2(\A[50] ), .ZN(new_n7652_));
  INV_X1     g06646(.I(\A[50] ), .ZN(new_n7653_));
  NOR2_X1    g06647(.A1(new_n7653_), .A2(\A[51] ), .ZN(new_n7654_));
  OAI21_X1   g06648(.A1(new_n7652_), .A2(new_n7654_), .B(\A[49] ), .ZN(new_n7655_));
  INV_X1     g06649(.I(\A[49] ), .ZN(new_n7656_));
  AND2_X2    g06650(.A1(\A[50] ), .A2(\A[51] ), .Z(new_n7657_));
  OAI21_X1   g06651(.A1(new_n7657_), .A2(new_n7224_), .B(new_n7656_), .ZN(new_n7658_));
  NAND2_X1   g06652(.A1(new_n7655_), .A2(new_n7658_), .ZN(new_n7659_));
  OAI22_X1   g06653(.A1(new_n7221_), .A2(new_n7222_), .B1(new_n7225_), .B2(new_n7224_), .ZN(new_n7660_));
  NOR2_X1    g06654(.A1(new_n7659_), .A2(new_n7660_), .ZN(new_n7661_));
  NAND2_X1   g06655(.A1(new_n7653_), .A2(\A[51] ), .ZN(new_n7662_));
  NAND2_X1   g06656(.A1(new_n7651_), .A2(\A[50] ), .ZN(new_n7663_));
  AOI21_X1   g06657(.A1(new_n7662_), .A2(new_n7663_), .B(new_n7656_), .ZN(new_n7664_));
  INV_X1     g06658(.I(new_n7224_), .ZN(new_n7665_));
  NAND2_X1   g06659(.A1(\A[50] ), .A2(\A[51] ), .ZN(new_n7666_));
  AOI21_X1   g06660(.A1(new_n7665_), .A2(new_n7666_), .B(\A[49] ), .ZN(new_n7667_));
  NOR2_X1    g06661(.A1(new_n7667_), .A2(new_n7664_), .ZN(new_n7668_));
  INV_X1     g06662(.I(new_n7660_), .ZN(new_n7669_));
  NOR2_X1    g06663(.A1(new_n7668_), .A2(new_n7669_), .ZN(new_n7670_));
  OAI21_X1   g06664(.A1(new_n7670_), .A2(new_n7661_), .B(new_n7650_), .ZN(new_n7671_));
  NOR2_X1    g06665(.A1(new_n7644_), .A2(\A[53] ), .ZN(new_n7672_));
  NOR2_X1    g06666(.A1(new_n7642_), .A2(\A[54] ), .ZN(new_n7673_));
  OAI21_X1   g06667(.A1(new_n7672_), .A2(new_n7673_), .B(\A[52] ), .ZN(new_n7674_));
  INV_X1     g06668(.I(new_n7648_), .ZN(new_n7675_));
  OAI21_X1   g06669(.A1(new_n7675_), .A2(new_n7221_), .B(new_n7641_), .ZN(new_n7676_));
  NAND2_X1   g06670(.A1(new_n7674_), .A2(new_n7676_), .ZN(new_n7677_));
  NAND3_X1   g06671(.A1(new_n7669_), .A2(new_n7655_), .A3(new_n7658_), .ZN(new_n7678_));
  NAND2_X1   g06672(.A1(new_n7659_), .A2(new_n7660_), .ZN(new_n7679_));
  NAND3_X1   g06673(.A1(new_n7679_), .A2(new_n7678_), .A3(new_n7677_), .ZN(new_n7680_));
  NAND2_X1   g06674(.A1(new_n7671_), .A2(new_n7680_), .ZN(new_n7681_));
  NAND2_X1   g06675(.A1(new_n7650_), .A2(new_n7635_), .ZN(new_n7682_));
  NAND2_X1   g06676(.A1(new_n7608_), .A2(new_n7677_), .ZN(new_n7683_));
  NAND2_X1   g06677(.A1(new_n7627_), .A2(new_n7659_), .ZN(new_n7684_));
  NAND2_X1   g06678(.A1(new_n7668_), .A2(new_n7618_), .ZN(new_n7685_));
  AOI22_X1   g06679(.A1(new_n7682_), .A2(new_n7683_), .B1(new_n7685_), .B2(new_n7684_), .ZN(new_n7686_));
  NOR3_X1    g06680(.A1(new_n7608_), .A2(new_n7620_), .A3(new_n7627_), .ZN(new_n7687_));
  NAND2_X1   g06681(.A1(new_n7223_), .A2(new_n7226_), .ZN(new_n7688_));
  NAND3_X1   g06682(.A1(new_n7677_), .A2(new_n7659_), .A3(new_n7688_), .ZN(new_n7689_));
  INV_X1     g06683(.I(new_n7689_), .ZN(new_n7690_));
  NAND4_X1   g06684(.A1(new_n7681_), .A2(new_n7686_), .A3(new_n7687_), .A4(new_n7690_), .ZN(new_n7691_));
  NOR2_X1    g06685(.A1(new_n7608_), .A2(new_n7677_), .ZN(new_n7692_));
  NOR2_X1    g06686(.A1(new_n7650_), .A2(new_n7635_), .ZN(new_n7693_));
  NOR2_X1    g06687(.A1(new_n7692_), .A2(new_n7693_), .ZN(new_n7694_));
  NOR2_X1    g06688(.A1(new_n7668_), .A2(new_n7618_), .ZN(new_n7695_));
  NOR2_X1    g06689(.A1(new_n7627_), .A2(new_n7659_), .ZN(new_n7696_));
  NOR2_X1    g06690(.A1(new_n7695_), .A2(new_n7696_), .ZN(new_n7697_));
  NAND3_X1   g06691(.A1(new_n7677_), .A2(new_n7659_), .A3(new_n7669_), .ZN(new_n7698_));
  OAI21_X1   g06692(.A1(new_n7694_), .A2(new_n7697_), .B(new_n7698_), .ZN(new_n7699_));
  OAI21_X1   g06693(.A1(new_n7699_), .A2(new_n7681_), .B(new_n7687_), .ZN(new_n7700_));
  AOI21_X1   g06694(.A1(new_n7700_), .A2(new_n7691_), .B(new_n7640_), .ZN(new_n7701_));
  AOI21_X1   g06695(.A1(new_n7679_), .A2(new_n7678_), .B(new_n7677_), .ZN(new_n7702_));
  NOR3_X1    g06696(.A1(new_n7670_), .A2(new_n7661_), .A3(new_n7650_), .ZN(new_n7703_));
  NOR2_X1    g06697(.A1(new_n7703_), .A2(new_n7702_), .ZN(new_n7704_));
  INV_X1     g06698(.I(new_n7698_), .ZN(new_n7705_));
  NOR2_X1    g06699(.A1(new_n7705_), .A2(new_n7687_), .ZN(new_n7706_));
  AOI21_X1   g06700(.A1(new_n7686_), .A2(new_n7706_), .B(new_n7704_), .ZN(new_n7707_));
  INV_X1     g06701(.I(new_n7686_), .ZN(new_n7708_));
  INV_X1     g06702(.I(new_n7687_), .ZN(new_n7709_));
  NAND2_X1   g06703(.A1(new_n7709_), .A2(new_n7698_), .ZN(new_n7710_));
  NOR3_X1    g06704(.A1(new_n7708_), .A2(new_n7681_), .A3(new_n7710_), .ZN(new_n7711_));
  OAI21_X1   g06705(.A1(new_n7707_), .A2(new_n7711_), .B(new_n7640_), .ZN(new_n7712_));
  INV_X1     g06706(.I(\A[40] ), .ZN(new_n7713_));
  INV_X1     g06707(.I(\A[41] ), .ZN(new_n7714_));
  NAND2_X1   g06708(.A1(new_n7714_), .A2(\A[42] ), .ZN(new_n7715_));
  INV_X1     g06709(.I(\A[42] ), .ZN(new_n7716_));
  NAND2_X1   g06710(.A1(new_n7716_), .A2(\A[41] ), .ZN(new_n7717_));
  AOI21_X1   g06711(.A1(new_n7715_), .A2(new_n7717_), .B(new_n7713_), .ZN(new_n7718_));
  INV_X1     g06712(.I(new_n7228_), .ZN(new_n7719_));
  NAND2_X1   g06713(.A1(\A[41] ), .A2(\A[42] ), .ZN(new_n7720_));
  AOI21_X1   g06714(.A1(new_n7719_), .A2(new_n7720_), .B(\A[40] ), .ZN(new_n7721_));
  NOR2_X1    g06715(.A1(new_n7721_), .A2(new_n7718_), .ZN(new_n7722_));
  INV_X1     g06716(.I(\A[37] ), .ZN(new_n7723_));
  INV_X1     g06717(.I(\A[38] ), .ZN(new_n7724_));
  NAND2_X1   g06718(.A1(new_n7724_), .A2(\A[39] ), .ZN(new_n7725_));
  INV_X1     g06719(.I(\A[39] ), .ZN(new_n7726_));
  NAND2_X1   g06720(.A1(new_n7726_), .A2(\A[38] ), .ZN(new_n7727_));
  AOI21_X1   g06721(.A1(new_n7725_), .A2(new_n7727_), .B(new_n7723_), .ZN(new_n7728_));
  INV_X1     g06722(.I(new_n7231_), .ZN(new_n7729_));
  NAND2_X1   g06723(.A1(\A[38] ), .A2(\A[39] ), .ZN(new_n7730_));
  AOI21_X1   g06724(.A1(new_n7729_), .A2(new_n7730_), .B(\A[37] ), .ZN(new_n7731_));
  OAI22_X1   g06725(.A1(new_n7228_), .A2(new_n7229_), .B1(new_n7232_), .B2(new_n7231_), .ZN(new_n7732_));
  NOR3_X1    g06726(.A1(new_n7731_), .A2(new_n7732_), .A3(new_n7728_), .ZN(new_n7733_));
  NOR2_X1    g06727(.A1(new_n7731_), .A2(new_n7728_), .ZN(new_n7734_));
  NOR2_X1    g06728(.A1(new_n7230_), .A2(new_n7233_), .ZN(new_n7735_));
  NOR2_X1    g06729(.A1(new_n7734_), .A2(new_n7735_), .ZN(new_n7736_));
  OAI21_X1   g06730(.A1(new_n7736_), .A2(new_n7733_), .B(new_n7722_), .ZN(new_n7737_));
  NOR2_X1    g06731(.A1(new_n7716_), .A2(\A[41] ), .ZN(new_n7738_));
  NOR2_X1    g06732(.A1(new_n7714_), .A2(\A[42] ), .ZN(new_n7739_));
  OAI21_X1   g06733(.A1(new_n7738_), .A2(new_n7739_), .B(\A[40] ), .ZN(new_n7740_));
  INV_X1     g06734(.I(new_n7720_), .ZN(new_n7741_));
  OAI21_X1   g06735(.A1(new_n7741_), .A2(new_n7228_), .B(new_n7713_), .ZN(new_n7742_));
  NAND2_X1   g06736(.A1(new_n7740_), .A2(new_n7742_), .ZN(new_n7743_));
  NOR2_X1    g06737(.A1(new_n7726_), .A2(\A[38] ), .ZN(new_n7744_));
  NOR2_X1    g06738(.A1(new_n7724_), .A2(\A[39] ), .ZN(new_n7745_));
  OAI21_X1   g06739(.A1(new_n7744_), .A2(new_n7745_), .B(\A[37] ), .ZN(new_n7746_));
  INV_X1     g06740(.I(new_n7730_), .ZN(new_n7747_));
  OAI21_X1   g06741(.A1(new_n7747_), .A2(new_n7231_), .B(new_n7723_), .ZN(new_n7748_));
  NAND3_X1   g06742(.A1(new_n7735_), .A2(new_n7746_), .A3(new_n7748_), .ZN(new_n7749_));
  OAI21_X1   g06743(.A1(new_n7728_), .A2(new_n7731_), .B(new_n7732_), .ZN(new_n7750_));
  NAND3_X1   g06744(.A1(new_n7749_), .A2(new_n7750_), .A3(new_n7743_), .ZN(new_n7751_));
  NAND2_X1   g06745(.A1(new_n7737_), .A2(new_n7751_), .ZN(new_n7752_));
  INV_X1     g06746(.I(\A[36] ), .ZN(new_n7753_));
  NOR2_X1    g06747(.A1(new_n7753_), .A2(\A[35] ), .ZN(new_n7754_));
  INV_X1     g06748(.I(\A[35] ), .ZN(new_n7755_));
  NOR2_X1    g06749(.A1(new_n7755_), .A2(\A[36] ), .ZN(new_n7756_));
  OAI21_X1   g06750(.A1(new_n7754_), .A2(new_n7756_), .B(\A[34] ), .ZN(new_n7757_));
  INV_X1     g06751(.I(new_n7206_), .ZN(new_n7758_));
  OAI21_X1   g06752(.A1(new_n7758_), .A2(new_n7205_), .B(new_n7204_), .ZN(new_n7759_));
  NAND2_X1   g06753(.A1(new_n7757_), .A2(new_n7759_), .ZN(new_n7760_));
  NOR2_X1    g06754(.A1(new_n7722_), .A2(new_n7760_), .ZN(new_n7761_));
  NAND2_X1   g06755(.A1(new_n7755_), .A2(\A[36] ), .ZN(new_n7762_));
  NAND2_X1   g06756(.A1(new_n7753_), .A2(\A[35] ), .ZN(new_n7763_));
  AOI21_X1   g06757(.A1(new_n7762_), .A2(new_n7763_), .B(new_n7204_), .ZN(new_n7764_));
  INV_X1     g06758(.I(new_n7205_), .ZN(new_n7765_));
  AOI21_X1   g06759(.A1(new_n7765_), .A2(new_n7206_), .B(\A[34] ), .ZN(new_n7766_));
  NOR2_X1    g06760(.A1(new_n7766_), .A2(new_n7764_), .ZN(new_n7767_));
  NOR2_X1    g06761(.A1(new_n7767_), .A2(new_n7743_), .ZN(new_n7768_));
  NAND2_X1   g06762(.A1(new_n7746_), .A2(new_n7748_), .ZN(new_n7769_));
  INV_X1     g06763(.I(\A[32] ), .ZN(new_n7770_));
  NAND2_X1   g06764(.A1(new_n7770_), .A2(\A[33] ), .ZN(new_n7771_));
  INV_X1     g06765(.I(\A[33] ), .ZN(new_n7772_));
  NAND2_X1   g06766(.A1(new_n7772_), .A2(\A[32] ), .ZN(new_n7773_));
  AOI21_X1   g06767(.A1(new_n7771_), .A2(new_n7773_), .B(new_n7208_), .ZN(new_n7774_));
  INV_X1     g06768(.I(new_n7209_), .ZN(new_n7775_));
  AOI21_X1   g06769(.A1(new_n7775_), .A2(new_n7210_), .B(\A[31] ), .ZN(new_n7776_));
  NOR2_X1    g06770(.A1(new_n7776_), .A2(new_n7774_), .ZN(new_n7777_));
  NOR2_X1    g06771(.A1(new_n7777_), .A2(new_n7769_), .ZN(new_n7778_));
  NOR2_X1    g06772(.A1(new_n7772_), .A2(\A[32] ), .ZN(new_n7779_));
  NOR2_X1    g06773(.A1(new_n7770_), .A2(\A[33] ), .ZN(new_n7780_));
  OAI21_X1   g06774(.A1(new_n7779_), .A2(new_n7780_), .B(\A[31] ), .ZN(new_n7781_));
  INV_X1     g06775(.I(new_n7210_), .ZN(new_n7782_));
  OAI21_X1   g06776(.A1(new_n7782_), .A2(new_n7209_), .B(new_n7208_), .ZN(new_n7783_));
  NAND2_X1   g06777(.A1(new_n7781_), .A2(new_n7783_), .ZN(new_n7784_));
  NOR2_X1    g06778(.A1(new_n7734_), .A2(new_n7784_), .ZN(new_n7785_));
  OAI22_X1   g06779(.A1(new_n7761_), .A2(new_n7768_), .B1(new_n7778_), .B2(new_n7785_), .ZN(new_n7786_));
  NAND2_X1   g06780(.A1(new_n7230_), .A2(new_n7233_), .ZN(new_n7787_));
  AOI22_X1   g06781(.A1(new_n7740_), .A2(new_n7742_), .B1(new_n7746_), .B2(new_n7748_), .ZN(new_n7788_));
  AOI21_X1   g06782(.A1(new_n7788_), .A2(new_n7787_), .B(new_n7735_), .ZN(new_n7789_));
  NOR3_X1    g06783(.A1(new_n7752_), .A2(new_n7786_), .A3(new_n7789_), .ZN(new_n7790_));
  NOR2_X1    g06784(.A1(new_n7207_), .A2(new_n7211_), .ZN(new_n7791_));
  NAND3_X1   g06785(.A1(new_n7760_), .A2(new_n7784_), .A3(new_n7791_), .ZN(new_n7792_));
  INV_X1     g06786(.I(new_n7792_), .ZN(new_n7793_));
  NOR4_X1    g06787(.A1(new_n7718_), .A2(new_n7721_), .A3(new_n7731_), .A4(new_n7728_), .ZN(new_n7794_));
  NOR2_X1    g06788(.A1(new_n7788_), .A2(new_n7794_), .ZN(new_n7795_));
  AOI21_X1   g06789(.A1(new_n7789_), .A2(new_n7795_), .B(new_n7793_), .ZN(new_n7796_));
  NAND2_X1   g06790(.A1(new_n7777_), .A2(new_n7791_), .ZN(new_n7797_));
  INV_X1     g06791(.I(new_n7791_), .ZN(new_n7798_));
  NAND2_X1   g06792(.A1(new_n7798_), .A2(new_n7784_), .ZN(new_n7799_));
  AOI21_X1   g06793(.A1(new_n7799_), .A2(new_n7797_), .B(new_n7760_), .ZN(new_n7800_));
  NOR2_X1    g06794(.A1(new_n7798_), .A2(new_n7784_), .ZN(new_n7801_));
  NOR2_X1    g06795(.A1(new_n7777_), .A2(new_n7791_), .ZN(new_n7802_));
  NOR3_X1    g06796(.A1(new_n7801_), .A2(new_n7802_), .A3(new_n7767_), .ZN(new_n7803_));
  NOR2_X1    g06797(.A1(new_n7803_), .A2(new_n7800_), .ZN(new_n7804_));
  NAND2_X1   g06798(.A1(new_n7767_), .A2(new_n7743_), .ZN(new_n7805_));
  NAND2_X1   g06799(.A1(new_n7722_), .A2(new_n7760_), .ZN(new_n7806_));
  NAND2_X1   g06800(.A1(new_n7734_), .A2(new_n7784_), .ZN(new_n7807_));
  NAND2_X1   g06801(.A1(new_n7777_), .A2(new_n7769_), .ZN(new_n7808_));
  AOI22_X1   g06802(.A1(new_n7805_), .A2(new_n7806_), .B1(new_n7807_), .B2(new_n7808_), .ZN(new_n7809_));
  NOR3_X1    g06803(.A1(new_n7722_), .A2(new_n7734_), .A3(new_n7732_), .ZN(new_n7810_));
  NOR3_X1    g06804(.A1(new_n7752_), .A2(new_n7809_), .A3(new_n7810_), .ZN(new_n7811_));
  NOR3_X1    g06805(.A1(new_n7811_), .A2(new_n7792_), .A3(new_n7804_), .ZN(new_n7812_));
  OAI21_X1   g06806(.A1(new_n7812_), .A2(new_n7796_), .B(new_n7790_), .ZN(new_n7813_));
  OR2_X2     g06807(.A1(new_n7803_), .A2(new_n7800_), .Z(new_n7814_));
  INV_X1     g06808(.I(new_n7810_), .ZN(new_n7815_));
  NAND2_X1   g06809(.A1(new_n7815_), .A2(new_n7792_), .ZN(new_n7816_));
  OAI21_X1   g06810(.A1(new_n7786_), .A2(new_n7816_), .B(new_n7752_), .ZN(new_n7817_));
  AOI21_X1   g06811(.A1(new_n7749_), .A2(new_n7750_), .B(new_n7743_), .ZN(new_n7818_));
  NOR3_X1    g06812(.A1(new_n7736_), .A2(new_n7722_), .A3(new_n7733_), .ZN(new_n7819_));
  NOR2_X1    g06813(.A1(new_n7819_), .A2(new_n7818_), .ZN(new_n7820_));
  NOR2_X1    g06814(.A1(new_n7793_), .A2(new_n7810_), .ZN(new_n7821_));
  NAND3_X1   g06815(.A1(new_n7820_), .A2(new_n7821_), .A3(new_n7809_), .ZN(new_n7822_));
  AOI21_X1   g06816(.A1(new_n7817_), .A2(new_n7822_), .B(new_n7814_), .ZN(new_n7823_));
  NOR2_X1    g06817(.A1(new_n7220_), .A2(new_n7212_), .ZN(new_n7824_));
  NOR2_X1    g06818(.A1(new_n7240_), .A2(new_n7219_), .ZN(new_n7825_));
  NOR2_X1    g06819(.A1(new_n7825_), .A2(new_n7824_), .ZN(new_n7826_));
  NOR2_X1    g06820(.A1(new_n7826_), .A2(new_n7237_), .ZN(new_n7827_));
  INV_X1     g06821(.I(new_n7827_), .ZN(new_n7828_));
  NOR2_X1    g06822(.A1(new_n7823_), .A2(new_n7828_), .ZN(new_n7829_));
  NAND3_X1   g06823(.A1(new_n7829_), .A2(new_n7813_), .A3(new_n7712_), .ZN(new_n7830_));
  OAI21_X1   g06824(.A1(new_n7708_), .A2(new_n7710_), .B(new_n7681_), .ZN(new_n7831_));
  NAND3_X1   g06825(.A1(new_n7704_), .A2(new_n7686_), .A3(new_n7706_), .ZN(new_n7832_));
  AOI21_X1   g06826(.A1(new_n7831_), .A2(new_n7832_), .B(new_n7639_), .ZN(new_n7833_));
  INV_X1     g06827(.I(new_n7790_), .ZN(new_n7834_));
  INV_X1     g06828(.I(new_n7796_), .ZN(new_n7835_));
  NAND3_X1   g06829(.A1(new_n7820_), .A2(new_n7786_), .A3(new_n7815_), .ZN(new_n7836_));
  NAND3_X1   g06830(.A1(new_n7836_), .A2(new_n7814_), .A3(new_n7793_), .ZN(new_n7837_));
  AOI21_X1   g06831(.A1(new_n7837_), .A2(new_n7835_), .B(new_n7834_), .ZN(new_n7838_));
  AOI21_X1   g06832(.A1(new_n7809_), .A2(new_n7821_), .B(new_n7820_), .ZN(new_n7839_));
  NOR3_X1    g06833(.A1(new_n7752_), .A2(new_n7816_), .A3(new_n7786_), .ZN(new_n7840_));
  OAI21_X1   g06834(.A1(new_n7839_), .A2(new_n7840_), .B(new_n7804_), .ZN(new_n7841_));
  NAND2_X1   g06835(.A1(new_n7841_), .A2(new_n7827_), .ZN(new_n7842_));
  OAI21_X1   g06836(.A1(new_n7842_), .A2(new_n7838_), .B(new_n7833_), .ZN(new_n7843_));
  AOI21_X1   g06837(.A1(new_n7843_), .A2(new_n7830_), .B(new_n7701_), .ZN(new_n7844_));
  NOR4_X1    g06838(.A1(new_n7708_), .A2(new_n7704_), .A3(new_n7709_), .A4(new_n7689_), .ZN(new_n7845_));
  NAND2_X1   g06839(.A1(new_n7682_), .A2(new_n7683_), .ZN(new_n7846_));
  NAND2_X1   g06840(.A1(new_n7685_), .A2(new_n7684_), .ZN(new_n7847_));
  AOI21_X1   g06841(.A1(new_n7846_), .A2(new_n7847_), .B(new_n7705_), .ZN(new_n7848_));
  AOI21_X1   g06842(.A1(new_n7848_), .A2(new_n7704_), .B(new_n7709_), .ZN(new_n7849_));
  OAI21_X1   g06843(.A1(new_n7845_), .A2(new_n7849_), .B(new_n7639_), .ZN(new_n7850_));
  NOR3_X1    g06844(.A1(new_n7842_), .A2(new_n7838_), .A3(new_n7833_), .ZN(new_n7851_));
  AOI21_X1   g06845(.A1(new_n7829_), .A2(new_n7813_), .B(new_n7712_), .ZN(new_n7852_));
  NOR3_X1    g06846(.A1(new_n7852_), .A2(new_n7851_), .A3(new_n7850_), .ZN(new_n7853_));
  OAI21_X1   g06847(.A1(new_n7853_), .A2(new_n7844_), .B(new_n7598_), .ZN(new_n7854_));
  NAND2_X1   g06848(.A1(new_n7854_), .A2(new_n7597_), .ZN(new_n7855_));
  NOR3_X1    g06849(.A1(new_n7251_), .A2(new_n7477_), .A3(new_n7485_), .ZN(new_n7856_));
  OAI21_X1   g06850(.A1(new_n7855_), .A2(new_n7856_), .B(new_n7486_), .ZN(new_n7857_));
  INV_X1     g06851(.I(new_n7597_), .ZN(new_n7858_));
  NOR3_X1    g06852(.A1(new_n7598_), .A2(new_n7853_), .A3(new_n7844_), .ZN(new_n7859_));
  OAI21_X1   g06853(.A1(new_n7858_), .A2(new_n7859_), .B(new_n7854_), .ZN(new_n7860_));
  XOR2_X1    g06854(.A1(new_n7212_), .A2(new_n7219_), .Z(new_n7861_));
  NAND3_X1   g06855(.A1(new_n7235_), .A2(new_n7861_), .A3(new_n7639_), .ZN(new_n7862_));
  AOI21_X1   g06856(.A1(new_n7862_), .A2(new_n7700_), .B(new_n7691_), .ZN(new_n7863_));
  NAND2_X1   g06857(.A1(new_n7838_), .A2(new_n7863_), .ZN(new_n7864_));
  NAND2_X1   g06858(.A1(new_n7833_), .A2(new_n7823_), .ZN(new_n7865_));
  NAND2_X1   g06859(.A1(new_n7864_), .A2(new_n7865_), .ZN(new_n7866_));
  OAI21_X1   g06860(.A1(new_n7833_), .A2(new_n7701_), .B(new_n7827_), .ZN(new_n7867_));
  OAI21_X1   g06861(.A1(new_n7811_), .A2(new_n7792_), .B(new_n7814_), .ZN(new_n7868_));
  NOR4_X1    g06862(.A1(new_n7752_), .A2(new_n7786_), .A3(new_n7789_), .A4(new_n7793_), .ZN(new_n7869_));
  NAND3_X1   g06863(.A1(new_n7737_), .A2(new_n7795_), .A3(new_n7751_), .ZN(new_n7870_));
  AND2_X2    g06864(.A1(new_n7207_), .A2(new_n7211_), .Z(new_n7871_));
  NAND2_X1   g06865(.A1(new_n7760_), .A2(new_n7784_), .ZN(new_n7872_));
  OAI21_X1   g06866(.A1(new_n7872_), .A2(new_n7871_), .B(new_n7798_), .ZN(new_n7873_));
  NAND3_X1   g06867(.A1(new_n7870_), .A2(new_n7789_), .A3(new_n7873_), .ZN(new_n7874_));
  NOR2_X1    g06868(.A1(new_n7869_), .A2(new_n7874_), .ZN(new_n7875_));
  INV_X1     g06869(.I(new_n7789_), .ZN(new_n7876_));
  NAND4_X1   g06870(.A1(new_n7820_), .A2(new_n7809_), .A3(new_n7876_), .A4(new_n7792_), .ZN(new_n7877_));
  NOR4_X1    g06871(.A1(new_n7819_), .A2(new_n7818_), .A3(new_n7788_), .A4(new_n7794_), .ZN(new_n7878_));
  INV_X1     g06872(.I(new_n7873_), .ZN(new_n7879_));
  NOR3_X1    g06873(.A1(new_n7878_), .A2(new_n7876_), .A3(new_n7879_), .ZN(new_n7880_));
  NOR2_X1    g06874(.A1(new_n7880_), .A2(new_n7877_), .ZN(new_n7881_));
  OAI21_X1   g06875(.A1(new_n7881_), .A2(new_n7875_), .B(new_n7868_), .ZN(new_n7882_));
  AOI21_X1   g06876(.A1(new_n7836_), .A2(new_n7793_), .B(new_n7804_), .ZN(new_n7883_));
  NAND2_X1   g06877(.A1(new_n7880_), .A2(new_n7877_), .ZN(new_n7884_));
  NAND2_X1   g06878(.A1(new_n7869_), .A2(new_n7874_), .ZN(new_n7885_));
  NAND3_X1   g06879(.A1(new_n7884_), .A2(new_n7885_), .A3(new_n7883_), .ZN(new_n7886_));
  NAND2_X1   g06880(.A1(new_n7882_), .A2(new_n7886_), .ZN(new_n7887_));
  NAND2_X1   g06881(.A1(new_n7689_), .A2(new_n7660_), .ZN(new_n7888_));
  NAND2_X1   g06882(.A1(new_n7215_), .A2(new_n7218_), .ZN(new_n7889_));
  NAND3_X1   g06883(.A1(new_n7635_), .A2(new_n7618_), .A3(new_n7889_), .ZN(new_n7890_));
  NAND2_X1   g06884(.A1(new_n7890_), .A2(new_n7620_), .ZN(new_n7891_));
  NAND2_X1   g06885(.A1(new_n7891_), .A2(new_n7888_), .ZN(new_n7892_));
  AOI21_X1   g06886(.A1(new_n7700_), .A2(new_n7639_), .B(new_n7892_), .ZN(new_n7893_));
  INV_X1     g06887(.I(new_n7892_), .ZN(new_n7894_));
  NOR3_X1    g06888(.A1(new_n7849_), .A2(new_n7640_), .A3(new_n7894_), .ZN(new_n7895_));
  OAI21_X1   g06889(.A1(new_n7893_), .A2(new_n7895_), .B(new_n7691_), .ZN(new_n7896_));
  OAI21_X1   g06890(.A1(new_n7849_), .A2(new_n7640_), .B(new_n7894_), .ZN(new_n7897_));
  NAND3_X1   g06891(.A1(new_n7700_), .A2(new_n7639_), .A3(new_n7892_), .ZN(new_n7898_));
  NAND3_X1   g06892(.A1(new_n7897_), .A2(new_n7898_), .A3(new_n7845_), .ZN(new_n7899_));
  NAND2_X1   g06893(.A1(new_n7896_), .A2(new_n7899_), .ZN(new_n7900_));
  NAND3_X1   g06894(.A1(new_n7900_), .A2(new_n7887_), .A3(new_n7867_), .ZN(new_n7901_));
  AOI21_X1   g06895(.A1(new_n7850_), .A2(new_n7712_), .B(new_n7828_), .ZN(new_n7902_));
  AOI21_X1   g06896(.A1(new_n7884_), .A2(new_n7885_), .B(new_n7883_), .ZN(new_n7903_));
  NOR3_X1    g06897(.A1(new_n7881_), .A2(new_n7868_), .A3(new_n7875_), .ZN(new_n7904_));
  NOR2_X1    g06898(.A1(new_n7904_), .A2(new_n7903_), .ZN(new_n7905_));
  AOI21_X1   g06899(.A1(new_n7897_), .A2(new_n7898_), .B(new_n7845_), .ZN(new_n7906_));
  NOR3_X1    g06900(.A1(new_n7893_), .A2(new_n7895_), .A3(new_n7691_), .ZN(new_n7907_));
  NOR2_X1    g06901(.A1(new_n7906_), .A2(new_n7907_), .ZN(new_n7908_));
  OAI21_X1   g06902(.A1(new_n7908_), .A2(new_n7905_), .B(new_n7902_), .ZN(new_n7909_));
  AOI21_X1   g06903(.A1(new_n7909_), .A2(new_n7901_), .B(new_n7866_), .ZN(new_n7910_));
  NOR3_X1    g06904(.A1(new_n7640_), .A2(new_n7237_), .A3(new_n7826_), .ZN(new_n7911_));
  OAI21_X1   g06905(.A1(new_n7911_), .A2(new_n7849_), .B(new_n7845_), .ZN(new_n7912_));
  NOR2_X1    g06906(.A1(new_n7813_), .A2(new_n7912_), .ZN(new_n7913_));
  INV_X1     g06907(.I(new_n7865_), .ZN(new_n7914_));
  NOR2_X1    g06908(.A1(new_n7913_), .A2(new_n7914_), .ZN(new_n7915_));
  NOR3_X1    g06909(.A1(new_n7908_), .A2(new_n7905_), .A3(new_n7902_), .ZN(new_n7916_));
  AOI21_X1   g06910(.A1(new_n7900_), .A2(new_n7887_), .B(new_n7867_), .ZN(new_n7917_));
  NOR3_X1    g06911(.A1(new_n7916_), .A2(new_n7917_), .A3(new_n7915_), .ZN(new_n7918_));
  XOR2_X1    g06912(.A1(new_n7109_), .A2(new_n7197_), .Z(new_n7919_));
  AOI21_X1   g06913(.A1(new_n7561_), .A2(new_n7562_), .B(new_n7560_), .ZN(new_n7920_));
  NOR3_X1    g06914(.A1(new_n7553_), .A2(new_n7548_), .A3(new_n7183_), .ZN(new_n7921_));
  NOR2_X1    g06915(.A1(new_n7921_), .A2(new_n7920_), .ZN(new_n7922_));
  NAND2_X1   g06916(.A1(new_n7183_), .A2(new_n7105_), .ZN(new_n7923_));
  NAND3_X1   g06917(.A1(new_n7560_), .A2(new_n7099_), .A3(new_n7104_), .ZN(new_n7924_));
  NAND2_X1   g06918(.A1(new_n7094_), .A2(new_n7172_), .ZN(new_n7925_));
  NAND3_X1   g06919(.A1(new_n7573_), .A2(new_n7167_), .A3(new_n7171_), .ZN(new_n7926_));
  AOI22_X1   g06920(.A1(new_n7923_), .A2(new_n7924_), .B1(new_n7926_), .B2(new_n7925_), .ZN(new_n7927_));
  INV_X1     g06921(.I(new_n7580_), .ZN(new_n7928_));
  NAND2_X1   g06922(.A1(new_n7928_), .A2(new_n7927_), .ZN(new_n7929_));
  INV_X1     g06923(.I(new_n7585_), .ZN(new_n7930_));
  NAND3_X1   g06924(.A1(new_n7584_), .A2(new_n7582_), .A3(new_n7105_), .ZN(new_n7931_));
  NAND2_X1   g06925(.A1(new_n7930_), .A2(new_n7931_), .ZN(new_n7932_));
  NAND3_X1   g06926(.A1(new_n7932_), .A2(new_n7929_), .A3(new_n7922_), .ZN(new_n7933_));
  NOR3_X1    g06927(.A1(new_n7919_), .A2(new_n7933_), .A3(new_n7198_), .ZN(new_n7934_));
  OAI21_X1   g06928(.A1(new_n7919_), .A2(new_n7198_), .B(new_n7933_), .ZN(new_n7935_));
  NOR4_X1    g06929(.A1(new_n7495_), .A2(new_n7506_), .A3(new_n7533_), .A4(new_n7537_), .ZN(new_n7936_));
  NAND4_X1   g06930(.A1(new_n7936_), .A2(new_n7495_), .A3(new_n7510_), .A4(new_n7533_), .ZN(new_n7937_));
  INV_X1     g06931(.I(new_n7937_), .ZN(new_n7938_));
  AOI21_X1   g06932(.A1(new_n7938_), .A2(new_n7935_), .B(new_n7934_), .ZN(new_n7939_));
  NOR3_X1    g06933(.A1(new_n7576_), .A2(new_n7592_), .A3(new_n7922_), .ZN(new_n7940_));
  AOI21_X1   g06934(.A1(new_n7928_), .A2(new_n7927_), .B(new_n7564_), .ZN(new_n7941_));
  NAND2_X1   g06935(.A1(new_n7106_), .A2(new_n7107_), .ZN(new_n7942_));
  NAND3_X1   g06936(.A1(new_n7573_), .A2(new_n7105_), .A3(new_n7942_), .ZN(new_n7943_));
  AOI22_X1   g06937(.A1(new_n7943_), .A2(new_n7583_), .B1(new_n7591_), .B2(new_n7186_), .ZN(new_n7944_));
  OAI21_X1   g06938(.A1(new_n7941_), .A2(new_n7589_), .B(new_n7944_), .ZN(new_n7945_));
  OAI21_X1   g06939(.A1(new_n7576_), .A2(new_n7580_), .B(new_n7922_), .ZN(new_n7946_));
  INV_X1     g06940(.I(new_n7944_), .ZN(new_n7947_));
  NAND3_X1   g06941(.A1(new_n7946_), .A2(new_n7932_), .A3(new_n7947_), .ZN(new_n7948_));
  AOI21_X1   g06942(.A1(new_n7948_), .A2(new_n7945_), .B(new_n7940_), .ZN(new_n7949_));
  INV_X1     g06943(.I(new_n7940_), .ZN(new_n7950_));
  AOI21_X1   g06944(.A1(new_n7946_), .A2(new_n7932_), .B(new_n7947_), .ZN(new_n7951_));
  NOR3_X1    g06945(.A1(new_n7941_), .A2(new_n7589_), .A3(new_n7944_), .ZN(new_n7952_));
  NOR3_X1    g06946(.A1(new_n7951_), .A2(new_n7952_), .A3(new_n7950_), .ZN(new_n7953_));
  NOR2_X1    g06947(.A1(new_n7953_), .A2(new_n7949_), .ZN(new_n7954_));
  INV_X1     g06948(.I(new_n7538_), .ZN(new_n7955_));
  OAI21_X1   g06949(.A1(new_n7506_), .A2(new_n7509_), .B(new_n7533_), .ZN(new_n7956_));
  NAND2_X1   g06950(.A1(new_n7133_), .A2(new_n7134_), .ZN(new_n7957_));
  NAND3_X1   g06951(.A1(new_n7196_), .A2(new_n7132_), .A3(new_n7957_), .ZN(new_n7958_));
  AOI22_X1   g06952(.A1(new_n7958_), .A2(new_n7488_), .B1(new_n7536_), .B2(new_n7160_), .ZN(new_n7959_));
  INV_X1     g06953(.I(new_n7959_), .ZN(new_n7960_));
  AOI21_X1   g06954(.A1(new_n7956_), .A2(new_n7534_), .B(new_n7960_), .ZN(new_n7961_));
  NAND2_X1   g06955(.A1(new_n7157_), .A2(new_n7132_), .ZN(new_n7962_));
  NAND3_X1   g06956(.A1(new_n7501_), .A2(new_n7126_), .A3(new_n7131_), .ZN(new_n7963_));
  NAND2_X1   g06957(.A1(new_n7121_), .A2(new_n7146_), .ZN(new_n7964_));
  NAND3_X1   g06958(.A1(new_n7196_), .A2(new_n7141_), .A3(new_n7145_), .ZN(new_n7965_));
  AOI22_X1   g06959(.A1(new_n7962_), .A2(new_n7963_), .B1(new_n7965_), .B2(new_n7964_), .ZN(new_n7966_));
  AND2_X2    g06960(.A1(new_n7507_), .A2(new_n7508_), .Z(new_n7967_));
  AOI21_X1   g06961(.A1(new_n7967_), .A2(new_n7966_), .B(new_n7527_), .ZN(new_n7968_));
  NOR3_X1    g06962(.A1(new_n7968_), .A2(new_n7959_), .A3(new_n7495_), .ZN(new_n7969_));
  OAI21_X1   g06963(.A1(new_n7961_), .A2(new_n7969_), .B(new_n7955_), .ZN(new_n7970_));
  OAI21_X1   g06964(.A1(new_n7968_), .A2(new_n7495_), .B(new_n7959_), .ZN(new_n7971_));
  NAND3_X1   g06965(.A1(new_n7956_), .A2(new_n7534_), .A3(new_n7960_), .ZN(new_n7972_));
  NAND3_X1   g06966(.A1(new_n7972_), .A2(new_n7971_), .A3(new_n7538_), .ZN(new_n7973_));
  NAND2_X1   g06967(.A1(new_n7970_), .A2(new_n7973_), .ZN(new_n7974_));
  NAND2_X1   g06968(.A1(new_n7954_), .A2(new_n7974_), .ZN(new_n7975_));
  OAI21_X1   g06969(.A1(new_n7951_), .A2(new_n7952_), .B(new_n7950_), .ZN(new_n7976_));
  NAND3_X1   g06970(.A1(new_n7948_), .A2(new_n7945_), .A3(new_n7940_), .ZN(new_n7977_));
  NAND2_X1   g06971(.A1(new_n7976_), .A2(new_n7977_), .ZN(new_n7978_));
  AOI21_X1   g06972(.A1(new_n7972_), .A2(new_n7971_), .B(new_n7538_), .ZN(new_n7979_));
  NOR3_X1    g06973(.A1(new_n7961_), .A2(new_n7969_), .A3(new_n7955_), .ZN(new_n7980_));
  NOR2_X1    g06974(.A1(new_n7979_), .A2(new_n7980_), .ZN(new_n7981_));
  NAND2_X1   g06975(.A1(new_n7981_), .A2(new_n7978_), .ZN(new_n7982_));
  AOI21_X1   g06976(.A1(new_n7975_), .A2(new_n7982_), .B(new_n7939_), .ZN(new_n7983_));
  AOI21_X1   g06977(.A1(new_n7189_), .A2(new_n7541_), .B(new_n7594_), .ZN(new_n7984_));
  OAI21_X1   g06978(.A1(new_n7984_), .A2(new_n7937_), .B(new_n7595_), .ZN(new_n7985_));
  NAND2_X1   g06979(.A1(new_n7978_), .A2(new_n7974_), .ZN(new_n7986_));
  NAND4_X1   g06980(.A1(new_n7976_), .A2(new_n7977_), .A3(new_n7970_), .A4(new_n7973_), .ZN(new_n7987_));
  AOI21_X1   g06981(.A1(new_n7986_), .A2(new_n7987_), .B(new_n7985_), .ZN(new_n7988_));
  NOR2_X1    g06982(.A1(new_n7983_), .A2(new_n7988_), .ZN(new_n7989_));
  NOR3_X1    g06983(.A1(new_n7989_), .A2(new_n7910_), .A3(new_n7918_), .ZN(new_n7990_));
  OAI21_X1   g06984(.A1(new_n7916_), .A2(new_n7917_), .B(new_n7915_), .ZN(new_n7991_));
  NAND3_X1   g06985(.A1(new_n7909_), .A2(new_n7901_), .A3(new_n7866_), .ZN(new_n7992_));
  NOR2_X1    g06986(.A1(new_n7981_), .A2(new_n7978_), .ZN(new_n7993_));
  NOR2_X1    g06987(.A1(new_n7954_), .A2(new_n7974_), .ZN(new_n7994_));
  OAI21_X1   g06988(.A1(new_n7993_), .A2(new_n7994_), .B(new_n7985_), .ZN(new_n7995_));
  AOI22_X1   g06989(.A1(new_n7976_), .A2(new_n7977_), .B1(new_n7970_), .B2(new_n7973_), .ZN(new_n7996_));
  NOR4_X1    g06990(.A1(new_n7949_), .A2(new_n7953_), .A3(new_n7979_), .A4(new_n7980_), .ZN(new_n7997_));
  OAI21_X1   g06991(.A1(new_n7997_), .A2(new_n7996_), .B(new_n7939_), .ZN(new_n7998_));
  NAND2_X1   g06992(.A1(new_n7995_), .A2(new_n7998_), .ZN(new_n7999_));
  AOI21_X1   g06993(.A1(new_n7991_), .A2(new_n7992_), .B(new_n7999_), .ZN(new_n8000_));
  OAI21_X1   g06994(.A1(new_n8000_), .A2(new_n7990_), .B(new_n7860_), .ZN(new_n8001_));
  OAI21_X1   g06995(.A1(new_n7852_), .A2(new_n7851_), .B(new_n7850_), .ZN(new_n8002_));
  NAND3_X1   g06996(.A1(new_n7843_), .A2(new_n7830_), .A3(new_n7701_), .ZN(new_n8003_));
  AOI21_X1   g06997(.A1(new_n8002_), .A2(new_n8003_), .B(new_n7249_), .ZN(new_n8004_));
  NAND3_X1   g06998(.A1(new_n8002_), .A2(new_n8003_), .A3(new_n7249_), .ZN(new_n8005_));
  AOI21_X1   g06999(.A1(new_n7597_), .A2(new_n8005_), .B(new_n8004_), .ZN(new_n8006_));
  AOI22_X1   g07000(.A1(new_n7991_), .A2(new_n7992_), .B1(new_n7995_), .B2(new_n7998_), .ZN(new_n8007_));
  NOR3_X1    g07001(.A1(new_n7999_), .A2(new_n7910_), .A3(new_n7918_), .ZN(new_n8008_));
  OAI21_X1   g07002(.A1(new_n8008_), .A2(new_n8007_), .B(new_n8006_), .ZN(new_n8009_));
  NAND2_X1   g07003(.A1(new_n7403_), .A2(new_n7380_), .ZN(new_n8010_));
  NOR4_X1    g07004(.A1(new_n7397_), .A2(new_n7394_), .A3(new_n7311_), .A4(new_n7314_), .ZN(new_n8011_));
  AOI21_X1   g07005(.A1(new_n8010_), .A2(new_n8011_), .B(new_n7482_), .ZN(new_n8012_));
  NOR4_X1    g07006(.A1(new_n7078_), .A2(new_n7428_), .A3(new_n7430_), .A4(new_n7457_), .ZN(new_n8013_));
  INV_X1     g07007(.I(new_n8013_), .ZN(new_n8014_));
  NAND2_X1   g07008(.A1(new_n7017_), .A2(new_n7021_), .ZN(new_n8015_));
  NOR2_X1    g07009(.A1(new_n7440_), .A2(new_n7449_), .ZN(new_n8016_));
  AOI21_X1   g07010(.A1(new_n8016_), .A2(new_n8015_), .B(new_n7450_), .ZN(new_n8017_));
  INV_X1     g07011(.I(new_n8017_), .ZN(new_n8018_));
  INV_X1     g07012(.I(new_n7414_), .ZN(new_n8019_));
  OAI22_X1   g07013(.A1(new_n7029_), .A2(new_n8019_), .B1(new_n7415_), .B2(new_n7416_), .ZN(new_n8020_));
  OAI22_X1   g07014(.A1(new_n8020_), .A2(new_n7412_), .B1(new_n7070_), .B2(new_n7414_), .ZN(new_n8021_));
  NAND3_X1   g07015(.A1(new_n7464_), .A2(new_n8021_), .A3(new_n7465_), .ZN(new_n8022_));
  AOI21_X1   g07016(.A1(new_n7070_), .A2(new_n7414_), .B(new_n7417_), .ZN(new_n8023_));
  AOI22_X1   g07017(.A1(new_n7461_), .A2(new_n8023_), .B1(new_n7029_), .B2(new_n8019_), .ZN(new_n8024_));
  NAND2_X1   g07018(.A1(new_n7428_), .A2(new_n7430_), .ZN(new_n8025_));
  NAND2_X1   g07019(.A1(new_n8022_), .A2(new_n8025_), .ZN(new_n8026_));
  NOR2_X1    g07020(.A1(new_n8026_), .A2(new_n8018_), .ZN(new_n8027_));
  NOR4_X1    g07021(.A1(new_n7428_), .A2(new_n8024_), .A3(new_n7465_), .A4(new_n8017_), .ZN(new_n8028_));
  NAND3_X1   g07022(.A1(new_n8027_), .A2(new_n8014_), .A3(new_n8028_), .ZN(new_n8029_));
  NOR3_X1    g07023(.A1(new_n7428_), .A2(new_n8024_), .A3(new_n7430_), .ZN(new_n8030_));
  NOR2_X1    g07024(.A1(new_n7464_), .A2(new_n7465_), .ZN(new_n8031_));
  NOR2_X1    g07025(.A1(new_n8030_), .A2(new_n8031_), .ZN(new_n8032_));
  NAND2_X1   g07026(.A1(new_n8032_), .A2(new_n8017_), .ZN(new_n8033_));
  INV_X1     g07027(.I(new_n8028_), .ZN(new_n8034_));
  OAI21_X1   g07028(.A1(new_n8033_), .A2(new_n8034_), .B(new_n8013_), .ZN(new_n8035_));
  NAND2_X1   g07029(.A1(new_n8035_), .A2(new_n8029_), .ZN(new_n8036_));
  NAND2_X1   g07030(.A1(new_n7464_), .A2(new_n7465_), .ZN(new_n8037_));
  NOR2_X1    g07031(.A1(new_n7470_), .A2(new_n7466_), .ZN(new_n8038_));
  NOR2_X1    g07032(.A1(new_n7458_), .A2(new_n7432_), .ZN(new_n8039_));
  OAI21_X1   g07033(.A1(new_n8039_), .A2(new_n8038_), .B(new_n8037_), .ZN(new_n8040_));
  INV_X1     g07034(.I(new_n7473_), .ZN(new_n8041_));
  NAND2_X1   g07035(.A1(new_n8040_), .A2(new_n8041_), .ZN(new_n8042_));
  OAI21_X1   g07036(.A1(new_n7410_), .A2(new_n8042_), .B(new_n7405_), .ZN(new_n8043_));
  NOR3_X1    g07037(.A1(new_n7340_), .A2(new_n7375_), .A3(new_n7378_), .ZN(new_n8044_));
  INV_X1     g07038(.I(new_n7370_), .ZN(new_n8045_));
  OAI21_X1   g07039(.A1(new_n7338_), .A2(new_n7337_), .B(new_n7336_), .ZN(new_n8046_));
  NAND3_X1   g07040(.A1(new_n7322_), .A2(new_n7329_), .A3(new_n6979_), .ZN(new_n8047_));
  NAND2_X1   g07041(.A1(new_n8046_), .A2(new_n8047_), .ZN(new_n8048_));
  AOI22_X1   g07042(.A1(new_n7341_), .A2(new_n7348_), .B1(new_n7356_), .B2(new_n7358_), .ZN(new_n8049_));
  AOI21_X1   g07043(.A1(new_n8049_), .A2(new_n7362_), .B(new_n8048_), .ZN(new_n8050_));
  NAND3_X1   g07044(.A1(new_n6968_), .A2(new_n6979_), .A3(new_n7376_), .ZN(new_n8051_));
  NAND2_X1   g07045(.A1(new_n8051_), .A2(new_n7328_), .ZN(new_n8052_));
  OR4_X2     g07046(.A1(new_n6992_), .A2(new_n7008_), .A3(new_n7009_), .A4(new_n7005_), .Z(new_n8053_));
  NAND3_X1   g07047(.A1(new_n6996_), .A2(new_n7007_), .A3(new_n8053_), .ZN(new_n8054_));
  NAND2_X1   g07048(.A1(new_n8054_), .A2(new_n7010_), .ZN(new_n8055_));
  NAND2_X1   g07049(.A1(new_n8052_), .A2(new_n8055_), .ZN(new_n8056_));
  INV_X1     g07050(.I(new_n8056_), .ZN(new_n8057_));
  OAI21_X1   g07051(.A1(new_n8050_), .A2(new_n8045_), .B(new_n8057_), .ZN(new_n8058_));
  NAND2_X1   g07052(.A1(new_n7363_), .A2(new_n7340_), .ZN(new_n8059_));
  NAND3_X1   g07053(.A1(new_n8059_), .A2(new_n7370_), .A3(new_n8056_), .ZN(new_n8060_));
  AOI21_X1   g07054(.A1(new_n8060_), .A2(new_n8058_), .B(new_n8044_), .ZN(new_n8061_));
  INV_X1     g07055(.I(new_n8044_), .ZN(new_n8062_));
  AOI21_X1   g07056(.A1(new_n8059_), .A2(new_n7370_), .B(new_n8056_), .ZN(new_n8063_));
  NOR3_X1    g07057(.A1(new_n8050_), .A2(new_n8057_), .A3(new_n8045_), .ZN(new_n8064_));
  NOR3_X1    g07058(.A1(new_n8063_), .A2(new_n8064_), .A3(new_n8062_), .ZN(new_n8065_));
  NAND3_X1   g07059(.A1(new_n7310_), .A2(new_n7314_), .A3(new_n7396_), .ZN(new_n8066_));
  INV_X1     g07060(.I(new_n8066_), .ZN(new_n8067_));
  AOI21_X1   g07061(.A1(new_n7310_), .A2(new_n7291_), .B(new_n7314_), .ZN(new_n8068_));
  NOR4_X1    g07062(.A1(new_n6952_), .A2(new_n6953_), .A3(new_n6936_), .A4(new_n6949_), .ZN(new_n8069_));
  OR3_X2     g07063(.A1(new_n6940_), .A2(new_n7265_), .A3(new_n8069_), .Z(new_n8070_));
  AOI22_X1   g07064(.A1(new_n8070_), .A2(new_n6954_), .B1(new_n7395_), .B2(new_n6927_), .ZN(new_n8071_));
  OAI21_X1   g07065(.A1(new_n8068_), .A2(new_n7269_), .B(new_n8071_), .ZN(new_n8072_));
  OAI21_X1   g07066(.A1(new_n7288_), .A2(new_n7292_), .B(new_n7304_), .ZN(new_n8073_));
  NAND2_X1   g07067(.A1(new_n7395_), .A2(new_n6927_), .ZN(new_n8074_));
  NAND2_X1   g07068(.A1(new_n8070_), .A2(new_n6954_), .ZN(new_n8075_));
  NAND2_X1   g07069(.A1(new_n8075_), .A2(new_n8074_), .ZN(new_n8076_));
  NAND3_X1   g07070(.A1(new_n8073_), .A2(new_n7394_), .A3(new_n8076_), .ZN(new_n8077_));
  AOI21_X1   g07071(.A1(new_n8077_), .A2(new_n8072_), .B(new_n8067_), .ZN(new_n8078_));
  AOI21_X1   g07072(.A1(new_n8073_), .A2(new_n7394_), .B(new_n8076_), .ZN(new_n8079_));
  NOR3_X1    g07073(.A1(new_n8068_), .A2(new_n7269_), .A3(new_n8071_), .ZN(new_n8080_));
  NOR3_X1    g07074(.A1(new_n8079_), .A2(new_n8080_), .A3(new_n8066_), .ZN(new_n8081_));
  OAI22_X1   g07075(.A1(new_n8061_), .A2(new_n8065_), .B1(new_n8078_), .B2(new_n8081_), .ZN(new_n8082_));
  OAI21_X1   g07076(.A1(new_n8063_), .A2(new_n8064_), .B(new_n8062_), .ZN(new_n8083_));
  NAND3_X1   g07077(.A1(new_n8060_), .A2(new_n8058_), .A3(new_n8044_), .ZN(new_n8084_));
  OAI21_X1   g07078(.A1(new_n8079_), .A2(new_n8080_), .B(new_n8066_), .ZN(new_n8085_));
  NAND3_X1   g07079(.A1(new_n8077_), .A2(new_n8072_), .A3(new_n8067_), .ZN(new_n8086_));
  NAND4_X1   g07080(.A1(new_n8083_), .A2(new_n8084_), .A3(new_n8085_), .A4(new_n8086_), .ZN(new_n8087_));
  NAND2_X1   g07081(.A1(new_n8082_), .A2(new_n8087_), .ZN(new_n8088_));
  NAND2_X1   g07082(.A1(new_n8043_), .A2(new_n8088_), .ZN(new_n8089_));
  AOI21_X1   g07083(.A1(new_n7411_), .A2(new_n7474_), .B(new_n7484_), .ZN(new_n8090_));
  AOI22_X1   g07084(.A1(new_n8083_), .A2(new_n8084_), .B1(new_n8085_), .B2(new_n8086_), .ZN(new_n8091_));
  NOR4_X1    g07085(.A1(new_n8061_), .A2(new_n8065_), .A3(new_n8078_), .A4(new_n8081_), .ZN(new_n8092_));
  NOR2_X1    g07086(.A1(new_n8092_), .A2(new_n8091_), .ZN(new_n8093_));
  NAND2_X1   g07087(.A1(new_n8090_), .A2(new_n8093_), .ZN(new_n8094_));
  AOI21_X1   g07088(.A1(new_n8094_), .A2(new_n8089_), .B(new_n8036_), .ZN(new_n8095_));
  NOR3_X1    g07089(.A1(new_n8033_), .A2(new_n8013_), .A3(new_n8034_), .ZN(new_n8096_));
  AOI21_X1   g07090(.A1(new_n8027_), .A2(new_n8028_), .B(new_n8014_), .ZN(new_n8097_));
  NOR2_X1    g07091(.A1(new_n8097_), .A2(new_n8096_), .ZN(new_n8098_));
  NOR2_X1    g07092(.A1(new_n8090_), .A2(new_n8093_), .ZN(new_n8099_));
  NOR2_X1    g07093(.A1(new_n8043_), .A2(new_n8088_), .ZN(new_n8100_));
  NOR3_X1    g07094(.A1(new_n8099_), .A2(new_n8100_), .A3(new_n8098_), .ZN(new_n8101_));
  OAI21_X1   g07095(.A1(new_n8095_), .A2(new_n8101_), .B(new_n8012_), .ZN(new_n8102_));
  INV_X1     g07096(.I(new_n8012_), .ZN(new_n8103_));
  OAI21_X1   g07097(.A1(new_n8099_), .A2(new_n8100_), .B(new_n8098_), .ZN(new_n8104_));
  NAND3_X1   g07098(.A1(new_n8094_), .A2(new_n8089_), .A3(new_n8036_), .ZN(new_n8105_));
  NAND3_X1   g07099(.A1(new_n8104_), .A2(new_n8105_), .A3(new_n8103_), .ZN(new_n8106_));
  NAND2_X1   g07100(.A1(new_n8102_), .A2(new_n8106_), .ZN(new_n8107_));
  NAND3_X1   g07101(.A1(new_n8107_), .A2(new_n8001_), .A3(new_n8009_), .ZN(new_n8108_));
  NAND2_X1   g07102(.A1(new_n8001_), .A2(new_n8009_), .ZN(new_n8109_));
  AOI21_X1   g07103(.A1(new_n8104_), .A2(new_n8105_), .B(new_n8103_), .ZN(new_n8110_));
  NOR3_X1    g07104(.A1(new_n8095_), .A2(new_n8101_), .A3(new_n8012_), .ZN(new_n8111_));
  NOR2_X1    g07105(.A1(new_n8111_), .A2(new_n8110_), .ZN(new_n8112_));
  NAND2_X1   g07106(.A1(new_n8109_), .A2(new_n8112_), .ZN(new_n8113_));
  AOI21_X1   g07107(.A1(new_n8113_), .A2(new_n8108_), .B(new_n7857_), .ZN(new_n8114_));
  INV_X1     g07108(.I(new_n7857_), .ZN(new_n8115_));
  NAND3_X1   g07109(.A1(new_n7999_), .A2(new_n7991_), .A3(new_n7992_), .ZN(new_n8116_));
  OAI21_X1   g07110(.A1(new_n7910_), .A2(new_n7918_), .B(new_n7989_), .ZN(new_n8117_));
  AOI21_X1   g07111(.A1(new_n8117_), .A2(new_n8116_), .B(new_n8006_), .ZN(new_n8118_));
  OAI22_X1   g07112(.A1(new_n7918_), .A2(new_n7910_), .B1(new_n7983_), .B2(new_n7988_), .ZN(new_n8119_));
  NAND4_X1   g07113(.A1(new_n7991_), .A2(new_n7992_), .A3(new_n7995_), .A4(new_n7998_), .ZN(new_n8120_));
  AOI21_X1   g07114(.A1(new_n8119_), .A2(new_n8120_), .B(new_n7860_), .ZN(new_n8121_));
  OAI22_X1   g07115(.A1(new_n8118_), .A2(new_n8121_), .B1(new_n8110_), .B2(new_n8111_), .ZN(new_n8122_));
  NAND4_X1   g07116(.A1(new_n8001_), .A2(new_n8009_), .A3(new_n8102_), .A4(new_n8106_), .ZN(new_n8123_));
  AOI21_X1   g07117(.A1(new_n8122_), .A2(new_n8123_), .B(new_n8115_), .ZN(new_n8124_));
  OAI21_X1   g07118(.A1(new_n8114_), .A2(new_n8124_), .B(new_n6903_), .ZN(new_n8125_));
  NOR3_X1    g07119(.A1(new_n8112_), .A2(new_n8118_), .A3(new_n8121_), .ZN(new_n8126_));
  AOI21_X1   g07120(.A1(new_n8001_), .A2(new_n8009_), .B(new_n8107_), .ZN(new_n8127_));
  OAI21_X1   g07121(.A1(new_n8127_), .A2(new_n8126_), .B(new_n8115_), .ZN(new_n8128_));
  AOI22_X1   g07122(.A1(new_n8001_), .A2(new_n8009_), .B1(new_n8102_), .B2(new_n8106_), .ZN(new_n8129_));
  NOR4_X1    g07123(.A1(new_n8118_), .A2(new_n8121_), .A3(new_n8110_), .A4(new_n8111_), .ZN(new_n8130_));
  OAI21_X1   g07124(.A1(new_n8129_), .A2(new_n8130_), .B(new_n7857_), .ZN(new_n8131_));
  NAND3_X1   g07125(.A1(new_n8128_), .A2(new_n6902_), .A3(new_n8131_), .ZN(new_n8132_));
  NAND2_X1   g07126(.A1(new_n8125_), .A2(new_n8132_), .ZN(new_n8133_));
  OAI21_X1   g07127(.A1(new_n5910_), .A2(new_n5912_), .B(new_n5797_), .ZN(new_n8134_));
  XNOR2_X1   g07128(.A1(new_n5795_), .A2(new_n5577_), .ZN(new_n8135_));
  INV_X1     g07129(.I(new_n6458_), .ZN(new_n8136_));
  OAI21_X1   g07130(.A1(new_n8136_), .A2(new_n6456_), .B(new_n6676_), .ZN(new_n8137_));
  INV_X1     g07131(.I(new_n6600_), .ZN(new_n8138_));
  AOI21_X1   g07132(.A1(new_n6460_), .A2(new_n8137_), .B(new_n8138_), .ZN(new_n8139_));
  NOR2_X1    g07133(.A1(new_n6601_), .A2(new_n8139_), .ZN(new_n8140_));
  NAND2_X1   g07134(.A1(new_n8140_), .A2(new_n7250_), .ZN(new_n8141_));
  INV_X1     g07135(.I(new_n7250_), .ZN(new_n8142_));
  NAND3_X1   g07136(.A1(new_n6460_), .A2(new_n8137_), .A3(new_n8138_), .ZN(new_n8143_));
  OAI21_X1   g07137(.A1(new_n6461_), .A2(new_n6459_), .B(new_n6600_), .ZN(new_n8144_));
  NAND2_X1   g07138(.A1(new_n8144_), .A2(new_n8143_), .ZN(new_n8145_));
  NAND2_X1   g07139(.A1(new_n8142_), .A2(new_n8145_), .ZN(new_n8146_));
  AOI21_X1   g07140(.A1(new_n8146_), .A2(new_n8141_), .B(new_n7083_), .ZN(new_n8147_));
  NOR2_X1    g07141(.A1(new_n7082_), .A2(new_n6957_), .ZN(new_n8148_));
  AOI21_X1   g07142(.A1(new_n6957_), .A2(new_n7080_), .B(new_n8148_), .ZN(new_n8149_));
  NOR2_X1    g07143(.A1(new_n8142_), .A2(new_n8145_), .ZN(new_n8150_));
  NOR2_X1    g07144(.A1(new_n8140_), .A2(new_n7250_), .ZN(new_n8151_));
  NOR3_X1    g07145(.A1(new_n8150_), .A2(new_n8151_), .A3(new_n8149_), .ZN(new_n8152_));
  OAI21_X1   g07146(.A1(new_n8152_), .A2(new_n8147_), .B(new_n8135_), .ZN(new_n8153_));
  NOR2_X1    g07147(.A1(new_n8153_), .A2(new_n8134_), .ZN(new_n8154_));
  NAND3_X1   g07148(.A1(new_n7486_), .A2(new_n7597_), .A3(new_n7854_), .ZN(new_n8155_));
  NAND2_X1   g07149(.A1(new_n8142_), .A2(new_n7083_), .ZN(new_n8156_));
  NAND2_X1   g07150(.A1(new_n8149_), .A2(new_n7250_), .ZN(new_n8157_));
  AOI21_X1   g07151(.A1(new_n8156_), .A2(new_n8157_), .B(new_n8145_), .ZN(new_n8158_));
  INV_X1     g07152(.I(new_n6686_), .ZN(new_n8159_));
  NAND3_X1   g07153(.A1(new_n8159_), .A2(new_n6787_), .A3(new_n6601_), .ZN(new_n8160_));
  NAND3_X1   g07154(.A1(new_n6787_), .A2(new_n6686_), .A3(new_n6601_), .ZN(new_n8161_));
  NAND2_X1   g07155(.A1(new_n8160_), .A2(new_n8161_), .ZN(new_n8162_));
  NAND2_X1   g07156(.A1(new_n8162_), .A2(new_n8158_), .ZN(new_n8163_));
  INV_X1     g07157(.I(new_n8163_), .ZN(new_n8164_));
  AOI21_X1   g07158(.A1(new_n6013_), .A2(new_n6014_), .B(new_n5796_), .ZN(new_n8165_));
  OAI21_X1   g07159(.A1(new_n8150_), .A2(new_n8151_), .B(new_n8149_), .ZN(new_n8166_));
  NAND3_X1   g07160(.A1(new_n8146_), .A2(new_n8141_), .A3(new_n7083_), .ZN(new_n8167_));
  NAND2_X1   g07161(.A1(new_n8166_), .A2(new_n8167_), .ZN(new_n8168_));
  AOI21_X1   g07162(.A1(new_n8168_), .A2(new_n8135_), .B(new_n8165_), .ZN(new_n8169_));
  NOR3_X1    g07163(.A1(new_n8169_), .A2(new_n8155_), .A3(new_n8164_), .ZN(new_n8170_));
  NOR2_X1    g07164(.A1(new_n8162_), .A2(new_n8158_), .ZN(new_n8171_));
  NOR2_X1    g07165(.A1(new_n8155_), .A2(new_n8171_), .ZN(new_n8172_));
  NOR2_X1    g07166(.A1(new_n8172_), .A2(new_n8164_), .ZN(new_n8173_));
  NOR3_X1    g07167(.A1(new_n8170_), .A2(new_n8173_), .A3(new_n8154_), .ZN(new_n8174_));
  INV_X1     g07168(.I(new_n8154_), .ZN(new_n8175_));
  INV_X1     g07169(.I(new_n8155_), .ZN(new_n8176_));
  NAND2_X1   g07170(.A1(new_n8153_), .A2(new_n8134_), .ZN(new_n8177_));
  NAND3_X1   g07171(.A1(new_n8177_), .A2(new_n8176_), .A3(new_n8163_), .ZN(new_n8178_));
  OAI21_X1   g07172(.A1(new_n8155_), .A2(new_n8171_), .B(new_n8163_), .ZN(new_n8179_));
  AOI21_X1   g07173(.A1(new_n8178_), .A2(new_n8175_), .B(new_n8179_), .ZN(new_n8180_));
  NOR2_X1    g07174(.A1(new_n8174_), .A2(new_n8180_), .ZN(new_n8181_));
  NOR2_X1    g07175(.A1(new_n8133_), .A2(new_n8181_), .ZN(new_n8182_));
  NAND3_X1   g07176(.A1(new_n8178_), .A2(new_n8175_), .A3(new_n8179_), .ZN(new_n8183_));
  OAI21_X1   g07177(.A1(new_n8170_), .A2(new_n8154_), .B(new_n8173_), .ZN(new_n8184_));
  NAND2_X1   g07178(.A1(new_n8184_), .A2(new_n8183_), .ZN(new_n8185_));
  AOI21_X1   g07179(.A1(new_n8125_), .A2(new_n8132_), .B(new_n8185_), .ZN(new_n8186_));
  OAI21_X1   g07180(.A1(new_n8182_), .A2(new_n8186_), .B(new_n6273_), .ZN(new_n8187_));
  NOR2_X1    g07181(.A1(new_n6267_), .A2(new_n6260_), .ZN(new_n8188_));
  NOR2_X1    g07182(.A1(new_n6253_), .A2(new_n6125_), .ZN(new_n8189_));
  OAI21_X1   g07183(.A1(new_n8189_), .A2(new_n8188_), .B(new_n6017_), .ZN(new_n8190_));
  NOR2_X1    g07184(.A1(new_n6267_), .A2(new_n6125_), .ZN(new_n8191_));
  NOR2_X1    g07185(.A1(new_n6253_), .A2(new_n6260_), .ZN(new_n8192_));
  OAI21_X1   g07186(.A1(new_n8191_), .A2(new_n8192_), .B(new_n6018_), .ZN(new_n8193_));
  NAND2_X1   g07187(.A1(new_n8190_), .A2(new_n8193_), .ZN(new_n8194_));
  NAND3_X1   g07188(.A1(new_n8185_), .A2(new_n8125_), .A3(new_n8132_), .ZN(new_n8195_));
  NAND2_X1   g07189(.A1(new_n8133_), .A2(new_n8181_), .ZN(new_n8196_));
  NAND3_X1   g07190(.A1(new_n8196_), .A2(new_n8195_), .A3(new_n8194_), .ZN(new_n8197_));
  NAND2_X1   g07191(.A1(new_n8187_), .A2(new_n8197_), .ZN(new_n8198_));
  NAND3_X1   g07192(.A1(new_n8168_), .A2(new_n8165_), .A3(new_n8135_), .ZN(new_n8199_));
  INV_X1     g07193(.I(\A[391] ), .ZN(new_n8200_));
  INV_X1     g07194(.I(\A[392] ), .ZN(new_n8201_));
  NAND2_X1   g07195(.A1(new_n8201_), .A2(\A[393] ), .ZN(new_n8202_));
  INV_X1     g07196(.I(\A[393] ), .ZN(new_n8203_));
  NAND2_X1   g07197(.A1(new_n8203_), .A2(\A[392] ), .ZN(new_n8204_));
  AOI21_X1   g07198(.A1(new_n8202_), .A2(new_n8204_), .B(new_n8200_), .ZN(new_n8205_));
  NAND2_X1   g07199(.A1(\A[392] ), .A2(\A[393] ), .ZN(new_n8206_));
  NOR2_X1    g07200(.A1(\A[392] ), .A2(\A[393] ), .ZN(new_n8207_));
  INV_X1     g07201(.I(new_n8207_), .ZN(new_n8208_));
  AOI21_X1   g07202(.A1(new_n8208_), .A2(new_n8206_), .B(\A[391] ), .ZN(new_n8209_));
  NOR2_X1    g07203(.A1(new_n8209_), .A2(new_n8205_), .ZN(new_n8210_));
  INV_X1     g07204(.I(\A[394] ), .ZN(new_n8211_));
  INV_X1     g07205(.I(\A[395] ), .ZN(new_n8212_));
  NAND2_X1   g07206(.A1(new_n8212_), .A2(\A[396] ), .ZN(new_n8213_));
  INV_X1     g07207(.I(\A[396] ), .ZN(new_n8214_));
  NAND2_X1   g07208(.A1(new_n8214_), .A2(\A[395] ), .ZN(new_n8215_));
  AOI21_X1   g07209(.A1(new_n8213_), .A2(new_n8215_), .B(new_n8211_), .ZN(new_n8216_));
  NAND2_X1   g07210(.A1(\A[395] ), .A2(\A[396] ), .ZN(new_n8217_));
  NOR2_X1    g07211(.A1(\A[395] ), .A2(\A[396] ), .ZN(new_n8218_));
  INV_X1     g07212(.I(new_n8218_), .ZN(new_n8219_));
  AOI21_X1   g07213(.A1(new_n8219_), .A2(new_n8217_), .B(\A[394] ), .ZN(new_n8220_));
  NOR2_X1    g07214(.A1(new_n8220_), .A2(new_n8216_), .ZN(new_n8221_));
  NOR2_X1    g07215(.A1(new_n8210_), .A2(new_n8221_), .ZN(new_n8222_));
  NOR4_X1    g07216(.A1(new_n8205_), .A2(new_n8209_), .A3(new_n8220_), .A4(new_n8216_), .ZN(new_n8223_));
  NOR2_X1    g07217(.A1(new_n8222_), .A2(new_n8223_), .ZN(new_n8224_));
  NOR2_X1    g07218(.A1(new_n8214_), .A2(\A[395] ), .ZN(new_n8225_));
  NOR2_X1    g07219(.A1(new_n8212_), .A2(\A[396] ), .ZN(new_n8226_));
  OAI21_X1   g07220(.A1(new_n8225_), .A2(new_n8226_), .B(\A[394] ), .ZN(new_n8227_));
  INV_X1     g07221(.I(new_n8217_), .ZN(new_n8228_));
  OAI21_X1   g07222(.A1(new_n8228_), .A2(new_n8218_), .B(new_n8211_), .ZN(new_n8229_));
  NAND2_X1   g07223(.A1(new_n8227_), .A2(new_n8229_), .ZN(new_n8230_));
  AOI21_X1   g07224(.A1(\A[395] ), .A2(\A[396] ), .B(\A[394] ), .ZN(new_n8231_));
  NOR2_X1    g07225(.A1(new_n8231_), .A2(new_n8218_), .ZN(new_n8232_));
  NOR4_X1    g07226(.A1(new_n8232_), .A2(\A[391] ), .A3(\A[392] ), .A4(\A[393] ), .ZN(new_n8233_));
  NAND2_X1   g07227(.A1(new_n8230_), .A2(new_n8233_), .ZN(new_n8234_));
  NAND2_X1   g07228(.A1(new_n8224_), .A2(new_n8234_), .ZN(new_n8235_));
  INV_X1     g07229(.I(\A[399] ), .ZN(new_n8236_));
  NOR2_X1    g07230(.A1(new_n8236_), .A2(\A[398] ), .ZN(new_n8237_));
  INV_X1     g07231(.I(\A[398] ), .ZN(new_n8238_));
  NOR2_X1    g07232(.A1(new_n8238_), .A2(\A[399] ), .ZN(new_n8239_));
  OAI21_X1   g07233(.A1(new_n8237_), .A2(new_n8239_), .B(\A[397] ), .ZN(new_n8240_));
  INV_X1     g07234(.I(\A[397] ), .ZN(new_n8241_));
  NOR2_X1    g07235(.A1(\A[398] ), .A2(\A[399] ), .ZN(new_n8242_));
  NAND2_X1   g07236(.A1(\A[398] ), .A2(\A[399] ), .ZN(new_n8243_));
  INV_X1     g07237(.I(new_n8243_), .ZN(new_n8244_));
  OAI21_X1   g07238(.A1(new_n8244_), .A2(new_n8242_), .B(new_n8241_), .ZN(new_n8245_));
  INV_X1     g07239(.I(\A[402] ), .ZN(new_n8246_));
  NOR2_X1    g07240(.A1(new_n8246_), .A2(\A[401] ), .ZN(new_n8247_));
  INV_X1     g07241(.I(\A[401] ), .ZN(new_n8248_));
  NOR2_X1    g07242(.A1(new_n8248_), .A2(\A[402] ), .ZN(new_n8249_));
  OAI21_X1   g07243(.A1(new_n8247_), .A2(new_n8249_), .B(\A[400] ), .ZN(new_n8250_));
  INV_X1     g07244(.I(\A[400] ), .ZN(new_n8251_));
  NOR2_X1    g07245(.A1(\A[401] ), .A2(\A[402] ), .ZN(new_n8252_));
  NAND2_X1   g07246(.A1(\A[401] ), .A2(\A[402] ), .ZN(new_n8253_));
  INV_X1     g07247(.I(new_n8253_), .ZN(new_n8254_));
  OAI21_X1   g07248(.A1(new_n8254_), .A2(new_n8252_), .B(new_n8251_), .ZN(new_n8255_));
  NAND4_X1   g07249(.A1(new_n8240_), .A2(new_n8245_), .A3(new_n8250_), .A4(new_n8255_), .ZN(new_n8256_));
  AOI21_X1   g07250(.A1(\A[401] ), .A2(\A[402] ), .B(\A[400] ), .ZN(new_n8257_));
  NOR2_X1    g07251(.A1(new_n8257_), .A2(new_n8252_), .ZN(new_n8258_));
  AOI21_X1   g07252(.A1(\A[398] ), .A2(\A[399] ), .B(\A[397] ), .ZN(new_n8259_));
  NOR2_X1    g07253(.A1(new_n8259_), .A2(new_n8242_), .ZN(new_n8260_));
  NAND2_X1   g07254(.A1(new_n8258_), .A2(new_n8260_), .ZN(new_n8261_));
  NOR2_X1    g07255(.A1(new_n8256_), .A2(new_n8261_), .ZN(new_n8262_));
  NAND2_X1   g07256(.A1(new_n8238_), .A2(\A[399] ), .ZN(new_n8263_));
  NAND2_X1   g07257(.A1(new_n8236_), .A2(\A[398] ), .ZN(new_n8264_));
  AOI21_X1   g07258(.A1(new_n8263_), .A2(new_n8264_), .B(new_n8241_), .ZN(new_n8265_));
  INV_X1     g07259(.I(new_n8242_), .ZN(new_n8266_));
  AOI21_X1   g07260(.A1(new_n8266_), .A2(new_n8243_), .B(\A[397] ), .ZN(new_n8267_));
  NAND2_X1   g07261(.A1(new_n8248_), .A2(\A[402] ), .ZN(new_n8268_));
  NAND2_X1   g07262(.A1(new_n8246_), .A2(\A[401] ), .ZN(new_n8269_));
  AOI21_X1   g07263(.A1(new_n8268_), .A2(new_n8269_), .B(new_n8251_), .ZN(new_n8270_));
  INV_X1     g07264(.I(new_n8252_), .ZN(new_n8271_));
  AOI21_X1   g07265(.A1(new_n8271_), .A2(new_n8253_), .B(\A[400] ), .ZN(new_n8272_));
  OAI22_X1   g07266(.A1(new_n8265_), .A2(new_n8267_), .B1(new_n8272_), .B2(new_n8270_), .ZN(new_n8273_));
  NAND2_X1   g07267(.A1(new_n8273_), .A2(new_n8256_), .ZN(new_n8274_));
  NOR2_X1    g07268(.A1(new_n8274_), .A2(new_n8262_), .ZN(new_n8275_));
  INV_X1     g07269(.I(\A[409] ), .ZN(new_n8276_));
  INV_X1     g07270(.I(\A[410] ), .ZN(new_n8277_));
  NAND2_X1   g07271(.A1(new_n8277_), .A2(\A[411] ), .ZN(new_n8278_));
  INV_X1     g07272(.I(\A[411] ), .ZN(new_n8279_));
  NAND2_X1   g07273(.A1(new_n8279_), .A2(\A[410] ), .ZN(new_n8280_));
  AOI21_X1   g07274(.A1(new_n8278_), .A2(new_n8280_), .B(new_n8276_), .ZN(new_n8281_));
  NOR2_X1    g07275(.A1(\A[410] ), .A2(\A[411] ), .ZN(new_n8282_));
  INV_X1     g07276(.I(new_n8282_), .ZN(new_n8283_));
  NAND2_X1   g07277(.A1(\A[410] ), .A2(\A[411] ), .ZN(new_n8284_));
  AOI21_X1   g07278(.A1(new_n8283_), .A2(new_n8284_), .B(\A[409] ), .ZN(new_n8285_));
  INV_X1     g07279(.I(\A[412] ), .ZN(new_n8286_));
  INV_X1     g07280(.I(\A[413] ), .ZN(new_n8287_));
  NAND2_X1   g07281(.A1(new_n8287_), .A2(\A[414] ), .ZN(new_n8288_));
  INV_X1     g07282(.I(\A[414] ), .ZN(new_n8289_));
  NAND2_X1   g07283(.A1(new_n8289_), .A2(\A[413] ), .ZN(new_n8290_));
  AOI21_X1   g07284(.A1(new_n8288_), .A2(new_n8290_), .B(new_n8286_), .ZN(new_n8291_));
  NOR2_X1    g07285(.A1(\A[413] ), .A2(\A[414] ), .ZN(new_n8292_));
  INV_X1     g07286(.I(new_n8292_), .ZN(new_n8293_));
  NAND2_X1   g07287(.A1(\A[413] ), .A2(\A[414] ), .ZN(new_n8294_));
  AOI21_X1   g07288(.A1(new_n8293_), .A2(new_n8294_), .B(\A[412] ), .ZN(new_n8295_));
  NOR4_X1    g07289(.A1(new_n8281_), .A2(new_n8285_), .A3(new_n8295_), .A4(new_n8291_), .ZN(new_n8296_));
  AOI21_X1   g07290(.A1(\A[413] ), .A2(\A[414] ), .B(\A[412] ), .ZN(new_n8297_));
  NOR2_X1    g07291(.A1(new_n8297_), .A2(new_n8292_), .ZN(new_n8298_));
  AOI21_X1   g07292(.A1(\A[410] ), .A2(\A[411] ), .B(\A[409] ), .ZN(new_n8299_));
  NOR2_X1    g07293(.A1(new_n8299_), .A2(new_n8282_), .ZN(new_n8300_));
  NAND2_X1   g07294(.A1(new_n8298_), .A2(new_n8300_), .ZN(new_n8301_));
  INV_X1     g07295(.I(new_n8301_), .ZN(new_n8302_));
  NAND2_X1   g07296(.A1(new_n8296_), .A2(new_n8302_), .ZN(new_n8303_));
  NOR2_X1    g07297(.A1(new_n8279_), .A2(\A[410] ), .ZN(new_n8304_));
  NOR2_X1    g07298(.A1(new_n8277_), .A2(\A[411] ), .ZN(new_n8305_));
  OAI21_X1   g07299(.A1(new_n8304_), .A2(new_n8305_), .B(\A[409] ), .ZN(new_n8306_));
  INV_X1     g07300(.I(new_n8284_), .ZN(new_n8307_));
  OAI21_X1   g07301(.A1(new_n8307_), .A2(new_n8282_), .B(new_n8276_), .ZN(new_n8308_));
  NOR2_X1    g07302(.A1(new_n8289_), .A2(\A[413] ), .ZN(new_n8309_));
  NOR2_X1    g07303(.A1(new_n8287_), .A2(\A[414] ), .ZN(new_n8310_));
  OAI21_X1   g07304(.A1(new_n8309_), .A2(new_n8310_), .B(\A[412] ), .ZN(new_n8311_));
  INV_X1     g07305(.I(new_n8294_), .ZN(new_n8312_));
  OAI21_X1   g07306(.A1(new_n8312_), .A2(new_n8292_), .B(new_n8286_), .ZN(new_n8313_));
  AOI22_X1   g07307(.A1(new_n8306_), .A2(new_n8308_), .B1(new_n8311_), .B2(new_n8313_), .ZN(new_n8314_));
  NOR2_X1    g07308(.A1(new_n8314_), .A2(new_n8296_), .ZN(new_n8315_));
  NAND2_X1   g07309(.A1(new_n8315_), .A2(new_n8303_), .ZN(new_n8316_));
  INV_X1     g07310(.I(\A[403] ), .ZN(new_n8317_));
  INV_X1     g07311(.I(\A[404] ), .ZN(new_n8318_));
  NAND2_X1   g07312(.A1(new_n8318_), .A2(\A[405] ), .ZN(new_n8319_));
  INV_X1     g07313(.I(\A[405] ), .ZN(new_n8320_));
  NAND2_X1   g07314(.A1(new_n8320_), .A2(\A[404] ), .ZN(new_n8321_));
  AOI21_X1   g07315(.A1(new_n8319_), .A2(new_n8321_), .B(new_n8317_), .ZN(new_n8322_));
  NAND2_X1   g07316(.A1(\A[404] ), .A2(\A[405] ), .ZN(new_n8323_));
  NOR2_X1    g07317(.A1(\A[404] ), .A2(\A[405] ), .ZN(new_n8324_));
  INV_X1     g07318(.I(new_n8324_), .ZN(new_n8325_));
  AOI21_X1   g07319(.A1(new_n8325_), .A2(new_n8323_), .B(\A[403] ), .ZN(new_n8326_));
  INV_X1     g07320(.I(\A[406] ), .ZN(new_n8327_));
  INV_X1     g07321(.I(\A[407] ), .ZN(new_n8328_));
  NAND2_X1   g07322(.A1(new_n8328_), .A2(\A[408] ), .ZN(new_n8329_));
  INV_X1     g07323(.I(\A[408] ), .ZN(new_n8330_));
  NAND2_X1   g07324(.A1(new_n8330_), .A2(\A[407] ), .ZN(new_n8331_));
  AOI21_X1   g07325(.A1(new_n8329_), .A2(new_n8331_), .B(new_n8327_), .ZN(new_n8332_));
  NAND2_X1   g07326(.A1(\A[407] ), .A2(\A[408] ), .ZN(new_n8333_));
  NOR2_X1    g07327(.A1(\A[407] ), .A2(\A[408] ), .ZN(new_n8334_));
  INV_X1     g07328(.I(new_n8334_), .ZN(new_n8335_));
  AOI21_X1   g07329(.A1(new_n8335_), .A2(new_n8333_), .B(\A[406] ), .ZN(new_n8336_));
  OAI22_X1   g07330(.A1(new_n8322_), .A2(new_n8326_), .B1(new_n8336_), .B2(new_n8332_), .ZN(new_n8337_));
  NOR2_X1    g07331(.A1(new_n8320_), .A2(\A[404] ), .ZN(new_n8338_));
  NOR2_X1    g07332(.A1(new_n8318_), .A2(\A[405] ), .ZN(new_n8339_));
  OAI21_X1   g07333(.A1(new_n8338_), .A2(new_n8339_), .B(\A[403] ), .ZN(new_n8340_));
  INV_X1     g07334(.I(new_n8323_), .ZN(new_n8341_));
  OAI21_X1   g07335(.A1(new_n8341_), .A2(new_n8324_), .B(new_n8317_), .ZN(new_n8342_));
  NOR2_X1    g07336(.A1(new_n8330_), .A2(\A[407] ), .ZN(new_n8343_));
  NOR2_X1    g07337(.A1(new_n8328_), .A2(\A[408] ), .ZN(new_n8344_));
  OAI21_X1   g07338(.A1(new_n8343_), .A2(new_n8344_), .B(\A[406] ), .ZN(new_n8345_));
  INV_X1     g07339(.I(new_n8333_), .ZN(new_n8346_));
  OAI21_X1   g07340(.A1(new_n8346_), .A2(new_n8334_), .B(new_n8327_), .ZN(new_n8347_));
  NAND4_X1   g07341(.A1(new_n8340_), .A2(new_n8342_), .A3(new_n8345_), .A4(new_n8347_), .ZN(new_n8348_));
  NAND2_X1   g07342(.A1(new_n8337_), .A2(new_n8348_), .ZN(new_n8349_));
  NOR2_X1    g07343(.A1(new_n8326_), .A2(new_n8322_), .ZN(new_n8350_));
  NOR2_X1    g07344(.A1(new_n8336_), .A2(new_n8332_), .ZN(new_n8351_));
  AOI21_X1   g07345(.A1(\A[404] ), .A2(\A[405] ), .B(\A[403] ), .ZN(new_n8352_));
  AOI21_X1   g07346(.A1(\A[407] ), .A2(\A[408] ), .B(\A[406] ), .ZN(new_n8353_));
  OAI22_X1   g07347(.A1(new_n8324_), .A2(new_n8352_), .B1(new_n8353_), .B2(new_n8334_), .ZN(new_n8354_));
  NOR3_X1    g07348(.A1(new_n8350_), .A2(new_n8351_), .A3(new_n8354_), .ZN(new_n8355_));
  NOR2_X1    g07349(.A1(new_n8349_), .A2(new_n8355_), .ZN(new_n8356_));
  NAND2_X1   g07350(.A1(new_n8316_), .A2(new_n8356_), .ZN(new_n8357_));
  NAND4_X1   g07351(.A1(new_n8306_), .A2(new_n8308_), .A3(new_n8311_), .A4(new_n8313_), .ZN(new_n8358_));
  NOR2_X1    g07352(.A1(new_n8358_), .A2(new_n8301_), .ZN(new_n8359_));
  OAI22_X1   g07353(.A1(new_n8281_), .A2(new_n8285_), .B1(new_n8295_), .B2(new_n8291_), .ZN(new_n8360_));
  NAND2_X1   g07354(.A1(new_n8360_), .A2(new_n8358_), .ZN(new_n8361_));
  NOR2_X1    g07355(.A1(new_n8361_), .A2(new_n8359_), .ZN(new_n8362_));
  AOI22_X1   g07356(.A1(new_n8340_), .A2(new_n8342_), .B1(new_n8345_), .B2(new_n8347_), .ZN(new_n8363_));
  NOR4_X1    g07357(.A1(new_n8322_), .A2(new_n8326_), .A3(new_n8336_), .A4(new_n8332_), .ZN(new_n8364_));
  NOR2_X1    g07358(.A1(new_n8363_), .A2(new_n8364_), .ZN(new_n8365_));
  NAND2_X1   g07359(.A1(new_n8340_), .A2(new_n8342_), .ZN(new_n8366_));
  NAND2_X1   g07360(.A1(new_n8345_), .A2(new_n8347_), .ZN(new_n8367_));
  NOR2_X1    g07361(.A1(new_n8352_), .A2(new_n8324_), .ZN(new_n8368_));
  NOR2_X1    g07362(.A1(new_n8353_), .A2(new_n8334_), .ZN(new_n8369_));
  NOR2_X1    g07363(.A1(new_n8368_), .A2(new_n8369_), .ZN(new_n8370_));
  NAND3_X1   g07364(.A1(new_n8366_), .A2(new_n8367_), .A3(new_n8370_), .ZN(new_n8371_));
  NAND2_X1   g07365(.A1(new_n8365_), .A2(new_n8371_), .ZN(new_n8372_));
  NAND2_X1   g07366(.A1(new_n8372_), .A2(new_n8362_), .ZN(new_n8373_));
  AOI21_X1   g07367(.A1(new_n8373_), .A2(new_n8357_), .B(new_n8275_), .ZN(new_n8374_));
  INV_X1     g07368(.I(new_n8374_), .ZN(new_n8375_));
  NAND3_X1   g07369(.A1(new_n8373_), .A2(new_n8357_), .A3(new_n8275_), .ZN(new_n8376_));
  NAND2_X1   g07370(.A1(new_n8375_), .A2(new_n8376_), .ZN(new_n8377_));
  NAND2_X1   g07371(.A1(new_n8377_), .A2(new_n8235_), .ZN(new_n8378_));
  OAI22_X1   g07372(.A1(new_n8205_), .A2(new_n8209_), .B1(new_n8220_), .B2(new_n8216_), .ZN(new_n8379_));
  NOR2_X1    g07373(.A1(new_n8203_), .A2(\A[392] ), .ZN(new_n8380_));
  NOR2_X1    g07374(.A1(new_n8201_), .A2(\A[393] ), .ZN(new_n8381_));
  OAI21_X1   g07375(.A1(new_n8380_), .A2(new_n8381_), .B(\A[391] ), .ZN(new_n8382_));
  INV_X1     g07376(.I(new_n8206_), .ZN(new_n8383_));
  OAI21_X1   g07377(.A1(new_n8383_), .A2(new_n8207_), .B(new_n8200_), .ZN(new_n8384_));
  NAND4_X1   g07378(.A1(new_n8382_), .A2(new_n8384_), .A3(new_n8227_), .A4(new_n8229_), .ZN(new_n8385_));
  NAND2_X1   g07379(.A1(new_n8379_), .A2(new_n8385_), .ZN(new_n8386_));
  AOI21_X1   g07380(.A1(\A[392] ), .A2(\A[393] ), .B(\A[391] ), .ZN(new_n8387_));
  OAI22_X1   g07381(.A1(new_n8207_), .A2(new_n8387_), .B1(new_n8231_), .B2(new_n8218_), .ZN(new_n8388_));
  NOR3_X1    g07382(.A1(new_n8210_), .A2(new_n8221_), .A3(new_n8388_), .ZN(new_n8389_));
  NOR2_X1    g07383(.A1(new_n8386_), .A2(new_n8389_), .ZN(new_n8390_));
  NAND3_X1   g07384(.A1(new_n8375_), .A2(new_n8390_), .A3(new_n8376_), .ZN(new_n8391_));
  INV_X1     g07385(.I(\A[385] ), .ZN(new_n8392_));
  INV_X1     g07386(.I(\A[386] ), .ZN(new_n8393_));
  NAND2_X1   g07387(.A1(new_n8393_), .A2(\A[387] ), .ZN(new_n8394_));
  INV_X1     g07388(.I(\A[387] ), .ZN(new_n8395_));
  NAND2_X1   g07389(.A1(new_n8395_), .A2(\A[386] ), .ZN(new_n8396_));
  AOI21_X1   g07390(.A1(new_n8394_), .A2(new_n8396_), .B(new_n8392_), .ZN(new_n8397_));
  NAND2_X1   g07391(.A1(\A[386] ), .A2(\A[387] ), .ZN(new_n8398_));
  NOR2_X1    g07392(.A1(\A[386] ), .A2(\A[387] ), .ZN(new_n8399_));
  INV_X1     g07393(.I(new_n8399_), .ZN(new_n8400_));
  AOI21_X1   g07394(.A1(new_n8400_), .A2(new_n8398_), .B(\A[385] ), .ZN(new_n8401_));
  NOR2_X1    g07395(.A1(new_n8401_), .A2(new_n8397_), .ZN(new_n8402_));
  INV_X1     g07396(.I(\A[388] ), .ZN(new_n8403_));
  INV_X1     g07397(.I(\A[389] ), .ZN(new_n8404_));
  NAND2_X1   g07398(.A1(new_n8404_), .A2(\A[390] ), .ZN(new_n8405_));
  INV_X1     g07399(.I(\A[390] ), .ZN(new_n8406_));
  NAND2_X1   g07400(.A1(new_n8406_), .A2(\A[389] ), .ZN(new_n8407_));
  AOI21_X1   g07401(.A1(new_n8405_), .A2(new_n8407_), .B(new_n8403_), .ZN(new_n8408_));
  NAND2_X1   g07402(.A1(\A[389] ), .A2(\A[390] ), .ZN(new_n8409_));
  NOR2_X1    g07403(.A1(\A[389] ), .A2(\A[390] ), .ZN(new_n8410_));
  INV_X1     g07404(.I(new_n8410_), .ZN(new_n8411_));
  AOI21_X1   g07405(.A1(new_n8411_), .A2(new_n8409_), .B(\A[388] ), .ZN(new_n8412_));
  NOR2_X1    g07406(.A1(new_n8412_), .A2(new_n8408_), .ZN(new_n8413_));
  AOI21_X1   g07407(.A1(\A[386] ), .A2(\A[387] ), .B(\A[385] ), .ZN(new_n8414_));
  AOI21_X1   g07408(.A1(\A[389] ), .A2(\A[390] ), .B(\A[388] ), .ZN(new_n8415_));
  OAI22_X1   g07409(.A1(new_n8399_), .A2(new_n8414_), .B1(new_n8415_), .B2(new_n8410_), .ZN(new_n8416_));
  NOR3_X1    g07410(.A1(new_n8402_), .A2(new_n8413_), .A3(new_n8416_), .ZN(new_n8417_));
  INV_X1     g07411(.I(\A[381] ), .ZN(new_n8418_));
  NOR2_X1    g07412(.A1(new_n8418_), .A2(\A[380] ), .ZN(new_n8419_));
  INV_X1     g07413(.I(\A[380] ), .ZN(new_n8420_));
  NOR2_X1    g07414(.A1(new_n8420_), .A2(\A[381] ), .ZN(new_n8421_));
  OAI21_X1   g07415(.A1(new_n8419_), .A2(new_n8421_), .B(\A[379] ), .ZN(new_n8422_));
  INV_X1     g07416(.I(\A[379] ), .ZN(new_n8423_));
  NAND2_X1   g07417(.A1(\A[380] ), .A2(\A[381] ), .ZN(new_n8424_));
  INV_X1     g07418(.I(new_n8424_), .ZN(new_n8425_));
  NOR2_X1    g07419(.A1(\A[380] ), .A2(\A[381] ), .ZN(new_n8426_));
  OAI21_X1   g07420(.A1(new_n8425_), .A2(new_n8426_), .B(new_n8423_), .ZN(new_n8427_));
  NAND2_X1   g07421(.A1(new_n8422_), .A2(new_n8427_), .ZN(new_n8428_));
  INV_X1     g07422(.I(\A[384] ), .ZN(new_n8429_));
  NOR2_X1    g07423(.A1(new_n8429_), .A2(\A[383] ), .ZN(new_n8430_));
  INV_X1     g07424(.I(\A[383] ), .ZN(new_n8431_));
  NOR2_X1    g07425(.A1(new_n8431_), .A2(\A[384] ), .ZN(new_n8432_));
  OAI21_X1   g07426(.A1(new_n8430_), .A2(new_n8432_), .B(\A[382] ), .ZN(new_n8433_));
  INV_X1     g07427(.I(\A[382] ), .ZN(new_n8434_));
  NAND2_X1   g07428(.A1(\A[383] ), .A2(\A[384] ), .ZN(new_n8435_));
  INV_X1     g07429(.I(new_n8435_), .ZN(new_n8436_));
  NOR2_X1    g07430(.A1(\A[383] ), .A2(\A[384] ), .ZN(new_n8437_));
  OAI21_X1   g07431(.A1(new_n8436_), .A2(new_n8437_), .B(new_n8434_), .ZN(new_n8438_));
  NAND2_X1   g07432(.A1(new_n8433_), .A2(new_n8438_), .ZN(new_n8439_));
  AOI21_X1   g07433(.A1(\A[380] ), .A2(\A[381] ), .B(\A[379] ), .ZN(new_n8440_));
  AOI21_X1   g07434(.A1(\A[383] ), .A2(\A[384] ), .B(\A[382] ), .ZN(new_n8441_));
  OAI22_X1   g07435(.A1(new_n8426_), .A2(new_n8440_), .B1(new_n8441_), .B2(new_n8437_), .ZN(new_n8442_));
  INV_X1     g07436(.I(new_n8442_), .ZN(new_n8443_));
  NAND3_X1   g07437(.A1(new_n8428_), .A2(new_n8439_), .A3(new_n8443_), .ZN(new_n8444_));
  NOR2_X1    g07438(.A1(new_n8417_), .A2(new_n8444_), .ZN(new_n8445_));
  NOR2_X1    g07439(.A1(new_n8395_), .A2(\A[386] ), .ZN(new_n8446_));
  NOR2_X1    g07440(.A1(new_n8393_), .A2(\A[387] ), .ZN(new_n8447_));
  OAI21_X1   g07441(.A1(new_n8446_), .A2(new_n8447_), .B(\A[385] ), .ZN(new_n8448_));
  INV_X1     g07442(.I(new_n8398_), .ZN(new_n8449_));
  OAI21_X1   g07443(.A1(new_n8449_), .A2(new_n8399_), .B(new_n8392_), .ZN(new_n8450_));
  NAND2_X1   g07444(.A1(new_n8448_), .A2(new_n8450_), .ZN(new_n8451_));
  NOR2_X1    g07445(.A1(new_n8406_), .A2(\A[389] ), .ZN(new_n8452_));
  NOR2_X1    g07446(.A1(new_n8404_), .A2(\A[390] ), .ZN(new_n8453_));
  OAI21_X1   g07447(.A1(new_n8452_), .A2(new_n8453_), .B(\A[388] ), .ZN(new_n8454_));
  INV_X1     g07448(.I(new_n8409_), .ZN(new_n8455_));
  OAI21_X1   g07449(.A1(new_n8455_), .A2(new_n8410_), .B(new_n8403_), .ZN(new_n8456_));
  NAND2_X1   g07450(.A1(new_n8454_), .A2(new_n8456_), .ZN(new_n8457_));
  NOR2_X1    g07451(.A1(new_n8414_), .A2(new_n8399_), .ZN(new_n8458_));
  NOR2_X1    g07452(.A1(new_n8415_), .A2(new_n8410_), .ZN(new_n8459_));
  NOR2_X1    g07453(.A1(new_n8458_), .A2(new_n8459_), .ZN(new_n8460_));
  NAND3_X1   g07454(.A1(new_n8451_), .A2(new_n8457_), .A3(new_n8460_), .ZN(new_n8461_));
  NAND2_X1   g07455(.A1(new_n8420_), .A2(\A[381] ), .ZN(new_n8462_));
  NAND2_X1   g07456(.A1(new_n8418_), .A2(\A[380] ), .ZN(new_n8463_));
  AOI21_X1   g07457(.A1(new_n8462_), .A2(new_n8463_), .B(new_n8423_), .ZN(new_n8464_));
  INV_X1     g07458(.I(new_n8426_), .ZN(new_n8465_));
  AOI21_X1   g07459(.A1(new_n8465_), .A2(new_n8424_), .B(\A[379] ), .ZN(new_n8466_));
  NOR2_X1    g07460(.A1(new_n8466_), .A2(new_n8464_), .ZN(new_n8467_));
  NAND2_X1   g07461(.A1(new_n8431_), .A2(\A[384] ), .ZN(new_n8468_));
  NAND2_X1   g07462(.A1(new_n8429_), .A2(\A[383] ), .ZN(new_n8469_));
  AOI21_X1   g07463(.A1(new_n8468_), .A2(new_n8469_), .B(new_n8434_), .ZN(new_n8470_));
  INV_X1     g07464(.I(new_n8437_), .ZN(new_n8471_));
  AOI21_X1   g07465(.A1(new_n8471_), .A2(new_n8435_), .B(\A[382] ), .ZN(new_n8472_));
  NOR2_X1    g07466(.A1(new_n8472_), .A2(new_n8470_), .ZN(new_n8473_));
  NOR3_X1    g07467(.A1(new_n8467_), .A2(new_n8473_), .A3(new_n8442_), .ZN(new_n8474_));
  NOR2_X1    g07468(.A1(new_n8474_), .A2(new_n8461_), .ZN(new_n8475_));
  INV_X1     g07469(.I(\A[373] ), .ZN(new_n8476_));
  INV_X1     g07470(.I(\A[374] ), .ZN(new_n8477_));
  NAND2_X1   g07471(.A1(new_n8477_), .A2(\A[375] ), .ZN(new_n8478_));
  INV_X1     g07472(.I(\A[375] ), .ZN(new_n8479_));
  NAND2_X1   g07473(.A1(new_n8479_), .A2(\A[374] ), .ZN(new_n8480_));
  AOI21_X1   g07474(.A1(new_n8478_), .A2(new_n8480_), .B(new_n8476_), .ZN(new_n8481_));
  NAND2_X1   g07475(.A1(\A[374] ), .A2(\A[375] ), .ZN(new_n8482_));
  NOR2_X1    g07476(.A1(\A[374] ), .A2(\A[375] ), .ZN(new_n8483_));
  INV_X1     g07477(.I(new_n8483_), .ZN(new_n8484_));
  AOI21_X1   g07478(.A1(new_n8484_), .A2(new_n8482_), .B(\A[373] ), .ZN(new_n8485_));
  NOR2_X1    g07479(.A1(new_n8485_), .A2(new_n8481_), .ZN(new_n8486_));
  INV_X1     g07480(.I(\A[376] ), .ZN(new_n8487_));
  INV_X1     g07481(.I(\A[377] ), .ZN(new_n8488_));
  NAND2_X1   g07482(.A1(new_n8488_), .A2(\A[378] ), .ZN(new_n8489_));
  INV_X1     g07483(.I(\A[378] ), .ZN(new_n8490_));
  NAND2_X1   g07484(.A1(new_n8490_), .A2(\A[377] ), .ZN(new_n8491_));
  AOI21_X1   g07485(.A1(new_n8489_), .A2(new_n8491_), .B(new_n8487_), .ZN(new_n8492_));
  NAND2_X1   g07486(.A1(\A[377] ), .A2(\A[378] ), .ZN(new_n8493_));
  NOR2_X1    g07487(.A1(\A[377] ), .A2(\A[378] ), .ZN(new_n8494_));
  INV_X1     g07488(.I(new_n8494_), .ZN(new_n8495_));
  AOI21_X1   g07489(.A1(new_n8495_), .A2(new_n8493_), .B(\A[376] ), .ZN(new_n8496_));
  NOR2_X1    g07490(.A1(new_n8496_), .A2(new_n8492_), .ZN(new_n8497_));
  AOI21_X1   g07491(.A1(\A[374] ), .A2(\A[375] ), .B(\A[373] ), .ZN(new_n8498_));
  AOI21_X1   g07492(.A1(\A[377] ), .A2(\A[378] ), .B(\A[376] ), .ZN(new_n8499_));
  OAI22_X1   g07493(.A1(new_n8483_), .A2(new_n8498_), .B1(new_n8499_), .B2(new_n8494_), .ZN(new_n8500_));
  NOR3_X1    g07494(.A1(new_n8486_), .A2(new_n8497_), .A3(new_n8500_), .ZN(new_n8501_));
  INV_X1     g07495(.I(\A[369] ), .ZN(new_n8502_));
  NOR2_X1    g07496(.A1(new_n8502_), .A2(\A[368] ), .ZN(new_n8503_));
  INV_X1     g07497(.I(\A[368] ), .ZN(new_n8504_));
  NOR2_X1    g07498(.A1(new_n8504_), .A2(\A[369] ), .ZN(new_n8505_));
  OAI21_X1   g07499(.A1(new_n8503_), .A2(new_n8505_), .B(\A[367] ), .ZN(new_n8506_));
  INV_X1     g07500(.I(\A[367] ), .ZN(new_n8507_));
  NAND2_X1   g07501(.A1(\A[368] ), .A2(\A[369] ), .ZN(new_n8508_));
  INV_X1     g07502(.I(new_n8508_), .ZN(new_n8509_));
  NOR2_X1    g07503(.A1(\A[368] ), .A2(\A[369] ), .ZN(new_n8510_));
  OAI21_X1   g07504(.A1(new_n8509_), .A2(new_n8510_), .B(new_n8507_), .ZN(new_n8511_));
  NAND2_X1   g07505(.A1(new_n8506_), .A2(new_n8511_), .ZN(new_n8512_));
  INV_X1     g07506(.I(\A[372] ), .ZN(new_n8513_));
  NOR2_X1    g07507(.A1(new_n8513_), .A2(\A[371] ), .ZN(new_n8514_));
  INV_X1     g07508(.I(\A[371] ), .ZN(new_n8515_));
  NOR2_X1    g07509(.A1(new_n8515_), .A2(\A[372] ), .ZN(new_n8516_));
  OAI21_X1   g07510(.A1(new_n8514_), .A2(new_n8516_), .B(\A[370] ), .ZN(new_n8517_));
  INV_X1     g07511(.I(\A[370] ), .ZN(new_n8518_));
  NAND2_X1   g07512(.A1(\A[371] ), .A2(\A[372] ), .ZN(new_n8519_));
  INV_X1     g07513(.I(new_n8519_), .ZN(new_n8520_));
  NOR2_X1    g07514(.A1(\A[371] ), .A2(\A[372] ), .ZN(new_n8521_));
  OAI21_X1   g07515(.A1(new_n8520_), .A2(new_n8521_), .B(new_n8518_), .ZN(new_n8522_));
  NAND2_X1   g07516(.A1(new_n8517_), .A2(new_n8522_), .ZN(new_n8523_));
  AOI21_X1   g07517(.A1(\A[368] ), .A2(\A[369] ), .B(\A[367] ), .ZN(new_n8524_));
  AOI21_X1   g07518(.A1(\A[371] ), .A2(\A[372] ), .B(\A[370] ), .ZN(new_n8525_));
  OAI22_X1   g07519(.A1(new_n8510_), .A2(new_n8524_), .B1(new_n8525_), .B2(new_n8521_), .ZN(new_n8526_));
  INV_X1     g07520(.I(new_n8526_), .ZN(new_n8527_));
  NAND3_X1   g07521(.A1(new_n8512_), .A2(new_n8523_), .A3(new_n8527_), .ZN(new_n8528_));
  NOR2_X1    g07522(.A1(new_n8501_), .A2(new_n8528_), .ZN(new_n8529_));
  NOR2_X1    g07523(.A1(new_n8479_), .A2(\A[374] ), .ZN(new_n8530_));
  NOR2_X1    g07524(.A1(new_n8477_), .A2(\A[375] ), .ZN(new_n8531_));
  OAI21_X1   g07525(.A1(new_n8530_), .A2(new_n8531_), .B(\A[373] ), .ZN(new_n8532_));
  INV_X1     g07526(.I(new_n8482_), .ZN(new_n8533_));
  OAI21_X1   g07527(.A1(new_n8533_), .A2(new_n8483_), .B(new_n8476_), .ZN(new_n8534_));
  NAND2_X1   g07528(.A1(new_n8532_), .A2(new_n8534_), .ZN(new_n8535_));
  NOR2_X1    g07529(.A1(new_n8490_), .A2(\A[377] ), .ZN(new_n8536_));
  NOR2_X1    g07530(.A1(new_n8488_), .A2(\A[378] ), .ZN(new_n8537_));
  OAI21_X1   g07531(.A1(new_n8536_), .A2(new_n8537_), .B(\A[376] ), .ZN(new_n8538_));
  INV_X1     g07532(.I(new_n8493_), .ZN(new_n8539_));
  OAI21_X1   g07533(.A1(new_n8539_), .A2(new_n8494_), .B(new_n8487_), .ZN(new_n8540_));
  NAND2_X1   g07534(.A1(new_n8538_), .A2(new_n8540_), .ZN(new_n8541_));
  NOR2_X1    g07535(.A1(new_n8498_), .A2(new_n8483_), .ZN(new_n8542_));
  NOR2_X1    g07536(.A1(new_n8499_), .A2(new_n8494_), .ZN(new_n8543_));
  NOR2_X1    g07537(.A1(new_n8542_), .A2(new_n8543_), .ZN(new_n8544_));
  NAND3_X1   g07538(.A1(new_n8535_), .A2(new_n8541_), .A3(new_n8544_), .ZN(new_n8545_));
  NAND2_X1   g07539(.A1(new_n8504_), .A2(\A[369] ), .ZN(new_n8546_));
  NAND2_X1   g07540(.A1(new_n8502_), .A2(\A[368] ), .ZN(new_n8547_));
  AOI21_X1   g07541(.A1(new_n8546_), .A2(new_n8547_), .B(new_n8507_), .ZN(new_n8548_));
  INV_X1     g07542(.I(new_n8510_), .ZN(new_n8549_));
  AOI21_X1   g07543(.A1(new_n8549_), .A2(new_n8508_), .B(\A[367] ), .ZN(new_n8550_));
  NOR2_X1    g07544(.A1(new_n8550_), .A2(new_n8548_), .ZN(new_n8551_));
  NAND2_X1   g07545(.A1(new_n8515_), .A2(\A[372] ), .ZN(new_n8552_));
  NAND2_X1   g07546(.A1(new_n8513_), .A2(\A[371] ), .ZN(new_n8553_));
  AOI21_X1   g07547(.A1(new_n8552_), .A2(new_n8553_), .B(new_n8518_), .ZN(new_n8554_));
  INV_X1     g07548(.I(new_n8521_), .ZN(new_n8555_));
  AOI21_X1   g07549(.A1(new_n8555_), .A2(new_n8519_), .B(\A[370] ), .ZN(new_n8556_));
  NOR2_X1    g07550(.A1(new_n8556_), .A2(new_n8554_), .ZN(new_n8557_));
  NOR3_X1    g07551(.A1(new_n8551_), .A2(new_n8557_), .A3(new_n8526_), .ZN(new_n8558_));
  NOR2_X1    g07552(.A1(new_n8558_), .A2(new_n8545_), .ZN(new_n8559_));
  OAI22_X1   g07553(.A1(new_n8445_), .A2(new_n8475_), .B1(new_n8529_), .B2(new_n8559_), .ZN(new_n8560_));
  NOR2_X1    g07554(.A1(new_n8445_), .A2(new_n8475_), .ZN(new_n8561_));
  NOR2_X1    g07555(.A1(new_n8529_), .A2(new_n8559_), .ZN(new_n8562_));
  NAND2_X1   g07556(.A1(new_n8561_), .A2(new_n8562_), .ZN(new_n8563_));
  AND2_X2    g07557(.A1(new_n8563_), .A2(new_n8560_), .Z(new_n8564_));
  AOI21_X1   g07558(.A1(new_n8378_), .A2(new_n8391_), .B(new_n8564_), .ZN(new_n8565_));
  AND3_X2    g07559(.A1(new_n8378_), .A2(new_n8391_), .A3(new_n8564_), .Z(new_n8566_));
  INV_X1     g07560(.I(\A[439] ), .ZN(new_n8567_));
  INV_X1     g07561(.I(\A[440] ), .ZN(new_n8568_));
  NAND2_X1   g07562(.A1(new_n8568_), .A2(\A[441] ), .ZN(new_n8569_));
  INV_X1     g07563(.I(\A[441] ), .ZN(new_n8570_));
  NAND2_X1   g07564(.A1(new_n8570_), .A2(\A[440] ), .ZN(new_n8571_));
  AOI21_X1   g07565(.A1(new_n8569_), .A2(new_n8571_), .B(new_n8567_), .ZN(new_n8572_));
  NOR2_X1    g07566(.A1(\A[440] ), .A2(\A[441] ), .ZN(new_n8573_));
  INV_X1     g07567(.I(new_n8573_), .ZN(new_n8574_));
  NAND2_X1   g07568(.A1(\A[440] ), .A2(\A[441] ), .ZN(new_n8575_));
  AOI21_X1   g07569(.A1(new_n8574_), .A2(new_n8575_), .B(\A[439] ), .ZN(new_n8576_));
  NOR2_X1    g07570(.A1(new_n8576_), .A2(new_n8572_), .ZN(new_n8577_));
  INV_X1     g07571(.I(\A[444] ), .ZN(new_n8578_));
  NOR2_X1    g07572(.A1(new_n8578_), .A2(\A[443] ), .ZN(new_n8579_));
  INV_X1     g07573(.I(\A[443] ), .ZN(new_n8580_));
  NOR2_X1    g07574(.A1(new_n8580_), .A2(\A[444] ), .ZN(new_n8581_));
  OAI21_X1   g07575(.A1(new_n8579_), .A2(new_n8581_), .B(\A[442] ), .ZN(new_n8582_));
  INV_X1     g07576(.I(\A[442] ), .ZN(new_n8583_));
  NAND2_X1   g07577(.A1(\A[443] ), .A2(\A[444] ), .ZN(new_n8584_));
  INV_X1     g07578(.I(new_n8584_), .ZN(new_n8585_));
  NOR2_X1    g07579(.A1(\A[443] ), .A2(\A[444] ), .ZN(new_n8586_));
  OAI21_X1   g07580(.A1(new_n8585_), .A2(new_n8586_), .B(new_n8583_), .ZN(new_n8587_));
  NAND2_X1   g07581(.A1(new_n8582_), .A2(new_n8587_), .ZN(new_n8588_));
  AOI21_X1   g07582(.A1(new_n8567_), .A2(new_n8575_), .B(new_n8573_), .ZN(new_n8589_));
  AOI21_X1   g07583(.A1(new_n8583_), .A2(new_n8584_), .B(new_n8586_), .ZN(new_n8590_));
  NOR2_X1    g07584(.A1(new_n8589_), .A2(new_n8590_), .ZN(new_n8591_));
  XOR2_X1    g07585(.A1(new_n8577_), .A2(new_n8588_), .Z(new_n8592_));
  INV_X1     g07586(.I(\A[453] ), .ZN(new_n8593_));
  NOR2_X1    g07587(.A1(new_n8593_), .A2(\A[452] ), .ZN(new_n8594_));
  INV_X1     g07588(.I(\A[452] ), .ZN(new_n8595_));
  NOR2_X1    g07589(.A1(new_n8595_), .A2(\A[453] ), .ZN(new_n8596_));
  OAI21_X1   g07590(.A1(new_n8594_), .A2(new_n8596_), .B(\A[451] ), .ZN(new_n8597_));
  INV_X1     g07591(.I(\A[451] ), .ZN(new_n8598_));
  NOR2_X1    g07592(.A1(\A[452] ), .A2(\A[453] ), .ZN(new_n8599_));
  NAND2_X1   g07593(.A1(\A[452] ), .A2(\A[453] ), .ZN(new_n8600_));
  INV_X1     g07594(.I(new_n8600_), .ZN(new_n8601_));
  OAI21_X1   g07595(.A1(new_n8601_), .A2(new_n8599_), .B(new_n8598_), .ZN(new_n8602_));
  NAND2_X1   g07596(.A1(new_n8597_), .A2(new_n8602_), .ZN(new_n8603_));
  INV_X1     g07597(.I(\A[456] ), .ZN(new_n8604_));
  NOR2_X1    g07598(.A1(new_n8604_), .A2(\A[455] ), .ZN(new_n8605_));
  INV_X1     g07599(.I(\A[455] ), .ZN(new_n8606_));
  NOR2_X1    g07600(.A1(new_n8606_), .A2(\A[456] ), .ZN(new_n8607_));
  OAI21_X1   g07601(.A1(new_n8605_), .A2(new_n8607_), .B(\A[454] ), .ZN(new_n8608_));
  INV_X1     g07602(.I(\A[454] ), .ZN(new_n8609_));
  NAND2_X1   g07603(.A1(\A[455] ), .A2(\A[456] ), .ZN(new_n8610_));
  INV_X1     g07604(.I(new_n8610_), .ZN(new_n8611_));
  NOR2_X1    g07605(.A1(\A[455] ), .A2(\A[456] ), .ZN(new_n8612_));
  OAI21_X1   g07606(.A1(new_n8611_), .A2(new_n8612_), .B(new_n8609_), .ZN(new_n8613_));
  NAND2_X1   g07607(.A1(new_n8608_), .A2(new_n8613_), .ZN(new_n8614_));
  AOI21_X1   g07608(.A1(new_n8598_), .A2(new_n8600_), .B(new_n8599_), .ZN(new_n8615_));
  AOI21_X1   g07609(.A1(new_n8609_), .A2(new_n8610_), .B(new_n8612_), .ZN(new_n8616_));
  NOR2_X1    g07610(.A1(new_n8615_), .A2(new_n8616_), .ZN(new_n8617_));
  XOR2_X1    g07611(.A1(new_n8603_), .A2(new_n8614_), .Z(new_n8618_));
  INV_X1     g07612(.I(\A[457] ), .ZN(new_n8619_));
  INV_X1     g07613(.I(\A[458] ), .ZN(new_n8620_));
  NAND2_X1   g07614(.A1(new_n8620_), .A2(\A[459] ), .ZN(new_n8621_));
  INV_X1     g07615(.I(\A[459] ), .ZN(new_n8622_));
  NAND2_X1   g07616(.A1(new_n8622_), .A2(\A[458] ), .ZN(new_n8623_));
  AOI21_X1   g07617(.A1(new_n8621_), .A2(new_n8623_), .B(new_n8619_), .ZN(new_n8624_));
  NOR2_X1    g07618(.A1(\A[458] ), .A2(\A[459] ), .ZN(new_n8625_));
  INV_X1     g07619(.I(new_n8625_), .ZN(new_n8626_));
  NAND2_X1   g07620(.A1(\A[458] ), .A2(\A[459] ), .ZN(new_n8627_));
  AOI21_X1   g07621(.A1(new_n8626_), .A2(new_n8627_), .B(\A[457] ), .ZN(new_n8628_));
  NOR2_X1    g07622(.A1(new_n8628_), .A2(new_n8624_), .ZN(new_n8629_));
  INV_X1     g07623(.I(\A[462] ), .ZN(new_n8630_));
  NOR2_X1    g07624(.A1(new_n8630_), .A2(\A[461] ), .ZN(new_n8631_));
  INV_X1     g07625(.I(\A[461] ), .ZN(new_n8632_));
  NOR2_X1    g07626(.A1(new_n8632_), .A2(\A[462] ), .ZN(new_n8633_));
  OAI21_X1   g07627(.A1(new_n8631_), .A2(new_n8633_), .B(\A[460] ), .ZN(new_n8634_));
  INV_X1     g07628(.I(\A[460] ), .ZN(new_n8635_));
  NAND2_X1   g07629(.A1(\A[461] ), .A2(\A[462] ), .ZN(new_n8636_));
  INV_X1     g07630(.I(new_n8636_), .ZN(new_n8637_));
  NOR2_X1    g07631(.A1(\A[461] ), .A2(\A[462] ), .ZN(new_n8638_));
  OAI21_X1   g07632(.A1(new_n8637_), .A2(new_n8638_), .B(new_n8635_), .ZN(new_n8639_));
  NAND2_X1   g07633(.A1(new_n8634_), .A2(new_n8639_), .ZN(new_n8640_));
  AOI21_X1   g07634(.A1(\A[458] ), .A2(\A[459] ), .B(\A[457] ), .ZN(new_n8641_));
  NOR2_X1    g07635(.A1(new_n8641_), .A2(new_n8625_), .ZN(new_n8642_));
  AOI21_X1   g07636(.A1(\A[461] ), .A2(\A[462] ), .B(\A[460] ), .ZN(new_n8643_));
  NOR2_X1    g07637(.A1(new_n8643_), .A2(new_n8638_), .ZN(new_n8644_));
  NOR2_X1    g07638(.A1(new_n8642_), .A2(new_n8644_), .ZN(new_n8645_));
  XOR2_X1    g07639(.A1(new_n8629_), .A2(new_n8640_), .Z(new_n8646_));
  INV_X1     g07640(.I(\A[447] ), .ZN(new_n8647_));
  NOR2_X1    g07641(.A1(new_n8647_), .A2(\A[446] ), .ZN(new_n8648_));
  INV_X1     g07642(.I(\A[446] ), .ZN(new_n8649_));
  NOR2_X1    g07643(.A1(new_n8649_), .A2(\A[447] ), .ZN(new_n8650_));
  OAI21_X1   g07644(.A1(new_n8648_), .A2(new_n8650_), .B(\A[445] ), .ZN(new_n8651_));
  INV_X1     g07645(.I(\A[445] ), .ZN(new_n8652_));
  NOR2_X1    g07646(.A1(\A[446] ), .A2(\A[447] ), .ZN(new_n8653_));
  NAND2_X1   g07647(.A1(\A[446] ), .A2(\A[447] ), .ZN(new_n8654_));
  INV_X1     g07648(.I(new_n8654_), .ZN(new_n8655_));
  OAI21_X1   g07649(.A1(new_n8655_), .A2(new_n8653_), .B(new_n8652_), .ZN(new_n8656_));
  NAND2_X1   g07650(.A1(new_n8651_), .A2(new_n8656_), .ZN(new_n8657_));
  INV_X1     g07651(.I(\A[450] ), .ZN(new_n8658_));
  NOR2_X1    g07652(.A1(new_n8658_), .A2(\A[449] ), .ZN(new_n8659_));
  INV_X1     g07653(.I(\A[449] ), .ZN(new_n8660_));
  NOR2_X1    g07654(.A1(new_n8660_), .A2(\A[450] ), .ZN(new_n8661_));
  OAI21_X1   g07655(.A1(new_n8659_), .A2(new_n8661_), .B(\A[448] ), .ZN(new_n8662_));
  INV_X1     g07656(.I(\A[448] ), .ZN(new_n8663_));
  NOR2_X1    g07657(.A1(new_n8660_), .A2(new_n8658_), .ZN(new_n8664_));
  NOR2_X1    g07658(.A1(\A[449] ), .A2(\A[450] ), .ZN(new_n8665_));
  OAI21_X1   g07659(.A1(new_n8664_), .A2(new_n8665_), .B(new_n8663_), .ZN(new_n8666_));
  NAND2_X1   g07660(.A1(new_n8666_), .A2(new_n8662_), .ZN(new_n8667_));
  AOI21_X1   g07661(.A1(\A[446] ), .A2(\A[447] ), .B(\A[445] ), .ZN(new_n8668_));
  NOR2_X1    g07662(.A1(new_n8668_), .A2(new_n8653_), .ZN(new_n8669_));
  AOI21_X1   g07663(.A1(\A[449] ), .A2(\A[450] ), .B(\A[448] ), .ZN(new_n8670_));
  NOR2_X1    g07664(.A1(new_n8670_), .A2(new_n8665_), .ZN(new_n8671_));
  NOR2_X1    g07665(.A1(new_n8669_), .A2(new_n8671_), .ZN(new_n8672_));
  XOR2_X1    g07666(.A1(new_n8667_), .A2(new_n8657_), .Z(new_n8673_));
  XOR2_X1    g07667(.A1(new_n8646_), .A2(new_n8673_), .Z(new_n8674_));
  NOR2_X1    g07668(.A1(new_n8674_), .A2(new_n8618_), .ZN(new_n8675_));
  NAND2_X1   g07669(.A1(new_n8646_), .A2(new_n8673_), .ZN(new_n8676_));
  NOR2_X1    g07670(.A1(new_n8622_), .A2(\A[458] ), .ZN(new_n8677_));
  NOR2_X1    g07671(.A1(new_n8620_), .A2(\A[459] ), .ZN(new_n8678_));
  OAI21_X1   g07672(.A1(new_n8677_), .A2(new_n8678_), .B(\A[457] ), .ZN(new_n8679_));
  INV_X1     g07673(.I(new_n8627_), .ZN(new_n8680_));
  OAI21_X1   g07674(.A1(new_n8680_), .A2(new_n8625_), .B(new_n8619_), .ZN(new_n8681_));
  NAND2_X1   g07675(.A1(new_n8679_), .A2(new_n8681_), .ZN(new_n8682_));
  XOR2_X1    g07676(.A1(new_n8682_), .A2(new_n8640_), .Z(new_n8683_));
  NAND2_X1   g07677(.A1(new_n8649_), .A2(\A[447] ), .ZN(new_n8684_));
  NAND2_X1   g07678(.A1(new_n8647_), .A2(\A[446] ), .ZN(new_n8685_));
  AOI21_X1   g07679(.A1(new_n8684_), .A2(new_n8685_), .B(new_n8652_), .ZN(new_n8686_));
  INV_X1     g07680(.I(new_n8653_), .ZN(new_n8687_));
  AOI21_X1   g07681(.A1(new_n8687_), .A2(new_n8654_), .B(\A[445] ), .ZN(new_n8688_));
  NOR2_X1    g07682(.A1(new_n8688_), .A2(new_n8686_), .ZN(new_n8689_));
  XOR2_X1    g07683(.A1(new_n8689_), .A2(new_n8667_), .Z(new_n8690_));
  NAND2_X1   g07684(.A1(new_n8690_), .A2(new_n8683_), .ZN(new_n8691_));
  NAND3_X1   g07685(.A1(new_n8676_), .A2(new_n8691_), .A3(new_n8618_), .ZN(new_n8692_));
  INV_X1     g07686(.I(new_n8692_), .ZN(new_n8693_));
  OAI21_X1   g07687(.A1(new_n8675_), .A2(new_n8693_), .B(new_n8592_), .ZN(new_n8694_));
  INV_X1     g07688(.I(new_n8592_), .ZN(new_n8695_));
  NAND2_X1   g07689(.A1(new_n8595_), .A2(\A[453] ), .ZN(new_n8696_));
  NAND2_X1   g07690(.A1(new_n8593_), .A2(\A[452] ), .ZN(new_n8697_));
  AOI21_X1   g07691(.A1(new_n8696_), .A2(new_n8697_), .B(new_n8598_), .ZN(new_n8698_));
  INV_X1     g07692(.I(new_n8599_), .ZN(new_n8699_));
  AOI21_X1   g07693(.A1(new_n8699_), .A2(new_n8600_), .B(\A[451] ), .ZN(new_n8700_));
  NOR2_X1    g07694(.A1(new_n8700_), .A2(new_n8698_), .ZN(new_n8701_));
  XOR2_X1    g07695(.A1(new_n8701_), .A2(new_n8614_), .Z(new_n8702_));
  NAND2_X1   g07696(.A1(new_n8676_), .A2(new_n8691_), .ZN(new_n8703_));
  NAND2_X1   g07697(.A1(new_n8703_), .A2(new_n8702_), .ZN(new_n8704_));
  NAND3_X1   g07698(.A1(new_n8704_), .A2(new_n8692_), .A3(new_n8695_), .ZN(new_n8705_));
  INV_X1     g07699(.I(\A[415] ), .ZN(new_n8706_));
  INV_X1     g07700(.I(\A[416] ), .ZN(new_n8707_));
  NAND2_X1   g07701(.A1(new_n8707_), .A2(\A[417] ), .ZN(new_n8708_));
  INV_X1     g07702(.I(\A[417] ), .ZN(new_n8709_));
  NAND2_X1   g07703(.A1(new_n8709_), .A2(\A[416] ), .ZN(new_n8710_));
  AOI21_X1   g07704(.A1(new_n8708_), .A2(new_n8710_), .B(new_n8706_), .ZN(new_n8711_));
  NAND2_X1   g07705(.A1(\A[416] ), .A2(\A[417] ), .ZN(new_n8712_));
  NOR2_X1    g07706(.A1(\A[416] ), .A2(\A[417] ), .ZN(new_n8713_));
  INV_X1     g07707(.I(new_n8713_), .ZN(new_n8714_));
  AOI21_X1   g07708(.A1(new_n8714_), .A2(new_n8712_), .B(\A[415] ), .ZN(new_n8715_));
  INV_X1     g07709(.I(\A[418] ), .ZN(new_n8716_));
  INV_X1     g07710(.I(\A[419] ), .ZN(new_n8717_));
  NAND2_X1   g07711(.A1(new_n8717_), .A2(\A[420] ), .ZN(new_n8718_));
  INV_X1     g07712(.I(\A[420] ), .ZN(new_n8719_));
  NAND2_X1   g07713(.A1(new_n8719_), .A2(\A[419] ), .ZN(new_n8720_));
  AOI21_X1   g07714(.A1(new_n8718_), .A2(new_n8720_), .B(new_n8716_), .ZN(new_n8721_));
  NAND2_X1   g07715(.A1(\A[419] ), .A2(\A[420] ), .ZN(new_n8722_));
  NOR2_X1    g07716(.A1(\A[419] ), .A2(\A[420] ), .ZN(new_n8723_));
  INV_X1     g07717(.I(new_n8723_), .ZN(new_n8724_));
  AOI21_X1   g07718(.A1(new_n8724_), .A2(new_n8722_), .B(\A[418] ), .ZN(new_n8725_));
  OAI22_X1   g07719(.A1(new_n8711_), .A2(new_n8715_), .B1(new_n8725_), .B2(new_n8721_), .ZN(new_n8726_));
  NOR2_X1    g07720(.A1(new_n8709_), .A2(\A[416] ), .ZN(new_n8727_));
  NOR2_X1    g07721(.A1(new_n8707_), .A2(\A[417] ), .ZN(new_n8728_));
  OAI21_X1   g07722(.A1(new_n8727_), .A2(new_n8728_), .B(\A[415] ), .ZN(new_n8729_));
  INV_X1     g07723(.I(new_n8712_), .ZN(new_n8730_));
  OAI21_X1   g07724(.A1(new_n8730_), .A2(new_n8713_), .B(new_n8706_), .ZN(new_n8731_));
  NOR2_X1    g07725(.A1(new_n8719_), .A2(\A[419] ), .ZN(new_n8732_));
  NOR2_X1    g07726(.A1(new_n8717_), .A2(\A[420] ), .ZN(new_n8733_));
  OAI21_X1   g07727(.A1(new_n8732_), .A2(new_n8733_), .B(\A[418] ), .ZN(new_n8734_));
  INV_X1     g07728(.I(new_n8722_), .ZN(new_n8735_));
  OAI21_X1   g07729(.A1(new_n8735_), .A2(new_n8723_), .B(new_n8716_), .ZN(new_n8736_));
  NAND4_X1   g07730(.A1(new_n8729_), .A2(new_n8731_), .A3(new_n8734_), .A4(new_n8736_), .ZN(new_n8737_));
  NAND2_X1   g07731(.A1(new_n8734_), .A2(new_n8736_), .ZN(new_n8738_));
  AOI21_X1   g07732(.A1(\A[419] ), .A2(\A[420] ), .B(\A[418] ), .ZN(new_n8739_));
  NOR2_X1    g07733(.A1(new_n8739_), .A2(new_n8723_), .ZN(new_n8740_));
  NOR4_X1    g07734(.A1(new_n8740_), .A2(\A[415] ), .A3(\A[416] ), .A4(\A[417] ), .ZN(new_n8741_));
  NAND2_X1   g07735(.A1(new_n8738_), .A2(new_n8741_), .ZN(new_n8742_));
  NAND3_X1   g07736(.A1(new_n8742_), .A2(new_n8726_), .A3(new_n8737_), .ZN(new_n8743_));
  INV_X1     g07737(.I(\A[429] ), .ZN(new_n8744_));
  NOR2_X1    g07738(.A1(new_n8744_), .A2(\A[428] ), .ZN(new_n8745_));
  INV_X1     g07739(.I(\A[428] ), .ZN(new_n8746_));
  NOR2_X1    g07740(.A1(new_n8746_), .A2(\A[429] ), .ZN(new_n8747_));
  OAI21_X1   g07741(.A1(new_n8745_), .A2(new_n8747_), .B(\A[427] ), .ZN(new_n8748_));
  INV_X1     g07742(.I(\A[427] ), .ZN(new_n8749_));
  NAND2_X1   g07743(.A1(\A[428] ), .A2(\A[429] ), .ZN(new_n8750_));
  INV_X1     g07744(.I(new_n8750_), .ZN(new_n8751_));
  NOR2_X1    g07745(.A1(\A[428] ), .A2(\A[429] ), .ZN(new_n8752_));
  OAI21_X1   g07746(.A1(new_n8751_), .A2(new_n8752_), .B(new_n8749_), .ZN(new_n8753_));
  NAND2_X1   g07747(.A1(new_n8748_), .A2(new_n8753_), .ZN(new_n8754_));
  INV_X1     g07748(.I(\A[432] ), .ZN(new_n8755_));
  NOR2_X1    g07749(.A1(new_n8755_), .A2(\A[431] ), .ZN(new_n8756_));
  INV_X1     g07750(.I(\A[431] ), .ZN(new_n8757_));
  NOR2_X1    g07751(.A1(new_n8757_), .A2(\A[432] ), .ZN(new_n8758_));
  OAI21_X1   g07752(.A1(new_n8756_), .A2(new_n8758_), .B(\A[430] ), .ZN(new_n8759_));
  INV_X1     g07753(.I(\A[430] ), .ZN(new_n8760_));
  NAND2_X1   g07754(.A1(\A[431] ), .A2(\A[432] ), .ZN(new_n8761_));
  INV_X1     g07755(.I(new_n8761_), .ZN(new_n8762_));
  NOR2_X1    g07756(.A1(\A[431] ), .A2(\A[432] ), .ZN(new_n8763_));
  OAI21_X1   g07757(.A1(new_n8762_), .A2(new_n8763_), .B(new_n8760_), .ZN(new_n8764_));
  NAND2_X1   g07758(.A1(new_n8759_), .A2(new_n8764_), .ZN(new_n8765_));
  AOI21_X1   g07759(.A1(new_n8749_), .A2(new_n8750_), .B(new_n8752_), .ZN(new_n8766_));
  AOI21_X1   g07760(.A1(new_n8760_), .A2(new_n8761_), .B(new_n8763_), .ZN(new_n8767_));
  NOR2_X1    g07761(.A1(new_n8766_), .A2(new_n8767_), .ZN(new_n8768_));
  XOR2_X1    g07762(.A1(new_n8754_), .A2(new_n8765_), .Z(new_n8769_));
  INV_X1     g07763(.I(\A[433] ), .ZN(new_n8770_));
  INV_X1     g07764(.I(\A[434] ), .ZN(new_n8771_));
  NAND2_X1   g07765(.A1(new_n8771_), .A2(\A[435] ), .ZN(new_n8772_));
  INV_X1     g07766(.I(\A[435] ), .ZN(new_n8773_));
  NAND2_X1   g07767(.A1(new_n8773_), .A2(\A[434] ), .ZN(new_n8774_));
  AOI21_X1   g07768(.A1(new_n8772_), .A2(new_n8774_), .B(new_n8770_), .ZN(new_n8775_));
  NOR2_X1    g07769(.A1(\A[434] ), .A2(\A[435] ), .ZN(new_n8776_));
  INV_X1     g07770(.I(new_n8776_), .ZN(new_n8777_));
  NAND2_X1   g07771(.A1(\A[434] ), .A2(\A[435] ), .ZN(new_n8778_));
  AOI21_X1   g07772(.A1(new_n8777_), .A2(new_n8778_), .B(\A[433] ), .ZN(new_n8779_));
  NOR2_X1    g07773(.A1(new_n8779_), .A2(new_n8775_), .ZN(new_n8780_));
  INV_X1     g07774(.I(\A[438] ), .ZN(new_n8781_));
  NOR2_X1    g07775(.A1(new_n8781_), .A2(\A[437] ), .ZN(new_n8782_));
  INV_X1     g07776(.I(\A[437] ), .ZN(new_n8783_));
  NOR2_X1    g07777(.A1(new_n8783_), .A2(\A[438] ), .ZN(new_n8784_));
  OAI21_X1   g07778(.A1(new_n8782_), .A2(new_n8784_), .B(\A[436] ), .ZN(new_n8785_));
  INV_X1     g07779(.I(\A[436] ), .ZN(new_n8786_));
  NAND2_X1   g07780(.A1(\A[437] ), .A2(\A[438] ), .ZN(new_n8787_));
  INV_X1     g07781(.I(new_n8787_), .ZN(new_n8788_));
  NOR2_X1    g07782(.A1(\A[437] ), .A2(\A[438] ), .ZN(new_n8789_));
  OAI21_X1   g07783(.A1(new_n8788_), .A2(new_n8789_), .B(new_n8786_), .ZN(new_n8790_));
  NAND2_X1   g07784(.A1(new_n8785_), .A2(new_n8790_), .ZN(new_n8791_));
  AOI21_X1   g07785(.A1(\A[434] ), .A2(\A[435] ), .B(\A[433] ), .ZN(new_n8792_));
  AOI21_X1   g07786(.A1(\A[437] ), .A2(\A[438] ), .B(\A[436] ), .ZN(new_n8793_));
  OAI22_X1   g07787(.A1(new_n8776_), .A2(new_n8792_), .B1(new_n8793_), .B2(new_n8789_), .ZN(new_n8794_));
  INV_X1     g07788(.I(new_n8794_), .ZN(new_n8795_));
  XOR2_X1    g07789(.A1(new_n8780_), .A2(new_n8791_), .Z(new_n8796_));
  INV_X1     g07790(.I(\A[421] ), .ZN(new_n8797_));
  INV_X1     g07791(.I(\A[422] ), .ZN(new_n8798_));
  NAND2_X1   g07792(.A1(new_n8798_), .A2(\A[423] ), .ZN(new_n8799_));
  INV_X1     g07793(.I(\A[423] ), .ZN(new_n8800_));
  NAND2_X1   g07794(.A1(new_n8800_), .A2(\A[422] ), .ZN(new_n8801_));
  AOI21_X1   g07795(.A1(new_n8799_), .A2(new_n8801_), .B(new_n8797_), .ZN(new_n8802_));
  NAND2_X1   g07796(.A1(\A[422] ), .A2(\A[423] ), .ZN(new_n8803_));
  NOR2_X1    g07797(.A1(\A[422] ), .A2(\A[423] ), .ZN(new_n8804_));
  INV_X1     g07798(.I(new_n8804_), .ZN(new_n8805_));
  AOI21_X1   g07799(.A1(new_n8805_), .A2(new_n8803_), .B(\A[421] ), .ZN(new_n8806_));
  INV_X1     g07800(.I(\A[424] ), .ZN(new_n8807_));
  INV_X1     g07801(.I(\A[425] ), .ZN(new_n8808_));
  NAND2_X1   g07802(.A1(new_n8808_), .A2(\A[426] ), .ZN(new_n8809_));
  INV_X1     g07803(.I(\A[426] ), .ZN(new_n8810_));
  NAND2_X1   g07804(.A1(new_n8810_), .A2(\A[425] ), .ZN(new_n8811_));
  AOI21_X1   g07805(.A1(new_n8809_), .A2(new_n8811_), .B(new_n8807_), .ZN(new_n8812_));
  NAND2_X1   g07806(.A1(\A[425] ), .A2(\A[426] ), .ZN(new_n8813_));
  NOR2_X1    g07807(.A1(\A[425] ), .A2(\A[426] ), .ZN(new_n8814_));
  INV_X1     g07808(.I(new_n8814_), .ZN(new_n8815_));
  AOI21_X1   g07809(.A1(new_n8815_), .A2(new_n8813_), .B(\A[424] ), .ZN(new_n8816_));
  OAI22_X1   g07810(.A1(new_n8802_), .A2(new_n8806_), .B1(new_n8816_), .B2(new_n8812_), .ZN(new_n8817_));
  NOR2_X1    g07811(.A1(new_n8800_), .A2(\A[422] ), .ZN(new_n8818_));
  NOR2_X1    g07812(.A1(new_n8798_), .A2(\A[423] ), .ZN(new_n8819_));
  OAI21_X1   g07813(.A1(new_n8818_), .A2(new_n8819_), .B(\A[421] ), .ZN(new_n8820_));
  INV_X1     g07814(.I(new_n8803_), .ZN(new_n8821_));
  OAI21_X1   g07815(.A1(new_n8821_), .A2(new_n8804_), .B(new_n8797_), .ZN(new_n8822_));
  NOR2_X1    g07816(.A1(new_n8810_), .A2(\A[425] ), .ZN(new_n8823_));
  NOR2_X1    g07817(.A1(new_n8808_), .A2(\A[426] ), .ZN(new_n8824_));
  OAI21_X1   g07818(.A1(new_n8823_), .A2(new_n8824_), .B(\A[424] ), .ZN(new_n8825_));
  INV_X1     g07819(.I(new_n8813_), .ZN(new_n8826_));
  OAI21_X1   g07820(.A1(new_n8826_), .A2(new_n8814_), .B(new_n8807_), .ZN(new_n8827_));
  NAND4_X1   g07821(.A1(new_n8820_), .A2(new_n8822_), .A3(new_n8825_), .A4(new_n8827_), .ZN(new_n8828_));
  NAND2_X1   g07822(.A1(new_n8817_), .A2(new_n8828_), .ZN(new_n8829_));
  NAND2_X1   g07823(.A1(new_n8825_), .A2(new_n8827_), .ZN(new_n8830_));
  AOI21_X1   g07824(.A1(\A[425] ), .A2(\A[426] ), .B(\A[424] ), .ZN(new_n8831_));
  NOR2_X1    g07825(.A1(new_n8831_), .A2(new_n8814_), .ZN(new_n8832_));
  NOR4_X1    g07826(.A1(new_n8832_), .A2(\A[421] ), .A3(\A[422] ), .A4(\A[423] ), .ZN(new_n8833_));
  NAND2_X1   g07827(.A1(new_n8830_), .A2(new_n8833_), .ZN(new_n8834_));
  INV_X1     g07828(.I(new_n8834_), .ZN(new_n8835_));
  NOR2_X1    g07829(.A1(new_n8835_), .A2(new_n8829_), .ZN(new_n8836_));
  NAND2_X1   g07830(.A1(new_n8836_), .A2(new_n8796_), .ZN(new_n8837_));
  NOR2_X1    g07831(.A1(new_n8773_), .A2(\A[434] ), .ZN(new_n8838_));
  NOR2_X1    g07832(.A1(new_n8771_), .A2(\A[435] ), .ZN(new_n8839_));
  OAI21_X1   g07833(.A1(new_n8838_), .A2(new_n8839_), .B(\A[433] ), .ZN(new_n8840_));
  INV_X1     g07834(.I(new_n8778_), .ZN(new_n8841_));
  OAI21_X1   g07835(.A1(new_n8841_), .A2(new_n8776_), .B(new_n8770_), .ZN(new_n8842_));
  NAND2_X1   g07836(.A1(new_n8840_), .A2(new_n8842_), .ZN(new_n8843_));
  XOR2_X1    g07837(.A1(new_n8843_), .A2(new_n8791_), .Z(new_n8844_));
  AOI22_X1   g07838(.A1(new_n8820_), .A2(new_n8822_), .B1(new_n8825_), .B2(new_n8827_), .ZN(new_n8845_));
  NOR4_X1    g07839(.A1(new_n8802_), .A2(new_n8806_), .A3(new_n8816_), .A4(new_n8812_), .ZN(new_n8846_));
  NOR2_X1    g07840(.A1(new_n8845_), .A2(new_n8846_), .ZN(new_n8847_));
  NAND2_X1   g07841(.A1(new_n8847_), .A2(new_n8834_), .ZN(new_n8848_));
  NAND2_X1   g07842(.A1(new_n8848_), .A2(new_n8844_), .ZN(new_n8849_));
  AOI21_X1   g07843(.A1(new_n8837_), .A2(new_n8849_), .B(new_n8769_), .ZN(new_n8850_));
  NAND2_X1   g07844(.A1(new_n8754_), .A2(new_n8765_), .ZN(new_n8851_));
  NAND2_X1   g07845(.A1(new_n8746_), .A2(\A[429] ), .ZN(new_n8852_));
  NAND2_X1   g07846(.A1(new_n8744_), .A2(\A[428] ), .ZN(new_n8853_));
  AOI21_X1   g07847(.A1(new_n8852_), .A2(new_n8853_), .B(new_n8749_), .ZN(new_n8854_));
  INV_X1     g07848(.I(new_n8752_), .ZN(new_n8855_));
  AOI21_X1   g07849(.A1(new_n8855_), .A2(new_n8750_), .B(\A[427] ), .ZN(new_n8856_));
  NOR2_X1    g07850(.A1(new_n8856_), .A2(new_n8854_), .ZN(new_n8857_));
  NAND2_X1   g07851(.A1(new_n8757_), .A2(\A[432] ), .ZN(new_n8858_));
  NAND2_X1   g07852(.A1(new_n8755_), .A2(\A[431] ), .ZN(new_n8859_));
  AOI21_X1   g07853(.A1(new_n8858_), .A2(new_n8859_), .B(new_n8760_), .ZN(new_n8860_));
  INV_X1     g07854(.I(new_n8763_), .ZN(new_n8861_));
  AOI21_X1   g07855(.A1(new_n8861_), .A2(new_n8761_), .B(\A[430] ), .ZN(new_n8862_));
  NOR2_X1    g07856(.A1(new_n8862_), .A2(new_n8860_), .ZN(new_n8863_));
  NAND2_X1   g07857(.A1(new_n8857_), .A2(new_n8863_), .ZN(new_n8864_));
  NOR4_X1    g07858(.A1(new_n8767_), .A2(\A[427] ), .A3(\A[428] ), .A4(\A[429] ), .ZN(new_n8865_));
  NAND2_X1   g07859(.A1(new_n8765_), .A2(new_n8865_), .ZN(new_n8866_));
  NAND3_X1   g07860(.A1(new_n8864_), .A2(new_n8851_), .A3(new_n8866_), .ZN(new_n8867_));
  NOR2_X1    g07861(.A1(new_n8848_), .A2(new_n8844_), .ZN(new_n8868_));
  NOR2_X1    g07862(.A1(new_n8836_), .A2(new_n8796_), .ZN(new_n8869_));
  NOR3_X1    g07863(.A1(new_n8869_), .A2(new_n8868_), .A3(new_n8867_), .ZN(new_n8870_));
  OAI21_X1   g07864(.A1(new_n8850_), .A2(new_n8870_), .B(new_n8743_), .ZN(new_n8871_));
  INV_X1     g07865(.I(new_n8743_), .ZN(new_n8872_));
  INV_X1     g07866(.I(new_n8850_), .ZN(new_n8873_));
  NAND3_X1   g07867(.A1(new_n8837_), .A2(new_n8849_), .A3(new_n8769_), .ZN(new_n8874_));
  NAND3_X1   g07868(.A1(new_n8873_), .A2(new_n8874_), .A3(new_n8872_), .ZN(new_n8875_));
  AOI22_X1   g07869(.A1(new_n8694_), .A2(new_n8705_), .B1(new_n8871_), .B2(new_n8875_), .ZN(new_n8876_));
  AOI21_X1   g07870(.A1(new_n8704_), .A2(new_n8692_), .B(new_n8695_), .ZN(new_n8877_));
  NOR3_X1    g07871(.A1(new_n8675_), .A2(new_n8693_), .A3(new_n8592_), .ZN(new_n8878_));
  AOI21_X1   g07872(.A1(new_n8873_), .A2(new_n8874_), .B(new_n8872_), .ZN(new_n8879_));
  NOR3_X1    g07873(.A1(new_n8850_), .A2(new_n8870_), .A3(new_n8743_), .ZN(new_n8880_));
  NOR4_X1    g07874(.A1(new_n8878_), .A2(new_n8877_), .A3(new_n8879_), .A4(new_n8880_), .ZN(new_n8881_));
  OAI22_X1   g07875(.A1(new_n8566_), .A2(new_n8565_), .B1(new_n8876_), .B2(new_n8881_), .ZN(new_n8882_));
  NOR2_X1    g07876(.A1(new_n8566_), .A2(new_n8565_), .ZN(new_n8883_));
  NOR2_X1    g07877(.A1(new_n8876_), .A2(new_n8881_), .ZN(new_n8884_));
  NAND2_X1   g07878(.A1(new_n8883_), .A2(new_n8884_), .ZN(new_n8885_));
  INV_X1     g07879(.I(\A[343] ), .ZN(new_n8886_));
  INV_X1     g07880(.I(\A[344] ), .ZN(new_n8887_));
  NAND2_X1   g07881(.A1(new_n8887_), .A2(\A[345] ), .ZN(new_n8888_));
  INV_X1     g07882(.I(\A[345] ), .ZN(new_n8889_));
  NAND2_X1   g07883(.A1(new_n8889_), .A2(\A[344] ), .ZN(new_n8890_));
  AOI21_X1   g07884(.A1(new_n8888_), .A2(new_n8890_), .B(new_n8886_), .ZN(new_n8891_));
  NOR2_X1    g07885(.A1(\A[344] ), .A2(\A[345] ), .ZN(new_n8892_));
  INV_X1     g07886(.I(new_n8892_), .ZN(new_n8893_));
  NAND2_X1   g07887(.A1(\A[344] ), .A2(\A[345] ), .ZN(new_n8894_));
  AOI21_X1   g07888(.A1(new_n8893_), .A2(new_n8894_), .B(\A[343] ), .ZN(new_n8895_));
  NOR2_X1    g07889(.A1(new_n8895_), .A2(new_n8891_), .ZN(new_n8896_));
  INV_X1     g07890(.I(\A[348] ), .ZN(new_n8897_));
  NOR2_X1    g07891(.A1(new_n8897_), .A2(\A[347] ), .ZN(new_n8898_));
  INV_X1     g07892(.I(\A[347] ), .ZN(new_n8899_));
  NOR2_X1    g07893(.A1(new_n8899_), .A2(\A[348] ), .ZN(new_n8900_));
  OAI21_X1   g07894(.A1(new_n8898_), .A2(new_n8900_), .B(\A[346] ), .ZN(new_n8901_));
  INV_X1     g07895(.I(\A[346] ), .ZN(new_n8902_));
  NAND2_X1   g07896(.A1(\A[347] ), .A2(\A[348] ), .ZN(new_n8903_));
  INV_X1     g07897(.I(new_n8903_), .ZN(new_n8904_));
  NOR2_X1    g07898(.A1(\A[347] ), .A2(\A[348] ), .ZN(new_n8905_));
  OAI21_X1   g07899(.A1(new_n8904_), .A2(new_n8905_), .B(new_n8902_), .ZN(new_n8906_));
  NAND2_X1   g07900(.A1(new_n8901_), .A2(new_n8906_), .ZN(new_n8907_));
  AOI21_X1   g07901(.A1(new_n8886_), .A2(new_n8894_), .B(new_n8892_), .ZN(new_n8908_));
  AOI21_X1   g07902(.A1(new_n8902_), .A2(new_n8903_), .B(new_n8905_), .ZN(new_n8909_));
  NOR2_X1    g07903(.A1(new_n8908_), .A2(new_n8909_), .ZN(new_n8910_));
  XOR2_X1    g07904(.A1(new_n8896_), .A2(new_n8907_), .Z(new_n8911_));
  INV_X1     g07905(.I(\A[357] ), .ZN(new_n8912_));
  NOR2_X1    g07906(.A1(new_n8912_), .A2(\A[356] ), .ZN(new_n8913_));
  INV_X1     g07907(.I(\A[356] ), .ZN(new_n8914_));
  NOR2_X1    g07908(.A1(new_n8914_), .A2(\A[357] ), .ZN(new_n8915_));
  OAI21_X1   g07909(.A1(new_n8913_), .A2(new_n8915_), .B(\A[355] ), .ZN(new_n8916_));
  INV_X1     g07910(.I(\A[355] ), .ZN(new_n8917_));
  NOR2_X1    g07911(.A1(\A[356] ), .A2(\A[357] ), .ZN(new_n8918_));
  NAND2_X1   g07912(.A1(\A[356] ), .A2(\A[357] ), .ZN(new_n8919_));
  INV_X1     g07913(.I(new_n8919_), .ZN(new_n8920_));
  OAI21_X1   g07914(.A1(new_n8920_), .A2(new_n8918_), .B(new_n8917_), .ZN(new_n8921_));
  NAND2_X1   g07915(.A1(new_n8916_), .A2(new_n8921_), .ZN(new_n8922_));
  INV_X1     g07916(.I(\A[360] ), .ZN(new_n8923_));
  NOR2_X1    g07917(.A1(new_n8923_), .A2(\A[359] ), .ZN(new_n8924_));
  INV_X1     g07918(.I(\A[359] ), .ZN(new_n8925_));
  NOR2_X1    g07919(.A1(new_n8925_), .A2(\A[360] ), .ZN(new_n8926_));
  OAI21_X1   g07920(.A1(new_n8924_), .A2(new_n8926_), .B(\A[358] ), .ZN(new_n8927_));
  INV_X1     g07921(.I(\A[358] ), .ZN(new_n8928_));
  NAND2_X1   g07922(.A1(\A[359] ), .A2(\A[360] ), .ZN(new_n8929_));
  INV_X1     g07923(.I(new_n8929_), .ZN(new_n8930_));
  NOR2_X1    g07924(.A1(\A[359] ), .A2(\A[360] ), .ZN(new_n8931_));
  OAI21_X1   g07925(.A1(new_n8930_), .A2(new_n8931_), .B(new_n8928_), .ZN(new_n8932_));
  NAND2_X1   g07926(.A1(new_n8927_), .A2(new_n8932_), .ZN(new_n8933_));
  AOI21_X1   g07927(.A1(new_n8917_), .A2(new_n8919_), .B(new_n8918_), .ZN(new_n8934_));
  AOI21_X1   g07928(.A1(new_n8928_), .A2(new_n8929_), .B(new_n8931_), .ZN(new_n8935_));
  NOR2_X1    g07929(.A1(new_n8934_), .A2(new_n8935_), .ZN(new_n8936_));
  XOR2_X1    g07930(.A1(new_n8922_), .A2(new_n8933_), .Z(new_n8937_));
  INV_X1     g07931(.I(\A[363] ), .ZN(new_n8938_));
  NOR2_X1    g07932(.A1(new_n8938_), .A2(\A[362] ), .ZN(new_n8939_));
  INV_X1     g07933(.I(\A[362] ), .ZN(new_n8940_));
  NOR2_X1    g07934(.A1(new_n8940_), .A2(\A[363] ), .ZN(new_n8941_));
  OAI21_X1   g07935(.A1(new_n8939_), .A2(new_n8941_), .B(\A[361] ), .ZN(new_n8942_));
  INV_X1     g07936(.I(\A[361] ), .ZN(new_n8943_));
  NOR2_X1    g07937(.A1(\A[362] ), .A2(\A[363] ), .ZN(new_n8944_));
  AND2_X2    g07938(.A1(\A[362] ), .A2(\A[363] ), .Z(new_n8945_));
  OAI21_X1   g07939(.A1(new_n8945_), .A2(new_n8944_), .B(new_n8943_), .ZN(new_n8946_));
  NAND2_X1   g07940(.A1(new_n8942_), .A2(new_n8946_), .ZN(new_n8947_));
  INV_X1     g07941(.I(\A[366] ), .ZN(new_n8948_));
  NOR2_X1    g07942(.A1(new_n8948_), .A2(\A[365] ), .ZN(new_n8949_));
  INV_X1     g07943(.I(\A[365] ), .ZN(new_n8950_));
  NOR2_X1    g07944(.A1(new_n8950_), .A2(\A[366] ), .ZN(new_n8951_));
  OAI21_X1   g07945(.A1(new_n8949_), .A2(new_n8951_), .B(\A[364] ), .ZN(new_n8952_));
  INV_X1     g07946(.I(\A[364] ), .ZN(new_n8953_));
  NAND2_X1   g07947(.A1(\A[365] ), .A2(\A[366] ), .ZN(new_n8954_));
  INV_X1     g07948(.I(new_n8954_), .ZN(new_n8955_));
  NOR2_X1    g07949(.A1(\A[365] ), .A2(\A[366] ), .ZN(new_n8956_));
  OAI21_X1   g07950(.A1(new_n8955_), .A2(new_n8956_), .B(new_n8953_), .ZN(new_n8957_));
  NAND2_X1   g07951(.A1(new_n8952_), .A2(new_n8957_), .ZN(new_n8958_));
  AOI21_X1   g07952(.A1(\A[362] ), .A2(\A[363] ), .B(\A[361] ), .ZN(new_n8959_));
  NOR2_X1    g07953(.A1(new_n8959_), .A2(new_n8944_), .ZN(new_n8960_));
  AOI21_X1   g07954(.A1(\A[365] ), .A2(\A[366] ), .B(\A[364] ), .ZN(new_n8961_));
  NOR2_X1    g07955(.A1(new_n8961_), .A2(new_n8956_), .ZN(new_n8962_));
  NOR2_X1    g07956(.A1(new_n8960_), .A2(new_n8962_), .ZN(new_n8963_));
  XOR2_X1    g07957(.A1(new_n8958_), .A2(new_n8947_), .Z(new_n8964_));
  INV_X1     g07958(.I(\A[349] ), .ZN(new_n8965_));
  INV_X1     g07959(.I(\A[350] ), .ZN(new_n8966_));
  NAND2_X1   g07960(.A1(new_n8966_), .A2(\A[351] ), .ZN(new_n8967_));
  INV_X1     g07961(.I(\A[351] ), .ZN(new_n8968_));
  NAND2_X1   g07962(.A1(new_n8968_), .A2(\A[350] ), .ZN(new_n8969_));
  AOI21_X1   g07963(.A1(new_n8967_), .A2(new_n8969_), .B(new_n8965_), .ZN(new_n8970_));
  NOR2_X1    g07964(.A1(\A[350] ), .A2(\A[351] ), .ZN(new_n8971_));
  INV_X1     g07965(.I(new_n8971_), .ZN(new_n8972_));
  NAND2_X1   g07966(.A1(\A[350] ), .A2(\A[351] ), .ZN(new_n8973_));
  AOI21_X1   g07967(.A1(new_n8972_), .A2(new_n8973_), .B(\A[349] ), .ZN(new_n8974_));
  NOR2_X1    g07968(.A1(new_n8974_), .A2(new_n8970_), .ZN(new_n8975_));
  INV_X1     g07969(.I(\A[354] ), .ZN(new_n8976_));
  NOR2_X1    g07970(.A1(new_n8976_), .A2(\A[353] ), .ZN(new_n8977_));
  INV_X1     g07971(.I(\A[353] ), .ZN(new_n8978_));
  NOR2_X1    g07972(.A1(new_n8978_), .A2(\A[354] ), .ZN(new_n8979_));
  OAI21_X1   g07973(.A1(new_n8977_), .A2(new_n8979_), .B(\A[352] ), .ZN(new_n8980_));
  INV_X1     g07974(.I(\A[352] ), .ZN(new_n8981_));
  NAND2_X1   g07975(.A1(\A[353] ), .A2(\A[354] ), .ZN(new_n8982_));
  INV_X1     g07976(.I(new_n8982_), .ZN(new_n8983_));
  NOR2_X1    g07977(.A1(\A[353] ), .A2(\A[354] ), .ZN(new_n8984_));
  OAI21_X1   g07978(.A1(new_n8983_), .A2(new_n8984_), .B(new_n8981_), .ZN(new_n8985_));
  NAND2_X1   g07979(.A1(new_n8980_), .A2(new_n8985_), .ZN(new_n8986_));
  AOI21_X1   g07980(.A1(\A[350] ), .A2(\A[351] ), .B(\A[349] ), .ZN(new_n8987_));
  NOR2_X1    g07981(.A1(new_n8987_), .A2(new_n8971_), .ZN(new_n8988_));
  AOI21_X1   g07982(.A1(\A[353] ), .A2(\A[354] ), .B(\A[352] ), .ZN(new_n8989_));
  NOR2_X1    g07983(.A1(new_n8989_), .A2(new_n8984_), .ZN(new_n8990_));
  NOR2_X1    g07984(.A1(new_n8988_), .A2(new_n8990_), .ZN(new_n8991_));
  XOR2_X1    g07985(.A1(new_n8975_), .A2(new_n8986_), .Z(new_n8992_));
  XOR2_X1    g07986(.A1(new_n8992_), .A2(new_n8964_), .Z(new_n8993_));
  NOR2_X1    g07987(.A1(new_n8993_), .A2(new_n8937_), .ZN(new_n8994_));
  NAND2_X1   g07988(.A1(new_n8914_), .A2(\A[357] ), .ZN(new_n8995_));
  NAND2_X1   g07989(.A1(new_n8912_), .A2(\A[356] ), .ZN(new_n8996_));
  AOI21_X1   g07990(.A1(new_n8995_), .A2(new_n8996_), .B(new_n8917_), .ZN(new_n8997_));
  INV_X1     g07991(.I(new_n8918_), .ZN(new_n8998_));
  AOI21_X1   g07992(.A1(new_n8998_), .A2(new_n8919_), .B(\A[355] ), .ZN(new_n8999_));
  NOR2_X1    g07993(.A1(new_n8999_), .A2(new_n8997_), .ZN(new_n9000_));
  XOR2_X1    g07994(.A1(new_n9000_), .A2(new_n8933_), .Z(new_n9001_));
  NAND2_X1   g07995(.A1(new_n8950_), .A2(\A[366] ), .ZN(new_n9002_));
  NAND2_X1   g07996(.A1(new_n8948_), .A2(\A[365] ), .ZN(new_n9003_));
  AOI21_X1   g07997(.A1(new_n9002_), .A2(new_n9003_), .B(new_n8953_), .ZN(new_n9004_));
  INV_X1     g07998(.I(new_n8956_), .ZN(new_n9005_));
  AOI21_X1   g07999(.A1(new_n9005_), .A2(new_n8954_), .B(\A[364] ), .ZN(new_n9006_));
  NOR2_X1    g08000(.A1(new_n9006_), .A2(new_n9004_), .ZN(new_n9007_));
  XOR2_X1    g08001(.A1(new_n9007_), .A2(new_n8947_), .Z(new_n9008_));
  NOR2_X1    g08002(.A1(new_n8968_), .A2(\A[350] ), .ZN(new_n9009_));
  NOR2_X1    g08003(.A1(new_n8966_), .A2(\A[351] ), .ZN(new_n9010_));
  OAI21_X1   g08004(.A1(new_n9009_), .A2(new_n9010_), .B(\A[349] ), .ZN(new_n9011_));
  INV_X1     g08005(.I(new_n8973_), .ZN(new_n9012_));
  OAI21_X1   g08006(.A1(new_n9012_), .A2(new_n8971_), .B(new_n8965_), .ZN(new_n9013_));
  NAND2_X1   g08007(.A1(new_n9011_), .A2(new_n9013_), .ZN(new_n9014_));
  XOR2_X1    g08008(.A1(new_n9014_), .A2(new_n8986_), .Z(new_n9015_));
  NAND2_X1   g08009(.A1(new_n9015_), .A2(new_n9008_), .ZN(new_n9016_));
  NAND2_X1   g08010(.A1(new_n8992_), .A2(new_n8964_), .ZN(new_n9017_));
  NAND2_X1   g08011(.A1(new_n9016_), .A2(new_n9017_), .ZN(new_n9018_));
  NOR2_X1    g08012(.A1(new_n9018_), .A2(new_n9001_), .ZN(new_n9019_));
  OAI21_X1   g08013(.A1(new_n8994_), .A2(new_n9019_), .B(new_n8911_), .ZN(new_n9020_));
  INV_X1     g08014(.I(new_n8911_), .ZN(new_n9021_));
  NAND2_X1   g08015(.A1(new_n9018_), .A2(new_n9001_), .ZN(new_n9022_));
  NAND2_X1   g08016(.A1(new_n8993_), .A2(new_n8937_), .ZN(new_n9023_));
  NAND3_X1   g08017(.A1(new_n9023_), .A2(new_n9022_), .A3(new_n9021_), .ZN(new_n9024_));
  INV_X1     g08018(.I(\A[319] ), .ZN(new_n9025_));
  INV_X1     g08019(.I(\A[320] ), .ZN(new_n9026_));
  NAND2_X1   g08020(.A1(new_n9026_), .A2(\A[321] ), .ZN(new_n9027_));
  INV_X1     g08021(.I(\A[321] ), .ZN(new_n9028_));
  NAND2_X1   g08022(.A1(new_n9028_), .A2(\A[320] ), .ZN(new_n9029_));
  AOI21_X1   g08023(.A1(new_n9027_), .A2(new_n9029_), .B(new_n9025_), .ZN(new_n9030_));
  NAND2_X1   g08024(.A1(\A[320] ), .A2(\A[321] ), .ZN(new_n9031_));
  NOR2_X1    g08025(.A1(\A[320] ), .A2(\A[321] ), .ZN(new_n9032_));
  INV_X1     g08026(.I(new_n9032_), .ZN(new_n9033_));
  AOI21_X1   g08027(.A1(new_n9033_), .A2(new_n9031_), .B(\A[319] ), .ZN(new_n9034_));
  INV_X1     g08028(.I(\A[322] ), .ZN(new_n9035_));
  INV_X1     g08029(.I(\A[323] ), .ZN(new_n9036_));
  NAND2_X1   g08030(.A1(new_n9036_), .A2(\A[324] ), .ZN(new_n9037_));
  INV_X1     g08031(.I(\A[324] ), .ZN(new_n9038_));
  NAND2_X1   g08032(.A1(new_n9038_), .A2(\A[323] ), .ZN(new_n9039_));
  AOI21_X1   g08033(.A1(new_n9037_), .A2(new_n9039_), .B(new_n9035_), .ZN(new_n9040_));
  NAND2_X1   g08034(.A1(\A[323] ), .A2(\A[324] ), .ZN(new_n9041_));
  NOR2_X1    g08035(.A1(\A[323] ), .A2(\A[324] ), .ZN(new_n9042_));
  INV_X1     g08036(.I(new_n9042_), .ZN(new_n9043_));
  AOI21_X1   g08037(.A1(new_n9043_), .A2(new_n9041_), .B(\A[322] ), .ZN(new_n9044_));
  OAI22_X1   g08038(.A1(new_n9030_), .A2(new_n9034_), .B1(new_n9044_), .B2(new_n9040_), .ZN(new_n9045_));
  NOR2_X1    g08039(.A1(new_n9028_), .A2(\A[320] ), .ZN(new_n9046_));
  NOR2_X1    g08040(.A1(new_n9026_), .A2(\A[321] ), .ZN(new_n9047_));
  OAI21_X1   g08041(.A1(new_n9046_), .A2(new_n9047_), .B(\A[319] ), .ZN(new_n9048_));
  INV_X1     g08042(.I(new_n9031_), .ZN(new_n9049_));
  OAI21_X1   g08043(.A1(new_n9049_), .A2(new_n9032_), .B(new_n9025_), .ZN(new_n9050_));
  NOR2_X1    g08044(.A1(new_n9038_), .A2(\A[323] ), .ZN(new_n9051_));
  NOR2_X1    g08045(.A1(new_n9036_), .A2(\A[324] ), .ZN(new_n9052_));
  OAI21_X1   g08046(.A1(new_n9051_), .A2(new_n9052_), .B(\A[322] ), .ZN(new_n9053_));
  INV_X1     g08047(.I(new_n9041_), .ZN(new_n9054_));
  OAI21_X1   g08048(.A1(new_n9054_), .A2(new_n9042_), .B(new_n9035_), .ZN(new_n9055_));
  NAND4_X1   g08049(.A1(new_n9048_), .A2(new_n9050_), .A3(new_n9053_), .A4(new_n9055_), .ZN(new_n9056_));
  NAND2_X1   g08050(.A1(new_n9045_), .A2(new_n9056_), .ZN(new_n9057_));
  NOR2_X1    g08051(.A1(new_n9034_), .A2(new_n9030_), .ZN(new_n9058_));
  NOR2_X1    g08052(.A1(new_n9044_), .A2(new_n9040_), .ZN(new_n9059_));
  AOI21_X1   g08053(.A1(\A[320] ), .A2(\A[321] ), .B(\A[319] ), .ZN(new_n9060_));
  AOI21_X1   g08054(.A1(\A[323] ), .A2(\A[324] ), .B(\A[322] ), .ZN(new_n9061_));
  OAI22_X1   g08055(.A1(new_n9032_), .A2(new_n9060_), .B1(new_n9061_), .B2(new_n9042_), .ZN(new_n9062_));
  NOR3_X1    g08056(.A1(new_n9058_), .A2(new_n9059_), .A3(new_n9062_), .ZN(new_n9063_));
  NOR2_X1    g08057(.A1(new_n9057_), .A2(new_n9063_), .ZN(new_n9064_));
  INV_X1     g08058(.I(\A[331] ), .ZN(new_n9065_));
  INV_X1     g08059(.I(\A[332] ), .ZN(new_n9066_));
  NAND2_X1   g08060(.A1(new_n9066_), .A2(\A[333] ), .ZN(new_n9067_));
  INV_X1     g08061(.I(\A[333] ), .ZN(new_n9068_));
  NAND2_X1   g08062(.A1(new_n9068_), .A2(\A[332] ), .ZN(new_n9069_));
  AOI21_X1   g08063(.A1(new_n9067_), .A2(new_n9069_), .B(new_n9065_), .ZN(new_n9070_));
  NAND2_X1   g08064(.A1(\A[332] ), .A2(\A[333] ), .ZN(new_n9071_));
  NOR2_X1    g08065(.A1(\A[332] ), .A2(\A[333] ), .ZN(new_n9072_));
  INV_X1     g08066(.I(new_n9072_), .ZN(new_n9073_));
  AOI21_X1   g08067(.A1(new_n9073_), .A2(new_n9071_), .B(\A[331] ), .ZN(new_n9074_));
  NOR2_X1    g08068(.A1(new_n9074_), .A2(new_n9070_), .ZN(new_n9075_));
  INV_X1     g08069(.I(\A[336] ), .ZN(new_n9076_));
  NOR2_X1    g08070(.A1(new_n9076_), .A2(\A[335] ), .ZN(new_n9077_));
  INV_X1     g08071(.I(\A[335] ), .ZN(new_n9078_));
  NOR2_X1    g08072(.A1(new_n9078_), .A2(\A[336] ), .ZN(new_n9079_));
  OAI21_X1   g08073(.A1(new_n9077_), .A2(new_n9079_), .B(\A[334] ), .ZN(new_n9080_));
  INV_X1     g08074(.I(\A[334] ), .ZN(new_n9081_));
  NAND2_X1   g08075(.A1(\A[335] ), .A2(\A[336] ), .ZN(new_n9082_));
  INV_X1     g08076(.I(new_n9082_), .ZN(new_n9083_));
  NOR2_X1    g08077(.A1(\A[335] ), .A2(\A[336] ), .ZN(new_n9084_));
  OAI21_X1   g08078(.A1(new_n9083_), .A2(new_n9084_), .B(new_n9081_), .ZN(new_n9085_));
  NAND2_X1   g08079(.A1(new_n9080_), .A2(new_n9085_), .ZN(new_n9086_));
  AOI21_X1   g08080(.A1(new_n9065_), .A2(new_n9071_), .B(new_n9072_), .ZN(new_n9087_));
  AOI21_X1   g08081(.A1(new_n9081_), .A2(new_n9082_), .B(new_n9084_), .ZN(new_n9088_));
  NOR2_X1    g08082(.A1(new_n9087_), .A2(new_n9088_), .ZN(new_n9089_));
  XOR2_X1    g08083(.A1(new_n9075_), .A2(new_n9086_), .Z(new_n9090_));
  INV_X1     g08084(.I(\A[339] ), .ZN(new_n9091_));
  NOR2_X1    g08085(.A1(new_n9091_), .A2(\A[338] ), .ZN(new_n9092_));
  INV_X1     g08086(.I(\A[338] ), .ZN(new_n9093_));
  NOR2_X1    g08087(.A1(new_n9093_), .A2(\A[339] ), .ZN(new_n9094_));
  OAI21_X1   g08088(.A1(new_n9092_), .A2(new_n9094_), .B(\A[337] ), .ZN(new_n9095_));
  INV_X1     g08089(.I(\A[337] ), .ZN(new_n9096_));
  NOR2_X1    g08090(.A1(\A[338] ), .A2(\A[339] ), .ZN(new_n9097_));
  NAND2_X1   g08091(.A1(\A[338] ), .A2(\A[339] ), .ZN(new_n9098_));
  INV_X1     g08092(.I(new_n9098_), .ZN(new_n9099_));
  OAI21_X1   g08093(.A1(new_n9099_), .A2(new_n9097_), .B(new_n9096_), .ZN(new_n9100_));
  NAND2_X1   g08094(.A1(new_n9095_), .A2(new_n9100_), .ZN(new_n9101_));
  INV_X1     g08095(.I(\A[342] ), .ZN(new_n9102_));
  NOR2_X1    g08096(.A1(new_n9102_), .A2(\A[341] ), .ZN(new_n9103_));
  INV_X1     g08097(.I(\A[341] ), .ZN(new_n9104_));
  NOR2_X1    g08098(.A1(new_n9104_), .A2(\A[342] ), .ZN(new_n9105_));
  OAI21_X1   g08099(.A1(new_n9103_), .A2(new_n9105_), .B(\A[340] ), .ZN(new_n9106_));
  INV_X1     g08100(.I(\A[340] ), .ZN(new_n9107_));
  NAND2_X1   g08101(.A1(\A[341] ), .A2(\A[342] ), .ZN(new_n9108_));
  INV_X1     g08102(.I(new_n9108_), .ZN(new_n9109_));
  NOR2_X1    g08103(.A1(\A[341] ), .A2(\A[342] ), .ZN(new_n9110_));
  OAI21_X1   g08104(.A1(new_n9109_), .A2(new_n9110_), .B(new_n9107_), .ZN(new_n9111_));
  NAND2_X1   g08105(.A1(new_n9106_), .A2(new_n9111_), .ZN(new_n9112_));
  AOI21_X1   g08106(.A1(\A[338] ), .A2(\A[339] ), .B(\A[337] ), .ZN(new_n9113_));
  AOI21_X1   g08107(.A1(\A[341] ), .A2(\A[342] ), .B(\A[340] ), .ZN(new_n9114_));
  OAI22_X1   g08108(.A1(new_n9097_), .A2(new_n9113_), .B1(new_n9114_), .B2(new_n9110_), .ZN(new_n9115_));
  INV_X1     g08109(.I(new_n9115_), .ZN(new_n9116_));
  XOR2_X1    g08110(.A1(new_n9101_), .A2(new_n9112_), .Z(new_n9117_));
  INV_X1     g08111(.I(\A[327] ), .ZN(new_n9118_));
  NOR2_X1    g08112(.A1(new_n9118_), .A2(\A[326] ), .ZN(new_n9119_));
  INV_X1     g08113(.I(\A[326] ), .ZN(new_n9120_));
  NOR2_X1    g08114(.A1(new_n9120_), .A2(\A[327] ), .ZN(new_n9121_));
  OAI21_X1   g08115(.A1(new_n9119_), .A2(new_n9121_), .B(\A[325] ), .ZN(new_n9122_));
  INV_X1     g08116(.I(\A[325] ), .ZN(new_n9123_));
  AND2_X2    g08117(.A1(\A[326] ), .A2(\A[327] ), .Z(new_n9124_));
  NOR2_X1    g08118(.A1(\A[326] ), .A2(\A[327] ), .ZN(new_n9125_));
  OAI21_X1   g08119(.A1(new_n9124_), .A2(new_n9125_), .B(new_n9123_), .ZN(new_n9126_));
  INV_X1     g08120(.I(\A[330] ), .ZN(new_n9127_));
  NOR2_X1    g08121(.A1(new_n9127_), .A2(\A[329] ), .ZN(new_n9128_));
  INV_X1     g08122(.I(\A[329] ), .ZN(new_n9129_));
  NOR2_X1    g08123(.A1(new_n9129_), .A2(\A[330] ), .ZN(new_n9130_));
  OAI21_X1   g08124(.A1(new_n9128_), .A2(new_n9130_), .B(\A[328] ), .ZN(new_n9131_));
  INV_X1     g08125(.I(\A[328] ), .ZN(new_n9132_));
  NAND2_X1   g08126(.A1(\A[329] ), .A2(\A[330] ), .ZN(new_n9133_));
  INV_X1     g08127(.I(new_n9133_), .ZN(new_n9134_));
  NOR2_X1    g08128(.A1(\A[329] ), .A2(\A[330] ), .ZN(new_n9135_));
  OAI21_X1   g08129(.A1(new_n9134_), .A2(new_n9135_), .B(new_n9132_), .ZN(new_n9136_));
  AOI22_X1   g08130(.A1(new_n9131_), .A2(new_n9136_), .B1(new_n9122_), .B2(new_n9126_), .ZN(new_n9137_));
  NAND2_X1   g08131(.A1(new_n9120_), .A2(\A[327] ), .ZN(new_n9138_));
  NAND2_X1   g08132(.A1(new_n9118_), .A2(\A[326] ), .ZN(new_n9139_));
  AOI21_X1   g08133(.A1(new_n9138_), .A2(new_n9139_), .B(new_n9123_), .ZN(new_n9140_));
  NAND2_X1   g08134(.A1(\A[326] ), .A2(\A[327] ), .ZN(new_n9141_));
  INV_X1     g08135(.I(new_n9125_), .ZN(new_n9142_));
  AOI21_X1   g08136(.A1(new_n9142_), .A2(new_n9141_), .B(\A[325] ), .ZN(new_n9143_));
  NAND2_X1   g08137(.A1(new_n9129_), .A2(\A[330] ), .ZN(new_n9144_));
  NAND2_X1   g08138(.A1(new_n9127_), .A2(\A[329] ), .ZN(new_n9145_));
  AOI21_X1   g08139(.A1(new_n9144_), .A2(new_n9145_), .B(new_n9132_), .ZN(new_n9146_));
  INV_X1     g08140(.I(new_n9135_), .ZN(new_n9147_));
  AOI21_X1   g08141(.A1(new_n9147_), .A2(new_n9133_), .B(\A[328] ), .ZN(new_n9148_));
  NOR4_X1    g08142(.A1(new_n9140_), .A2(new_n9143_), .A3(new_n9148_), .A4(new_n9146_), .ZN(new_n9149_));
  NOR2_X1    g08143(.A1(new_n9149_), .A2(new_n9137_), .ZN(new_n9150_));
  NAND2_X1   g08144(.A1(new_n9131_), .A2(new_n9136_), .ZN(new_n9151_));
  AOI21_X1   g08145(.A1(\A[329] ), .A2(\A[330] ), .B(\A[328] ), .ZN(new_n9152_));
  NOR2_X1    g08146(.A1(new_n9152_), .A2(new_n9135_), .ZN(new_n9153_));
  NOR4_X1    g08147(.A1(new_n9153_), .A2(\A[325] ), .A3(\A[326] ), .A4(\A[327] ), .ZN(new_n9154_));
  NAND2_X1   g08148(.A1(new_n9151_), .A2(new_n9154_), .ZN(new_n9155_));
  NAND2_X1   g08149(.A1(new_n9150_), .A2(new_n9155_), .ZN(new_n9156_));
  NOR2_X1    g08150(.A1(new_n9156_), .A2(new_n9117_), .ZN(new_n9157_));
  NAND2_X1   g08151(.A1(new_n9093_), .A2(\A[339] ), .ZN(new_n9158_));
  NAND2_X1   g08152(.A1(new_n9091_), .A2(\A[338] ), .ZN(new_n9159_));
  AOI21_X1   g08153(.A1(new_n9158_), .A2(new_n9159_), .B(new_n9096_), .ZN(new_n9160_));
  INV_X1     g08154(.I(new_n9097_), .ZN(new_n9161_));
  AOI21_X1   g08155(.A1(new_n9161_), .A2(new_n9098_), .B(\A[337] ), .ZN(new_n9162_));
  NOR2_X1    g08156(.A1(new_n9162_), .A2(new_n9160_), .ZN(new_n9163_));
  XOR2_X1    g08157(.A1(new_n9163_), .A2(new_n9112_), .Z(new_n9164_));
  OAI22_X1   g08158(.A1(new_n9140_), .A2(new_n9143_), .B1(new_n9148_), .B2(new_n9146_), .ZN(new_n9165_));
  NAND4_X1   g08159(.A1(new_n9122_), .A2(new_n9131_), .A3(new_n9136_), .A4(new_n9126_), .ZN(new_n9166_));
  NAND2_X1   g08160(.A1(new_n9165_), .A2(new_n9166_), .ZN(new_n9167_));
  NOR2_X1    g08161(.A1(new_n9143_), .A2(new_n9140_), .ZN(new_n9168_));
  NOR2_X1    g08162(.A1(new_n9148_), .A2(new_n9146_), .ZN(new_n9169_));
  AOI21_X1   g08163(.A1(\A[326] ), .A2(\A[327] ), .B(\A[325] ), .ZN(new_n9170_));
  OAI22_X1   g08164(.A1(new_n9125_), .A2(new_n9170_), .B1(new_n9152_), .B2(new_n9135_), .ZN(new_n9171_));
  NOR3_X1    g08165(.A1(new_n9168_), .A2(new_n9169_), .A3(new_n9171_), .ZN(new_n9172_));
  NOR2_X1    g08166(.A1(new_n9167_), .A2(new_n9172_), .ZN(new_n9173_));
  NOR2_X1    g08167(.A1(new_n9164_), .A2(new_n9173_), .ZN(new_n9174_));
  OAI21_X1   g08168(.A1(new_n9157_), .A2(new_n9174_), .B(new_n9090_), .ZN(new_n9175_));
  NOR2_X1    g08169(.A1(new_n9068_), .A2(\A[332] ), .ZN(new_n9176_));
  NOR2_X1    g08170(.A1(new_n9066_), .A2(\A[333] ), .ZN(new_n9177_));
  OAI21_X1   g08171(.A1(new_n9176_), .A2(new_n9177_), .B(\A[331] ), .ZN(new_n9178_));
  INV_X1     g08172(.I(new_n9071_), .ZN(new_n9179_));
  OAI21_X1   g08173(.A1(new_n9179_), .A2(new_n9072_), .B(new_n9065_), .ZN(new_n9180_));
  NAND2_X1   g08174(.A1(new_n9178_), .A2(new_n9180_), .ZN(new_n9181_));
  XOR2_X1    g08175(.A1(new_n9181_), .A2(new_n9086_), .Z(new_n9182_));
  NAND2_X1   g08176(.A1(new_n9164_), .A2(new_n9173_), .ZN(new_n9183_));
  NAND2_X1   g08177(.A1(new_n9156_), .A2(new_n9117_), .ZN(new_n9184_));
  NAND3_X1   g08178(.A1(new_n9184_), .A2(new_n9183_), .A3(new_n9182_), .ZN(new_n9185_));
  AOI21_X1   g08179(.A1(new_n9175_), .A2(new_n9185_), .B(new_n9064_), .ZN(new_n9186_));
  INV_X1     g08180(.I(new_n9186_), .ZN(new_n9187_));
  NAND3_X1   g08181(.A1(new_n9175_), .A2(new_n9185_), .A3(new_n9064_), .ZN(new_n9188_));
  AOI22_X1   g08182(.A1(new_n9020_), .A2(new_n9024_), .B1(new_n9187_), .B2(new_n9188_), .ZN(new_n9189_));
  AOI21_X1   g08183(.A1(new_n9023_), .A2(new_n9022_), .B(new_n9021_), .ZN(new_n9190_));
  NOR3_X1    g08184(.A1(new_n8994_), .A2(new_n9019_), .A3(new_n8911_), .ZN(new_n9191_));
  INV_X1     g08185(.I(new_n9188_), .ZN(new_n9192_));
  NOR4_X1    g08186(.A1(new_n9191_), .A2(new_n9190_), .A3(new_n9192_), .A4(new_n9186_), .ZN(new_n9193_));
  INV_X1     g08187(.I(\A[315] ), .ZN(new_n9194_));
  NOR2_X1    g08188(.A1(new_n9194_), .A2(\A[314] ), .ZN(new_n9195_));
  INV_X1     g08189(.I(\A[314] ), .ZN(new_n9196_));
  NOR2_X1    g08190(.A1(new_n9196_), .A2(\A[315] ), .ZN(new_n9197_));
  OAI21_X1   g08191(.A1(new_n9195_), .A2(new_n9197_), .B(\A[313] ), .ZN(new_n9198_));
  INV_X1     g08192(.I(\A[313] ), .ZN(new_n9199_));
  NAND2_X1   g08193(.A1(\A[314] ), .A2(\A[315] ), .ZN(new_n9200_));
  INV_X1     g08194(.I(new_n9200_), .ZN(new_n9201_));
  NOR2_X1    g08195(.A1(\A[314] ), .A2(\A[315] ), .ZN(new_n9202_));
  OAI21_X1   g08196(.A1(new_n9201_), .A2(new_n9202_), .B(new_n9199_), .ZN(new_n9203_));
  NAND2_X1   g08197(.A1(new_n9198_), .A2(new_n9203_), .ZN(new_n9204_));
  INV_X1     g08198(.I(\A[318] ), .ZN(new_n9205_));
  NOR2_X1    g08199(.A1(new_n9205_), .A2(\A[317] ), .ZN(new_n9206_));
  INV_X1     g08200(.I(\A[317] ), .ZN(new_n9207_));
  NOR2_X1    g08201(.A1(new_n9207_), .A2(\A[318] ), .ZN(new_n9208_));
  OAI21_X1   g08202(.A1(new_n9206_), .A2(new_n9208_), .B(\A[316] ), .ZN(new_n9209_));
  INV_X1     g08203(.I(\A[316] ), .ZN(new_n9210_));
  NAND2_X1   g08204(.A1(\A[317] ), .A2(\A[318] ), .ZN(new_n9211_));
  INV_X1     g08205(.I(new_n9211_), .ZN(new_n9212_));
  NOR2_X1    g08206(.A1(\A[317] ), .A2(\A[318] ), .ZN(new_n9213_));
  OAI21_X1   g08207(.A1(new_n9212_), .A2(new_n9213_), .B(new_n9210_), .ZN(new_n9214_));
  NAND2_X1   g08208(.A1(new_n9209_), .A2(new_n9214_), .ZN(new_n9215_));
  AOI21_X1   g08209(.A1(\A[314] ), .A2(\A[315] ), .B(\A[313] ), .ZN(new_n9216_));
  AOI21_X1   g08210(.A1(\A[317] ), .A2(\A[318] ), .B(\A[316] ), .ZN(new_n9217_));
  OAI22_X1   g08211(.A1(new_n9202_), .A2(new_n9216_), .B1(new_n9217_), .B2(new_n9213_), .ZN(new_n9218_));
  INV_X1     g08212(.I(new_n9218_), .ZN(new_n9219_));
  NAND3_X1   g08213(.A1(new_n9204_), .A2(new_n9215_), .A3(new_n9219_), .ZN(new_n9220_));
  INV_X1     g08214(.I(\A[307] ), .ZN(new_n9221_));
  INV_X1     g08215(.I(\A[308] ), .ZN(new_n9222_));
  NAND2_X1   g08216(.A1(new_n9222_), .A2(\A[309] ), .ZN(new_n9223_));
  INV_X1     g08217(.I(\A[309] ), .ZN(new_n9224_));
  NAND2_X1   g08218(.A1(new_n9224_), .A2(\A[308] ), .ZN(new_n9225_));
  AOI21_X1   g08219(.A1(new_n9223_), .A2(new_n9225_), .B(new_n9221_), .ZN(new_n9226_));
  NAND2_X1   g08220(.A1(\A[308] ), .A2(\A[309] ), .ZN(new_n9227_));
  NOR2_X1    g08221(.A1(\A[308] ), .A2(\A[309] ), .ZN(new_n9228_));
  INV_X1     g08222(.I(new_n9228_), .ZN(new_n9229_));
  AOI21_X1   g08223(.A1(new_n9229_), .A2(new_n9227_), .B(\A[307] ), .ZN(new_n9230_));
  NOR2_X1    g08224(.A1(new_n9230_), .A2(new_n9226_), .ZN(new_n9231_));
  INV_X1     g08225(.I(\A[310] ), .ZN(new_n9232_));
  INV_X1     g08226(.I(\A[311] ), .ZN(new_n9233_));
  NAND2_X1   g08227(.A1(new_n9233_), .A2(\A[312] ), .ZN(new_n9234_));
  INV_X1     g08228(.I(\A[312] ), .ZN(new_n9235_));
  NAND2_X1   g08229(.A1(new_n9235_), .A2(\A[311] ), .ZN(new_n9236_));
  AOI21_X1   g08230(.A1(new_n9234_), .A2(new_n9236_), .B(new_n9232_), .ZN(new_n9237_));
  NAND2_X1   g08231(.A1(\A[311] ), .A2(\A[312] ), .ZN(new_n9238_));
  NOR2_X1    g08232(.A1(\A[311] ), .A2(\A[312] ), .ZN(new_n9239_));
  INV_X1     g08233(.I(new_n9239_), .ZN(new_n9240_));
  AOI21_X1   g08234(.A1(new_n9240_), .A2(new_n9238_), .B(\A[310] ), .ZN(new_n9241_));
  NOR2_X1    g08235(.A1(new_n9241_), .A2(new_n9237_), .ZN(new_n9242_));
  AOI21_X1   g08236(.A1(\A[308] ), .A2(\A[309] ), .B(\A[307] ), .ZN(new_n9243_));
  AOI21_X1   g08237(.A1(\A[311] ), .A2(\A[312] ), .B(\A[310] ), .ZN(new_n9244_));
  OAI22_X1   g08238(.A1(new_n9228_), .A2(new_n9243_), .B1(new_n9244_), .B2(new_n9239_), .ZN(new_n9245_));
  NOR3_X1    g08239(.A1(new_n9231_), .A2(new_n9242_), .A3(new_n9245_), .ZN(new_n9246_));
  NAND2_X1   g08240(.A1(new_n9246_), .A2(new_n9220_), .ZN(new_n9247_));
  NAND2_X1   g08241(.A1(new_n9196_), .A2(\A[315] ), .ZN(new_n9248_));
  NAND2_X1   g08242(.A1(new_n9194_), .A2(\A[314] ), .ZN(new_n9249_));
  AOI21_X1   g08243(.A1(new_n9248_), .A2(new_n9249_), .B(new_n9199_), .ZN(new_n9250_));
  INV_X1     g08244(.I(new_n9202_), .ZN(new_n9251_));
  AOI21_X1   g08245(.A1(new_n9251_), .A2(new_n9200_), .B(\A[313] ), .ZN(new_n9252_));
  NOR2_X1    g08246(.A1(new_n9252_), .A2(new_n9250_), .ZN(new_n9253_));
  NAND2_X1   g08247(.A1(new_n9207_), .A2(\A[318] ), .ZN(new_n9254_));
  NAND2_X1   g08248(.A1(new_n9205_), .A2(\A[317] ), .ZN(new_n9255_));
  AOI21_X1   g08249(.A1(new_n9254_), .A2(new_n9255_), .B(new_n9210_), .ZN(new_n9256_));
  INV_X1     g08250(.I(new_n9213_), .ZN(new_n9257_));
  AOI21_X1   g08251(.A1(new_n9257_), .A2(new_n9211_), .B(\A[316] ), .ZN(new_n9258_));
  NOR2_X1    g08252(.A1(new_n9258_), .A2(new_n9256_), .ZN(new_n9259_));
  NOR3_X1    g08253(.A1(new_n9253_), .A2(new_n9259_), .A3(new_n9218_), .ZN(new_n9260_));
  NOR2_X1    g08254(.A1(new_n9224_), .A2(\A[308] ), .ZN(new_n9261_));
  NOR2_X1    g08255(.A1(new_n9222_), .A2(\A[309] ), .ZN(new_n9262_));
  OAI21_X1   g08256(.A1(new_n9261_), .A2(new_n9262_), .B(\A[307] ), .ZN(new_n9263_));
  INV_X1     g08257(.I(new_n9227_), .ZN(new_n9264_));
  OAI21_X1   g08258(.A1(new_n9264_), .A2(new_n9228_), .B(new_n9221_), .ZN(new_n9265_));
  NAND2_X1   g08259(.A1(new_n9263_), .A2(new_n9265_), .ZN(new_n9266_));
  NOR2_X1    g08260(.A1(new_n9235_), .A2(\A[311] ), .ZN(new_n9267_));
  NOR2_X1    g08261(.A1(new_n9233_), .A2(\A[312] ), .ZN(new_n9268_));
  OAI21_X1   g08262(.A1(new_n9267_), .A2(new_n9268_), .B(\A[310] ), .ZN(new_n9269_));
  INV_X1     g08263(.I(new_n9238_), .ZN(new_n9270_));
  OAI21_X1   g08264(.A1(new_n9270_), .A2(new_n9239_), .B(new_n9232_), .ZN(new_n9271_));
  NAND2_X1   g08265(.A1(new_n9269_), .A2(new_n9271_), .ZN(new_n9272_));
  NOR2_X1    g08266(.A1(new_n9243_), .A2(new_n9228_), .ZN(new_n9273_));
  NOR2_X1    g08267(.A1(new_n9244_), .A2(new_n9239_), .ZN(new_n9274_));
  NOR2_X1    g08268(.A1(new_n9273_), .A2(new_n9274_), .ZN(new_n9275_));
  NAND3_X1   g08269(.A1(new_n9266_), .A2(new_n9272_), .A3(new_n9275_), .ZN(new_n9276_));
  NAND2_X1   g08270(.A1(new_n9260_), .A2(new_n9276_), .ZN(new_n9277_));
  NAND2_X1   g08271(.A1(new_n9247_), .A2(new_n9277_), .ZN(new_n9278_));
  INV_X1     g08272(.I(\A[303] ), .ZN(new_n9279_));
  NOR2_X1    g08273(.A1(new_n9279_), .A2(\A[302] ), .ZN(new_n9280_));
  INV_X1     g08274(.I(\A[302] ), .ZN(new_n9281_));
  NOR2_X1    g08275(.A1(new_n9281_), .A2(\A[303] ), .ZN(new_n9282_));
  OAI21_X1   g08276(.A1(new_n9280_), .A2(new_n9282_), .B(\A[301] ), .ZN(new_n9283_));
  INV_X1     g08277(.I(\A[301] ), .ZN(new_n9284_));
  NAND2_X1   g08278(.A1(\A[302] ), .A2(\A[303] ), .ZN(new_n9285_));
  INV_X1     g08279(.I(new_n9285_), .ZN(new_n9286_));
  NOR2_X1    g08280(.A1(\A[302] ), .A2(\A[303] ), .ZN(new_n9287_));
  OAI21_X1   g08281(.A1(new_n9286_), .A2(new_n9287_), .B(new_n9284_), .ZN(new_n9288_));
  NAND2_X1   g08282(.A1(new_n9283_), .A2(new_n9288_), .ZN(new_n9289_));
  INV_X1     g08283(.I(\A[306] ), .ZN(new_n9290_));
  NOR2_X1    g08284(.A1(new_n9290_), .A2(\A[305] ), .ZN(new_n9291_));
  INV_X1     g08285(.I(\A[305] ), .ZN(new_n9292_));
  NOR2_X1    g08286(.A1(new_n9292_), .A2(\A[306] ), .ZN(new_n9293_));
  OAI21_X1   g08287(.A1(new_n9291_), .A2(new_n9293_), .B(\A[304] ), .ZN(new_n9294_));
  INV_X1     g08288(.I(\A[304] ), .ZN(new_n9295_));
  NAND2_X1   g08289(.A1(\A[305] ), .A2(\A[306] ), .ZN(new_n9296_));
  INV_X1     g08290(.I(new_n9296_), .ZN(new_n9297_));
  NOR2_X1    g08291(.A1(\A[305] ), .A2(\A[306] ), .ZN(new_n9298_));
  OAI21_X1   g08292(.A1(new_n9297_), .A2(new_n9298_), .B(new_n9295_), .ZN(new_n9299_));
  NAND2_X1   g08293(.A1(new_n9294_), .A2(new_n9299_), .ZN(new_n9300_));
  AOI21_X1   g08294(.A1(\A[302] ), .A2(\A[303] ), .B(\A[301] ), .ZN(new_n9301_));
  AOI21_X1   g08295(.A1(\A[305] ), .A2(\A[306] ), .B(\A[304] ), .ZN(new_n9302_));
  OAI22_X1   g08296(.A1(new_n9287_), .A2(new_n9301_), .B1(new_n9302_), .B2(new_n9298_), .ZN(new_n9303_));
  INV_X1     g08297(.I(new_n9303_), .ZN(new_n9304_));
  NAND3_X1   g08298(.A1(new_n9289_), .A2(new_n9300_), .A3(new_n9304_), .ZN(new_n9305_));
  INV_X1     g08299(.I(\A[295] ), .ZN(new_n9306_));
  INV_X1     g08300(.I(\A[296] ), .ZN(new_n9307_));
  NAND2_X1   g08301(.A1(new_n9307_), .A2(\A[297] ), .ZN(new_n9308_));
  INV_X1     g08302(.I(\A[297] ), .ZN(new_n9309_));
  NAND2_X1   g08303(.A1(new_n9309_), .A2(\A[296] ), .ZN(new_n9310_));
  AOI21_X1   g08304(.A1(new_n9308_), .A2(new_n9310_), .B(new_n9306_), .ZN(new_n9311_));
  NAND2_X1   g08305(.A1(\A[296] ), .A2(\A[297] ), .ZN(new_n9312_));
  NOR2_X1    g08306(.A1(\A[296] ), .A2(\A[297] ), .ZN(new_n9313_));
  INV_X1     g08307(.I(new_n9313_), .ZN(new_n9314_));
  AOI21_X1   g08308(.A1(new_n9314_), .A2(new_n9312_), .B(\A[295] ), .ZN(new_n9315_));
  NOR2_X1    g08309(.A1(new_n9315_), .A2(new_n9311_), .ZN(new_n9316_));
  INV_X1     g08310(.I(\A[298] ), .ZN(new_n9317_));
  INV_X1     g08311(.I(\A[299] ), .ZN(new_n9318_));
  NAND2_X1   g08312(.A1(new_n9318_), .A2(\A[300] ), .ZN(new_n9319_));
  INV_X1     g08313(.I(\A[300] ), .ZN(new_n9320_));
  NAND2_X1   g08314(.A1(new_n9320_), .A2(\A[299] ), .ZN(new_n9321_));
  AOI21_X1   g08315(.A1(new_n9319_), .A2(new_n9321_), .B(new_n9317_), .ZN(new_n9322_));
  NAND2_X1   g08316(.A1(\A[299] ), .A2(\A[300] ), .ZN(new_n9323_));
  NOR2_X1    g08317(.A1(\A[299] ), .A2(\A[300] ), .ZN(new_n9324_));
  INV_X1     g08318(.I(new_n9324_), .ZN(new_n9325_));
  AOI21_X1   g08319(.A1(new_n9325_), .A2(new_n9323_), .B(\A[298] ), .ZN(new_n9326_));
  NOR2_X1    g08320(.A1(new_n9326_), .A2(new_n9322_), .ZN(new_n9327_));
  AOI21_X1   g08321(.A1(\A[296] ), .A2(\A[297] ), .B(\A[295] ), .ZN(new_n9328_));
  AOI21_X1   g08322(.A1(\A[299] ), .A2(\A[300] ), .B(\A[298] ), .ZN(new_n9329_));
  OAI22_X1   g08323(.A1(new_n9313_), .A2(new_n9328_), .B1(new_n9329_), .B2(new_n9324_), .ZN(new_n9330_));
  NOR3_X1    g08324(.A1(new_n9316_), .A2(new_n9327_), .A3(new_n9330_), .ZN(new_n9331_));
  NAND2_X1   g08325(.A1(new_n9331_), .A2(new_n9305_), .ZN(new_n9332_));
  NAND2_X1   g08326(.A1(new_n9281_), .A2(\A[303] ), .ZN(new_n9333_));
  NAND2_X1   g08327(.A1(new_n9279_), .A2(\A[302] ), .ZN(new_n9334_));
  AOI21_X1   g08328(.A1(new_n9333_), .A2(new_n9334_), .B(new_n9284_), .ZN(new_n9335_));
  INV_X1     g08329(.I(new_n9287_), .ZN(new_n9336_));
  AOI21_X1   g08330(.A1(new_n9336_), .A2(new_n9285_), .B(\A[301] ), .ZN(new_n9337_));
  NOR2_X1    g08331(.A1(new_n9337_), .A2(new_n9335_), .ZN(new_n9338_));
  NAND2_X1   g08332(.A1(new_n9292_), .A2(\A[306] ), .ZN(new_n9339_));
  NAND2_X1   g08333(.A1(new_n9290_), .A2(\A[305] ), .ZN(new_n9340_));
  AOI21_X1   g08334(.A1(new_n9339_), .A2(new_n9340_), .B(new_n9295_), .ZN(new_n9341_));
  INV_X1     g08335(.I(new_n9298_), .ZN(new_n9342_));
  AOI21_X1   g08336(.A1(new_n9342_), .A2(new_n9296_), .B(\A[304] ), .ZN(new_n9343_));
  NOR2_X1    g08337(.A1(new_n9343_), .A2(new_n9341_), .ZN(new_n9344_));
  NOR3_X1    g08338(.A1(new_n9338_), .A2(new_n9344_), .A3(new_n9303_), .ZN(new_n9345_));
  NOR2_X1    g08339(.A1(new_n9309_), .A2(\A[296] ), .ZN(new_n9346_));
  NOR2_X1    g08340(.A1(new_n9307_), .A2(\A[297] ), .ZN(new_n9347_));
  OAI21_X1   g08341(.A1(new_n9346_), .A2(new_n9347_), .B(\A[295] ), .ZN(new_n9348_));
  INV_X1     g08342(.I(new_n9312_), .ZN(new_n9349_));
  OAI21_X1   g08343(.A1(new_n9349_), .A2(new_n9313_), .B(new_n9306_), .ZN(new_n9350_));
  NAND2_X1   g08344(.A1(new_n9348_), .A2(new_n9350_), .ZN(new_n9351_));
  NOR2_X1    g08345(.A1(new_n9320_), .A2(\A[299] ), .ZN(new_n9352_));
  NOR2_X1    g08346(.A1(new_n9318_), .A2(\A[300] ), .ZN(new_n9353_));
  OAI21_X1   g08347(.A1(new_n9352_), .A2(new_n9353_), .B(\A[298] ), .ZN(new_n9354_));
  INV_X1     g08348(.I(new_n9323_), .ZN(new_n9355_));
  OAI21_X1   g08349(.A1(new_n9355_), .A2(new_n9324_), .B(new_n9317_), .ZN(new_n9356_));
  NAND2_X1   g08350(.A1(new_n9354_), .A2(new_n9356_), .ZN(new_n9357_));
  INV_X1     g08351(.I(new_n9330_), .ZN(new_n9358_));
  NAND3_X1   g08352(.A1(new_n9351_), .A2(new_n9357_), .A3(new_n9358_), .ZN(new_n9359_));
  NAND2_X1   g08353(.A1(new_n9345_), .A2(new_n9359_), .ZN(new_n9360_));
  NAND2_X1   g08354(.A1(new_n9332_), .A2(new_n9360_), .ZN(new_n9361_));
  NAND2_X1   g08355(.A1(new_n9278_), .A2(new_n9361_), .ZN(new_n9362_));
  NAND4_X1   g08356(.A1(new_n9247_), .A2(new_n9277_), .A3(new_n9332_), .A4(new_n9360_), .ZN(new_n9363_));
  NAND2_X1   g08357(.A1(new_n9362_), .A2(new_n9363_), .ZN(new_n9364_));
  INV_X1     g08358(.I(\A[289] ), .ZN(new_n9365_));
  INV_X1     g08359(.I(\A[290] ), .ZN(new_n9366_));
  NAND2_X1   g08360(.A1(new_n9366_), .A2(\A[291] ), .ZN(new_n9367_));
  INV_X1     g08361(.I(\A[291] ), .ZN(new_n9368_));
  NAND2_X1   g08362(.A1(new_n9368_), .A2(\A[290] ), .ZN(new_n9369_));
  AOI21_X1   g08363(.A1(new_n9367_), .A2(new_n9369_), .B(new_n9365_), .ZN(new_n9370_));
  NAND2_X1   g08364(.A1(\A[290] ), .A2(\A[291] ), .ZN(new_n9371_));
  NOR2_X1    g08365(.A1(\A[290] ), .A2(\A[291] ), .ZN(new_n9372_));
  INV_X1     g08366(.I(new_n9372_), .ZN(new_n9373_));
  AOI21_X1   g08367(.A1(new_n9373_), .A2(new_n9371_), .B(\A[289] ), .ZN(new_n9374_));
  NOR2_X1    g08368(.A1(new_n9374_), .A2(new_n9370_), .ZN(new_n9375_));
  INV_X1     g08369(.I(\A[292] ), .ZN(new_n9376_));
  INV_X1     g08370(.I(\A[293] ), .ZN(new_n9377_));
  NAND2_X1   g08371(.A1(new_n9377_), .A2(\A[294] ), .ZN(new_n9378_));
  INV_X1     g08372(.I(\A[294] ), .ZN(new_n9379_));
  NAND2_X1   g08373(.A1(new_n9379_), .A2(\A[293] ), .ZN(new_n9380_));
  AOI21_X1   g08374(.A1(new_n9378_), .A2(new_n9380_), .B(new_n9376_), .ZN(new_n9381_));
  NAND2_X1   g08375(.A1(\A[293] ), .A2(\A[294] ), .ZN(new_n9382_));
  NOR2_X1    g08376(.A1(\A[293] ), .A2(\A[294] ), .ZN(new_n9383_));
  INV_X1     g08377(.I(new_n9383_), .ZN(new_n9384_));
  AOI21_X1   g08378(.A1(new_n9384_), .A2(new_n9382_), .B(\A[292] ), .ZN(new_n9385_));
  NOR2_X1    g08379(.A1(new_n9385_), .A2(new_n9381_), .ZN(new_n9386_));
  AOI21_X1   g08380(.A1(\A[290] ), .A2(\A[291] ), .B(\A[289] ), .ZN(new_n9387_));
  AOI21_X1   g08381(.A1(\A[293] ), .A2(\A[294] ), .B(\A[292] ), .ZN(new_n9388_));
  OAI22_X1   g08382(.A1(new_n9372_), .A2(new_n9387_), .B1(new_n9388_), .B2(new_n9383_), .ZN(new_n9389_));
  NOR3_X1    g08383(.A1(new_n9375_), .A2(new_n9386_), .A3(new_n9389_), .ZN(new_n9390_));
  INV_X1     g08384(.I(\A[285] ), .ZN(new_n9391_));
  NOR2_X1    g08385(.A1(new_n9391_), .A2(\A[284] ), .ZN(new_n9392_));
  INV_X1     g08386(.I(\A[284] ), .ZN(new_n9393_));
  NOR2_X1    g08387(.A1(new_n9393_), .A2(\A[285] ), .ZN(new_n9394_));
  OAI21_X1   g08388(.A1(new_n9392_), .A2(new_n9394_), .B(\A[283] ), .ZN(new_n9395_));
  INV_X1     g08389(.I(\A[283] ), .ZN(new_n9396_));
  NAND2_X1   g08390(.A1(\A[284] ), .A2(\A[285] ), .ZN(new_n9397_));
  INV_X1     g08391(.I(new_n9397_), .ZN(new_n9398_));
  NOR2_X1    g08392(.A1(\A[284] ), .A2(\A[285] ), .ZN(new_n9399_));
  OAI21_X1   g08393(.A1(new_n9398_), .A2(new_n9399_), .B(new_n9396_), .ZN(new_n9400_));
  NAND2_X1   g08394(.A1(new_n9395_), .A2(new_n9400_), .ZN(new_n9401_));
  INV_X1     g08395(.I(\A[288] ), .ZN(new_n9402_));
  NOR2_X1    g08396(.A1(new_n9402_), .A2(\A[287] ), .ZN(new_n9403_));
  INV_X1     g08397(.I(\A[287] ), .ZN(new_n9404_));
  NOR2_X1    g08398(.A1(new_n9404_), .A2(\A[288] ), .ZN(new_n9405_));
  OAI21_X1   g08399(.A1(new_n9403_), .A2(new_n9405_), .B(\A[286] ), .ZN(new_n9406_));
  INV_X1     g08400(.I(\A[286] ), .ZN(new_n9407_));
  NAND2_X1   g08401(.A1(\A[287] ), .A2(\A[288] ), .ZN(new_n9408_));
  INV_X1     g08402(.I(new_n9408_), .ZN(new_n9409_));
  NOR2_X1    g08403(.A1(\A[287] ), .A2(\A[288] ), .ZN(new_n9410_));
  OAI21_X1   g08404(.A1(new_n9409_), .A2(new_n9410_), .B(new_n9407_), .ZN(new_n9411_));
  NAND2_X1   g08405(.A1(new_n9406_), .A2(new_n9411_), .ZN(new_n9412_));
  AOI21_X1   g08406(.A1(\A[284] ), .A2(\A[285] ), .B(\A[283] ), .ZN(new_n9413_));
  NOR2_X1    g08407(.A1(new_n9413_), .A2(new_n9399_), .ZN(new_n9414_));
  AOI21_X1   g08408(.A1(\A[287] ), .A2(\A[288] ), .B(\A[286] ), .ZN(new_n9415_));
  NOR2_X1    g08409(.A1(new_n9415_), .A2(new_n9410_), .ZN(new_n9416_));
  NOR2_X1    g08410(.A1(new_n9414_), .A2(new_n9416_), .ZN(new_n9417_));
  NAND3_X1   g08411(.A1(new_n9401_), .A2(new_n9412_), .A3(new_n9417_), .ZN(new_n9418_));
  NOR2_X1    g08412(.A1(new_n9390_), .A2(new_n9418_), .ZN(new_n9419_));
  NOR2_X1    g08413(.A1(new_n9368_), .A2(\A[290] ), .ZN(new_n9420_));
  NOR2_X1    g08414(.A1(new_n9366_), .A2(\A[291] ), .ZN(new_n9421_));
  OAI21_X1   g08415(.A1(new_n9420_), .A2(new_n9421_), .B(\A[289] ), .ZN(new_n9422_));
  INV_X1     g08416(.I(new_n9371_), .ZN(new_n9423_));
  OAI21_X1   g08417(.A1(new_n9423_), .A2(new_n9372_), .B(new_n9365_), .ZN(new_n9424_));
  NAND2_X1   g08418(.A1(new_n9422_), .A2(new_n9424_), .ZN(new_n9425_));
  NOR2_X1    g08419(.A1(new_n9379_), .A2(\A[293] ), .ZN(new_n9426_));
  NOR2_X1    g08420(.A1(new_n9377_), .A2(\A[294] ), .ZN(new_n9427_));
  OAI21_X1   g08421(.A1(new_n9426_), .A2(new_n9427_), .B(\A[292] ), .ZN(new_n9428_));
  INV_X1     g08422(.I(new_n9382_), .ZN(new_n9429_));
  OAI21_X1   g08423(.A1(new_n9429_), .A2(new_n9383_), .B(new_n9376_), .ZN(new_n9430_));
  NAND2_X1   g08424(.A1(new_n9428_), .A2(new_n9430_), .ZN(new_n9431_));
  NOR2_X1    g08425(.A1(new_n9387_), .A2(new_n9372_), .ZN(new_n9432_));
  NOR2_X1    g08426(.A1(new_n9388_), .A2(new_n9383_), .ZN(new_n9433_));
  NOR2_X1    g08427(.A1(new_n9432_), .A2(new_n9433_), .ZN(new_n9434_));
  NAND3_X1   g08428(.A1(new_n9425_), .A2(new_n9431_), .A3(new_n9434_), .ZN(new_n9435_));
  NAND2_X1   g08429(.A1(new_n9393_), .A2(\A[285] ), .ZN(new_n9436_));
  NAND2_X1   g08430(.A1(new_n9391_), .A2(\A[284] ), .ZN(new_n9437_));
  AOI21_X1   g08431(.A1(new_n9436_), .A2(new_n9437_), .B(new_n9396_), .ZN(new_n9438_));
  INV_X1     g08432(.I(new_n9399_), .ZN(new_n9439_));
  AOI21_X1   g08433(.A1(new_n9439_), .A2(new_n9397_), .B(\A[283] ), .ZN(new_n9440_));
  NOR2_X1    g08434(.A1(new_n9440_), .A2(new_n9438_), .ZN(new_n9441_));
  NAND2_X1   g08435(.A1(new_n9404_), .A2(\A[288] ), .ZN(new_n9442_));
  NAND2_X1   g08436(.A1(new_n9402_), .A2(\A[287] ), .ZN(new_n9443_));
  AOI21_X1   g08437(.A1(new_n9442_), .A2(new_n9443_), .B(new_n9407_), .ZN(new_n9444_));
  INV_X1     g08438(.I(new_n9410_), .ZN(new_n9445_));
  AOI21_X1   g08439(.A1(new_n9445_), .A2(new_n9408_), .B(\A[286] ), .ZN(new_n9446_));
  NOR2_X1    g08440(.A1(new_n9446_), .A2(new_n9444_), .ZN(new_n9447_));
  OAI22_X1   g08441(.A1(new_n9399_), .A2(new_n9413_), .B1(new_n9415_), .B2(new_n9410_), .ZN(new_n9448_));
  NOR3_X1    g08442(.A1(new_n9441_), .A2(new_n9447_), .A3(new_n9448_), .ZN(new_n9449_));
  NOR2_X1    g08443(.A1(new_n9449_), .A2(new_n9435_), .ZN(new_n9450_));
  INV_X1     g08444(.I(\A[277] ), .ZN(new_n9451_));
  INV_X1     g08445(.I(\A[278] ), .ZN(new_n9452_));
  NAND2_X1   g08446(.A1(new_n9452_), .A2(\A[279] ), .ZN(new_n9453_));
  INV_X1     g08447(.I(\A[279] ), .ZN(new_n9454_));
  NAND2_X1   g08448(.A1(new_n9454_), .A2(\A[278] ), .ZN(new_n9455_));
  AOI21_X1   g08449(.A1(new_n9453_), .A2(new_n9455_), .B(new_n9451_), .ZN(new_n9456_));
  NAND2_X1   g08450(.A1(\A[278] ), .A2(\A[279] ), .ZN(new_n9457_));
  NOR2_X1    g08451(.A1(\A[278] ), .A2(\A[279] ), .ZN(new_n9458_));
  INV_X1     g08452(.I(new_n9458_), .ZN(new_n9459_));
  AOI21_X1   g08453(.A1(new_n9459_), .A2(new_n9457_), .B(\A[277] ), .ZN(new_n9460_));
  NOR2_X1    g08454(.A1(new_n9460_), .A2(new_n9456_), .ZN(new_n9461_));
  INV_X1     g08455(.I(\A[280] ), .ZN(new_n9462_));
  INV_X1     g08456(.I(\A[281] ), .ZN(new_n9463_));
  NAND2_X1   g08457(.A1(new_n9463_), .A2(\A[282] ), .ZN(new_n9464_));
  INV_X1     g08458(.I(\A[282] ), .ZN(new_n9465_));
  NAND2_X1   g08459(.A1(new_n9465_), .A2(\A[281] ), .ZN(new_n9466_));
  AOI21_X1   g08460(.A1(new_n9464_), .A2(new_n9466_), .B(new_n9462_), .ZN(new_n9467_));
  NAND2_X1   g08461(.A1(\A[281] ), .A2(\A[282] ), .ZN(new_n9468_));
  NOR2_X1    g08462(.A1(\A[281] ), .A2(\A[282] ), .ZN(new_n9469_));
  INV_X1     g08463(.I(new_n9469_), .ZN(new_n9470_));
  AOI21_X1   g08464(.A1(new_n9470_), .A2(new_n9468_), .B(\A[280] ), .ZN(new_n9471_));
  NOR2_X1    g08465(.A1(new_n9471_), .A2(new_n9467_), .ZN(new_n9472_));
  AOI21_X1   g08466(.A1(\A[278] ), .A2(\A[279] ), .B(\A[277] ), .ZN(new_n9473_));
  AOI21_X1   g08467(.A1(\A[281] ), .A2(\A[282] ), .B(\A[280] ), .ZN(new_n9474_));
  OAI22_X1   g08468(.A1(new_n9458_), .A2(new_n9473_), .B1(new_n9474_), .B2(new_n9469_), .ZN(new_n9475_));
  NOR3_X1    g08469(.A1(new_n9461_), .A2(new_n9472_), .A3(new_n9475_), .ZN(new_n9476_));
  INV_X1     g08470(.I(\A[273] ), .ZN(new_n9477_));
  NOR2_X1    g08471(.A1(new_n9477_), .A2(\A[272] ), .ZN(new_n9478_));
  INV_X1     g08472(.I(\A[272] ), .ZN(new_n9479_));
  NOR2_X1    g08473(.A1(new_n9479_), .A2(\A[273] ), .ZN(new_n9480_));
  OAI21_X1   g08474(.A1(new_n9478_), .A2(new_n9480_), .B(\A[271] ), .ZN(new_n9481_));
  INV_X1     g08475(.I(\A[271] ), .ZN(new_n9482_));
  NAND2_X1   g08476(.A1(\A[272] ), .A2(\A[273] ), .ZN(new_n9483_));
  INV_X1     g08477(.I(new_n9483_), .ZN(new_n9484_));
  NOR2_X1    g08478(.A1(\A[272] ), .A2(\A[273] ), .ZN(new_n9485_));
  OAI21_X1   g08479(.A1(new_n9484_), .A2(new_n9485_), .B(new_n9482_), .ZN(new_n9486_));
  NAND2_X1   g08480(.A1(new_n9481_), .A2(new_n9486_), .ZN(new_n9487_));
  INV_X1     g08481(.I(\A[276] ), .ZN(new_n9488_));
  NOR2_X1    g08482(.A1(new_n9488_), .A2(\A[275] ), .ZN(new_n9489_));
  INV_X1     g08483(.I(\A[275] ), .ZN(new_n9490_));
  NOR2_X1    g08484(.A1(new_n9490_), .A2(\A[276] ), .ZN(new_n9491_));
  OAI21_X1   g08485(.A1(new_n9489_), .A2(new_n9491_), .B(\A[274] ), .ZN(new_n9492_));
  INV_X1     g08486(.I(\A[274] ), .ZN(new_n9493_));
  NAND2_X1   g08487(.A1(\A[275] ), .A2(\A[276] ), .ZN(new_n9494_));
  INV_X1     g08488(.I(new_n9494_), .ZN(new_n9495_));
  NOR2_X1    g08489(.A1(\A[275] ), .A2(\A[276] ), .ZN(new_n9496_));
  OAI21_X1   g08490(.A1(new_n9495_), .A2(new_n9496_), .B(new_n9493_), .ZN(new_n9497_));
  NAND2_X1   g08491(.A1(new_n9492_), .A2(new_n9497_), .ZN(new_n9498_));
  AOI21_X1   g08492(.A1(\A[272] ), .A2(\A[273] ), .B(\A[271] ), .ZN(new_n9499_));
  AOI21_X1   g08493(.A1(\A[275] ), .A2(\A[276] ), .B(\A[274] ), .ZN(new_n9500_));
  OAI22_X1   g08494(.A1(new_n9485_), .A2(new_n9499_), .B1(new_n9500_), .B2(new_n9496_), .ZN(new_n9501_));
  INV_X1     g08495(.I(new_n9501_), .ZN(new_n9502_));
  NAND3_X1   g08496(.A1(new_n9487_), .A2(new_n9498_), .A3(new_n9502_), .ZN(new_n9503_));
  NOR2_X1    g08497(.A1(new_n9476_), .A2(new_n9503_), .ZN(new_n9504_));
  NOR2_X1    g08498(.A1(new_n9454_), .A2(\A[278] ), .ZN(new_n9505_));
  NOR2_X1    g08499(.A1(new_n9452_), .A2(\A[279] ), .ZN(new_n9506_));
  OAI21_X1   g08500(.A1(new_n9505_), .A2(new_n9506_), .B(\A[277] ), .ZN(new_n9507_));
  INV_X1     g08501(.I(new_n9457_), .ZN(new_n9508_));
  OAI21_X1   g08502(.A1(new_n9508_), .A2(new_n9458_), .B(new_n9451_), .ZN(new_n9509_));
  NAND2_X1   g08503(.A1(new_n9507_), .A2(new_n9509_), .ZN(new_n9510_));
  NOR2_X1    g08504(.A1(new_n9465_), .A2(\A[281] ), .ZN(new_n9511_));
  NOR2_X1    g08505(.A1(new_n9463_), .A2(\A[282] ), .ZN(new_n9512_));
  OAI21_X1   g08506(.A1(new_n9511_), .A2(new_n9512_), .B(\A[280] ), .ZN(new_n9513_));
  INV_X1     g08507(.I(new_n9468_), .ZN(new_n9514_));
  OAI21_X1   g08508(.A1(new_n9514_), .A2(new_n9469_), .B(new_n9462_), .ZN(new_n9515_));
  NAND2_X1   g08509(.A1(new_n9513_), .A2(new_n9515_), .ZN(new_n9516_));
  NOR2_X1    g08510(.A1(new_n9473_), .A2(new_n9458_), .ZN(new_n9517_));
  NOR2_X1    g08511(.A1(new_n9474_), .A2(new_n9469_), .ZN(new_n9518_));
  NOR2_X1    g08512(.A1(new_n9517_), .A2(new_n9518_), .ZN(new_n9519_));
  NAND3_X1   g08513(.A1(new_n9510_), .A2(new_n9516_), .A3(new_n9519_), .ZN(new_n9520_));
  NAND2_X1   g08514(.A1(new_n9479_), .A2(\A[273] ), .ZN(new_n9521_));
  NAND2_X1   g08515(.A1(new_n9477_), .A2(\A[272] ), .ZN(new_n9522_));
  AOI21_X1   g08516(.A1(new_n9521_), .A2(new_n9522_), .B(new_n9482_), .ZN(new_n9523_));
  INV_X1     g08517(.I(new_n9485_), .ZN(new_n9524_));
  AOI21_X1   g08518(.A1(new_n9524_), .A2(new_n9483_), .B(\A[271] ), .ZN(new_n9525_));
  NOR2_X1    g08519(.A1(new_n9525_), .A2(new_n9523_), .ZN(new_n9526_));
  NAND2_X1   g08520(.A1(new_n9490_), .A2(\A[276] ), .ZN(new_n9527_));
  NAND2_X1   g08521(.A1(new_n9488_), .A2(\A[275] ), .ZN(new_n9528_));
  AOI21_X1   g08522(.A1(new_n9527_), .A2(new_n9528_), .B(new_n9493_), .ZN(new_n9529_));
  INV_X1     g08523(.I(new_n9496_), .ZN(new_n9530_));
  AOI21_X1   g08524(.A1(new_n9530_), .A2(new_n9494_), .B(\A[274] ), .ZN(new_n9531_));
  NOR2_X1    g08525(.A1(new_n9531_), .A2(new_n9529_), .ZN(new_n9532_));
  NOR3_X1    g08526(.A1(new_n9526_), .A2(new_n9532_), .A3(new_n9501_), .ZN(new_n9533_));
  NOR2_X1    g08527(.A1(new_n9533_), .A2(new_n9520_), .ZN(new_n9534_));
  OAI22_X1   g08528(.A1(new_n9419_), .A2(new_n9450_), .B1(new_n9504_), .B2(new_n9534_), .ZN(new_n9535_));
  NAND2_X1   g08529(.A1(new_n9449_), .A2(new_n9435_), .ZN(new_n9536_));
  NAND2_X1   g08530(.A1(new_n9390_), .A2(new_n9418_), .ZN(new_n9537_));
  NAND2_X1   g08531(.A1(new_n9533_), .A2(new_n9520_), .ZN(new_n9538_));
  NAND2_X1   g08532(.A1(new_n9476_), .A2(new_n9503_), .ZN(new_n9539_));
  NAND4_X1   g08533(.A1(new_n9536_), .A2(new_n9537_), .A3(new_n9538_), .A4(new_n9539_), .ZN(new_n9540_));
  NAND2_X1   g08534(.A1(new_n9535_), .A2(new_n9540_), .ZN(new_n9541_));
  NAND2_X1   g08535(.A1(new_n9364_), .A2(new_n9541_), .ZN(new_n9542_));
  NOR2_X1    g08536(.A1(new_n9364_), .A2(new_n9541_), .ZN(new_n9543_));
  INV_X1     g08537(.I(new_n9543_), .ZN(new_n9544_));
  NAND2_X1   g08538(.A1(new_n9544_), .A2(new_n9542_), .ZN(new_n9545_));
  OAI21_X1   g08539(.A1(new_n9189_), .A2(new_n9193_), .B(new_n9545_), .ZN(new_n9546_));
  NOR3_X1    g08540(.A1(new_n9189_), .A2(new_n9193_), .A3(new_n9545_), .ZN(new_n9547_));
  INV_X1     g08541(.I(new_n9547_), .ZN(new_n9548_));
  AOI22_X1   g08542(.A1(new_n8885_), .A2(new_n8882_), .B1(new_n9546_), .B2(new_n9548_), .ZN(new_n9549_));
  NAND4_X1   g08543(.A1(new_n8885_), .A2(new_n8882_), .A3(new_n9548_), .A4(new_n9546_), .ZN(new_n9550_));
  INV_X1     g08544(.I(new_n9550_), .ZN(new_n9551_));
  INV_X1     g08545(.I(\A[201] ), .ZN(new_n9552_));
  NOR2_X1    g08546(.A1(new_n9552_), .A2(\A[200] ), .ZN(new_n9553_));
  INV_X1     g08547(.I(\A[200] ), .ZN(new_n9554_));
  NOR2_X1    g08548(.A1(new_n9554_), .A2(\A[201] ), .ZN(new_n9555_));
  OAI21_X1   g08549(.A1(new_n9553_), .A2(new_n9555_), .B(\A[199] ), .ZN(new_n9556_));
  INV_X1     g08550(.I(\A[199] ), .ZN(new_n9557_));
  NOR2_X1    g08551(.A1(\A[200] ), .A2(\A[201] ), .ZN(new_n9558_));
  AND2_X2    g08552(.A1(\A[200] ), .A2(\A[201] ), .Z(new_n9559_));
  OAI21_X1   g08553(.A1(new_n9559_), .A2(new_n9558_), .B(new_n9557_), .ZN(new_n9560_));
  NAND2_X1   g08554(.A1(new_n9556_), .A2(new_n9560_), .ZN(new_n9561_));
  INV_X1     g08555(.I(\A[204] ), .ZN(new_n9562_));
  NOR2_X1    g08556(.A1(new_n9562_), .A2(\A[203] ), .ZN(new_n9563_));
  INV_X1     g08557(.I(\A[203] ), .ZN(new_n9564_));
  NOR2_X1    g08558(.A1(new_n9564_), .A2(\A[204] ), .ZN(new_n9565_));
  OAI21_X1   g08559(.A1(new_n9563_), .A2(new_n9565_), .B(\A[202] ), .ZN(new_n9566_));
  INV_X1     g08560(.I(\A[202] ), .ZN(new_n9567_));
  NAND2_X1   g08561(.A1(\A[203] ), .A2(\A[204] ), .ZN(new_n9568_));
  INV_X1     g08562(.I(new_n9568_), .ZN(new_n9569_));
  NOR2_X1    g08563(.A1(\A[203] ), .A2(\A[204] ), .ZN(new_n9570_));
  OAI21_X1   g08564(.A1(new_n9569_), .A2(new_n9570_), .B(new_n9567_), .ZN(new_n9571_));
  NAND2_X1   g08565(.A1(new_n9566_), .A2(new_n9571_), .ZN(new_n9572_));
  AOI21_X1   g08566(.A1(\A[200] ), .A2(\A[201] ), .B(\A[199] ), .ZN(new_n9573_));
  OR2_X2     g08567(.A1(new_n9573_), .A2(new_n9558_), .Z(new_n9574_));
  OR2_X2     g08568(.A1(\A[203] ), .A2(\A[204] ), .Z(new_n9575_));
  OAI21_X1   g08569(.A1(new_n9569_), .A2(\A[202] ), .B(new_n9575_), .ZN(new_n9576_));
  NAND4_X1   g08570(.A1(new_n9572_), .A2(new_n9561_), .A3(new_n9574_), .A4(new_n9576_), .ZN(new_n9577_));
  AOI22_X1   g08571(.A1(new_n9566_), .A2(new_n9571_), .B1(new_n9556_), .B2(new_n9560_), .ZN(new_n9578_));
  NAND2_X1   g08572(.A1(new_n9554_), .A2(\A[201] ), .ZN(new_n9579_));
  NAND2_X1   g08573(.A1(new_n9552_), .A2(\A[200] ), .ZN(new_n9580_));
  AOI21_X1   g08574(.A1(new_n9579_), .A2(new_n9580_), .B(new_n9557_), .ZN(new_n9581_));
  INV_X1     g08575(.I(new_n9558_), .ZN(new_n9582_));
  NAND2_X1   g08576(.A1(\A[200] ), .A2(\A[201] ), .ZN(new_n9583_));
  AOI21_X1   g08577(.A1(new_n9582_), .A2(new_n9583_), .B(\A[199] ), .ZN(new_n9584_));
  NAND2_X1   g08578(.A1(new_n9564_), .A2(\A[204] ), .ZN(new_n9585_));
  NAND2_X1   g08579(.A1(new_n9562_), .A2(\A[203] ), .ZN(new_n9586_));
  AOI21_X1   g08580(.A1(new_n9585_), .A2(new_n9586_), .B(new_n9567_), .ZN(new_n9587_));
  AOI21_X1   g08581(.A1(new_n9575_), .A2(new_n9568_), .B(\A[202] ), .ZN(new_n9588_));
  NOR4_X1    g08582(.A1(new_n9581_), .A2(new_n9584_), .A3(new_n9587_), .A4(new_n9588_), .ZN(new_n9589_));
  NOR2_X1    g08583(.A1(new_n9578_), .A2(new_n9589_), .ZN(new_n9590_));
  NAND2_X1   g08584(.A1(new_n9590_), .A2(new_n9577_), .ZN(new_n9591_));
  INV_X1     g08585(.I(\A[208] ), .ZN(new_n9592_));
  INV_X1     g08586(.I(\A[209] ), .ZN(new_n9593_));
  NAND2_X1   g08587(.A1(new_n9593_), .A2(\A[210] ), .ZN(new_n9594_));
  INV_X1     g08588(.I(\A[210] ), .ZN(new_n9595_));
  NAND2_X1   g08589(.A1(new_n9595_), .A2(\A[209] ), .ZN(new_n9596_));
  AOI21_X1   g08590(.A1(new_n9594_), .A2(new_n9596_), .B(new_n9592_), .ZN(new_n9597_));
  NOR2_X1    g08591(.A1(\A[209] ), .A2(\A[210] ), .ZN(new_n9598_));
  INV_X1     g08592(.I(new_n9598_), .ZN(new_n9599_));
  NAND2_X1   g08593(.A1(\A[209] ), .A2(\A[210] ), .ZN(new_n9600_));
  AOI21_X1   g08594(.A1(new_n9599_), .A2(new_n9600_), .B(\A[208] ), .ZN(new_n9601_));
  NOR2_X1    g08595(.A1(new_n9601_), .A2(new_n9597_), .ZN(new_n9602_));
  INV_X1     g08596(.I(\A[205] ), .ZN(new_n9603_));
  INV_X1     g08597(.I(\A[206] ), .ZN(new_n9604_));
  NAND2_X1   g08598(.A1(new_n9604_), .A2(\A[207] ), .ZN(new_n9605_));
  INV_X1     g08599(.I(\A[207] ), .ZN(new_n9606_));
  NAND2_X1   g08600(.A1(new_n9606_), .A2(\A[206] ), .ZN(new_n9607_));
  AOI21_X1   g08601(.A1(new_n9605_), .A2(new_n9607_), .B(new_n9603_), .ZN(new_n9608_));
  OR2_X2     g08602(.A1(\A[206] ), .A2(\A[207] ), .Z(new_n9609_));
  NAND2_X1   g08603(.A1(\A[206] ), .A2(\A[207] ), .ZN(new_n9610_));
  AOI21_X1   g08604(.A1(new_n9609_), .A2(new_n9610_), .B(\A[205] ), .ZN(new_n9611_));
  NOR2_X1    g08605(.A1(new_n9608_), .A2(new_n9611_), .ZN(new_n9612_));
  NOR2_X1    g08606(.A1(new_n9602_), .A2(new_n9612_), .ZN(new_n9613_));
  NOR4_X1    g08607(.A1(new_n9597_), .A2(new_n9601_), .A3(new_n9608_), .A4(new_n9611_), .ZN(new_n9614_));
  AOI21_X1   g08608(.A1(\A[209] ), .A2(\A[210] ), .B(\A[208] ), .ZN(new_n9615_));
  NOR2_X1    g08609(.A1(new_n9615_), .A2(new_n9598_), .ZN(new_n9616_));
  NOR2_X1    g08610(.A1(\A[206] ), .A2(\A[207] ), .ZN(new_n9617_));
  AOI21_X1   g08611(.A1(\A[206] ), .A2(\A[207] ), .B(\A[205] ), .ZN(new_n9618_));
  NOR2_X1    g08612(.A1(new_n9618_), .A2(new_n9617_), .ZN(new_n9619_));
  NAND2_X1   g08613(.A1(new_n9616_), .A2(new_n9619_), .ZN(new_n9620_));
  INV_X1     g08614(.I(new_n9620_), .ZN(new_n9621_));
  NOR2_X1    g08615(.A1(new_n9613_), .A2(new_n9614_), .ZN(new_n9622_));
  INV_X1     g08616(.I(\A[211] ), .ZN(new_n9623_));
  INV_X1     g08617(.I(\A[212] ), .ZN(new_n9624_));
  NAND2_X1   g08618(.A1(new_n9624_), .A2(\A[213] ), .ZN(new_n9625_));
  INV_X1     g08619(.I(\A[213] ), .ZN(new_n9626_));
  NAND2_X1   g08620(.A1(new_n9626_), .A2(\A[212] ), .ZN(new_n9627_));
  AOI21_X1   g08621(.A1(new_n9625_), .A2(new_n9627_), .B(new_n9623_), .ZN(new_n9628_));
  NOR2_X1    g08622(.A1(\A[212] ), .A2(\A[213] ), .ZN(new_n9629_));
  INV_X1     g08623(.I(new_n9629_), .ZN(new_n9630_));
  NAND2_X1   g08624(.A1(\A[212] ), .A2(\A[213] ), .ZN(new_n9631_));
  AOI21_X1   g08625(.A1(new_n9630_), .A2(new_n9631_), .B(\A[211] ), .ZN(new_n9632_));
  NOR2_X1    g08626(.A1(new_n9632_), .A2(new_n9628_), .ZN(new_n9633_));
  INV_X1     g08627(.I(\A[214] ), .ZN(new_n9634_));
  INV_X1     g08628(.I(\A[215] ), .ZN(new_n9635_));
  NAND2_X1   g08629(.A1(new_n9635_), .A2(\A[216] ), .ZN(new_n9636_));
  INV_X1     g08630(.I(\A[216] ), .ZN(new_n9637_));
  NAND2_X1   g08631(.A1(new_n9637_), .A2(\A[215] ), .ZN(new_n9638_));
  AOI21_X1   g08632(.A1(new_n9636_), .A2(new_n9638_), .B(new_n9634_), .ZN(new_n9639_));
  NAND2_X1   g08633(.A1(\A[215] ), .A2(\A[216] ), .ZN(new_n9640_));
  NOR2_X1    g08634(.A1(\A[215] ), .A2(\A[216] ), .ZN(new_n9641_));
  INV_X1     g08635(.I(new_n9641_), .ZN(new_n9642_));
  AOI21_X1   g08636(.A1(new_n9642_), .A2(new_n9640_), .B(\A[214] ), .ZN(new_n9643_));
  NOR2_X1    g08637(.A1(new_n9643_), .A2(new_n9639_), .ZN(new_n9644_));
  AOI21_X1   g08638(.A1(\A[212] ), .A2(\A[213] ), .B(\A[211] ), .ZN(new_n9645_));
  AOI21_X1   g08639(.A1(\A[215] ), .A2(\A[216] ), .B(\A[214] ), .ZN(new_n9646_));
  OAI22_X1   g08640(.A1(new_n9629_), .A2(new_n9645_), .B1(new_n9646_), .B2(new_n9641_), .ZN(new_n9647_));
  NOR3_X1    g08641(.A1(new_n9633_), .A2(new_n9644_), .A3(new_n9647_), .ZN(new_n9648_));
  OAI22_X1   g08642(.A1(new_n9628_), .A2(new_n9632_), .B1(new_n9643_), .B2(new_n9639_), .ZN(new_n9649_));
  NOR2_X1    g08643(.A1(new_n9626_), .A2(\A[212] ), .ZN(new_n9650_));
  NOR2_X1    g08644(.A1(new_n9624_), .A2(\A[213] ), .ZN(new_n9651_));
  OAI21_X1   g08645(.A1(new_n9650_), .A2(new_n9651_), .B(\A[211] ), .ZN(new_n9652_));
  INV_X1     g08646(.I(new_n9631_), .ZN(new_n9653_));
  OAI21_X1   g08647(.A1(new_n9653_), .A2(new_n9629_), .B(new_n9623_), .ZN(new_n9654_));
  NOR2_X1    g08648(.A1(new_n9637_), .A2(\A[215] ), .ZN(new_n9655_));
  NOR2_X1    g08649(.A1(new_n9635_), .A2(\A[216] ), .ZN(new_n9656_));
  OAI21_X1   g08650(.A1(new_n9655_), .A2(new_n9656_), .B(\A[214] ), .ZN(new_n9657_));
  INV_X1     g08651(.I(new_n9640_), .ZN(new_n9658_));
  OAI21_X1   g08652(.A1(new_n9658_), .A2(new_n9641_), .B(new_n9634_), .ZN(new_n9659_));
  NAND4_X1   g08653(.A1(new_n9652_), .A2(new_n9659_), .A3(new_n9657_), .A4(new_n9654_), .ZN(new_n9660_));
  NAND2_X1   g08654(.A1(new_n9649_), .A2(new_n9660_), .ZN(new_n9661_));
  NOR2_X1    g08655(.A1(new_n9661_), .A2(new_n9648_), .ZN(new_n9662_));
  INV_X1     g08656(.I(\A[217] ), .ZN(new_n9663_));
  INV_X1     g08657(.I(\A[218] ), .ZN(new_n9664_));
  NAND2_X1   g08658(.A1(new_n9664_), .A2(\A[219] ), .ZN(new_n9665_));
  INV_X1     g08659(.I(\A[219] ), .ZN(new_n9666_));
  NAND2_X1   g08660(.A1(new_n9666_), .A2(\A[218] ), .ZN(new_n9667_));
  AOI21_X1   g08661(.A1(new_n9665_), .A2(new_n9667_), .B(new_n9663_), .ZN(new_n9668_));
  NOR2_X1    g08662(.A1(\A[218] ), .A2(\A[219] ), .ZN(new_n9669_));
  INV_X1     g08663(.I(new_n9669_), .ZN(new_n9670_));
  NAND2_X1   g08664(.A1(\A[218] ), .A2(\A[219] ), .ZN(new_n9671_));
  AOI21_X1   g08665(.A1(new_n9670_), .A2(new_n9671_), .B(\A[217] ), .ZN(new_n9672_));
  INV_X1     g08666(.I(\A[220] ), .ZN(new_n9673_));
  INV_X1     g08667(.I(\A[221] ), .ZN(new_n9674_));
  NAND2_X1   g08668(.A1(new_n9674_), .A2(\A[222] ), .ZN(new_n9675_));
  INV_X1     g08669(.I(\A[222] ), .ZN(new_n9676_));
  NAND2_X1   g08670(.A1(new_n9676_), .A2(\A[221] ), .ZN(new_n9677_));
  AOI21_X1   g08671(.A1(new_n9675_), .A2(new_n9677_), .B(new_n9673_), .ZN(new_n9678_));
  NOR2_X1    g08672(.A1(\A[221] ), .A2(\A[222] ), .ZN(new_n9679_));
  INV_X1     g08673(.I(new_n9679_), .ZN(new_n9680_));
  NAND2_X1   g08674(.A1(\A[221] ), .A2(\A[222] ), .ZN(new_n9681_));
  AOI21_X1   g08675(.A1(new_n9680_), .A2(new_n9681_), .B(\A[220] ), .ZN(new_n9682_));
  NOR4_X1    g08676(.A1(new_n9668_), .A2(new_n9672_), .A3(new_n9682_), .A4(new_n9678_), .ZN(new_n9683_));
  AOI21_X1   g08677(.A1(\A[221] ), .A2(\A[222] ), .B(\A[220] ), .ZN(new_n9684_));
  NOR2_X1    g08678(.A1(new_n9684_), .A2(new_n9679_), .ZN(new_n9685_));
  AOI21_X1   g08679(.A1(\A[218] ), .A2(\A[219] ), .B(\A[217] ), .ZN(new_n9686_));
  NOR2_X1    g08680(.A1(new_n9686_), .A2(new_n9669_), .ZN(new_n9687_));
  NAND2_X1   g08681(.A1(new_n9685_), .A2(new_n9687_), .ZN(new_n9688_));
  INV_X1     g08682(.I(new_n9688_), .ZN(new_n9689_));
  NAND2_X1   g08683(.A1(new_n9683_), .A2(new_n9689_), .ZN(new_n9690_));
  NOR2_X1    g08684(.A1(new_n9666_), .A2(\A[218] ), .ZN(new_n9691_));
  NOR2_X1    g08685(.A1(new_n9664_), .A2(\A[219] ), .ZN(new_n9692_));
  OAI21_X1   g08686(.A1(new_n9691_), .A2(new_n9692_), .B(\A[217] ), .ZN(new_n9693_));
  INV_X1     g08687(.I(new_n9671_), .ZN(new_n9694_));
  OAI21_X1   g08688(.A1(new_n9694_), .A2(new_n9669_), .B(new_n9663_), .ZN(new_n9695_));
  NOR2_X1    g08689(.A1(new_n9676_), .A2(\A[221] ), .ZN(new_n9696_));
  NOR2_X1    g08690(.A1(new_n9674_), .A2(\A[222] ), .ZN(new_n9697_));
  OAI21_X1   g08691(.A1(new_n9696_), .A2(new_n9697_), .B(\A[220] ), .ZN(new_n9698_));
  AND2_X2    g08692(.A1(\A[221] ), .A2(\A[222] ), .Z(new_n9699_));
  OAI21_X1   g08693(.A1(new_n9699_), .A2(new_n9679_), .B(new_n9673_), .ZN(new_n9700_));
  AOI22_X1   g08694(.A1(new_n9693_), .A2(new_n9695_), .B1(new_n9698_), .B2(new_n9700_), .ZN(new_n9701_));
  NOR2_X1    g08695(.A1(new_n9683_), .A2(new_n9701_), .ZN(new_n9702_));
  NAND2_X1   g08696(.A1(new_n9702_), .A2(new_n9690_), .ZN(new_n9703_));
  XOR2_X1    g08697(.A1(new_n9703_), .A2(new_n9662_), .Z(new_n9704_));
  NOR2_X1    g08698(.A1(new_n9704_), .A2(new_n9622_), .ZN(new_n9705_));
  NOR2_X1    g08699(.A1(new_n9595_), .A2(\A[209] ), .ZN(new_n9706_));
  NOR2_X1    g08700(.A1(new_n9593_), .A2(\A[210] ), .ZN(new_n9707_));
  OAI21_X1   g08701(.A1(new_n9706_), .A2(new_n9707_), .B(\A[208] ), .ZN(new_n9708_));
  INV_X1     g08702(.I(new_n9600_), .ZN(new_n9709_));
  OAI21_X1   g08703(.A1(new_n9709_), .A2(new_n9598_), .B(new_n9592_), .ZN(new_n9710_));
  NAND2_X1   g08704(.A1(new_n9708_), .A2(new_n9710_), .ZN(new_n9711_));
  NOR2_X1    g08705(.A1(new_n9606_), .A2(\A[206] ), .ZN(new_n9712_));
  NOR2_X1    g08706(.A1(new_n9604_), .A2(\A[207] ), .ZN(new_n9713_));
  OAI21_X1   g08707(.A1(new_n9712_), .A2(new_n9713_), .B(\A[205] ), .ZN(new_n9714_));
  AND2_X2    g08708(.A1(\A[206] ), .A2(\A[207] ), .Z(new_n9715_));
  OAI21_X1   g08709(.A1(new_n9715_), .A2(new_n9617_), .B(new_n9603_), .ZN(new_n9716_));
  NAND2_X1   g08710(.A1(new_n9714_), .A2(new_n9716_), .ZN(new_n9717_));
  NAND2_X1   g08711(.A1(new_n9711_), .A2(new_n9717_), .ZN(new_n9718_));
  NAND2_X1   g08712(.A1(new_n9602_), .A2(new_n9612_), .ZN(new_n9719_));
  NAND2_X1   g08713(.A1(new_n9719_), .A2(new_n9718_), .ZN(new_n9720_));
  NAND2_X1   g08714(.A1(new_n9652_), .A2(new_n9654_), .ZN(new_n9721_));
  NAND2_X1   g08715(.A1(new_n9657_), .A2(new_n9659_), .ZN(new_n9722_));
  INV_X1     g08716(.I(new_n9647_), .ZN(new_n9723_));
  NAND3_X1   g08717(.A1(new_n9722_), .A2(new_n9721_), .A3(new_n9723_), .ZN(new_n9724_));
  NAND3_X1   g08718(.A1(new_n9724_), .A2(new_n9649_), .A3(new_n9660_), .ZN(new_n9725_));
  XOR2_X1    g08719(.A1(new_n9703_), .A2(new_n9725_), .Z(new_n9726_));
  NOR2_X1    g08720(.A1(new_n9726_), .A2(new_n9720_), .ZN(new_n9727_));
  OAI21_X1   g08721(.A1(new_n9705_), .A2(new_n9727_), .B(new_n9591_), .ZN(new_n9728_));
  NOR2_X1    g08722(.A1(new_n9584_), .A2(new_n9581_), .ZN(new_n9729_));
  NOR2_X1    g08723(.A1(new_n9587_), .A2(new_n9588_), .ZN(new_n9730_));
  AOI21_X1   g08724(.A1(\A[203] ), .A2(\A[204] ), .B(\A[202] ), .ZN(new_n9731_));
  OAI22_X1   g08725(.A1(new_n9558_), .A2(new_n9573_), .B1(new_n9731_), .B2(new_n9570_), .ZN(new_n9732_));
  NOR3_X1    g08726(.A1(new_n9729_), .A2(new_n9730_), .A3(new_n9732_), .ZN(new_n9733_));
  OAI22_X1   g08727(.A1(new_n9581_), .A2(new_n9584_), .B1(new_n9587_), .B2(new_n9588_), .ZN(new_n9734_));
  NAND4_X1   g08728(.A1(new_n9556_), .A2(new_n9566_), .A3(new_n9571_), .A4(new_n9560_), .ZN(new_n9735_));
  NAND2_X1   g08729(.A1(new_n9734_), .A2(new_n9735_), .ZN(new_n9736_));
  NOR2_X1    g08730(.A1(new_n9736_), .A2(new_n9733_), .ZN(new_n9737_));
  NAND2_X1   g08731(.A1(new_n9726_), .A2(new_n9720_), .ZN(new_n9738_));
  NAND2_X1   g08732(.A1(new_n9704_), .A2(new_n9622_), .ZN(new_n9739_));
  NAND3_X1   g08733(.A1(new_n9739_), .A2(new_n9738_), .A3(new_n9737_), .ZN(new_n9740_));
  INV_X1     g08734(.I(\A[195] ), .ZN(new_n9741_));
  NOR2_X1    g08735(.A1(new_n9741_), .A2(\A[194] ), .ZN(new_n9742_));
  INV_X1     g08736(.I(\A[194] ), .ZN(new_n9743_));
  NOR2_X1    g08737(.A1(new_n9743_), .A2(\A[195] ), .ZN(new_n9744_));
  OAI21_X1   g08738(.A1(new_n9742_), .A2(new_n9744_), .B(\A[193] ), .ZN(new_n9745_));
  INV_X1     g08739(.I(\A[193] ), .ZN(new_n9746_));
  NAND2_X1   g08740(.A1(\A[194] ), .A2(\A[195] ), .ZN(new_n9747_));
  INV_X1     g08741(.I(new_n9747_), .ZN(new_n9748_));
  NOR2_X1    g08742(.A1(\A[194] ), .A2(\A[195] ), .ZN(new_n9749_));
  OAI21_X1   g08743(.A1(new_n9748_), .A2(new_n9749_), .B(new_n9746_), .ZN(new_n9750_));
  NAND2_X1   g08744(.A1(new_n9745_), .A2(new_n9750_), .ZN(new_n9751_));
  INV_X1     g08745(.I(\A[198] ), .ZN(new_n9752_));
  NOR2_X1    g08746(.A1(new_n9752_), .A2(\A[197] ), .ZN(new_n9753_));
  INV_X1     g08747(.I(\A[197] ), .ZN(new_n9754_));
  NOR2_X1    g08748(.A1(new_n9754_), .A2(\A[198] ), .ZN(new_n9755_));
  OAI21_X1   g08749(.A1(new_n9753_), .A2(new_n9755_), .B(\A[196] ), .ZN(new_n9756_));
  INV_X1     g08750(.I(\A[196] ), .ZN(new_n9757_));
  AND2_X2    g08751(.A1(\A[197] ), .A2(\A[198] ), .Z(new_n9758_));
  NOR2_X1    g08752(.A1(\A[197] ), .A2(\A[198] ), .ZN(new_n9759_));
  OAI21_X1   g08753(.A1(new_n9758_), .A2(new_n9759_), .B(new_n9757_), .ZN(new_n9760_));
  NAND2_X1   g08754(.A1(new_n9756_), .A2(new_n9760_), .ZN(new_n9761_));
  AOI21_X1   g08755(.A1(\A[194] ), .A2(\A[195] ), .B(\A[193] ), .ZN(new_n9762_));
  NOR2_X1    g08756(.A1(new_n9762_), .A2(new_n9749_), .ZN(new_n9763_));
  AOI21_X1   g08757(.A1(\A[197] ), .A2(\A[198] ), .B(\A[196] ), .ZN(new_n9764_));
  NOR2_X1    g08758(.A1(new_n9764_), .A2(new_n9759_), .ZN(new_n9765_));
  NOR2_X1    g08759(.A1(new_n9763_), .A2(new_n9765_), .ZN(new_n9766_));
  NAND3_X1   g08760(.A1(new_n9751_), .A2(new_n9761_), .A3(new_n9766_), .ZN(new_n9767_));
  INV_X1     g08761(.I(\A[187] ), .ZN(new_n9768_));
  INV_X1     g08762(.I(\A[188] ), .ZN(new_n9769_));
  NAND2_X1   g08763(.A1(new_n9769_), .A2(\A[189] ), .ZN(new_n9770_));
  INV_X1     g08764(.I(\A[189] ), .ZN(new_n9771_));
  NAND2_X1   g08765(.A1(new_n9771_), .A2(\A[188] ), .ZN(new_n9772_));
  AOI21_X1   g08766(.A1(new_n9770_), .A2(new_n9772_), .B(new_n9768_), .ZN(new_n9773_));
  NAND2_X1   g08767(.A1(\A[188] ), .A2(\A[189] ), .ZN(new_n9774_));
  NOR2_X1    g08768(.A1(\A[188] ), .A2(\A[189] ), .ZN(new_n9775_));
  INV_X1     g08769(.I(new_n9775_), .ZN(new_n9776_));
  AOI21_X1   g08770(.A1(new_n9776_), .A2(new_n9774_), .B(\A[187] ), .ZN(new_n9777_));
  NOR2_X1    g08771(.A1(new_n9777_), .A2(new_n9773_), .ZN(new_n9778_));
  INV_X1     g08772(.I(\A[190] ), .ZN(new_n9779_));
  INV_X1     g08773(.I(\A[191] ), .ZN(new_n9780_));
  NAND2_X1   g08774(.A1(new_n9780_), .A2(\A[192] ), .ZN(new_n9781_));
  INV_X1     g08775(.I(\A[192] ), .ZN(new_n9782_));
  NAND2_X1   g08776(.A1(new_n9782_), .A2(\A[191] ), .ZN(new_n9783_));
  AOI21_X1   g08777(.A1(new_n9781_), .A2(new_n9783_), .B(new_n9779_), .ZN(new_n9784_));
  NAND2_X1   g08778(.A1(\A[191] ), .A2(\A[192] ), .ZN(new_n9785_));
  NOR2_X1    g08779(.A1(\A[191] ), .A2(\A[192] ), .ZN(new_n9786_));
  INV_X1     g08780(.I(new_n9786_), .ZN(new_n9787_));
  AOI21_X1   g08781(.A1(new_n9787_), .A2(new_n9785_), .B(\A[190] ), .ZN(new_n9788_));
  NOR2_X1    g08782(.A1(new_n9788_), .A2(new_n9784_), .ZN(new_n9789_));
  AOI21_X1   g08783(.A1(\A[188] ), .A2(\A[189] ), .B(\A[187] ), .ZN(new_n9790_));
  AOI21_X1   g08784(.A1(\A[191] ), .A2(\A[192] ), .B(\A[190] ), .ZN(new_n9791_));
  OAI22_X1   g08785(.A1(new_n9775_), .A2(new_n9790_), .B1(new_n9791_), .B2(new_n9786_), .ZN(new_n9792_));
  NOR3_X1    g08786(.A1(new_n9778_), .A2(new_n9789_), .A3(new_n9792_), .ZN(new_n9793_));
  NAND2_X1   g08787(.A1(new_n9793_), .A2(new_n9767_), .ZN(new_n9794_));
  INV_X1     g08788(.I(new_n9767_), .ZN(new_n9795_));
  NOR2_X1    g08789(.A1(new_n9771_), .A2(\A[188] ), .ZN(new_n9796_));
  NOR2_X1    g08790(.A1(new_n9769_), .A2(\A[189] ), .ZN(new_n9797_));
  OAI21_X1   g08791(.A1(new_n9796_), .A2(new_n9797_), .B(\A[187] ), .ZN(new_n9798_));
  INV_X1     g08792(.I(new_n9774_), .ZN(new_n9799_));
  OAI21_X1   g08793(.A1(new_n9799_), .A2(new_n9775_), .B(new_n9768_), .ZN(new_n9800_));
  NAND2_X1   g08794(.A1(new_n9798_), .A2(new_n9800_), .ZN(new_n9801_));
  NOR2_X1    g08795(.A1(new_n9782_), .A2(\A[191] ), .ZN(new_n9802_));
  NOR2_X1    g08796(.A1(new_n9780_), .A2(\A[192] ), .ZN(new_n9803_));
  OAI21_X1   g08797(.A1(new_n9802_), .A2(new_n9803_), .B(\A[190] ), .ZN(new_n9804_));
  INV_X1     g08798(.I(new_n9785_), .ZN(new_n9805_));
  OAI21_X1   g08799(.A1(new_n9805_), .A2(new_n9786_), .B(new_n9779_), .ZN(new_n9806_));
  NAND2_X1   g08800(.A1(new_n9804_), .A2(new_n9806_), .ZN(new_n9807_));
  INV_X1     g08801(.I(new_n9792_), .ZN(new_n9808_));
  NAND3_X1   g08802(.A1(new_n9801_), .A2(new_n9807_), .A3(new_n9808_), .ZN(new_n9809_));
  NAND2_X1   g08803(.A1(new_n9795_), .A2(new_n9809_), .ZN(new_n9810_));
  INV_X1     g08804(.I(\A[183] ), .ZN(new_n9811_));
  NOR2_X1    g08805(.A1(new_n9811_), .A2(\A[182] ), .ZN(new_n9812_));
  INV_X1     g08806(.I(\A[182] ), .ZN(new_n9813_));
  NOR2_X1    g08807(.A1(new_n9813_), .A2(\A[183] ), .ZN(new_n9814_));
  OAI21_X1   g08808(.A1(new_n9812_), .A2(new_n9814_), .B(\A[181] ), .ZN(new_n9815_));
  INV_X1     g08809(.I(\A[181] ), .ZN(new_n9816_));
  NAND2_X1   g08810(.A1(\A[182] ), .A2(\A[183] ), .ZN(new_n9817_));
  INV_X1     g08811(.I(new_n9817_), .ZN(new_n9818_));
  NOR2_X1    g08812(.A1(\A[182] ), .A2(\A[183] ), .ZN(new_n9819_));
  OAI21_X1   g08813(.A1(new_n9818_), .A2(new_n9819_), .B(new_n9816_), .ZN(new_n9820_));
  NAND2_X1   g08814(.A1(new_n9815_), .A2(new_n9820_), .ZN(new_n9821_));
  INV_X1     g08815(.I(\A[186] ), .ZN(new_n9822_));
  NOR2_X1    g08816(.A1(new_n9822_), .A2(\A[185] ), .ZN(new_n9823_));
  INV_X1     g08817(.I(\A[185] ), .ZN(new_n9824_));
  NOR2_X1    g08818(.A1(new_n9824_), .A2(\A[186] ), .ZN(new_n9825_));
  OAI21_X1   g08819(.A1(new_n9823_), .A2(new_n9825_), .B(\A[184] ), .ZN(new_n9826_));
  INV_X1     g08820(.I(\A[184] ), .ZN(new_n9827_));
  NAND2_X1   g08821(.A1(\A[185] ), .A2(\A[186] ), .ZN(new_n9828_));
  INV_X1     g08822(.I(new_n9828_), .ZN(new_n9829_));
  NOR2_X1    g08823(.A1(\A[185] ), .A2(\A[186] ), .ZN(new_n9830_));
  OAI21_X1   g08824(.A1(new_n9829_), .A2(new_n9830_), .B(new_n9827_), .ZN(new_n9831_));
  NAND2_X1   g08825(.A1(new_n9826_), .A2(new_n9831_), .ZN(new_n9832_));
  AOI21_X1   g08826(.A1(\A[182] ), .A2(\A[183] ), .B(\A[181] ), .ZN(new_n9833_));
  NOR2_X1    g08827(.A1(new_n9833_), .A2(new_n9819_), .ZN(new_n9834_));
  AOI21_X1   g08828(.A1(\A[185] ), .A2(\A[186] ), .B(\A[184] ), .ZN(new_n9835_));
  NOR2_X1    g08829(.A1(new_n9835_), .A2(new_n9830_), .ZN(new_n9836_));
  NOR2_X1    g08830(.A1(new_n9834_), .A2(new_n9836_), .ZN(new_n9837_));
  NAND3_X1   g08831(.A1(new_n9821_), .A2(new_n9832_), .A3(new_n9837_), .ZN(new_n9838_));
  INV_X1     g08832(.I(\A[175] ), .ZN(new_n9839_));
  INV_X1     g08833(.I(\A[176] ), .ZN(new_n9840_));
  NAND2_X1   g08834(.A1(new_n9840_), .A2(\A[177] ), .ZN(new_n9841_));
  INV_X1     g08835(.I(\A[177] ), .ZN(new_n9842_));
  NAND2_X1   g08836(.A1(new_n9842_), .A2(\A[176] ), .ZN(new_n9843_));
  AOI21_X1   g08837(.A1(new_n9841_), .A2(new_n9843_), .B(new_n9839_), .ZN(new_n9844_));
  NAND2_X1   g08838(.A1(\A[176] ), .A2(\A[177] ), .ZN(new_n9845_));
  NOR2_X1    g08839(.A1(\A[176] ), .A2(\A[177] ), .ZN(new_n9846_));
  INV_X1     g08840(.I(new_n9846_), .ZN(new_n9847_));
  AOI21_X1   g08841(.A1(new_n9847_), .A2(new_n9845_), .B(\A[175] ), .ZN(new_n9848_));
  NOR2_X1    g08842(.A1(new_n9848_), .A2(new_n9844_), .ZN(new_n9849_));
  INV_X1     g08843(.I(\A[178] ), .ZN(new_n9850_));
  INV_X1     g08844(.I(\A[179] ), .ZN(new_n9851_));
  NAND2_X1   g08845(.A1(new_n9851_), .A2(\A[180] ), .ZN(new_n9852_));
  INV_X1     g08846(.I(\A[180] ), .ZN(new_n9853_));
  NAND2_X1   g08847(.A1(new_n9853_), .A2(\A[179] ), .ZN(new_n9854_));
  AOI21_X1   g08848(.A1(new_n9852_), .A2(new_n9854_), .B(new_n9850_), .ZN(new_n9855_));
  NAND2_X1   g08849(.A1(\A[179] ), .A2(\A[180] ), .ZN(new_n9856_));
  NOR2_X1    g08850(.A1(\A[179] ), .A2(\A[180] ), .ZN(new_n9857_));
  INV_X1     g08851(.I(new_n9857_), .ZN(new_n9858_));
  AOI21_X1   g08852(.A1(new_n9858_), .A2(new_n9856_), .B(\A[178] ), .ZN(new_n9859_));
  NOR2_X1    g08853(.A1(new_n9859_), .A2(new_n9855_), .ZN(new_n9860_));
  AOI21_X1   g08854(.A1(\A[176] ), .A2(\A[177] ), .B(\A[175] ), .ZN(new_n9861_));
  AOI21_X1   g08855(.A1(\A[179] ), .A2(\A[180] ), .B(\A[178] ), .ZN(new_n9862_));
  OAI22_X1   g08856(.A1(new_n9846_), .A2(new_n9861_), .B1(new_n9862_), .B2(new_n9857_), .ZN(new_n9863_));
  NOR3_X1    g08857(.A1(new_n9849_), .A2(new_n9860_), .A3(new_n9863_), .ZN(new_n9864_));
  NAND2_X1   g08858(.A1(new_n9864_), .A2(new_n9838_), .ZN(new_n9865_));
  NAND2_X1   g08859(.A1(new_n9813_), .A2(\A[183] ), .ZN(new_n9866_));
  NAND2_X1   g08860(.A1(new_n9811_), .A2(\A[182] ), .ZN(new_n9867_));
  AOI21_X1   g08861(.A1(new_n9866_), .A2(new_n9867_), .B(new_n9816_), .ZN(new_n9868_));
  INV_X1     g08862(.I(new_n9819_), .ZN(new_n9869_));
  AOI21_X1   g08863(.A1(new_n9869_), .A2(new_n9817_), .B(\A[181] ), .ZN(new_n9870_));
  NOR2_X1    g08864(.A1(new_n9870_), .A2(new_n9868_), .ZN(new_n9871_));
  NAND2_X1   g08865(.A1(new_n9824_), .A2(\A[186] ), .ZN(new_n9872_));
  NAND2_X1   g08866(.A1(new_n9822_), .A2(\A[185] ), .ZN(new_n9873_));
  AOI21_X1   g08867(.A1(new_n9872_), .A2(new_n9873_), .B(new_n9827_), .ZN(new_n9874_));
  INV_X1     g08868(.I(new_n9830_), .ZN(new_n9875_));
  AOI21_X1   g08869(.A1(new_n9875_), .A2(new_n9828_), .B(\A[184] ), .ZN(new_n9876_));
  NOR2_X1    g08870(.A1(new_n9876_), .A2(new_n9874_), .ZN(new_n9877_));
  OAI22_X1   g08871(.A1(new_n9819_), .A2(new_n9833_), .B1(new_n9835_), .B2(new_n9830_), .ZN(new_n9878_));
  NOR3_X1    g08872(.A1(new_n9871_), .A2(new_n9877_), .A3(new_n9878_), .ZN(new_n9879_));
  NOR2_X1    g08873(.A1(new_n9842_), .A2(\A[176] ), .ZN(new_n9880_));
  NOR2_X1    g08874(.A1(new_n9840_), .A2(\A[177] ), .ZN(new_n9881_));
  OAI21_X1   g08875(.A1(new_n9880_), .A2(new_n9881_), .B(\A[175] ), .ZN(new_n9882_));
  INV_X1     g08876(.I(new_n9845_), .ZN(new_n9883_));
  OAI21_X1   g08877(.A1(new_n9883_), .A2(new_n9846_), .B(new_n9839_), .ZN(new_n9884_));
  NAND2_X1   g08878(.A1(new_n9882_), .A2(new_n9884_), .ZN(new_n9885_));
  NOR2_X1    g08879(.A1(new_n9853_), .A2(\A[179] ), .ZN(new_n9886_));
  NOR2_X1    g08880(.A1(new_n9851_), .A2(\A[180] ), .ZN(new_n9887_));
  OAI21_X1   g08881(.A1(new_n9886_), .A2(new_n9887_), .B(\A[178] ), .ZN(new_n9888_));
  INV_X1     g08882(.I(new_n9856_), .ZN(new_n9889_));
  OAI21_X1   g08883(.A1(new_n9889_), .A2(new_n9857_), .B(new_n9850_), .ZN(new_n9890_));
  NAND2_X1   g08884(.A1(new_n9888_), .A2(new_n9890_), .ZN(new_n9891_));
  INV_X1     g08885(.I(new_n9863_), .ZN(new_n9892_));
  NAND3_X1   g08886(.A1(new_n9885_), .A2(new_n9891_), .A3(new_n9892_), .ZN(new_n9893_));
  NAND2_X1   g08887(.A1(new_n9879_), .A2(new_n9893_), .ZN(new_n9894_));
  AOI22_X1   g08888(.A1(new_n9865_), .A2(new_n9894_), .B1(new_n9810_), .B2(new_n9794_), .ZN(new_n9895_));
  INV_X1     g08889(.I(new_n9794_), .ZN(new_n9896_));
  NOR2_X1    g08890(.A1(new_n9793_), .A2(new_n9767_), .ZN(new_n9897_));
  NOR2_X1    g08891(.A1(new_n9879_), .A2(new_n9893_), .ZN(new_n9898_));
  NOR2_X1    g08892(.A1(new_n9864_), .A2(new_n9838_), .ZN(new_n9899_));
  NOR4_X1    g08893(.A1(new_n9896_), .A2(new_n9898_), .A3(new_n9899_), .A4(new_n9897_), .ZN(new_n9900_));
  NOR2_X1    g08894(.A1(new_n9895_), .A2(new_n9900_), .ZN(new_n9901_));
  NAND3_X1   g08895(.A1(new_n9728_), .A2(new_n9740_), .A3(new_n9901_), .ZN(new_n9902_));
  INV_X1     g08896(.I(new_n9902_), .ZN(new_n9903_));
  AOI21_X1   g08897(.A1(new_n9728_), .A2(new_n9740_), .B(new_n9901_), .ZN(new_n9904_));
  NOR2_X1    g08898(.A1(new_n9903_), .A2(new_n9904_), .ZN(new_n9905_));
  INV_X1     g08899(.I(\A[247] ), .ZN(new_n9906_));
  INV_X1     g08900(.I(\A[248] ), .ZN(new_n9907_));
  NAND2_X1   g08901(.A1(new_n9907_), .A2(\A[249] ), .ZN(new_n9908_));
  INV_X1     g08902(.I(\A[249] ), .ZN(new_n9909_));
  NAND2_X1   g08903(.A1(new_n9909_), .A2(\A[248] ), .ZN(new_n9910_));
  AOI21_X1   g08904(.A1(new_n9908_), .A2(new_n9910_), .B(new_n9906_), .ZN(new_n9911_));
  NOR2_X1    g08905(.A1(\A[248] ), .A2(\A[249] ), .ZN(new_n9912_));
  INV_X1     g08906(.I(new_n9912_), .ZN(new_n9913_));
  NAND2_X1   g08907(.A1(\A[248] ), .A2(\A[249] ), .ZN(new_n9914_));
  AOI21_X1   g08908(.A1(new_n9913_), .A2(new_n9914_), .B(\A[247] ), .ZN(new_n9915_));
  NOR2_X1    g08909(.A1(new_n9915_), .A2(new_n9911_), .ZN(new_n9916_));
  INV_X1     g08910(.I(\A[252] ), .ZN(new_n9917_));
  NOR2_X1    g08911(.A1(new_n9917_), .A2(\A[251] ), .ZN(new_n9918_));
  INV_X1     g08912(.I(\A[251] ), .ZN(new_n9919_));
  NOR2_X1    g08913(.A1(new_n9919_), .A2(\A[252] ), .ZN(new_n9920_));
  OAI21_X1   g08914(.A1(new_n9918_), .A2(new_n9920_), .B(\A[250] ), .ZN(new_n9921_));
  INV_X1     g08915(.I(\A[250] ), .ZN(new_n9922_));
  NAND2_X1   g08916(.A1(\A[251] ), .A2(\A[252] ), .ZN(new_n9923_));
  INV_X1     g08917(.I(new_n9923_), .ZN(new_n9924_));
  NOR2_X1    g08918(.A1(\A[251] ), .A2(\A[252] ), .ZN(new_n9925_));
  OAI21_X1   g08919(.A1(new_n9924_), .A2(new_n9925_), .B(new_n9922_), .ZN(new_n9926_));
  NAND2_X1   g08920(.A1(new_n9921_), .A2(new_n9926_), .ZN(new_n9927_));
  AOI21_X1   g08921(.A1(new_n9906_), .A2(new_n9914_), .B(new_n9912_), .ZN(new_n9928_));
  AOI21_X1   g08922(.A1(new_n9922_), .A2(new_n9923_), .B(new_n9925_), .ZN(new_n9929_));
  NOR2_X1    g08923(.A1(new_n9928_), .A2(new_n9929_), .ZN(new_n9930_));
  XOR2_X1    g08924(.A1(new_n9916_), .A2(new_n9927_), .Z(new_n9931_));
  INV_X1     g08925(.I(new_n9931_), .ZN(new_n9932_));
  INV_X1     g08926(.I(\A[259] ), .ZN(new_n9933_));
  INV_X1     g08927(.I(\A[260] ), .ZN(new_n9934_));
  NAND2_X1   g08928(.A1(new_n9934_), .A2(\A[261] ), .ZN(new_n9935_));
  INV_X1     g08929(.I(\A[261] ), .ZN(new_n9936_));
  NAND2_X1   g08930(.A1(new_n9936_), .A2(\A[260] ), .ZN(new_n9937_));
  AOI21_X1   g08931(.A1(new_n9935_), .A2(new_n9937_), .B(new_n9933_), .ZN(new_n9938_));
  NOR2_X1    g08932(.A1(\A[260] ), .A2(\A[261] ), .ZN(new_n9939_));
  INV_X1     g08933(.I(new_n9939_), .ZN(new_n9940_));
  NAND2_X1   g08934(.A1(\A[260] ), .A2(\A[261] ), .ZN(new_n9941_));
  AOI21_X1   g08935(.A1(new_n9940_), .A2(new_n9941_), .B(\A[259] ), .ZN(new_n9942_));
  NOR2_X1    g08936(.A1(new_n9942_), .A2(new_n9938_), .ZN(new_n9943_));
  INV_X1     g08937(.I(\A[264] ), .ZN(new_n9944_));
  NOR2_X1    g08938(.A1(new_n9944_), .A2(\A[263] ), .ZN(new_n9945_));
  INV_X1     g08939(.I(\A[263] ), .ZN(new_n9946_));
  NOR2_X1    g08940(.A1(new_n9946_), .A2(\A[264] ), .ZN(new_n9947_));
  OAI21_X1   g08941(.A1(new_n9945_), .A2(new_n9947_), .B(\A[262] ), .ZN(new_n9948_));
  INV_X1     g08942(.I(\A[262] ), .ZN(new_n9949_));
  NAND2_X1   g08943(.A1(\A[263] ), .A2(\A[264] ), .ZN(new_n9950_));
  INV_X1     g08944(.I(new_n9950_), .ZN(new_n9951_));
  NOR2_X1    g08945(.A1(\A[263] ), .A2(\A[264] ), .ZN(new_n9952_));
  OAI21_X1   g08946(.A1(new_n9951_), .A2(new_n9952_), .B(new_n9949_), .ZN(new_n9953_));
  NAND2_X1   g08947(.A1(new_n9948_), .A2(new_n9953_), .ZN(new_n9954_));
  AOI21_X1   g08948(.A1(new_n9933_), .A2(new_n9941_), .B(new_n9939_), .ZN(new_n9955_));
  AOI21_X1   g08949(.A1(new_n9949_), .A2(new_n9950_), .B(new_n9952_), .ZN(new_n9956_));
  NOR2_X1    g08950(.A1(new_n9955_), .A2(new_n9956_), .ZN(new_n9957_));
  XOR2_X1    g08951(.A1(new_n9943_), .A2(new_n9954_), .Z(new_n9958_));
  INV_X1     g08952(.I(\A[267] ), .ZN(new_n9959_));
  NOR2_X1    g08953(.A1(new_n9959_), .A2(\A[266] ), .ZN(new_n9960_));
  INV_X1     g08954(.I(\A[266] ), .ZN(new_n9961_));
  NOR2_X1    g08955(.A1(new_n9961_), .A2(\A[267] ), .ZN(new_n9962_));
  OAI21_X1   g08956(.A1(new_n9960_), .A2(new_n9962_), .B(\A[265] ), .ZN(new_n9963_));
  INV_X1     g08957(.I(\A[265] ), .ZN(new_n9964_));
  NOR2_X1    g08958(.A1(\A[266] ), .A2(\A[267] ), .ZN(new_n9965_));
  AND2_X2    g08959(.A1(\A[266] ), .A2(\A[267] ), .Z(new_n9966_));
  OAI21_X1   g08960(.A1(new_n9966_), .A2(new_n9965_), .B(new_n9964_), .ZN(new_n9967_));
  NAND2_X1   g08961(.A1(new_n9963_), .A2(new_n9967_), .ZN(new_n9968_));
  INV_X1     g08962(.I(\A[268] ), .ZN(new_n9969_));
  INV_X1     g08963(.I(\A[269] ), .ZN(new_n9970_));
  NAND2_X1   g08964(.A1(new_n9970_), .A2(\A[270] ), .ZN(new_n9971_));
  INV_X1     g08965(.I(\A[270] ), .ZN(new_n9972_));
  NAND2_X1   g08966(.A1(new_n9972_), .A2(\A[269] ), .ZN(new_n9973_));
  AOI21_X1   g08967(.A1(new_n9971_), .A2(new_n9973_), .B(new_n9969_), .ZN(new_n9974_));
  NAND2_X1   g08968(.A1(\A[269] ), .A2(\A[270] ), .ZN(new_n9975_));
  NOR2_X1    g08969(.A1(\A[269] ), .A2(\A[270] ), .ZN(new_n9976_));
  INV_X1     g08970(.I(new_n9976_), .ZN(new_n9977_));
  AOI21_X1   g08971(.A1(new_n9977_), .A2(new_n9975_), .B(\A[268] ), .ZN(new_n9978_));
  NOR2_X1    g08972(.A1(new_n9978_), .A2(new_n9974_), .ZN(new_n9979_));
  AOI21_X1   g08973(.A1(\A[266] ), .A2(\A[267] ), .B(\A[265] ), .ZN(new_n9980_));
  NOR2_X1    g08974(.A1(new_n9980_), .A2(new_n9965_), .ZN(new_n9981_));
  AOI21_X1   g08975(.A1(\A[269] ), .A2(\A[270] ), .B(\A[268] ), .ZN(new_n9982_));
  NOR2_X1    g08976(.A1(new_n9982_), .A2(new_n9976_), .ZN(new_n9983_));
  NOR2_X1    g08977(.A1(new_n9981_), .A2(new_n9983_), .ZN(new_n9984_));
  XOR2_X1    g08978(.A1(new_n9979_), .A2(new_n9968_), .Z(new_n9985_));
  INV_X1     g08979(.I(\A[255] ), .ZN(new_n9986_));
  NOR2_X1    g08980(.A1(new_n9986_), .A2(\A[254] ), .ZN(new_n9987_));
  INV_X1     g08981(.I(\A[254] ), .ZN(new_n9988_));
  NOR2_X1    g08982(.A1(new_n9988_), .A2(\A[255] ), .ZN(new_n9989_));
  OAI21_X1   g08983(.A1(new_n9987_), .A2(new_n9989_), .B(\A[253] ), .ZN(new_n9990_));
  INV_X1     g08984(.I(\A[253] ), .ZN(new_n9991_));
  NOR2_X1    g08985(.A1(\A[254] ), .A2(\A[255] ), .ZN(new_n9992_));
  NAND2_X1   g08986(.A1(\A[254] ), .A2(\A[255] ), .ZN(new_n9993_));
  INV_X1     g08987(.I(new_n9993_), .ZN(new_n9994_));
  OAI21_X1   g08988(.A1(new_n9994_), .A2(new_n9992_), .B(new_n9991_), .ZN(new_n9995_));
  NAND2_X1   g08989(.A1(new_n9990_), .A2(new_n9995_), .ZN(new_n9996_));
  INV_X1     g08990(.I(\A[258] ), .ZN(new_n9997_));
  NOR2_X1    g08991(.A1(new_n9997_), .A2(\A[257] ), .ZN(new_n9998_));
  INV_X1     g08992(.I(\A[257] ), .ZN(new_n9999_));
  NOR2_X1    g08993(.A1(new_n9999_), .A2(\A[258] ), .ZN(new_n10000_));
  OAI21_X1   g08994(.A1(new_n9998_), .A2(new_n10000_), .B(\A[256] ), .ZN(new_n10001_));
  INV_X1     g08995(.I(\A[256] ), .ZN(new_n10002_));
  NAND2_X1   g08996(.A1(\A[257] ), .A2(\A[258] ), .ZN(new_n10003_));
  INV_X1     g08997(.I(new_n10003_), .ZN(new_n10004_));
  NOR2_X1    g08998(.A1(\A[257] ), .A2(\A[258] ), .ZN(new_n10005_));
  OAI21_X1   g08999(.A1(new_n10004_), .A2(new_n10005_), .B(new_n10002_), .ZN(new_n10006_));
  NAND2_X1   g09000(.A1(new_n10001_), .A2(new_n10006_), .ZN(new_n10007_));
  AOI21_X1   g09001(.A1(\A[254] ), .A2(\A[255] ), .B(\A[253] ), .ZN(new_n10008_));
  NOR2_X1    g09002(.A1(new_n10008_), .A2(new_n9992_), .ZN(new_n10009_));
  AOI21_X1   g09003(.A1(\A[257] ), .A2(\A[258] ), .B(\A[256] ), .ZN(new_n10010_));
  NOR2_X1    g09004(.A1(new_n10010_), .A2(new_n10005_), .ZN(new_n10011_));
  NOR2_X1    g09005(.A1(new_n10009_), .A2(new_n10011_), .ZN(new_n10012_));
  XOR2_X1    g09006(.A1(new_n9996_), .A2(new_n10007_), .Z(new_n10013_));
  NAND2_X1   g09007(.A1(new_n10013_), .A2(new_n9985_), .ZN(new_n10014_));
  NOR2_X1    g09008(.A1(new_n9972_), .A2(\A[269] ), .ZN(new_n10015_));
  NOR2_X1    g09009(.A1(new_n9970_), .A2(\A[270] ), .ZN(new_n10016_));
  OAI21_X1   g09010(.A1(new_n10015_), .A2(new_n10016_), .B(\A[268] ), .ZN(new_n10017_));
  INV_X1     g09011(.I(new_n9975_), .ZN(new_n10018_));
  OAI21_X1   g09012(.A1(new_n10018_), .A2(new_n9976_), .B(new_n9969_), .ZN(new_n10019_));
  NAND2_X1   g09013(.A1(new_n10017_), .A2(new_n10019_), .ZN(new_n10020_));
  XOR2_X1    g09014(.A1(new_n10020_), .A2(new_n9968_), .Z(new_n10021_));
  NAND2_X1   g09015(.A1(new_n9988_), .A2(\A[255] ), .ZN(new_n10022_));
  NAND2_X1   g09016(.A1(new_n9986_), .A2(\A[254] ), .ZN(new_n10023_));
  AOI21_X1   g09017(.A1(new_n10022_), .A2(new_n10023_), .B(new_n9991_), .ZN(new_n10024_));
  INV_X1     g09018(.I(new_n9992_), .ZN(new_n10025_));
  AOI21_X1   g09019(.A1(new_n10025_), .A2(new_n9993_), .B(\A[253] ), .ZN(new_n10026_));
  NOR2_X1    g09020(.A1(new_n10026_), .A2(new_n10024_), .ZN(new_n10027_));
  XOR2_X1    g09021(.A1(new_n10027_), .A2(new_n10007_), .Z(new_n10028_));
  NAND2_X1   g09022(.A1(new_n10028_), .A2(new_n10021_), .ZN(new_n10029_));
  NAND2_X1   g09023(.A1(new_n10014_), .A2(new_n10029_), .ZN(new_n10030_));
  NAND2_X1   g09024(.A1(new_n10030_), .A2(new_n9958_), .ZN(new_n10031_));
  NOR2_X1    g09025(.A1(new_n9936_), .A2(\A[260] ), .ZN(new_n10032_));
  NOR2_X1    g09026(.A1(new_n9934_), .A2(\A[261] ), .ZN(new_n10033_));
  OAI21_X1   g09027(.A1(new_n10032_), .A2(new_n10033_), .B(\A[259] ), .ZN(new_n10034_));
  INV_X1     g09028(.I(new_n9941_), .ZN(new_n10035_));
  OAI21_X1   g09029(.A1(new_n10035_), .A2(new_n9939_), .B(new_n9933_), .ZN(new_n10036_));
  NAND2_X1   g09030(.A1(new_n10034_), .A2(new_n10036_), .ZN(new_n10037_));
  XOR2_X1    g09031(.A1(new_n10037_), .A2(new_n9954_), .Z(new_n10038_));
  NOR2_X1    g09032(.A1(new_n10028_), .A2(new_n10021_), .ZN(new_n10039_));
  NOR2_X1    g09033(.A1(new_n10013_), .A2(new_n9985_), .ZN(new_n10040_));
  NOR2_X1    g09034(.A1(new_n10040_), .A2(new_n10039_), .ZN(new_n10041_));
  NAND2_X1   g09035(.A1(new_n10041_), .A2(new_n10038_), .ZN(new_n10042_));
  AOI21_X1   g09036(.A1(new_n10042_), .A2(new_n10031_), .B(new_n9932_), .ZN(new_n10043_));
  NOR2_X1    g09037(.A1(new_n10041_), .A2(new_n10038_), .ZN(new_n10044_));
  NOR2_X1    g09038(.A1(new_n10030_), .A2(new_n9958_), .ZN(new_n10045_));
  NOR3_X1    g09039(.A1(new_n10044_), .A2(new_n10045_), .A3(new_n9931_), .ZN(new_n10046_));
  INV_X1     g09040(.I(\A[223] ), .ZN(new_n10047_));
  INV_X1     g09041(.I(\A[224] ), .ZN(new_n10048_));
  NAND2_X1   g09042(.A1(new_n10048_), .A2(\A[225] ), .ZN(new_n10049_));
  INV_X1     g09043(.I(\A[225] ), .ZN(new_n10050_));
  NAND2_X1   g09044(.A1(new_n10050_), .A2(\A[224] ), .ZN(new_n10051_));
  AOI21_X1   g09045(.A1(new_n10049_), .A2(new_n10051_), .B(new_n10047_), .ZN(new_n10052_));
  NAND2_X1   g09046(.A1(\A[224] ), .A2(\A[225] ), .ZN(new_n10053_));
  NOR2_X1    g09047(.A1(\A[224] ), .A2(\A[225] ), .ZN(new_n10054_));
  INV_X1     g09048(.I(new_n10054_), .ZN(new_n10055_));
  AOI21_X1   g09049(.A1(new_n10055_), .A2(new_n10053_), .B(\A[223] ), .ZN(new_n10056_));
  INV_X1     g09050(.I(\A[226] ), .ZN(new_n10057_));
  INV_X1     g09051(.I(\A[227] ), .ZN(new_n10058_));
  NAND2_X1   g09052(.A1(new_n10058_), .A2(\A[228] ), .ZN(new_n10059_));
  INV_X1     g09053(.I(\A[228] ), .ZN(new_n10060_));
  NAND2_X1   g09054(.A1(new_n10060_), .A2(\A[227] ), .ZN(new_n10061_));
  AOI21_X1   g09055(.A1(new_n10059_), .A2(new_n10061_), .B(new_n10057_), .ZN(new_n10062_));
  NAND2_X1   g09056(.A1(\A[227] ), .A2(\A[228] ), .ZN(new_n10063_));
  NOR2_X1    g09057(.A1(\A[227] ), .A2(\A[228] ), .ZN(new_n10064_));
  INV_X1     g09058(.I(new_n10064_), .ZN(new_n10065_));
  AOI21_X1   g09059(.A1(new_n10065_), .A2(new_n10063_), .B(\A[226] ), .ZN(new_n10066_));
  OAI22_X1   g09060(.A1(new_n10052_), .A2(new_n10056_), .B1(new_n10066_), .B2(new_n10062_), .ZN(new_n10067_));
  NOR2_X1    g09061(.A1(new_n10050_), .A2(\A[224] ), .ZN(new_n10068_));
  NOR2_X1    g09062(.A1(new_n10048_), .A2(\A[225] ), .ZN(new_n10069_));
  OAI21_X1   g09063(.A1(new_n10068_), .A2(new_n10069_), .B(\A[223] ), .ZN(new_n10070_));
  INV_X1     g09064(.I(new_n10053_), .ZN(new_n10071_));
  OAI21_X1   g09065(.A1(new_n10071_), .A2(new_n10054_), .B(new_n10047_), .ZN(new_n10072_));
  NOR2_X1    g09066(.A1(new_n10060_), .A2(\A[227] ), .ZN(new_n10073_));
  NOR2_X1    g09067(.A1(new_n10058_), .A2(\A[228] ), .ZN(new_n10074_));
  OAI21_X1   g09068(.A1(new_n10073_), .A2(new_n10074_), .B(\A[226] ), .ZN(new_n10075_));
  INV_X1     g09069(.I(new_n10063_), .ZN(new_n10076_));
  OAI21_X1   g09070(.A1(new_n10076_), .A2(new_n10064_), .B(new_n10057_), .ZN(new_n10077_));
  NAND4_X1   g09071(.A1(new_n10070_), .A2(new_n10072_), .A3(new_n10075_), .A4(new_n10077_), .ZN(new_n10078_));
  NAND2_X1   g09072(.A1(new_n10067_), .A2(new_n10078_), .ZN(new_n10079_));
  NOR2_X1    g09073(.A1(new_n10056_), .A2(new_n10052_), .ZN(new_n10080_));
  NOR2_X1    g09074(.A1(new_n10066_), .A2(new_n10062_), .ZN(new_n10081_));
  AOI21_X1   g09075(.A1(\A[224] ), .A2(\A[225] ), .B(\A[223] ), .ZN(new_n10082_));
  AOI21_X1   g09076(.A1(\A[227] ), .A2(\A[228] ), .B(\A[226] ), .ZN(new_n10083_));
  OAI22_X1   g09077(.A1(new_n10054_), .A2(new_n10082_), .B1(new_n10083_), .B2(new_n10064_), .ZN(new_n10084_));
  NOR3_X1    g09078(.A1(new_n10080_), .A2(new_n10081_), .A3(new_n10084_), .ZN(new_n10085_));
  NOR2_X1    g09079(.A1(new_n10079_), .A2(new_n10085_), .ZN(new_n10086_));
  INV_X1     g09080(.I(\A[237] ), .ZN(new_n10087_));
  NOR2_X1    g09081(.A1(new_n10087_), .A2(\A[236] ), .ZN(new_n10088_));
  INV_X1     g09082(.I(\A[236] ), .ZN(new_n10089_));
  NOR2_X1    g09083(.A1(new_n10089_), .A2(\A[237] ), .ZN(new_n10090_));
  OAI21_X1   g09084(.A1(new_n10088_), .A2(new_n10090_), .B(\A[235] ), .ZN(new_n10091_));
  INV_X1     g09085(.I(\A[235] ), .ZN(new_n10092_));
  NAND2_X1   g09086(.A1(\A[236] ), .A2(\A[237] ), .ZN(new_n10093_));
  INV_X1     g09087(.I(new_n10093_), .ZN(new_n10094_));
  NOR2_X1    g09088(.A1(\A[236] ), .A2(\A[237] ), .ZN(new_n10095_));
  OAI21_X1   g09089(.A1(new_n10094_), .A2(new_n10095_), .B(new_n10092_), .ZN(new_n10096_));
  NAND2_X1   g09090(.A1(new_n10091_), .A2(new_n10096_), .ZN(new_n10097_));
  INV_X1     g09091(.I(\A[240] ), .ZN(new_n10098_));
  NOR2_X1    g09092(.A1(new_n10098_), .A2(\A[239] ), .ZN(new_n10099_));
  INV_X1     g09093(.I(\A[239] ), .ZN(new_n10100_));
  NOR2_X1    g09094(.A1(new_n10100_), .A2(\A[240] ), .ZN(new_n10101_));
  OAI21_X1   g09095(.A1(new_n10099_), .A2(new_n10101_), .B(\A[238] ), .ZN(new_n10102_));
  INV_X1     g09096(.I(\A[238] ), .ZN(new_n10103_));
  NAND2_X1   g09097(.A1(\A[239] ), .A2(\A[240] ), .ZN(new_n10104_));
  INV_X1     g09098(.I(new_n10104_), .ZN(new_n10105_));
  NOR2_X1    g09099(.A1(\A[239] ), .A2(\A[240] ), .ZN(new_n10106_));
  OAI21_X1   g09100(.A1(new_n10105_), .A2(new_n10106_), .B(new_n10103_), .ZN(new_n10107_));
  NAND2_X1   g09101(.A1(new_n10102_), .A2(new_n10107_), .ZN(new_n10108_));
  NAND2_X1   g09102(.A1(new_n10097_), .A2(new_n10108_), .ZN(new_n10109_));
  NAND2_X1   g09103(.A1(new_n10089_), .A2(\A[237] ), .ZN(new_n10110_));
  NAND2_X1   g09104(.A1(new_n10087_), .A2(\A[236] ), .ZN(new_n10111_));
  AOI21_X1   g09105(.A1(new_n10110_), .A2(new_n10111_), .B(new_n10092_), .ZN(new_n10112_));
  INV_X1     g09106(.I(new_n10095_), .ZN(new_n10113_));
  AOI21_X1   g09107(.A1(new_n10113_), .A2(new_n10093_), .B(\A[235] ), .ZN(new_n10114_));
  NOR2_X1    g09108(.A1(new_n10114_), .A2(new_n10112_), .ZN(new_n10115_));
  NAND2_X1   g09109(.A1(new_n10100_), .A2(\A[240] ), .ZN(new_n10116_));
  NAND2_X1   g09110(.A1(new_n10098_), .A2(\A[239] ), .ZN(new_n10117_));
  AOI21_X1   g09111(.A1(new_n10116_), .A2(new_n10117_), .B(new_n10103_), .ZN(new_n10118_));
  INV_X1     g09112(.I(new_n10106_), .ZN(new_n10119_));
  AOI21_X1   g09113(.A1(new_n10119_), .A2(new_n10104_), .B(\A[238] ), .ZN(new_n10120_));
  NOR2_X1    g09114(.A1(new_n10120_), .A2(new_n10118_), .ZN(new_n10121_));
  NAND2_X1   g09115(.A1(new_n10115_), .A2(new_n10121_), .ZN(new_n10122_));
  AOI21_X1   g09116(.A1(new_n10092_), .A2(new_n10093_), .B(new_n10095_), .ZN(new_n10123_));
  AOI21_X1   g09117(.A1(new_n10103_), .A2(new_n10104_), .B(new_n10106_), .ZN(new_n10124_));
  NOR2_X1    g09118(.A1(new_n10123_), .A2(new_n10124_), .ZN(new_n10125_));
  NAND3_X1   g09119(.A1(new_n10097_), .A2(new_n10108_), .A3(new_n10125_), .ZN(new_n10126_));
  NAND3_X1   g09120(.A1(new_n10122_), .A2(new_n10126_), .A3(new_n10109_), .ZN(new_n10127_));
  INV_X1     g09121(.I(\A[243] ), .ZN(new_n10128_));
  NOR2_X1    g09122(.A1(new_n10128_), .A2(\A[242] ), .ZN(new_n10129_));
  INV_X1     g09123(.I(\A[242] ), .ZN(new_n10130_));
  NOR2_X1    g09124(.A1(new_n10130_), .A2(\A[243] ), .ZN(new_n10131_));
  OAI21_X1   g09125(.A1(new_n10129_), .A2(new_n10131_), .B(\A[241] ), .ZN(new_n10132_));
  INV_X1     g09126(.I(\A[241] ), .ZN(new_n10133_));
  NOR2_X1    g09127(.A1(\A[242] ), .A2(\A[243] ), .ZN(new_n10134_));
  NAND2_X1   g09128(.A1(\A[242] ), .A2(\A[243] ), .ZN(new_n10135_));
  INV_X1     g09129(.I(new_n10135_), .ZN(new_n10136_));
  OAI21_X1   g09130(.A1(new_n10136_), .A2(new_n10134_), .B(new_n10133_), .ZN(new_n10137_));
  NAND2_X1   g09131(.A1(new_n10132_), .A2(new_n10137_), .ZN(new_n10138_));
  INV_X1     g09132(.I(\A[246] ), .ZN(new_n10139_));
  NOR2_X1    g09133(.A1(new_n10139_), .A2(\A[245] ), .ZN(new_n10140_));
  INV_X1     g09134(.I(\A[245] ), .ZN(new_n10141_));
  NOR2_X1    g09135(.A1(new_n10141_), .A2(\A[246] ), .ZN(new_n10142_));
  OAI21_X1   g09136(.A1(new_n10140_), .A2(new_n10142_), .B(\A[244] ), .ZN(new_n10143_));
  INV_X1     g09137(.I(\A[244] ), .ZN(new_n10144_));
  NAND2_X1   g09138(.A1(\A[245] ), .A2(\A[246] ), .ZN(new_n10145_));
  INV_X1     g09139(.I(new_n10145_), .ZN(new_n10146_));
  NOR2_X1    g09140(.A1(\A[245] ), .A2(\A[246] ), .ZN(new_n10147_));
  OAI21_X1   g09141(.A1(new_n10146_), .A2(new_n10147_), .B(new_n10144_), .ZN(new_n10148_));
  NAND2_X1   g09142(.A1(new_n10143_), .A2(new_n10148_), .ZN(new_n10149_));
  AOI21_X1   g09143(.A1(\A[242] ), .A2(\A[243] ), .B(\A[241] ), .ZN(new_n10150_));
  AOI21_X1   g09144(.A1(\A[245] ), .A2(\A[246] ), .B(\A[244] ), .ZN(new_n10151_));
  OAI22_X1   g09145(.A1(new_n10134_), .A2(new_n10150_), .B1(new_n10151_), .B2(new_n10147_), .ZN(new_n10152_));
  INV_X1     g09146(.I(new_n10152_), .ZN(new_n10153_));
  XOR2_X1    g09147(.A1(new_n10138_), .A2(new_n10149_), .Z(new_n10154_));
  INV_X1     g09148(.I(\A[231] ), .ZN(new_n10155_));
  NOR2_X1    g09149(.A1(new_n10155_), .A2(\A[230] ), .ZN(new_n10156_));
  INV_X1     g09150(.I(\A[230] ), .ZN(new_n10157_));
  NOR2_X1    g09151(.A1(new_n10157_), .A2(\A[231] ), .ZN(new_n10158_));
  OAI21_X1   g09152(.A1(new_n10156_), .A2(new_n10158_), .B(\A[229] ), .ZN(new_n10159_));
  INV_X1     g09153(.I(\A[229] ), .ZN(new_n10160_));
  AND2_X2    g09154(.A1(\A[230] ), .A2(\A[231] ), .Z(new_n10161_));
  NOR2_X1    g09155(.A1(\A[230] ), .A2(\A[231] ), .ZN(new_n10162_));
  OAI21_X1   g09156(.A1(new_n10161_), .A2(new_n10162_), .B(new_n10160_), .ZN(new_n10163_));
  INV_X1     g09157(.I(\A[234] ), .ZN(new_n10164_));
  NOR2_X1    g09158(.A1(new_n10164_), .A2(\A[233] ), .ZN(new_n10165_));
  INV_X1     g09159(.I(\A[233] ), .ZN(new_n10166_));
  NOR2_X1    g09160(.A1(new_n10166_), .A2(\A[234] ), .ZN(new_n10167_));
  OAI21_X1   g09161(.A1(new_n10165_), .A2(new_n10167_), .B(\A[232] ), .ZN(new_n10168_));
  INV_X1     g09162(.I(\A[232] ), .ZN(new_n10169_));
  AND2_X2    g09163(.A1(\A[233] ), .A2(\A[234] ), .Z(new_n10170_));
  NOR2_X1    g09164(.A1(\A[233] ), .A2(\A[234] ), .ZN(new_n10171_));
  OAI21_X1   g09165(.A1(new_n10170_), .A2(new_n10171_), .B(new_n10169_), .ZN(new_n10172_));
  AOI22_X1   g09166(.A1(new_n10159_), .A2(new_n10163_), .B1(new_n10168_), .B2(new_n10172_), .ZN(new_n10173_));
  NAND2_X1   g09167(.A1(new_n10157_), .A2(\A[231] ), .ZN(new_n10174_));
  NAND2_X1   g09168(.A1(new_n10155_), .A2(\A[230] ), .ZN(new_n10175_));
  AOI21_X1   g09169(.A1(new_n10174_), .A2(new_n10175_), .B(new_n10160_), .ZN(new_n10176_));
  NAND2_X1   g09170(.A1(\A[230] ), .A2(\A[231] ), .ZN(new_n10177_));
  OR2_X2     g09171(.A1(\A[230] ), .A2(\A[231] ), .Z(new_n10178_));
  AOI21_X1   g09172(.A1(new_n10178_), .A2(new_n10177_), .B(\A[229] ), .ZN(new_n10179_));
  NAND2_X1   g09173(.A1(new_n10166_), .A2(\A[234] ), .ZN(new_n10180_));
  NAND2_X1   g09174(.A1(new_n10164_), .A2(\A[233] ), .ZN(new_n10181_));
  AOI21_X1   g09175(.A1(new_n10180_), .A2(new_n10181_), .B(new_n10169_), .ZN(new_n10182_));
  NAND2_X1   g09176(.A1(\A[233] ), .A2(\A[234] ), .ZN(new_n10183_));
  INV_X1     g09177(.I(new_n10171_), .ZN(new_n10184_));
  AOI21_X1   g09178(.A1(new_n10184_), .A2(new_n10183_), .B(\A[232] ), .ZN(new_n10185_));
  NOR4_X1    g09179(.A1(new_n10176_), .A2(new_n10185_), .A3(new_n10182_), .A4(new_n10179_), .ZN(new_n10186_));
  NOR2_X1    g09180(.A1(new_n10173_), .A2(new_n10186_), .ZN(new_n10187_));
  NAND2_X1   g09181(.A1(new_n10168_), .A2(new_n10172_), .ZN(new_n10188_));
  AOI21_X1   g09182(.A1(\A[233] ), .A2(\A[234] ), .B(\A[232] ), .ZN(new_n10189_));
  NOR2_X1    g09183(.A1(new_n10189_), .A2(new_n10171_), .ZN(new_n10190_));
  NOR4_X1    g09184(.A1(new_n10190_), .A2(\A[229] ), .A3(\A[230] ), .A4(\A[231] ), .ZN(new_n10191_));
  NAND2_X1   g09185(.A1(new_n10188_), .A2(new_n10191_), .ZN(new_n10192_));
  NAND2_X1   g09186(.A1(new_n10187_), .A2(new_n10192_), .ZN(new_n10193_));
  NOR2_X1    g09187(.A1(new_n10154_), .A2(new_n10193_), .ZN(new_n10194_));
  NAND2_X1   g09188(.A1(new_n10130_), .A2(\A[243] ), .ZN(new_n10195_));
  NAND2_X1   g09189(.A1(new_n10128_), .A2(\A[242] ), .ZN(new_n10196_));
  AOI21_X1   g09190(.A1(new_n10195_), .A2(new_n10196_), .B(new_n10133_), .ZN(new_n10197_));
  INV_X1     g09191(.I(new_n10134_), .ZN(new_n10198_));
  AOI21_X1   g09192(.A1(new_n10198_), .A2(new_n10135_), .B(\A[241] ), .ZN(new_n10199_));
  NOR2_X1    g09193(.A1(new_n10199_), .A2(new_n10197_), .ZN(new_n10200_));
  XOR2_X1    g09194(.A1(new_n10200_), .A2(new_n10149_), .Z(new_n10201_));
  OAI22_X1   g09195(.A1(new_n10182_), .A2(new_n10185_), .B1(new_n10176_), .B2(new_n10179_), .ZN(new_n10202_));
  NAND4_X1   g09196(.A1(new_n10159_), .A2(new_n10168_), .A3(new_n10163_), .A4(new_n10172_), .ZN(new_n10203_));
  NAND2_X1   g09197(.A1(new_n10202_), .A2(new_n10203_), .ZN(new_n10204_));
  NOR2_X1    g09198(.A1(new_n10176_), .A2(new_n10179_), .ZN(new_n10205_));
  NOR2_X1    g09199(.A1(new_n10185_), .A2(new_n10182_), .ZN(new_n10206_));
  AOI21_X1   g09200(.A1(\A[230] ), .A2(\A[231] ), .B(\A[229] ), .ZN(new_n10207_));
  OAI22_X1   g09201(.A1(new_n10162_), .A2(new_n10207_), .B1(new_n10189_), .B2(new_n10171_), .ZN(new_n10208_));
  NOR3_X1    g09202(.A1(new_n10206_), .A2(new_n10205_), .A3(new_n10208_), .ZN(new_n10209_));
  NOR2_X1    g09203(.A1(new_n10204_), .A2(new_n10209_), .ZN(new_n10210_));
  NOR2_X1    g09204(.A1(new_n10201_), .A2(new_n10210_), .ZN(new_n10211_));
  OAI21_X1   g09205(.A1(new_n10194_), .A2(new_n10211_), .B(new_n10127_), .ZN(new_n10212_));
  XOR2_X1    g09206(.A1(new_n10097_), .A2(new_n10108_), .Z(new_n10213_));
  NAND2_X1   g09207(.A1(new_n10201_), .A2(new_n10210_), .ZN(new_n10214_));
  NAND2_X1   g09208(.A1(new_n10154_), .A2(new_n10193_), .ZN(new_n10215_));
  NAND3_X1   g09209(.A1(new_n10215_), .A2(new_n10214_), .A3(new_n10213_), .ZN(new_n10216_));
  AOI21_X1   g09210(.A1(new_n10212_), .A2(new_n10216_), .B(new_n10086_), .ZN(new_n10217_));
  NAND3_X1   g09211(.A1(new_n10212_), .A2(new_n10216_), .A3(new_n10086_), .ZN(new_n10218_));
  INV_X1     g09212(.I(new_n10218_), .ZN(new_n10219_));
  NOR4_X1    g09213(.A1(new_n10043_), .A2(new_n10046_), .A3(new_n10219_), .A4(new_n10217_), .ZN(new_n10220_));
  OAI21_X1   g09214(.A1(new_n10044_), .A2(new_n10045_), .B(new_n9931_), .ZN(new_n10221_));
  NAND3_X1   g09215(.A1(new_n10042_), .A2(new_n10031_), .A3(new_n9932_), .ZN(new_n10222_));
  INV_X1     g09216(.I(new_n10217_), .ZN(new_n10223_));
  AOI22_X1   g09217(.A1(new_n10221_), .A2(new_n10222_), .B1(new_n10223_), .B2(new_n10218_), .ZN(new_n10224_));
  NOR2_X1    g09218(.A1(new_n10224_), .A2(new_n10220_), .ZN(new_n10225_));
  NAND2_X1   g09219(.A1(new_n9905_), .A2(new_n10225_), .ZN(new_n10226_));
  OAI22_X1   g09220(.A1(new_n9903_), .A2(new_n9904_), .B1(new_n10220_), .B2(new_n10224_), .ZN(new_n10227_));
  INV_X1     g09221(.I(\A[169] ), .ZN(new_n10228_));
  INV_X1     g09222(.I(\A[170] ), .ZN(new_n10229_));
  NAND2_X1   g09223(.A1(new_n10229_), .A2(\A[171] ), .ZN(new_n10230_));
  INV_X1     g09224(.I(\A[171] ), .ZN(new_n10231_));
  NAND2_X1   g09225(.A1(new_n10231_), .A2(\A[170] ), .ZN(new_n10232_));
  AOI21_X1   g09226(.A1(new_n10230_), .A2(new_n10232_), .B(new_n10228_), .ZN(new_n10233_));
  NAND2_X1   g09227(.A1(\A[170] ), .A2(\A[171] ), .ZN(new_n10234_));
  NOR2_X1    g09228(.A1(\A[170] ), .A2(\A[171] ), .ZN(new_n10235_));
  INV_X1     g09229(.I(new_n10235_), .ZN(new_n10236_));
  AOI21_X1   g09230(.A1(new_n10236_), .A2(new_n10234_), .B(\A[169] ), .ZN(new_n10237_));
  NOR2_X1    g09231(.A1(new_n10237_), .A2(new_n10233_), .ZN(new_n10238_));
  INV_X1     g09232(.I(\A[172] ), .ZN(new_n10239_));
  INV_X1     g09233(.I(\A[173] ), .ZN(new_n10240_));
  NAND2_X1   g09234(.A1(new_n10240_), .A2(\A[174] ), .ZN(new_n10241_));
  INV_X1     g09235(.I(\A[174] ), .ZN(new_n10242_));
  NAND2_X1   g09236(.A1(new_n10242_), .A2(\A[173] ), .ZN(new_n10243_));
  AOI21_X1   g09237(.A1(new_n10241_), .A2(new_n10243_), .B(new_n10239_), .ZN(new_n10244_));
  NAND2_X1   g09238(.A1(\A[173] ), .A2(\A[174] ), .ZN(new_n10245_));
  NOR2_X1    g09239(.A1(\A[173] ), .A2(\A[174] ), .ZN(new_n10246_));
  INV_X1     g09240(.I(new_n10246_), .ZN(new_n10247_));
  AOI21_X1   g09241(.A1(new_n10247_), .A2(new_n10245_), .B(\A[172] ), .ZN(new_n10248_));
  NOR2_X1    g09242(.A1(new_n10248_), .A2(new_n10244_), .ZN(new_n10249_));
  AOI21_X1   g09243(.A1(\A[170] ), .A2(\A[171] ), .B(\A[169] ), .ZN(new_n10250_));
  AOI21_X1   g09244(.A1(\A[173] ), .A2(\A[174] ), .B(\A[172] ), .ZN(new_n10251_));
  OAI22_X1   g09245(.A1(new_n10235_), .A2(new_n10250_), .B1(new_n10251_), .B2(new_n10246_), .ZN(new_n10252_));
  NOR3_X1    g09246(.A1(new_n10238_), .A2(new_n10249_), .A3(new_n10252_), .ZN(new_n10253_));
  INV_X1     g09247(.I(\A[165] ), .ZN(new_n10254_));
  NOR2_X1    g09248(.A1(new_n10254_), .A2(\A[164] ), .ZN(new_n10255_));
  INV_X1     g09249(.I(\A[164] ), .ZN(new_n10256_));
  NOR2_X1    g09250(.A1(new_n10256_), .A2(\A[165] ), .ZN(new_n10257_));
  OAI21_X1   g09251(.A1(new_n10255_), .A2(new_n10257_), .B(\A[163] ), .ZN(new_n10258_));
  INV_X1     g09252(.I(\A[163] ), .ZN(new_n10259_));
  NAND2_X1   g09253(.A1(\A[164] ), .A2(\A[165] ), .ZN(new_n10260_));
  INV_X1     g09254(.I(new_n10260_), .ZN(new_n10261_));
  NOR2_X1    g09255(.A1(\A[164] ), .A2(\A[165] ), .ZN(new_n10262_));
  OAI21_X1   g09256(.A1(new_n10261_), .A2(new_n10262_), .B(new_n10259_), .ZN(new_n10263_));
  NAND2_X1   g09257(.A1(new_n10258_), .A2(new_n10263_), .ZN(new_n10264_));
  INV_X1     g09258(.I(\A[168] ), .ZN(new_n10265_));
  NOR2_X1    g09259(.A1(new_n10265_), .A2(\A[167] ), .ZN(new_n10266_));
  INV_X1     g09260(.I(\A[167] ), .ZN(new_n10267_));
  NOR2_X1    g09261(.A1(new_n10267_), .A2(\A[168] ), .ZN(new_n10268_));
  OAI21_X1   g09262(.A1(new_n10266_), .A2(new_n10268_), .B(\A[166] ), .ZN(new_n10269_));
  INV_X1     g09263(.I(\A[166] ), .ZN(new_n10270_));
  NAND2_X1   g09264(.A1(\A[167] ), .A2(\A[168] ), .ZN(new_n10271_));
  INV_X1     g09265(.I(new_n10271_), .ZN(new_n10272_));
  NOR2_X1    g09266(.A1(\A[167] ), .A2(\A[168] ), .ZN(new_n10273_));
  OAI21_X1   g09267(.A1(new_n10272_), .A2(new_n10273_), .B(new_n10270_), .ZN(new_n10274_));
  NAND2_X1   g09268(.A1(new_n10269_), .A2(new_n10274_), .ZN(new_n10275_));
  AOI21_X1   g09269(.A1(\A[164] ), .A2(\A[165] ), .B(\A[163] ), .ZN(new_n10276_));
  AOI21_X1   g09270(.A1(\A[167] ), .A2(\A[168] ), .B(\A[166] ), .ZN(new_n10277_));
  OAI22_X1   g09271(.A1(new_n10262_), .A2(new_n10276_), .B1(new_n10277_), .B2(new_n10273_), .ZN(new_n10278_));
  INV_X1     g09272(.I(new_n10278_), .ZN(new_n10279_));
  NAND3_X1   g09273(.A1(new_n10275_), .A2(new_n10264_), .A3(new_n10279_), .ZN(new_n10280_));
  NOR2_X1    g09274(.A1(new_n10253_), .A2(new_n10280_), .ZN(new_n10281_));
  NAND2_X1   g09275(.A1(new_n10253_), .A2(new_n10280_), .ZN(new_n10282_));
  INV_X1     g09276(.I(new_n10282_), .ZN(new_n10283_));
  INV_X1     g09277(.I(\A[157] ), .ZN(new_n10284_));
  INV_X1     g09278(.I(\A[158] ), .ZN(new_n10285_));
  NAND2_X1   g09279(.A1(new_n10285_), .A2(\A[159] ), .ZN(new_n10286_));
  INV_X1     g09280(.I(\A[159] ), .ZN(new_n10287_));
  NAND2_X1   g09281(.A1(new_n10287_), .A2(\A[158] ), .ZN(new_n10288_));
  AOI21_X1   g09282(.A1(new_n10286_), .A2(new_n10288_), .B(new_n10284_), .ZN(new_n10289_));
  NAND2_X1   g09283(.A1(\A[158] ), .A2(\A[159] ), .ZN(new_n10290_));
  NOR2_X1    g09284(.A1(\A[158] ), .A2(\A[159] ), .ZN(new_n10291_));
  INV_X1     g09285(.I(new_n10291_), .ZN(new_n10292_));
  AOI21_X1   g09286(.A1(new_n10292_), .A2(new_n10290_), .B(\A[157] ), .ZN(new_n10293_));
  NOR2_X1    g09287(.A1(new_n10293_), .A2(new_n10289_), .ZN(new_n10294_));
  INV_X1     g09288(.I(\A[160] ), .ZN(new_n10295_));
  INV_X1     g09289(.I(\A[161] ), .ZN(new_n10296_));
  NAND2_X1   g09290(.A1(new_n10296_), .A2(\A[162] ), .ZN(new_n10297_));
  INV_X1     g09291(.I(\A[162] ), .ZN(new_n10298_));
  NAND2_X1   g09292(.A1(new_n10298_), .A2(\A[161] ), .ZN(new_n10299_));
  AOI21_X1   g09293(.A1(new_n10297_), .A2(new_n10299_), .B(new_n10295_), .ZN(new_n10300_));
  NAND2_X1   g09294(.A1(\A[161] ), .A2(\A[162] ), .ZN(new_n10301_));
  NOR2_X1    g09295(.A1(\A[161] ), .A2(\A[162] ), .ZN(new_n10302_));
  INV_X1     g09296(.I(new_n10302_), .ZN(new_n10303_));
  AOI21_X1   g09297(.A1(new_n10303_), .A2(new_n10301_), .B(\A[160] ), .ZN(new_n10304_));
  NOR2_X1    g09298(.A1(new_n10304_), .A2(new_n10300_), .ZN(new_n10305_));
  AOI21_X1   g09299(.A1(\A[158] ), .A2(\A[159] ), .B(\A[157] ), .ZN(new_n10306_));
  AOI21_X1   g09300(.A1(\A[161] ), .A2(\A[162] ), .B(\A[160] ), .ZN(new_n10307_));
  OAI22_X1   g09301(.A1(new_n10291_), .A2(new_n10306_), .B1(new_n10307_), .B2(new_n10302_), .ZN(new_n10308_));
  NOR3_X1    g09302(.A1(new_n10294_), .A2(new_n10305_), .A3(new_n10308_), .ZN(new_n10309_));
  INV_X1     g09303(.I(\A[153] ), .ZN(new_n10310_));
  NOR2_X1    g09304(.A1(new_n10310_), .A2(\A[152] ), .ZN(new_n10311_));
  INV_X1     g09305(.I(\A[152] ), .ZN(new_n10312_));
  NOR2_X1    g09306(.A1(new_n10312_), .A2(\A[153] ), .ZN(new_n10313_));
  OAI21_X1   g09307(.A1(new_n10311_), .A2(new_n10313_), .B(\A[151] ), .ZN(new_n10314_));
  INV_X1     g09308(.I(\A[151] ), .ZN(new_n10315_));
  NAND2_X1   g09309(.A1(\A[152] ), .A2(\A[153] ), .ZN(new_n10316_));
  INV_X1     g09310(.I(new_n10316_), .ZN(new_n10317_));
  NOR2_X1    g09311(.A1(\A[152] ), .A2(\A[153] ), .ZN(new_n10318_));
  OAI21_X1   g09312(.A1(new_n10317_), .A2(new_n10318_), .B(new_n10315_), .ZN(new_n10319_));
  NAND2_X1   g09313(.A1(new_n10314_), .A2(new_n10319_), .ZN(new_n10320_));
  INV_X1     g09314(.I(\A[156] ), .ZN(new_n10321_));
  NOR2_X1    g09315(.A1(new_n10321_), .A2(\A[155] ), .ZN(new_n10322_));
  INV_X1     g09316(.I(\A[155] ), .ZN(new_n10323_));
  NOR2_X1    g09317(.A1(new_n10323_), .A2(\A[156] ), .ZN(new_n10324_));
  OAI21_X1   g09318(.A1(new_n10322_), .A2(new_n10324_), .B(\A[154] ), .ZN(new_n10325_));
  INV_X1     g09319(.I(\A[154] ), .ZN(new_n10326_));
  NAND2_X1   g09320(.A1(\A[155] ), .A2(\A[156] ), .ZN(new_n10327_));
  INV_X1     g09321(.I(new_n10327_), .ZN(new_n10328_));
  NOR2_X1    g09322(.A1(\A[155] ), .A2(\A[156] ), .ZN(new_n10329_));
  OAI21_X1   g09323(.A1(new_n10328_), .A2(new_n10329_), .B(new_n10326_), .ZN(new_n10330_));
  NAND2_X1   g09324(.A1(new_n10325_), .A2(new_n10330_), .ZN(new_n10331_));
  AOI21_X1   g09325(.A1(\A[152] ), .A2(\A[153] ), .B(\A[151] ), .ZN(new_n10332_));
  AOI21_X1   g09326(.A1(\A[155] ), .A2(\A[156] ), .B(\A[154] ), .ZN(new_n10333_));
  OAI22_X1   g09327(.A1(new_n10318_), .A2(new_n10332_), .B1(new_n10333_), .B2(new_n10329_), .ZN(new_n10334_));
  INV_X1     g09328(.I(new_n10334_), .ZN(new_n10335_));
  NAND3_X1   g09329(.A1(new_n10320_), .A2(new_n10331_), .A3(new_n10335_), .ZN(new_n10336_));
  NOR2_X1    g09330(.A1(new_n10309_), .A2(new_n10336_), .ZN(new_n10337_));
  NOR2_X1    g09331(.A1(new_n10287_), .A2(\A[158] ), .ZN(new_n10338_));
  NOR2_X1    g09332(.A1(new_n10285_), .A2(\A[159] ), .ZN(new_n10339_));
  OAI21_X1   g09333(.A1(new_n10338_), .A2(new_n10339_), .B(\A[157] ), .ZN(new_n10340_));
  INV_X1     g09334(.I(new_n10290_), .ZN(new_n10341_));
  OAI21_X1   g09335(.A1(new_n10341_), .A2(new_n10291_), .B(new_n10284_), .ZN(new_n10342_));
  NAND2_X1   g09336(.A1(new_n10340_), .A2(new_n10342_), .ZN(new_n10343_));
  NOR2_X1    g09337(.A1(new_n10298_), .A2(\A[161] ), .ZN(new_n10344_));
  NOR2_X1    g09338(.A1(new_n10296_), .A2(\A[162] ), .ZN(new_n10345_));
  OAI21_X1   g09339(.A1(new_n10344_), .A2(new_n10345_), .B(\A[160] ), .ZN(new_n10346_));
  INV_X1     g09340(.I(new_n10301_), .ZN(new_n10347_));
  OAI21_X1   g09341(.A1(new_n10347_), .A2(new_n10302_), .B(new_n10295_), .ZN(new_n10348_));
  NAND2_X1   g09342(.A1(new_n10346_), .A2(new_n10348_), .ZN(new_n10349_));
  INV_X1     g09343(.I(new_n10308_), .ZN(new_n10350_));
  NAND3_X1   g09344(.A1(new_n10343_), .A2(new_n10349_), .A3(new_n10350_), .ZN(new_n10351_));
  NAND2_X1   g09345(.A1(new_n10312_), .A2(\A[153] ), .ZN(new_n10352_));
  NAND2_X1   g09346(.A1(new_n10310_), .A2(\A[152] ), .ZN(new_n10353_));
  AOI21_X1   g09347(.A1(new_n10352_), .A2(new_n10353_), .B(new_n10315_), .ZN(new_n10354_));
  INV_X1     g09348(.I(new_n10318_), .ZN(new_n10355_));
  AOI21_X1   g09349(.A1(new_n10355_), .A2(new_n10316_), .B(\A[151] ), .ZN(new_n10356_));
  NOR2_X1    g09350(.A1(new_n10356_), .A2(new_n10354_), .ZN(new_n10357_));
  NAND2_X1   g09351(.A1(new_n10323_), .A2(\A[156] ), .ZN(new_n10358_));
  NAND2_X1   g09352(.A1(new_n10321_), .A2(\A[155] ), .ZN(new_n10359_));
  AOI21_X1   g09353(.A1(new_n10358_), .A2(new_n10359_), .B(new_n10326_), .ZN(new_n10360_));
  INV_X1     g09354(.I(new_n10329_), .ZN(new_n10361_));
  AOI21_X1   g09355(.A1(new_n10361_), .A2(new_n10327_), .B(\A[154] ), .ZN(new_n10362_));
  NOR2_X1    g09356(.A1(new_n10362_), .A2(new_n10360_), .ZN(new_n10363_));
  NOR3_X1    g09357(.A1(new_n10357_), .A2(new_n10363_), .A3(new_n10334_), .ZN(new_n10364_));
  NOR2_X1    g09358(.A1(new_n10364_), .A2(new_n10351_), .ZN(new_n10365_));
  OAI22_X1   g09359(.A1(new_n10281_), .A2(new_n10283_), .B1(new_n10337_), .B2(new_n10365_), .ZN(new_n10366_));
  NOR2_X1    g09360(.A1(new_n10231_), .A2(\A[170] ), .ZN(new_n10367_));
  NOR2_X1    g09361(.A1(new_n10229_), .A2(\A[171] ), .ZN(new_n10368_));
  OAI21_X1   g09362(.A1(new_n10367_), .A2(new_n10368_), .B(\A[169] ), .ZN(new_n10369_));
  INV_X1     g09363(.I(new_n10234_), .ZN(new_n10370_));
  OAI21_X1   g09364(.A1(new_n10370_), .A2(new_n10235_), .B(new_n10228_), .ZN(new_n10371_));
  NAND2_X1   g09365(.A1(new_n10369_), .A2(new_n10371_), .ZN(new_n10372_));
  NOR2_X1    g09366(.A1(new_n10242_), .A2(\A[173] ), .ZN(new_n10373_));
  NOR2_X1    g09367(.A1(new_n10240_), .A2(\A[174] ), .ZN(new_n10374_));
  OAI21_X1   g09368(.A1(new_n10373_), .A2(new_n10374_), .B(\A[172] ), .ZN(new_n10375_));
  INV_X1     g09369(.I(new_n10245_), .ZN(new_n10376_));
  OAI21_X1   g09370(.A1(new_n10376_), .A2(new_n10246_), .B(new_n10239_), .ZN(new_n10377_));
  NAND2_X1   g09371(.A1(new_n10375_), .A2(new_n10377_), .ZN(new_n10378_));
  INV_X1     g09372(.I(new_n10252_), .ZN(new_n10379_));
  NAND3_X1   g09373(.A1(new_n10372_), .A2(new_n10378_), .A3(new_n10379_), .ZN(new_n10380_));
  INV_X1     g09374(.I(new_n10280_), .ZN(new_n10381_));
  NAND2_X1   g09375(.A1(new_n10381_), .A2(new_n10380_), .ZN(new_n10382_));
  NAND2_X1   g09376(.A1(new_n10364_), .A2(new_n10351_), .ZN(new_n10383_));
  NAND2_X1   g09377(.A1(new_n10309_), .A2(new_n10336_), .ZN(new_n10384_));
  NAND4_X1   g09378(.A1(new_n10382_), .A2(new_n10383_), .A3(new_n10384_), .A4(new_n10282_), .ZN(new_n10385_));
  NAND2_X1   g09379(.A1(new_n10366_), .A2(new_n10385_), .ZN(new_n10386_));
  INV_X1     g09380(.I(\A[145] ), .ZN(new_n10387_));
  INV_X1     g09381(.I(\A[146] ), .ZN(new_n10388_));
  NAND2_X1   g09382(.A1(new_n10388_), .A2(\A[147] ), .ZN(new_n10389_));
  INV_X1     g09383(.I(\A[147] ), .ZN(new_n10390_));
  NAND2_X1   g09384(.A1(new_n10390_), .A2(\A[146] ), .ZN(new_n10391_));
  AOI21_X1   g09385(.A1(new_n10389_), .A2(new_n10391_), .B(new_n10387_), .ZN(new_n10392_));
  NAND2_X1   g09386(.A1(\A[146] ), .A2(\A[147] ), .ZN(new_n10393_));
  NOR2_X1    g09387(.A1(\A[146] ), .A2(\A[147] ), .ZN(new_n10394_));
  INV_X1     g09388(.I(new_n10394_), .ZN(new_n10395_));
  AOI21_X1   g09389(.A1(new_n10395_), .A2(new_n10393_), .B(\A[145] ), .ZN(new_n10396_));
  NOR2_X1    g09390(.A1(new_n10396_), .A2(new_n10392_), .ZN(new_n10397_));
  INV_X1     g09391(.I(\A[148] ), .ZN(new_n10398_));
  INV_X1     g09392(.I(\A[149] ), .ZN(new_n10399_));
  NAND2_X1   g09393(.A1(new_n10399_), .A2(\A[150] ), .ZN(new_n10400_));
  INV_X1     g09394(.I(\A[150] ), .ZN(new_n10401_));
  NAND2_X1   g09395(.A1(new_n10401_), .A2(\A[149] ), .ZN(new_n10402_));
  AOI21_X1   g09396(.A1(new_n10400_), .A2(new_n10402_), .B(new_n10398_), .ZN(new_n10403_));
  NAND2_X1   g09397(.A1(\A[149] ), .A2(\A[150] ), .ZN(new_n10404_));
  NOR2_X1    g09398(.A1(\A[149] ), .A2(\A[150] ), .ZN(new_n10405_));
  INV_X1     g09399(.I(new_n10405_), .ZN(new_n10406_));
  AOI21_X1   g09400(.A1(new_n10406_), .A2(new_n10404_), .B(\A[148] ), .ZN(new_n10407_));
  NOR2_X1    g09401(.A1(new_n10407_), .A2(new_n10403_), .ZN(new_n10408_));
  AOI21_X1   g09402(.A1(\A[146] ), .A2(\A[147] ), .B(\A[145] ), .ZN(new_n10409_));
  AOI21_X1   g09403(.A1(\A[149] ), .A2(\A[150] ), .B(\A[148] ), .ZN(new_n10410_));
  OAI22_X1   g09404(.A1(new_n10394_), .A2(new_n10409_), .B1(new_n10410_), .B2(new_n10405_), .ZN(new_n10411_));
  NOR3_X1    g09405(.A1(new_n10397_), .A2(new_n10408_), .A3(new_n10411_), .ZN(new_n10412_));
  INV_X1     g09406(.I(\A[141] ), .ZN(new_n10413_));
  NOR2_X1    g09407(.A1(new_n10413_), .A2(\A[140] ), .ZN(new_n10414_));
  INV_X1     g09408(.I(\A[140] ), .ZN(new_n10415_));
  NOR2_X1    g09409(.A1(new_n10415_), .A2(\A[141] ), .ZN(new_n10416_));
  OAI21_X1   g09410(.A1(new_n10414_), .A2(new_n10416_), .B(\A[139] ), .ZN(new_n10417_));
  INV_X1     g09411(.I(\A[139] ), .ZN(new_n10418_));
  NAND2_X1   g09412(.A1(\A[140] ), .A2(\A[141] ), .ZN(new_n10419_));
  INV_X1     g09413(.I(new_n10419_), .ZN(new_n10420_));
  NOR2_X1    g09414(.A1(\A[140] ), .A2(\A[141] ), .ZN(new_n10421_));
  OAI21_X1   g09415(.A1(new_n10420_), .A2(new_n10421_), .B(new_n10418_), .ZN(new_n10422_));
  NAND2_X1   g09416(.A1(new_n10417_), .A2(new_n10422_), .ZN(new_n10423_));
  INV_X1     g09417(.I(\A[144] ), .ZN(new_n10424_));
  NOR2_X1    g09418(.A1(new_n10424_), .A2(\A[143] ), .ZN(new_n10425_));
  INV_X1     g09419(.I(\A[143] ), .ZN(new_n10426_));
  NOR2_X1    g09420(.A1(new_n10426_), .A2(\A[144] ), .ZN(new_n10427_));
  OAI21_X1   g09421(.A1(new_n10425_), .A2(new_n10427_), .B(\A[142] ), .ZN(new_n10428_));
  INV_X1     g09422(.I(\A[142] ), .ZN(new_n10429_));
  NAND2_X1   g09423(.A1(\A[143] ), .A2(\A[144] ), .ZN(new_n10430_));
  INV_X1     g09424(.I(new_n10430_), .ZN(new_n10431_));
  NOR2_X1    g09425(.A1(\A[143] ), .A2(\A[144] ), .ZN(new_n10432_));
  OAI21_X1   g09426(.A1(new_n10431_), .A2(new_n10432_), .B(new_n10429_), .ZN(new_n10433_));
  NAND2_X1   g09427(.A1(new_n10428_), .A2(new_n10433_), .ZN(new_n10434_));
  AOI21_X1   g09428(.A1(\A[140] ), .A2(\A[141] ), .B(\A[139] ), .ZN(new_n10435_));
  NOR2_X1    g09429(.A1(new_n10435_), .A2(new_n10421_), .ZN(new_n10436_));
  AOI21_X1   g09430(.A1(\A[143] ), .A2(\A[144] ), .B(\A[142] ), .ZN(new_n10437_));
  NOR2_X1    g09431(.A1(new_n10437_), .A2(new_n10432_), .ZN(new_n10438_));
  NOR2_X1    g09432(.A1(new_n10436_), .A2(new_n10438_), .ZN(new_n10439_));
  NAND3_X1   g09433(.A1(new_n10423_), .A2(new_n10434_), .A3(new_n10439_), .ZN(new_n10440_));
  NOR2_X1    g09434(.A1(new_n10412_), .A2(new_n10440_), .ZN(new_n10441_));
  NOR2_X1    g09435(.A1(new_n10390_), .A2(\A[146] ), .ZN(new_n10442_));
  NOR2_X1    g09436(.A1(new_n10388_), .A2(\A[147] ), .ZN(new_n10443_));
  OAI21_X1   g09437(.A1(new_n10442_), .A2(new_n10443_), .B(\A[145] ), .ZN(new_n10444_));
  INV_X1     g09438(.I(new_n10393_), .ZN(new_n10445_));
  OAI21_X1   g09439(.A1(new_n10445_), .A2(new_n10394_), .B(new_n10387_), .ZN(new_n10446_));
  NAND2_X1   g09440(.A1(new_n10444_), .A2(new_n10446_), .ZN(new_n10447_));
  NOR2_X1    g09441(.A1(new_n10401_), .A2(\A[149] ), .ZN(new_n10448_));
  NOR2_X1    g09442(.A1(new_n10399_), .A2(\A[150] ), .ZN(new_n10449_));
  OAI21_X1   g09443(.A1(new_n10448_), .A2(new_n10449_), .B(\A[148] ), .ZN(new_n10450_));
  INV_X1     g09444(.I(new_n10404_), .ZN(new_n10451_));
  OAI21_X1   g09445(.A1(new_n10451_), .A2(new_n10405_), .B(new_n10398_), .ZN(new_n10452_));
  NAND2_X1   g09446(.A1(new_n10450_), .A2(new_n10452_), .ZN(new_n10453_));
  NOR2_X1    g09447(.A1(new_n10409_), .A2(new_n10394_), .ZN(new_n10454_));
  NOR2_X1    g09448(.A1(new_n10410_), .A2(new_n10405_), .ZN(new_n10455_));
  NOR2_X1    g09449(.A1(new_n10454_), .A2(new_n10455_), .ZN(new_n10456_));
  NAND3_X1   g09450(.A1(new_n10453_), .A2(new_n10447_), .A3(new_n10456_), .ZN(new_n10457_));
  NAND2_X1   g09451(.A1(new_n10415_), .A2(\A[141] ), .ZN(new_n10458_));
  NAND2_X1   g09452(.A1(new_n10413_), .A2(\A[140] ), .ZN(new_n10459_));
  AOI21_X1   g09453(.A1(new_n10458_), .A2(new_n10459_), .B(new_n10418_), .ZN(new_n10460_));
  INV_X1     g09454(.I(new_n10421_), .ZN(new_n10461_));
  AOI21_X1   g09455(.A1(new_n10461_), .A2(new_n10419_), .B(\A[139] ), .ZN(new_n10462_));
  NOR2_X1    g09456(.A1(new_n10462_), .A2(new_n10460_), .ZN(new_n10463_));
  NAND2_X1   g09457(.A1(new_n10426_), .A2(\A[144] ), .ZN(new_n10464_));
  NAND2_X1   g09458(.A1(new_n10424_), .A2(\A[143] ), .ZN(new_n10465_));
  AOI21_X1   g09459(.A1(new_n10464_), .A2(new_n10465_), .B(new_n10429_), .ZN(new_n10466_));
  INV_X1     g09460(.I(new_n10432_), .ZN(new_n10467_));
  AOI21_X1   g09461(.A1(new_n10467_), .A2(new_n10430_), .B(\A[142] ), .ZN(new_n10468_));
  NOR2_X1    g09462(.A1(new_n10468_), .A2(new_n10466_), .ZN(new_n10469_));
  OAI22_X1   g09463(.A1(new_n10421_), .A2(new_n10435_), .B1(new_n10437_), .B2(new_n10432_), .ZN(new_n10470_));
  NOR3_X1    g09464(.A1(new_n10463_), .A2(new_n10469_), .A3(new_n10470_), .ZN(new_n10471_));
  NOR2_X1    g09465(.A1(new_n10471_), .A2(new_n10457_), .ZN(new_n10472_));
  INV_X1     g09466(.I(\A[133] ), .ZN(new_n10473_));
  INV_X1     g09467(.I(\A[134] ), .ZN(new_n10474_));
  NAND2_X1   g09468(.A1(new_n10474_), .A2(\A[135] ), .ZN(new_n10475_));
  INV_X1     g09469(.I(\A[135] ), .ZN(new_n10476_));
  NAND2_X1   g09470(.A1(new_n10476_), .A2(\A[134] ), .ZN(new_n10477_));
  AOI21_X1   g09471(.A1(new_n10475_), .A2(new_n10477_), .B(new_n10473_), .ZN(new_n10478_));
  NAND2_X1   g09472(.A1(\A[134] ), .A2(\A[135] ), .ZN(new_n10479_));
  NOR2_X1    g09473(.A1(\A[134] ), .A2(\A[135] ), .ZN(new_n10480_));
  INV_X1     g09474(.I(new_n10480_), .ZN(new_n10481_));
  AOI21_X1   g09475(.A1(new_n10481_), .A2(new_n10479_), .B(\A[133] ), .ZN(new_n10482_));
  NOR2_X1    g09476(.A1(new_n10482_), .A2(new_n10478_), .ZN(new_n10483_));
  INV_X1     g09477(.I(\A[136] ), .ZN(new_n10484_));
  INV_X1     g09478(.I(\A[137] ), .ZN(new_n10485_));
  NAND2_X1   g09479(.A1(new_n10485_), .A2(\A[138] ), .ZN(new_n10486_));
  INV_X1     g09480(.I(\A[138] ), .ZN(new_n10487_));
  NAND2_X1   g09481(.A1(new_n10487_), .A2(\A[137] ), .ZN(new_n10488_));
  AOI21_X1   g09482(.A1(new_n10486_), .A2(new_n10488_), .B(new_n10484_), .ZN(new_n10489_));
  NAND2_X1   g09483(.A1(\A[137] ), .A2(\A[138] ), .ZN(new_n10490_));
  NOR2_X1    g09484(.A1(\A[137] ), .A2(\A[138] ), .ZN(new_n10491_));
  INV_X1     g09485(.I(new_n10491_), .ZN(new_n10492_));
  AOI21_X1   g09486(.A1(new_n10492_), .A2(new_n10490_), .B(\A[136] ), .ZN(new_n10493_));
  NOR2_X1    g09487(.A1(new_n10493_), .A2(new_n10489_), .ZN(new_n10494_));
  AOI21_X1   g09488(.A1(\A[134] ), .A2(\A[135] ), .B(\A[133] ), .ZN(new_n10495_));
  AOI21_X1   g09489(.A1(\A[137] ), .A2(\A[138] ), .B(\A[136] ), .ZN(new_n10496_));
  OAI22_X1   g09490(.A1(new_n10480_), .A2(new_n10495_), .B1(new_n10496_), .B2(new_n10491_), .ZN(new_n10497_));
  NOR3_X1    g09491(.A1(new_n10483_), .A2(new_n10494_), .A3(new_n10497_), .ZN(new_n10498_));
  INV_X1     g09492(.I(\A[129] ), .ZN(new_n10499_));
  NOR2_X1    g09493(.A1(new_n10499_), .A2(\A[128] ), .ZN(new_n10500_));
  INV_X1     g09494(.I(\A[128] ), .ZN(new_n10501_));
  NOR2_X1    g09495(.A1(new_n10501_), .A2(\A[129] ), .ZN(new_n10502_));
  OAI21_X1   g09496(.A1(new_n10500_), .A2(new_n10502_), .B(\A[127] ), .ZN(new_n10503_));
  INV_X1     g09497(.I(\A[127] ), .ZN(new_n10504_));
  NAND2_X1   g09498(.A1(\A[128] ), .A2(\A[129] ), .ZN(new_n10505_));
  INV_X1     g09499(.I(new_n10505_), .ZN(new_n10506_));
  NOR2_X1    g09500(.A1(\A[128] ), .A2(\A[129] ), .ZN(new_n10507_));
  OAI21_X1   g09501(.A1(new_n10506_), .A2(new_n10507_), .B(new_n10504_), .ZN(new_n10508_));
  NAND2_X1   g09502(.A1(new_n10503_), .A2(new_n10508_), .ZN(new_n10509_));
  INV_X1     g09503(.I(\A[132] ), .ZN(new_n10510_));
  NOR2_X1    g09504(.A1(new_n10510_), .A2(\A[131] ), .ZN(new_n10511_));
  INV_X1     g09505(.I(\A[131] ), .ZN(new_n10512_));
  NOR2_X1    g09506(.A1(new_n10512_), .A2(\A[132] ), .ZN(new_n10513_));
  OAI21_X1   g09507(.A1(new_n10511_), .A2(new_n10513_), .B(\A[130] ), .ZN(new_n10514_));
  INV_X1     g09508(.I(\A[130] ), .ZN(new_n10515_));
  NAND2_X1   g09509(.A1(\A[131] ), .A2(\A[132] ), .ZN(new_n10516_));
  INV_X1     g09510(.I(new_n10516_), .ZN(new_n10517_));
  NOR2_X1    g09511(.A1(\A[131] ), .A2(\A[132] ), .ZN(new_n10518_));
  OAI21_X1   g09512(.A1(new_n10517_), .A2(new_n10518_), .B(new_n10515_), .ZN(new_n10519_));
  NAND2_X1   g09513(.A1(new_n10514_), .A2(new_n10519_), .ZN(new_n10520_));
  AOI21_X1   g09514(.A1(\A[128] ), .A2(\A[129] ), .B(\A[127] ), .ZN(new_n10521_));
  AOI21_X1   g09515(.A1(\A[131] ), .A2(\A[132] ), .B(\A[130] ), .ZN(new_n10522_));
  OAI22_X1   g09516(.A1(new_n10507_), .A2(new_n10521_), .B1(new_n10522_), .B2(new_n10518_), .ZN(new_n10523_));
  INV_X1     g09517(.I(new_n10523_), .ZN(new_n10524_));
  NAND3_X1   g09518(.A1(new_n10509_), .A2(new_n10520_), .A3(new_n10524_), .ZN(new_n10525_));
  NOR2_X1    g09519(.A1(new_n10498_), .A2(new_n10525_), .ZN(new_n10526_));
  NOR2_X1    g09520(.A1(new_n10476_), .A2(\A[134] ), .ZN(new_n10527_));
  NOR2_X1    g09521(.A1(new_n10474_), .A2(\A[135] ), .ZN(new_n10528_));
  OAI21_X1   g09522(.A1(new_n10527_), .A2(new_n10528_), .B(\A[133] ), .ZN(new_n10529_));
  INV_X1     g09523(.I(new_n10479_), .ZN(new_n10530_));
  OAI21_X1   g09524(.A1(new_n10530_), .A2(new_n10480_), .B(new_n10473_), .ZN(new_n10531_));
  NAND2_X1   g09525(.A1(new_n10529_), .A2(new_n10531_), .ZN(new_n10532_));
  NOR2_X1    g09526(.A1(new_n10487_), .A2(\A[137] ), .ZN(new_n10533_));
  NOR2_X1    g09527(.A1(new_n10485_), .A2(\A[138] ), .ZN(new_n10534_));
  OAI21_X1   g09528(.A1(new_n10533_), .A2(new_n10534_), .B(\A[136] ), .ZN(new_n10535_));
  AND2_X2    g09529(.A1(\A[137] ), .A2(\A[138] ), .Z(new_n10536_));
  OAI21_X1   g09530(.A1(new_n10536_), .A2(new_n10491_), .B(new_n10484_), .ZN(new_n10537_));
  NAND2_X1   g09531(.A1(new_n10535_), .A2(new_n10537_), .ZN(new_n10538_));
  NOR2_X1    g09532(.A1(new_n10495_), .A2(new_n10480_), .ZN(new_n10539_));
  NOR2_X1    g09533(.A1(new_n10496_), .A2(new_n10491_), .ZN(new_n10540_));
  NOR2_X1    g09534(.A1(new_n10539_), .A2(new_n10540_), .ZN(new_n10541_));
  NAND3_X1   g09535(.A1(new_n10532_), .A2(new_n10538_), .A3(new_n10541_), .ZN(new_n10542_));
  NAND2_X1   g09536(.A1(new_n10501_), .A2(\A[129] ), .ZN(new_n10543_));
  NAND2_X1   g09537(.A1(new_n10499_), .A2(\A[128] ), .ZN(new_n10544_));
  AOI21_X1   g09538(.A1(new_n10543_), .A2(new_n10544_), .B(new_n10504_), .ZN(new_n10545_));
  INV_X1     g09539(.I(new_n10507_), .ZN(new_n10546_));
  AOI21_X1   g09540(.A1(new_n10546_), .A2(new_n10505_), .B(\A[127] ), .ZN(new_n10547_));
  NOR2_X1    g09541(.A1(new_n10547_), .A2(new_n10545_), .ZN(new_n10548_));
  NAND2_X1   g09542(.A1(new_n10512_), .A2(\A[132] ), .ZN(new_n10549_));
  NAND2_X1   g09543(.A1(new_n10510_), .A2(\A[131] ), .ZN(new_n10550_));
  AOI21_X1   g09544(.A1(new_n10549_), .A2(new_n10550_), .B(new_n10515_), .ZN(new_n10551_));
  INV_X1     g09545(.I(new_n10518_), .ZN(new_n10552_));
  AOI21_X1   g09546(.A1(new_n10552_), .A2(new_n10516_), .B(\A[130] ), .ZN(new_n10553_));
  NOR2_X1    g09547(.A1(new_n10553_), .A2(new_n10551_), .ZN(new_n10554_));
  NOR3_X1    g09548(.A1(new_n10548_), .A2(new_n10554_), .A3(new_n10523_), .ZN(new_n10555_));
  NOR2_X1    g09549(.A1(new_n10555_), .A2(new_n10542_), .ZN(new_n10556_));
  OAI22_X1   g09550(.A1(new_n10441_), .A2(new_n10472_), .B1(new_n10526_), .B2(new_n10556_), .ZN(new_n10557_));
  NAND2_X1   g09551(.A1(new_n10471_), .A2(new_n10457_), .ZN(new_n10558_));
  NAND2_X1   g09552(.A1(new_n10412_), .A2(new_n10440_), .ZN(new_n10559_));
  NAND2_X1   g09553(.A1(new_n10555_), .A2(new_n10542_), .ZN(new_n10560_));
  NAND2_X1   g09554(.A1(new_n10498_), .A2(new_n10525_), .ZN(new_n10561_));
  NAND4_X1   g09555(.A1(new_n10558_), .A2(new_n10559_), .A3(new_n10561_), .A4(new_n10560_), .ZN(new_n10562_));
  NAND2_X1   g09556(.A1(new_n10557_), .A2(new_n10562_), .ZN(new_n10563_));
  NAND2_X1   g09557(.A1(new_n10386_), .A2(new_n10563_), .ZN(new_n10564_));
  NOR2_X1    g09558(.A1(new_n10386_), .A2(new_n10563_), .ZN(new_n10565_));
  INV_X1     g09559(.I(new_n10565_), .ZN(new_n10566_));
  NAND2_X1   g09560(.A1(new_n10566_), .A2(new_n10564_), .ZN(new_n10567_));
  INV_X1     g09561(.I(\A[123] ), .ZN(new_n10568_));
  NOR2_X1    g09562(.A1(new_n10568_), .A2(\A[122] ), .ZN(new_n10569_));
  INV_X1     g09563(.I(\A[122] ), .ZN(new_n10570_));
  NOR2_X1    g09564(.A1(new_n10570_), .A2(\A[123] ), .ZN(new_n10571_));
  OAI21_X1   g09565(.A1(new_n10569_), .A2(new_n10571_), .B(\A[121] ), .ZN(new_n10572_));
  INV_X1     g09566(.I(\A[121] ), .ZN(new_n10573_));
  NAND2_X1   g09567(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n10574_));
  INV_X1     g09568(.I(new_n10574_), .ZN(new_n10575_));
  NOR2_X1    g09569(.A1(\A[122] ), .A2(\A[123] ), .ZN(new_n10576_));
  OAI21_X1   g09570(.A1(new_n10575_), .A2(new_n10576_), .B(new_n10573_), .ZN(new_n10577_));
  NAND2_X1   g09571(.A1(new_n10572_), .A2(new_n10577_), .ZN(new_n10578_));
  INV_X1     g09572(.I(\A[126] ), .ZN(new_n10579_));
  NOR2_X1    g09573(.A1(new_n10579_), .A2(\A[125] ), .ZN(new_n10580_));
  INV_X1     g09574(.I(\A[125] ), .ZN(new_n10581_));
  NOR2_X1    g09575(.A1(new_n10581_), .A2(\A[126] ), .ZN(new_n10582_));
  OAI21_X1   g09576(.A1(new_n10580_), .A2(new_n10582_), .B(\A[124] ), .ZN(new_n10583_));
  INV_X1     g09577(.I(\A[124] ), .ZN(new_n10584_));
  NAND2_X1   g09578(.A1(\A[125] ), .A2(\A[126] ), .ZN(new_n10585_));
  INV_X1     g09579(.I(new_n10585_), .ZN(new_n10586_));
  NOR2_X1    g09580(.A1(\A[125] ), .A2(\A[126] ), .ZN(new_n10587_));
  OAI21_X1   g09581(.A1(new_n10586_), .A2(new_n10587_), .B(new_n10584_), .ZN(new_n10588_));
  NAND2_X1   g09582(.A1(new_n10583_), .A2(new_n10588_), .ZN(new_n10589_));
  AOI21_X1   g09583(.A1(\A[122] ), .A2(\A[123] ), .B(\A[121] ), .ZN(new_n10590_));
  NOR2_X1    g09584(.A1(new_n10590_), .A2(new_n10576_), .ZN(new_n10591_));
  AOI21_X1   g09585(.A1(\A[125] ), .A2(\A[126] ), .B(\A[124] ), .ZN(new_n10592_));
  NOR2_X1    g09586(.A1(new_n10592_), .A2(new_n10587_), .ZN(new_n10593_));
  NOR2_X1    g09587(.A1(new_n10591_), .A2(new_n10593_), .ZN(new_n10594_));
  NAND3_X1   g09588(.A1(new_n10578_), .A2(new_n10589_), .A3(new_n10594_), .ZN(new_n10595_));
  INV_X1     g09589(.I(\A[115] ), .ZN(new_n10596_));
  INV_X1     g09590(.I(\A[116] ), .ZN(new_n10597_));
  NAND2_X1   g09591(.A1(new_n10597_), .A2(\A[117] ), .ZN(new_n10598_));
  INV_X1     g09592(.I(\A[117] ), .ZN(new_n10599_));
  NAND2_X1   g09593(.A1(new_n10599_), .A2(\A[116] ), .ZN(new_n10600_));
  AOI21_X1   g09594(.A1(new_n10598_), .A2(new_n10600_), .B(new_n10596_), .ZN(new_n10601_));
  NAND2_X1   g09595(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n10602_));
  OR2_X2     g09596(.A1(\A[116] ), .A2(\A[117] ), .Z(new_n10603_));
  AOI21_X1   g09597(.A1(new_n10603_), .A2(new_n10602_), .B(\A[115] ), .ZN(new_n10604_));
  NOR2_X1    g09598(.A1(new_n10601_), .A2(new_n10604_), .ZN(new_n10605_));
  INV_X1     g09599(.I(\A[118] ), .ZN(new_n10606_));
  INV_X1     g09600(.I(\A[119] ), .ZN(new_n10607_));
  NAND2_X1   g09601(.A1(new_n10607_), .A2(\A[120] ), .ZN(new_n10608_));
  INV_X1     g09602(.I(\A[120] ), .ZN(new_n10609_));
  NAND2_X1   g09603(.A1(new_n10609_), .A2(\A[119] ), .ZN(new_n10610_));
  AOI21_X1   g09604(.A1(new_n10608_), .A2(new_n10610_), .B(new_n10606_), .ZN(new_n10611_));
  NAND2_X1   g09605(.A1(\A[119] ), .A2(\A[120] ), .ZN(new_n10612_));
  NOR2_X1    g09606(.A1(\A[119] ), .A2(\A[120] ), .ZN(new_n10613_));
  INV_X1     g09607(.I(new_n10613_), .ZN(new_n10614_));
  AOI21_X1   g09608(.A1(new_n10614_), .A2(new_n10612_), .B(\A[118] ), .ZN(new_n10615_));
  NOR2_X1    g09609(.A1(new_n10615_), .A2(new_n10611_), .ZN(new_n10616_));
  NOR2_X1    g09610(.A1(\A[116] ), .A2(\A[117] ), .ZN(new_n10617_));
  AOI21_X1   g09611(.A1(\A[116] ), .A2(\A[117] ), .B(\A[115] ), .ZN(new_n10618_));
  AOI21_X1   g09612(.A1(\A[119] ), .A2(\A[120] ), .B(\A[118] ), .ZN(new_n10619_));
  OAI22_X1   g09613(.A1(new_n10617_), .A2(new_n10618_), .B1(new_n10619_), .B2(new_n10613_), .ZN(new_n10620_));
  NOR3_X1    g09614(.A1(new_n10616_), .A2(new_n10605_), .A3(new_n10620_), .ZN(new_n10621_));
  NAND2_X1   g09615(.A1(new_n10595_), .A2(new_n10621_), .ZN(new_n10622_));
  NAND2_X1   g09616(.A1(new_n10570_), .A2(\A[123] ), .ZN(new_n10623_));
  NAND2_X1   g09617(.A1(new_n10568_), .A2(\A[122] ), .ZN(new_n10624_));
  AOI21_X1   g09618(.A1(new_n10623_), .A2(new_n10624_), .B(new_n10573_), .ZN(new_n10625_));
  INV_X1     g09619(.I(new_n10576_), .ZN(new_n10626_));
  AOI21_X1   g09620(.A1(new_n10626_), .A2(new_n10574_), .B(\A[121] ), .ZN(new_n10627_));
  NOR2_X1    g09621(.A1(new_n10627_), .A2(new_n10625_), .ZN(new_n10628_));
  NAND2_X1   g09622(.A1(new_n10581_), .A2(\A[126] ), .ZN(new_n10629_));
  NAND2_X1   g09623(.A1(new_n10579_), .A2(\A[125] ), .ZN(new_n10630_));
  AOI21_X1   g09624(.A1(new_n10629_), .A2(new_n10630_), .B(new_n10584_), .ZN(new_n10631_));
  INV_X1     g09625(.I(new_n10587_), .ZN(new_n10632_));
  AOI21_X1   g09626(.A1(new_n10632_), .A2(new_n10585_), .B(\A[124] ), .ZN(new_n10633_));
  NOR2_X1    g09627(.A1(new_n10633_), .A2(new_n10631_), .ZN(new_n10634_));
  OAI22_X1   g09628(.A1(new_n10576_), .A2(new_n10590_), .B1(new_n10592_), .B2(new_n10587_), .ZN(new_n10635_));
  NOR3_X1    g09629(.A1(new_n10628_), .A2(new_n10634_), .A3(new_n10635_), .ZN(new_n10636_));
  NOR2_X1    g09630(.A1(new_n10599_), .A2(\A[116] ), .ZN(new_n10637_));
  NOR2_X1    g09631(.A1(new_n10597_), .A2(\A[117] ), .ZN(new_n10638_));
  OAI21_X1   g09632(.A1(new_n10637_), .A2(new_n10638_), .B(\A[115] ), .ZN(new_n10639_));
  AND2_X2    g09633(.A1(\A[116] ), .A2(\A[117] ), .Z(new_n10640_));
  OAI21_X1   g09634(.A1(new_n10640_), .A2(new_n10617_), .B(new_n10596_), .ZN(new_n10641_));
  NAND2_X1   g09635(.A1(new_n10639_), .A2(new_n10641_), .ZN(new_n10642_));
  NOR2_X1    g09636(.A1(new_n10609_), .A2(\A[119] ), .ZN(new_n10643_));
  NOR2_X1    g09637(.A1(new_n10607_), .A2(\A[120] ), .ZN(new_n10644_));
  OAI21_X1   g09638(.A1(new_n10643_), .A2(new_n10644_), .B(\A[118] ), .ZN(new_n10645_));
  INV_X1     g09639(.I(new_n10612_), .ZN(new_n10646_));
  OAI21_X1   g09640(.A1(new_n10646_), .A2(new_n10613_), .B(new_n10606_), .ZN(new_n10647_));
  NAND2_X1   g09641(.A1(new_n10645_), .A2(new_n10647_), .ZN(new_n10648_));
  INV_X1     g09642(.I(new_n10620_), .ZN(new_n10649_));
  NAND3_X1   g09643(.A1(new_n10648_), .A2(new_n10642_), .A3(new_n10649_), .ZN(new_n10650_));
  NAND2_X1   g09644(.A1(new_n10636_), .A2(new_n10650_), .ZN(new_n10651_));
  NAND2_X1   g09645(.A1(new_n10622_), .A2(new_n10651_), .ZN(new_n10652_));
  INV_X1     g09646(.I(\A[111] ), .ZN(new_n10653_));
  NOR2_X1    g09647(.A1(new_n10653_), .A2(\A[110] ), .ZN(new_n10654_));
  INV_X1     g09648(.I(\A[110] ), .ZN(new_n10655_));
  NOR2_X1    g09649(.A1(new_n10655_), .A2(\A[111] ), .ZN(new_n10656_));
  OAI21_X1   g09650(.A1(new_n10654_), .A2(new_n10656_), .B(\A[109] ), .ZN(new_n10657_));
  INV_X1     g09651(.I(\A[109] ), .ZN(new_n10658_));
  NAND2_X1   g09652(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n10659_));
  INV_X1     g09653(.I(new_n10659_), .ZN(new_n10660_));
  NOR2_X1    g09654(.A1(\A[110] ), .A2(\A[111] ), .ZN(new_n10661_));
  OAI21_X1   g09655(.A1(new_n10660_), .A2(new_n10661_), .B(new_n10658_), .ZN(new_n10662_));
  NAND2_X1   g09656(.A1(new_n10657_), .A2(new_n10662_), .ZN(new_n10663_));
  INV_X1     g09657(.I(\A[114] ), .ZN(new_n10664_));
  NOR2_X1    g09658(.A1(new_n10664_), .A2(\A[113] ), .ZN(new_n10665_));
  INV_X1     g09659(.I(\A[113] ), .ZN(new_n10666_));
  NOR2_X1    g09660(.A1(new_n10666_), .A2(\A[114] ), .ZN(new_n10667_));
  OAI21_X1   g09661(.A1(new_n10665_), .A2(new_n10667_), .B(\A[112] ), .ZN(new_n10668_));
  INV_X1     g09662(.I(\A[112] ), .ZN(new_n10669_));
  AND2_X2    g09663(.A1(\A[113] ), .A2(\A[114] ), .Z(new_n10670_));
  NOR2_X1    g09664(.A1(\A[113] ), .A2(\A[114] ), .ZN(new_n10671_));
  OAI21_X1   g09665(.A1(new_n10670_), .A2(new_n10671_), .B(new_n10669_), .ZN(new_n10672_));
  NAND2_X1   g09666(.A1(new_n10668_), .A2(new_n10672_), .ZN(new_n10673_));
  AOI21_X1   g09667(.A1(\A[110] ), .A2(\A[111] ), .B(\A[109] ), .ZN(new_n10674_));
  NOR2_X1    g09668(.A1(new_n10674_), .A2(new_n10661_), .ZN(new_n10675_));
  AOI21_X1   g09669(.A1(\A[113] ), .A2(\A[114] ), .B(\A[112] ), .ZN(new_n10676_));
  NOR2_X1    g09670(.A1(new_n10676_), .A2(new_n10671_), .ZN(new_n10677_));
  NOR2_X1    g09671(.A1(new_n10675_), .A2(new_n10677_), .ZN(new_n10678_));
  NAND3_X1   g09672(.A1(new_n10663_), .A2(new_n10673_), .A3(new_n10678_), .ZN(new_n10679_));
  INV_X1     g09673(.I(\A[103] ), .ZN(new_n10680_));
  INV_X1     g09674(.I(\A[104] ), .ZN(new_n10681_));
  NAND2_X1   g09675(.A1(new_n10681_), .A2(\A[105] ), .ZN(new_n10682_));
  INV_X1     g09676(.I(\A[105] ), .ZN(new_n10683_));
  NAND2_X1   g09677(.A1(new_n10683_), .A2(\A[104] ), .ZN(new_n10684_));
  AOI21_X1   g09678(.A1(new_n10682_), .A2(new_n10684_), .B(new_n10680_), .ZN(new_n10685_));
  NAND2_X1   g09679(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n10686_));
  NOR2_X1    g09680(.A1(\A[104] ), .A2(\A[105] ), .ZN(new_n10687_));
  INV_X1     g09681(.I(new_n10687_), .ZN(new_n10688_));
  AOI21_X1   g09682(.A1(new_n10688_), .A2(new_n10686_), .B(\A[103] ), .ZN(new_n10689_));
  NOR2_X1    g09683(.A1(new_n10689_), .A2(new_n10685_), .ZN(new_n10690_));
  INV_X1     g09684(.I(\A[106] ), .ZN(new_n10691_));
  INV_X1     g09685(.I(\A[107] ), .ZN(new_n10692_));
  NAND2_X1   g09686(.A1(new_n10692_), .A2(\A[108] ), .ZN(new_n10693_));
  INV_X1     g09687(.I(\A[108] ), .ZN(new_n10694_));
  NAND2_X1   g09688(.A1(new_n10694_), .A2(\A[107] ), .ZN(new_n10695_));
  AOI21_X1   g09689(.A1(new_n10693_), .A2(new_n10695_), .B(new_n10691_), .ZN(new_n10696_));
  NAND2_X1   g09690(.A1(\A[107] ), .A2(\A[108] ), .ZN(new_n10697_));
  NOR2_X1    g09691(.A1(\A[107] ), .A2(\A[108] ), .ZN(new_n10698_));
  INV_X1     g09692(.I(new_n10698_), .ZN(new_n10699_));
  AOI21_X1   g09693(.A1(new_n10699_), .A2(new_n10697_), .B(\A[106] ), .ZN(new_n10700_));
  NOR2_X1    g09694(.A1(new_n10700_), .A2(new_n10696_), .ZN(new_n10701_));
  AOI21_X1   g09695(.A1(\A[104] ), .A2(\A[105] ), .B(\A[103] ), .ZN(new_n10702_));
  AOI21_X1   g09696(.A1(\A[107] ), .A2(\A[108] ), .B(\A[106] ), .ZN(new_n10703_));
  OAI22_X1   g09697(.A1(new_n10687_), .A2(new_n10702_), .B1(new_n10703_), .B2(new_n10698_), .ZN(new_n10704_));
  NOR3_X1    g09698(.A1(new_n10690_), .A2(new_n10701_), .A3(new_n10704_), .ZN(new_n10705_));
  NAND2_X1   g09699(.A1(new_n10705_), .A2(new_n10679_), .ZN(new_n10706_));
  NAND2_X1   g09700(.A1(new_n10655_), .A2(\A[111] ), .ZN(new_n10707_));
  NAND2_X1   g09701(.A1(new_n10653_), .A2(\A[110] ), .ZN(new_n10708_));
  AOI21_X1   g09702(.A1(new_n10707_), .A2(new_n10708_), .B(new_n10658_), .ZN(new_n10709_));
  INV_X1     g09703(.I(new_n10661_), .ZN(new_n10710_));
  AOI21_X1   g09704(.A1(new_n10710_), .A2(new_n10659_), .B(\A[109] ), .ZN(new_n10711_));
  NOR2_X1    g09705(.A1(new_n10711_), .A2(new_n10709_), .ZN(new_n10712_));
  NAND2_X1   g09706(.A1(new_n10666_), .A2(\A[114] ), .ZN(new_n10713_));
  NAND2_X1   g09707(.A1(new_n10664_), .A2(\A[113] ), .ZN(new_n10714_));
  AOI21_X1   g09708(.A1(new_n10713_), .A2(new_n10714_), .B(new_n10669_), .ZN(new_n10715_));
  NAND2_X1   g09709(.A1(\A[113] ), .A2(\A[114] ), .ZN(new_n10716_));
  INV_X1     g09710(.I(new_n10671_), .ZN(new_n10717_));
  AOI21_X1   g09711(.A1(new_n10717_), .A2(new_n10716_), .B(\A[112] ), .ZN(new_n10718_));
  NOR2_X1    g09712(.A1(new_n10718_), .A2(new_n10715_), .ZN(new_n10719_));
  OAI22_X1   g09713(.A1(new_n10661_), .A2(new_n10674_), .B1(new_n10676_), .B2(new_n10671_), .ZN(new_n10720_));
  NOR3_X1    g09714(.A1(new_n10712_), .A2(new_n10719_), .A3(new_n10720_), .ZN(new_n10721_));
  NOR2_X1    g09715(.A1(new_n10683_), .A2(\A[104] ), .ZN(new_n10722_));
  NOR2_X1    g09716(.A1(new_n10681_), .A2(\A[105] ), .ZN(new_n10723_));
  OAI21_X1   g09717(.A1(new_n10722_), .A2(new_n10723_), .B(\A[103] ), .ZN(new_n10724_));
  INV_X1     g09718(.I(new_n10686_), .ZN(new_n10725_));
  OAI21_X1   g09719(.A1(new_n10725_), .A2(new_n10687_), .B(new_n10680_), .ZN(new_n10726_));
  NAND2_X1   g09720(.A1(new_n10724_), .A2(new_n10726_), .ZN(new_n10727_));
  NOR2_X1    g09721(.A1(new_n10694_), .A2(\A[107] ), .ZN(new_n10728_));
  NOR2_X1    g09722(.A1(new_n10692_), .A2(\A[108] ), .ZN(new_n10729_));
  OAI21_X1   g09723(.A1(new_n10728_), .A2(new_n10729_), .B(\A[106] ), .ZN(new_n10730_));
  INV_X1     g09724(.I(new_n10697_), .ZN(new_n10731_));
  OAI21_X1   g09725(.A1(new_n10731_), .A2(new_n10698_), .B(new_n10691_), .ZN(new_n10732_));
  NAND2_X1   g09726(.A1(new_n10730_), .A2(new_n10732_), .ZN(new_n10733_));
  INV_X1     g09727(.I(new_n10704_), .ZN(new_n10734_));
  NAND3_X1   g09728(.A1(new_n10727_), .A2(new_n10733_), .A3(new_n10734_), .ZN(new_n10735_));
  NAND2_X1   g09729(.A1(new_n10721_), .A2(new_n10735_), .ZN(new_n10736_));
  NAND2_X1   g09730(.A1(new_n10736_), .A2(new_n10706_), .ZN(new_n10737_));
  NAND2_X1   g09731(.A1(new_n10652_), .A2(new_n10737_), .ZN(new_n10738_));
  NAND4_X1   g09732(.A1(new_n10622_), .A2(new_n10651_), .A3(new_n10736_), .A4(new_n10706_), .ZN(new_n10739_));
  NAND2_X1   g09733(.A1(new_n10738_), .A2(new_n10739_), .ZN(new_n10740_));
  INV_X1     g09734(.I(\A[97] ), .ZN(new_n10741_));
  INV_X1     g09735(.I(\A[98] ), .ZN(new_n10742_));
  NAND2_X1   g09736(.A1(new_n10742_), .A2(\A[99] ), .ZN(new_n10743_));
  INV_X1     g09737(.I(\A[99] ), .ZN(new_n10744_));
  NAND2_X1   g09738(.A1(new_n10744_), .A2(\A[98] ), .ZN(new_n10745_));
  AOI21_X1   g09739(.A1(new_n10743_), .A2(new_n10745_), .B(new_n10741_), .ZN(new_n10746_));
  NAND2_X1   g09740(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n10747_));
  NOR2_X1    g09741(.A1(\A[98] ), .A2(\A[99] ), .ZN(new_n10748_));
  INV_X1     g09742(.I(new_n10748_), .ZN(new_n10749_));
  AOI21_X1   g09743(.A1(new_n10749_), .A2(new_n10747_), .B(\A[97] ), .ZN(new_n10750_));
  NOR2_X1    g09744(.A1(new_n10750_), .A2(new_n10746_), .ZN(new_n10751_));
  INV_X1     g09745(.I(\A[100] ), .ZN(new_n10752_));
  INV_X1     g09746(.I(\A[101] ), .ZN(new_n10753_));
  NAND2_X1   g09747(.A1(new_n10753_), .A2(\A[102] ), .ZN(new_n10754_));
  INV_X1     g09748(.I(\A[102] ), .ZN(new_n10755_));
  NAND2_X1   g09749(.A1(new_n10755_), .A2(\A[101] ), .ZN(new_n10756_));
  AOI21_X1   g09750(.A1(new_n10754_), .A2(new_n10756_), .B(new_n10752_), .ZN(new_n10757_));
  NAND2_X1   g09751(.A1(\A[101] ), .A2(\A[102] ), .ZN(new_n10758_));
  NOR2_X1    g09752(.A1(\A[101] ), .A2(\A[102] ), .ZN(new_n10759_));
  INV_X1     g09753(.I(new_n10759_), .ZN(new_n10760_));
  AOI21_X1   g09754(.A1(new_n10760_), .A2(new_n10758_), .B(\A[100] ), .ZN(new_n10761_));
  NOR2_X1    g09755(.A1(new_n10761_), .A2(new_n10757_), .ZN(new_n10762_));
  AOI21_X1   g09756(.A1(\A[98] ), .A2(\A[99] ), .B(\A[97] ), .ZN(new_n10763_));
  AOI21_X1   g09757(.A1(\A[101] ), .A2(\A[102] ), .B(\A[100] ), .ZN(new_n10764_));
  OAI22_X1   g09758(.A1(new_n10748_), .A2(new_n10763_), .B1(new_n10764_), .B2(new_n10759_), .ZN(new_n10765_));
  NOR3_X1    g09759(.A1(new_n10751_), .A2(new_n10762_), .A3(new_n10765_), .ZN(new_n10766_));
  INV_X1     g09760(.I(\A[93] ), .ZN(new_n10767_));
  NOR2_X1    g09761(.A1(new_n10767_), .A2(\A[92] ), .ZN(new_n10768_));
  INV_X1     g09762(.I(\A[92] ), .ZN(new_n10769_));
  NOR2_X1    g09763(.A1(new_n10769_), .A2(\A[93] ), .ZN(new_n10770_));
  OAI21_X1   g09764(.A1(new_n10768_), .A2(new_n10770_), .B(\A[91] ), .ZN(new_n10771_));
  INV_X1     g09765(.I(\A[91] ), .ZN(new_n10772_));
  NAND2_X1   g09766(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n10773_));
  INV_X1     g09767(.I(new_n10773_), .ZN(new_n10774_));
  NOR2_X1    g09768(.A1(\A[92] ), .A2(\A[93] ), .ZN(new_n10775_));
  OAI21_X1   g09769(.A1(new_n10774_), .A2(new_n10775_), .B(new_n10772_), .ZN(new_n10776_));
  NAND2_X1   g09770(.A1(new_n10771_), .A2(new_n10776_), .ZN(new_n10777_));
  INV_X1     g09771(.I(\A[96] ), .ZN(new_n10778_));
  NOR2_X1    g09772(.A1(new_n10778_), .A2(\A[95] ), .ZN(new_n10779_));
  INV_X1     g09773(.I(\A[95] ), .ZN(new_n10780_));
  NOR2_X1    g09774(.A1(new_n10780_), .A2(\A[96] ), .ZN(new_n10781_));
  OAI21_X1   g09775(.A1(new_n10779_), .A2(new_n10781_), .B(\A[94] ), .ZN(new_n10782_));
  INV_X1     g09776(.I(\A[94] ), .ZN(new_n10783_));
  AND2_X2    g09777(.A1(\A[95] ), .A2(\A[96] ), .Z(new_n10784_));
  NOR2_X1    g09778(.A1(\A[95] ), .A2(\A[96] ), .ZN(new_n10785_));
  OAI21_X1   g09779(.A1(new_n10784_), .A2(new_n10785_), .B(new_n10783_), .ZN(new_n10786_));
  NAND2_X1   g09780(.A1(new_n10782_), .A2(new_n10786_), .ZN(new_n10787_));
  AOI21_X1   g09781(.A1(\A[92] ), .A2(\A[93] ), .B(\A[91] ), .ZN(new_n10788_));
  NOR2_X1    g09782(.A1(new_n10788_), .A2(new_n10775_), .ZN(new_n10789_));
  AOI21_X1   g09783(.A1(\A[95] ), .A2(\A[96] ), .B(\A[94] ), .ZN(new_n10790_));
  NOR2_X1    g09784(.A1(new_n10790_), .A2(new_n10785_), .ZN(new_n10791_));
  NOR2_X1    g09785(.A1(new_n10789_), .A2(new_n10791_), .ZN(new_n10792_));
  NAND3_X1   g09786(.A1(new_n10777_), .A2(new_n10787_), .A3(new_n10792_), .ZN(new_n10793_));
  NOR2_X1    g09787(.A1(new_n10766_), .A2(new_n10793_), .ZN(new_n10794_));
  NOR2_X1    g09788(.A1(new_n10744_), .A2(\A[98] ), .ZN(new_n10795_));
  NOR2_X1    g09789(.A1(new_n10742_), .A2(\A[99] ), .ZN(new_n10796_));
  OAI21_X1   g09790(.A1(new_n10795_), .A2(new_n10796_), .B(\A[97] ), .ZN(new_n10797_));
  INV_X1     g09791(.I(new_n10747_), .ZN(new_n10798_));
  OAI21_X1   g09792(.A1(new_n10798_), .A2(new_n10748_), .B(new_n10741_), .ZN(new_n10799_));
  NAND2_X1   g09793(.A1(new_n10797_), .A2(new_n10799_), .ZN(new_n10800_));
  NOR2_X1    g09794(.A1(new_n10755_), .A2(\A[101] ), .ZN(new_n10801_));
  NOR2_X1    g09795(.A1(new_n10753_), .A2(\A[102] ), .ZN(new_n10802_));
  OAI21_X1   g09796(.A1(new_n10801_), .A2(new_n10802_), .B(\A[100] ), .ZN(new_n10803_));
  INV_X1     g09797(.I(new_n10758_), .ZN(new_n10804_));
  OAI21_X1   g09798(.A1(new_n10804_), .A2(new_n10759_), .B(new_n10752_), .ZN(new_n10805_));
  NAND2_X1   g09799(.A1(new_n10803_), .A2(new_n10805_), .ZN(new_n10806_));
  NOR2_X1    g09800(.A1(new_n10763_), .A2(new_n10748_), .ZN(new_n10807_));
  NOR2_X1    g09801(.A1(new_n10764_), .A2(new_n10759_), .ZN(new_n10808_));
  NOR2_X1    g09802(.A1(new_n10807_), .A2(new_n10808_), .ZN(new_n10809_));
  NAND3_X1   g09803(.A1(new_n10800_), .A2(new_n10806_), .A3(new_n10809_), .ZN(new_n10810_));
  NAND2_X1   g09804(.A1(new_n10769_), .A2(\A[93] ), .ZN(new_n10811_));
  NAND2_X1   g09805(.A1(new_n10767_), .A2(\A[92] ), .ZN(new_n10812_));
  AOI21_X1   g09806(.A1(new_n10811_), .A2(new_n10812_), .B(new_n10772_), .ZN(new_n10813_));
  INV_X1     g09807(.I(new_n10775_), .ZN(new_n10814_));
  AOI21_X1   g09808(.A1(new_n10814_), .A2(new_n10773_), .B(\A[91] ), .ZN(new_n10815_));
  NOR2_X1    g09809(.A1(new_n10815_), .A2(new_n10813_), .ZN(new_n10816_));
  NAND2_X1   g09810(.A1(new_n10780_), .A2(\A[96] ), .ZN(new_n10817_));
  NAND2_X1   g09811(.A1(new_n10778_), .A2(\A[95] ), .ZN(new_n10818_));
  AOI21_X1   g09812(.A1(new_n10817_), .A2(new_n10818_), .B(new_n10783_), .ZN(new_n10819_));
  NAND2_X1   g09813(.A1(\A[95] ), .A2(\A[96] ), .ZN(new_n10820_));
  INV_X1     g09814(.I(new_n10785_), .ZN(new_n10821_));
  AOI21_X1   g09815(.A1(new_n10821_), .A2(new_n10820_), .B(\A[94] ), .ZN(new_n10822_));
  NOR2_X1    g09816(.A1(new_n10822_), .A2(new_n10819_), .ZN(new_n10823_));
  OAI22_X1   g09817(.A1(new_n10775_), .A2(new_n10788_), .B1(new_n10790_), .B2(new_n10785_), .ZN(new_n10824_));
  NOR3_X1    g09818(.A1(new_n10816_), .A2(new_n10823_), .A3(new_n10824_), .ZN(new_n10825_));
  NOR2_X1    g09819(.A1(new_n10825_), .A2(new_n10810_), .ZN(new_n10826_));
  INV_X1     g09820(.I(\A[85] ), .ZN(new_n10827_));
  INV_X1     g09821(.I(\A[86] ), .ZN(new_n10828_));
  NAND2_X1   g09822(.A1(new_n10828_), .A2(\A[87] ), .ZN(new_n10829_));
  INV_X1     g09823(.I(\A[87] ), .ZN(new_n10830_));
  NAND2_X1   g09824(.A1(new_n10830_), .A2(\A[86] ), .ZN(new_n10831_));
  AOI21_X1   g09825(.A1(new_n10829_), .A2(new_n10831_), .B(new_n10827_), .ZN(new_n10832_));
  NAND2_X1   g09826(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n10833_));
  NOR2_X1    g09827(.A1(\A[86] ), .A2(\A[87] ), .ZN(new_n10834_));
  INV_X1     g09828(.I(new_n10834_), .ZN(new_n10835_));
  AOI21_X1   g09829(.A1(new_n10835_), .A2(new_n10833_), .B(\A[85] ), .ZN(new_n10836_));
  NOR2_X1    g09830(.A1(new_n10836_), .A2(new_n10832_), .ZN(new_n10837_));
  INV_X1     g09831(.I(\A[88] ), .ZN(new_n10838_));
  INV_X1     g09832(.I(\A[89] ), .ZN(new_n10839_));
  NAND2_X1   g09833(.A1(new_n10839_), .A2(\A[90] ), .ZN(new_n10840_));
  INV_X1     g09834(.I(\A[90] ), .ZN(new_n10841_));
  NAND2_X1   g09835(.A1(new_n10841_), .A2(\A[89] ), .ZN(new_n10842_));
  AOI21_X1   g09836(.A1(new_n10840_), .A2(new_n10842_), .B(new_n10838_), .ZN(new_n10843_));
  NAND2_X1   g09837(.A1(\A[89] ), .A2(\A[90] ), .ZN(new_n10844_));
  NOR2_X1    g09838(.A1(\A[89] ), .A2(\A[90] ), .ZN(new_n10845_));
  INV_X1     g09839(.I(new_n10845_), .ZN(new_n10846_));
  AOI21_X1   g09840(.A1(new_n10846_), .A2(new_n10844_), .B(\A[88] ), .ZN(new_n10847_));
  NOR2_X1    g09841(.A1(new_n10847_), .A2(new_n10843_), .ZN(new_n10848_));
  AOI21_X1   g09842(.A1(\A[86] ), .A2(\A[87] ), .B(\A[85] ), .ZN(new_n10849_));
  AOI21_X1   g09843(.A1(\A[89] ), .A2(\A[90] ), .B(\A[88] ), .ZN(new_n10850_));
  OAI22_X1   g09844(.A1(new_n10834_), .A2(new_n10849_), .B1(new_n10850_), .B2(new_n10845_), .ZN(new_n10851_));
  NOR3_X1    g09845(.A1(new_n10837_), .A2(new_n10848_), .A3(new_n10851_), .ZN(new_n10852_));
  INV_X1     g09846(.I(\A[81] ), .ZN(new_n10853_));
  NOR2_X1    g09847(.A1(new_n10853_), .A2(\A[80] ), .ZN(new_n10854_));
  INV_X1     g09848(.I(\A[80] ), .ZN(new_n10855_));
  NOR2_X1    g09849(.A1(new_n10855_), .A2(\A[81] ), .ZN(new_n10856_));
  OAI21_X1   g09850(.A1(new_n10854_), .A2(new_n10856_), .B(\A[79] ), .ZN(new_n10857_));
  INV_X1     g09851(.I(\A[79] ), .ZN(new_n10858_));
  NAND2_X1   g09852(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n10859_));
  INV_X1     g09853(.I(new_n10859_), .ZN(new_n10860_));
  NOR2_X1    g09854(.A1(\A[80] ), .A2(\A[81] ), .ZN(new_n10861_));
  OAI21_X1   g09855(.A1(new_n10860_), .A2(new_n10861_), .B(new_n10858_), .ZN(new_n10862_));
  NAND2_X1   g09856(.A1(new_n10857_), .A2(new_n10862_), .ZN(new_n10863_));
  INV_X1     g09857(.I(\A[84] ), .ZN(new_n10864_));
  NOR2_X1    g09858(.A1(new_n10864_), .A2(\A[83] ), .ZN(new_n10865_));
  INV_X1     g09859(.I(\A[83] ), .ZN(new_n10866_));
  NOR2_X1    g09860(.A1(new_n10866_), .A2(\A[84] ), .ZN(new_n10867_));
  OAI21_X1   g09861(.A1(new_n10865_), .A2(new_n10867_), .B(\A[82] ), .ZN(new_n10868_));
  INV_X1     g09862(.I(\A[82] ), .ZN(new_n10869_));
  AND2_X2    g09863(.A1(\A[83] ), .A2(\A[84] ), .Z(new_n10870_));
  NOR2_X1    g09864(.A1(\A[83] ), .A2(\A[84] ), .ZN(new_n10871_));
  OAI21_X1   g09865(.A1(new_n10870_), .A2(new_n10871_), .B(new_n10869_), .ZN(new_n10872_));
  NAND2_X1   g09866(.A1(new_n10868_), .A2(new_n10872_), .ZN(new_n10873_));
  AOI21_X1   g09867(.A1(\A[80] ), .A2(\A[81] ), .B(\A[79] ), .ZN(new_n10874_));
  AOI21_X1   g09868(.A1(\A[83] ), .A2(\A[84] ), .B(\A[82] ), .ZN(new_n10875_));
  OAI22_X1   g09869(.A1(new_n10861_), .A2(new_n10874_), .B1(new_n10875_), .B2(new_n10871_), .ZN(new_n10876_));
  INV_X1     g09870(.I(new_n10876_), .ZN(new_n10877_));
  NAND3_X1   g09871(.A1(new_n10863_), .A2(new_n10873_), .A3(new_n10877_), .ZN(new_n10878_));
  NOR2_X1    g09872(.A1(new_n10852_), .A2(new_n10878_), .ZN(new_n10879_));
  NOR2_X1    g09873(.A1(new_n10830_), .A2(\A[86] ), .ZN(new_n10880_));
  NOR2_X1    g09874(.A1(new_n10828_), .A2(\A[87] ), .ZN(new_n10881_));
  OAI21_X1   g09875(.A1(new_n10880_), .A2(new_n10881_), .B(\A[85] ), .ZN(new_n10882_));
  AND2_X2    g09876(.A1(\A[86] ), .A2(\A[87] ), .Z(new_n10883_));
  OAI21_X1   g09877(.A1(new_n10883_), .A2(new_n10834_), .B(new_n10827_), .ZN(new_n10884_));
  NAND2_X1   g09878(.A1(new_n10882_), .A2(new_n10884_), .ZN(new_n10885_));
  NOR2_X1    g09879(.A1(new_n10841_), .A2(\A[89] ), .ZN(new_n10886_));
  NOR2_X1    g09880(.A1(new_n10839_), .A2(\A[90] ), .ZN(new_n10887_));
  OAI21_X1   g09881(.A1(new_n10886_), .A2(new_n10887_), .B(\A[88] ), .ZN(new_n10888_));
  AND2_X2    g09882(.A1(\A[89] ), .A2(\A[90] ), .Z(new_n10889_));
  OAI21_X1   g09883(.A1(new_n10889_), .A2(new_n10845_), .B(new_n10838_), .ZN(new_n10890_));
  NAND2_X1   g09884(.A1(new_n10888_), .A2(new_n10890_), .ZN(new_n10891_));
  NOR2_X1    g09885(.A1(new_n10849_), .A2(new_n10834_), .ZN(new_n10892_));
  NOR2_X1    g09886(.A1(new_n10850_), .A2(new_n10845_), .ZN(new_n10893_));
  NOR2_X1    g09887(.A1(new_n10892_), .A2(new_n10893_), .ZN(new_n10894_));
  NAND3_X1   g09888(.A1(new_n10885_), .A2(new_n10891_), .A3(new_n10894_), .ZN(new_n10895_));
  NAND2_X1   g09889(.A1(new_n10855_), .A2(\A[81] ), .ZN(new_n10896_));
  NAND2_X1   g09890(.A1(new_n10853_), .A2(\A[80] ), .ZN(new_n10897_));
  AOI21_X1   g09891(.A1(new_n10896_), .A2(new_n10897_), .B(new_n10858_), .ZN(new_n10898_));
  INV_X1     g09892(.I(new_n10861_), .ZN(new_n10899_));
  AOI21_X1   g09893(.A1(new_n10899_), .A2(new_n10859_), .B(\A[79] ), .ZN(new_n10900_));
  NOR2_X1    g09894(.A1(new_n10900_), .A2(new_n10898_), .ZN(new_n10901_));
  NAND2_X1   g09895(.A1(new_n10866_), .A2(\A[84] ), .ZN(new_n10902_));
  NAND2_X1   g09896(.A1(new_n10864_), .A2(\A[83] ), .ZN(new_n10903_));
  AOI21_X1   g09897(.A1(new_n10902_), .A2(new_n10903_), .B(new_n10869_), .ZN(new_n10904_));
  NAND2_X1   g09898(.A1(\A[83] ), .A2(\A[84] ), .ZN(new_n10905_));
  OR2_X2     g09899(.A1(\A[83] ), .A2(\A[84] ), .Z(new_n10906_));
  AOI21_X1   g09900(.A1(new_n10906_), .A2(new_n10905_), .B(\A[82] ), .ZN(new_n10907_));
  NOR2_X1    g09901(.A1(new_n10904_), .A2(new_n10907_), .ZN(new_n10908_));
  NOR3_X1    g09902(.A1(new_n10901_), .A2(new_n10908_), .A3(new_n10876_), .ZN(new_n10909_));
  NOR2_X1    g09903(.A1(new_n10909_), .A2(new_n10895_), .ZN(new_n10910_));
  OAI22_X1   g09904(.A1(new_n10794_), .A2(new_n10826_), .B1(new_n10879_), .B2(new_n10910_), .ZN(new_n10911_));
  NAND2_X1   g09905(.A1(new_n10825_), .A2(new_n10810_), .ZN(new_n10912_));
  NAND2_X1   g09906(.A1(new_n10766_), .A2(new_n10793_), .ZN(new_n10913_));
  NAND2_X1   g09907(.A1(new_n10909_), .A2(new_n10895_), .ZN(new_n10914_));
  NAND2_X1   g09908(.A1(new_n10852_), .A2(new_n10878_), .ZN(new_n10915_));
  NAND4_X1   g09909(.A1(new_n10912_), .A2(new_n10913_), .A3(new_n10915_), .A4(new_n10914_), .ZN(new_n10916_));
  NAND2_X1   g09910(.A1(new_n10911_), .A2(new_n10916_), .ZN(new_n10917_));
  NAND2_X1   g09911(.A1(new_n10740_), .A2(new_n10917_), .ZN(new_n10918_));
  NOR2_X1    g09912(.A1(new_n10740_), .A2(new_n10917_), .ZN(new_n10919_));
  INV_X1     g09913(.I(new_n10919_), .ZN(new_n10920_));
  NAND2_X1   g09914(.A1(new_n10920_), .A2(new_n10918_), .ZN(new_n10921_));
  XOR2_X1    g09915(.A1(new_n10567_), .A2(new_n10921_), .Z(new_n10922_));
  NAND3_X1   g09916(.A1(new_n10226_), .A2(new_n10227_), .A3(new_n10922_), .ZN(new_n10923_));
  INV_X1     g09917(.I(new_n10923_), .ZN(new_n10924_));
  AOI21_X1   g09918(.A1(new_n10226_), .A2(new_n10227_), .B(new_n10922_), .ZN(new_n10925_));
  NOR4_X1    g09919(.A1(new_n9551_), .A2(new_n9549_), .A3(new_n10924_), .A4(new_n10925_), .ZN(new_n10926_));
  INV_X1     g09920(.I(new_n10926_), .ZN(new_n10927_));
  OAI22_X1   g09921(.A1(new_n9551_), .A2(new_n9549_), .B1(new_n10924_), .B2(new_n10925_), .ZN(new_n10928_));
  NOR2_X1    g09922(.A1(new_n8150_), .A2(new_n8151_), .ZN(new_n10929_));
  XOR2_X1    g09923(.A1(new_n10929_), .A2(new_n8135_), .Z(new_n10930_));
  XOR2_X1    g09924(.A1(new_n10930_), .A2(new_n7083_), .Z(new_n10931_));
  NAND3_X1   g09925(.A1(new_n10931_), .A2(new_n10927_), .A3(new_n10928_), .ZN(new_n10932_));
  NOR2_X1    g09926(.A1(new_n10932_), .A2(new_n8199_), .ZN(new_n10933_));
  NAND2_X1   g09927(.A1(new_n8701_), .A2(new_n8617_), .ZN(new_n10934_));
  INV_X1     g09928(.I(new_n8617_), .ZN(new_n10935_));
  NAND2_X1   g09929(.A1(new_n10935_), .A2(new_n8603_), .ZN(new_n10936_));
  AOI21_X1   g09930(.A1(new_n10936_), .A2(new_n10934_), .B(new_n8614_), .ZN(new_n10937_));
  AND2_X2    g09931(.A1(new_n8608_), .A2(new_n8613_), .Z(new_n10938_));
  NOR2_X1    g09932(.A1(new_n10935_), .A2(new_n8603_), .ZN(new_n10939_));
  NOR2_X1    g09933(.A1(new_n8701_), .A2(new_n8617_), .ZN(new_n10940_));
  NOR3_X1    g09934(.A1(new_n10939_), .A2(new_n10940_), .A3(new_n10938_), .ZN(new_n10941_));
  OR2_X2     g09935(.A1(new_n10941_), .A2(new_n10937_), .Z(new_n10942_));
  NOR2_X1    g09936(.A1(new_n10938_), .A2(new_n8640_), .ZN(new_n10943_));
  NAND2_X1   g09937(.A1(new_n8632_), .A2(\A[462] ), .ZN(new_n10944_));
  NAND2_X1   g09938(.A1(new_n8630_), .A2(\A[461] ), .ZN(new_n10945_));
  AOI21_X1   g09939(.A1(new_n10944_), .A2(new_n10945_), .B(new_n8635_), .ZN(new_n10946_));
  INV_X1     g09940(.I(new_n8638_), .ZN(new_n10947_));
  AOI21_X1   g09941(.A1(new_n10947_), .A2(new_n8636_), .B(\A[460] ), .ZN(new_n10948_));
  NOR2_X1    g09942(.A1(new_n10948_), .A2(new_n10946_), .ZN(new_n10949_));
  NOR2_X1    g09943(.A1(new_n10949_), .A2(new_n8614_), .ZN(new_n10950_));
  NOR2_X1    g09944(.A1(new_n8629_), .A2(new_n8603_), .ZN(new_n10951_));
  NOR2_X1    g09945(.A1(new_n8701_), .A2(new_n8682_), .ZN(new_n10952_));
  OAI22_X1   g09946(.A1(new_n10943_), .A2(new_n10950_), .B1(new_n10951_), .B2(new_n10952_), .ZN(new_n10953_));
  NAND3_X1   g09947(.A1(new_n8603_), .A2(new_n8614_), .A3(new_n8617_), .ZN(new_n10954_));
  NAND3_X1   g09948(.A1(new_n8682_), .A2(new_n8640_), .A3(new_n8645_), .ZN(new_n10955_));
  NAND2_X1   g09949(.A1(new_n10955_), .A2(new_n10954_), .ZN(new_n10956_));
  NOR2_X1    g09950(.A1(new_n10953_), .A2(new_n10956_), .ZN(new_n10957_));
  NAND3_X1   g09951(.A1(new_n8645_), .A2(new_n8679_), .A3(new_n8681_), .ZN(new_n10958_));
  OAI22_X1   g09952(.A1(new_n8625_), .A2(new_n8641_), .B1(new_n8643_), .B2(new_n8638_), .ZN(new_n10959_));
  OAI21_X1   g09953(.A1(new_n8624_), .A2(new_n8628_), .B(new_n10959_), .ZN(new_n10960_));
  AOI21_X1   g09954(.A1(new_n10958_), .A2(new_n10960_), .B(new_n8640_), .ZN(new_n10961_));
  NOR3_X1    g09955(.A1(new_n8628_), .A2(new_n10959_), .A3(new_n8624_), .ZN(new_n10962_));
  AOI21_X1   g09956(.A1(new_n8679_), .A2(new_n8681_), .B(new_n8645_), .ZN(new_n10963_));
  NOR3_X1    g09957(.A1(new_n10963_), .A2(new_n10949_), .A3(new_n10962_), .ZN(new_n10964_));
  NOR2_X1    g09958(.A1(new_n10964_), .A2(new_n10961_), .ZN(new_n10965_));
  XOR2_X1    g09959(.A1(new_n10957_), .A2(new_n10965_), .Z(new_n10966_));
  NOR2_X1    g09960(.A1(new_n10966_), .A2(new_n10942_), .ZN(new_n10967_));
  INV_X1     g09961(.I(new_n10967_), .ZN(new_n10968_));
  OAI21_X1   g09962(.A1(new_n10963_), .A2(new_n10962_), .B(new_n10949_), .ZN(new_n10969_));
  NAND3_X1   g09963(.A1(new_n10958_), .A2(new_n10960_), .A3(new_n8640_), .ZN(new_n10970_));
  NAND2_X1   g09964(.A1(new_n10969_), .A2(new_n10970_), .ZN(new_n10971_));
  NOR2_X1    g09965(.A1(new_n10941_), .A2(new_n10937_), .ZN(new_n10972_));
  NAND2_X1   g09966(.A1(new_n10949_), .A2(new_n8614_), .ZN(new_n10973_));
  NAND2_X1   g09967(.A1(new_n10938_), .A2(new_n8640_), .ZN(new_n10974_));
  NAND2_X1   g09968(.A1(new_n8701_), .A2(new_n8682_), .ZN(new_n10975_));
  NAND2_X1   g09969(.A1(new_n8629_), .A2(new_n8603_), .ZN(new_n10976_));
  AOI22_X1   g09970(.A1(new_n10974_), .A2(new_n10973_), .B1(new_n10975_), .B2(new_n10976_), .ZN(new_n10977_));
  NAND2_X1   g09971(.A1(new_n8642_), .A2(new_n8644_), .ZN(new_n10978_));
  NAND3_X1   g09972(.A1(new_n8682_), .A2(new_n8640_), .A3(new_n10978_), .ZN(new_n10979_));
  NOR2_X1    g09973(.A1(new_n10979_), .A2(new_n10954_), .ZN(new_n10980_));
  NAND3_X1   g09974(.A1(new_n10977_), .A2(new_n10971_), .A3(new_n10980_), .ZN(new_n10981_));
  NOR2_X1    g09975(.A1(new_n10981_), .A2(new_n10972_), .ZN(new_n10982_));
  OAI21_X1   g09976(.A1(new_n10982_), .A2(new_n10971_), .B(new_n10957_), .ZN(new_n10983_));
  XOR2_X1    g09977(.A1(new_n8592_), .A2(new_n8618_), .Z(new_n10984_));
  NAND3_X1   g09978(.A1(new_n8672_), .A2(new_n8651_), .A3(new_n8656_), .ZN(new_n10985_));
  OAI22_X1   g09979(.A1(new_n8653_), .A2(new_n8668_), .B1(new_n8670_), .B2(new_n8665_), .ZN(new_n10986_));
  OAI21_X1   g09980(.A1(new_n8686_), .A2(new_n8688_), .B(new_n10986_), .ZN(new_n10987_));
  AOI21_X1   g09981(.A1(new_n10985_), .A2(new_n10987_), .B(new_n8667_), .ZN(new_n10988_));
  AND2_X2    g09982(.A1(new_n8666_), .A2(new_n8662_), .Z(new_n10989_));
  NOR3_X1    g09983(.A1(new_n8688_), .A2(new_n10986_), .A3(new_n8686_), .ZN(new_n10990_));
  AOI21_X1   g09984(.A1(new_n8651_), .A2(new_n8656_), .B(new_n8672_), .ZN(new_n10991_));
  NOR3_X1    g09985(.A1(new_n10991_), .A2(new_n10989_), .A3(new_n10990_), .ZN(new_n10992_));
  NOR2_X1    g09986(.A1(new_n10992_), .A2(new_n10988_), .ZN(new_n10993_));
  NAND2_X1   g09987(.A1(new_n10989_), .A2(new_n8588_), .ZN(new_n10994_));
  INV_X1     g09988(.I(new_n8588_), .ZN(new_n10995_));
  NAND2_X1   g09989(.A1(new_n10995_), .A2(new_n8667_), .ZN(new_n10996_));
  NAND2_X1   g09990(.A1(new_n8577_), .A2(new_n8657_), .ZN(new_n10997_));
  NOR2_X1    g09991(.A1(new_n8570_), .A2(\A[440] ), .ZN(new_n10998_));
  NOR2_X1    g09992(.A1(new_n8568_), .A2(\A[441] ), .ZN(new_n10999_));
  OAI21_X1   g09993(.A1(new_n10998_), .A2(new_n10999_), .B(\A[439] ), .ZN(new_n11000_));
  INV_X1     g09994(.I(new_n8575_), .ZN(new_n11001_));
  OAI21_X1   g09995(.A1(new_n11001_), .A2(new_n8573_), .B(new_n8567_), .ZN(new_n11002_));
  NAND2_X1   g09996(.A1(new_n11000_), .A2(new_n11002_), .ZN(new_n11003_));
  NAND2_X1   g09997(.A1(new_n8689_), .A2(new_n11003_), .ZN(new_n11004_));
  AOI22_X1   g09998(.A1(new_n10996_), .A2(new_n10994_), .B1(new_n10997_), .B2(new_n11004_), .ZN(new_n11005_));
  NOR4_X1    g09999(.A1(new_n8589_), .A2(\A[442] ), .A3(\A[443] ), .A4(\A[444] ), .ZN(new_n11006_));
  AOI21_X1   g10000(.A1(new_n8662_), .A2(new_n8666_), .B(new_n10986_), .ZN(new_n11007_));
  AOI22_X1   g10001(.A1(new_n11007_), .A2(new_n8657_), .B1(new_n11003_), .B2(new_n11006_), .ZN(new_n11008_));
  NAND2_X1   g10002(.A1(new_n11005_), .A2(new_n11008_), .ZN(new_n11009_));
  NAND2_X1   g10003(.A1(new_n8577_), .A2(new_n8591_), .ZN(new_n11010_));
  INV_X1     g10004(.I(new_n11010_), .ZN(new_n11011_));
  NOR2_X1    g10005(.A1(new_n8577_), .A2(new_n8591_), .ZN(new_n11012_));
  OAI21_X1   g10006(.A1(new_n11011_), .A2(new_n11012_), .B(new_n10995_), .ZN(new_n11013_));
  INV_X1     g10007(.I(new_n8591_), .ZN(new_n11014_));
  NAND2_X1   g10008(.A1(new_n11014_), .A2(new_n11003_), .ZN(new_n11015_));
  NAND3_X1   g10009(.A1(new_n11015_), .A2(new_n11010_), .A3(new_n8588_), .ZN(new_n11016_));
  NAND2_X1   g10010(.A1(new_n11013_), .A2(new_n11016_), .ZN(new_n11017_));
  NOR2_X1    g10011(.A1(new_n10995_), .A2(new_n8667_), .ZN(new_n11018_));
  NOR2_X1    g10012(.A1(new_n10989_), .A2(new_n8588_), .ZN(new_n11019_));
  NOR2_X1    g10013(.A1(new_n8689_), .A2(new_n11003_), .ZN(new_n11020_));
  NOR2_X1    g10014(.A1(new_n8577_), .A2(new_n8657_), .ZN(new_n11021_));
  OAI22_X1   g10015(.A1(new_n11018_), .A2(new_n11019_), .B1(new_n11020_), .B2(new_n11021_), .ZN(new_n11022_));
  NAND2_X1   g10016(.A1(new_n8669_), .A2(new_n8671_), .ZN(new_n11023_));
  NOR2_X1    g10017(.A1(new_n10989_), .A2(new_n8689_), .ZN(new_n11024_));
  NAND4_X1   g10018(.A1(new_n11024_), .A2(new_n11003_), .A3(new_n11006_), .A4(new_n11023_), .ZN(new_n11025_));
  NAND3_X1   g10019(.A1(new_n11009_), .A2(new_n11017_), .A3(new_n10993_), .ZN(new_n11027_));
  NOR3_X1    g10020(.A1(new_n8674_), .A2(new_n10984_), .A3(new_n11027_), .ZN(new_n11028_));
  NAND2_X1   g10021(.A1(new_n11028_), .A2(new_n10983_), .ZN(new_n11029_));
  OR2_X2     g10022(.A1(new_n11028_), .A2(new_n10983_), .Z(new_n11030_));
  AOI21_X1   g10023(.A1(new_n11030_), .A2(new_n11029_), .B(new_n10968_), .ZN(new_n11031_));
  INV_X1     g10024(.I(new_n11031_), .ZN(new_n11032_));
  NAND4_X1   g10025(.A1(new_n8694_), .A2(new_n8705_), .A3(new_n8875_), .A4(new_n8871_), .ZN(new_n11033_));
  NAND2_X1   g10026(.A1(new_n8857_), .A2(new_n8768_), .ZN(new_n11034_));
  OR2_X2     g10027(.A1(new_n8766_), .A2(new_n8767_), .Z(new_n11035_));
  NAND2_X1   g10028(.A1(new_n11035_), .A2(new_n8754_), .ZN(new_n11036_));
  AOI21_X1   g10029(.A1(new_n11036_), .A2(new_n11034_), .B(new_n8765_), .ZN(new_n11037_));
  NOR2_X1    g10030(.A1(new_n11035_), .A2(new_n8754_), .ZN(new_n11038_));
  NOR2_X1    g10031(.A1(new_n8857_), .A2(new_n8768_), .ZN(new_n11039_));
  NOR3_X1    g10032(.A1(new_n11038_), .A2(new_n11039_), .A3(new_n8863_), .ZN(new_n11040_));
  NOR2_X1    g10033(.A1(new_n11040_), .A2(new_n11037_), .ZN(new_n11041_));
  NAND2_X1   g10034(.A1(new_n8783_), .A2(\A[438] ), .ZN(new_n11042_));
  NAND2_X1   g10035(.A1(new_n8781_), .A2(\A[437] ), .ZN(new_n11043_));
  AOI21_X1   g10036(.A1(new_n11042_), .A2(new_n11043_), .B(new_n8786_), .ZN(new_n11044_));
  INV_X1     g10037(.I(new_n8789_), .ZN(new_n11045_));
  AOI21_X1   g10038(.A1(new_n11045_), .A2(new_n8787_), .B(\A[436] ), .ZN(new_n11046_));
  NOR2_X1    g10039(.A1(new_n11046_), .A2(new_n11044_), .ZN(new_n11047_));
  NAND3_X1   g10040(.A1(new_n8754_), .A2(new_n8765_), .A3(new_n8768_), .ZN(new_n11048_));
  NOR4_X1    g10041(.A1(new_n11048_), .A2(new_n8780_), .A3(new_n11047_), .A4(new_n8794_), .ZN(new_n11049_));
  NOR2_X1    g10042(.A1(new_n8843_), .A2(new_n8794_), .ZN(new_n11050_));
  NOR2_X1    g10043(.A1(new_n8780_), .A2(new_n8795_), .ZN(new_n11051_));
  OAI21_X1   g10044(.A1(new_n11051_), .A2(new_n11050_), .B(new_n11047_), .ZN(new_n11052_));
  NAND2_X1   g10045(.A1(new_n8780_), .A2(new_n8795_), .ZN(new_n11053_));
  NAND2_X1   g10046(.A1(new_n8843_), .A2(new_n8794_), .ZN(new_n11054_));
  NAND3_X1   g10047(.A1(new_n11053_), .A2(new_n11054_), .A3(new_n8791_), .ZN(new_n11055_));
  AOI21_X1   g10048(.A1(new_n11052_), .A2(new_n11055_), .B(new_n11049_), .ZN(new_n11056_));
  NOR3_X1    g10049(.A1(new_n11035_), .A2(new_n8857_), .A3(new_n8863_), .ZN(new_n11057_));
  NAND4_X1   g10050(.A1(new_n11057_), .A2(new_n8843_), .A3(new_n8791_), .A4(new_n8795_), .ZN(new_n11058_));
  AOI21_X1   g10051(.A1(new_n11053_), .A2(new_n11054_), .B(new_n8791_), .ZN(new_n11059_));
  NOR3_X1    g10052(.A1(new_n11051_), .A2(new_n11050_), .A3(new_n11047_), .ZN(new_n11060_));
  NOR3_X1    g10053(.A1(new_n11058_), .A2(new_n11059_), .A3(new_n11060_), .ZN(new_n11061_));
  OAI21_X1   g10054(.A1(new_n11056_), .A2(new_n11061_), .B(new_n11041_), .ZN(new_n11062_));
  NAND2_X1   g10055(.A1(new_n11052_), .A2(new_n11055_), .ZN(new_n11063_));
  NAND2_X1   g10056(.A1(new_n8864_), .A2(new_n8851_), .ZN(new_n11064_));
  OR4_X2     g10057(.A1(new_n8776_), .A2(new_n8792_), .A3(new_n8793_), .A4(new_n8789_), .Z(new_n11065_));
  NAND3_X1   g10058(.A1(new_n8843_), .A2(new_n8791_), .A3(new_n11065_), .ZN(new_n11066_));
  NOR2_X1    g10059(.A1(new_n11064_), .A2(new_n11066_), .ZN(new_n11067_));
  NOR2_X1    g10060(.A1(new_n8780_), .A2(new_n11047_), .ZN(new_n11068_));
  NOR2_X1    g10061(.A1(new_n8843_), .A2(new_n8791_), .ZN(new_n11069_));
  NOR3_X1    g10062(.A1(new_n11068_), .A2(new_n11069_), .A3(new_n8866_), .ZN(new_n11070_));
  NAND3_X1   g10063(.A1(new_n11063_), .A2(new_n11067_), .A3(new_n11070_), .ZN(new_n11071_));
  NOR4_X1    g10064(.A1(new_n11048_), .A2(new_n8780_), .A3(new_n11047_), .A4(new_n8794_), .ZN(new_n11073_));
  AOI22_X1   g10065(.A1(new_n8729_), .A2(new_n8731_), .B1(new_n8734_), .B2(new_n8736_), .ZN(new_n11074_));
  NOR4_X1    g10066(.A1(new_n8711_), .A2(new_n8715_), .A3(new_n8725_), .A4(new_n8721_), .ZN(new_n11075_));
  NOR2_X1    g10067(.A1(new_n11074_), .A2(new_n11075_), .ZN(new_n11076_));
  NAND4_X1   g10068(.A1(new_n8738_), .A2(new_n8830_), .A3(new_n8741_), .A4(new_n8833_), .ZN(new_n11077_));
  NOR3_X1    g10069(.A1(new_n11076_), .A2(new_n8847_), .A3(new_n11077_), .ZN(new_n11078_));
  NOR2_X1    g10070(.A1(new_n8816_), .A2(new_n8812_), .ZN(new_n11079_));
  AOI21_X1   g10071(.A1(\A[422] ), .A2(\A[423] ), .B(\A[421] ), .ZN(new_n11080_));
  OAI22_X1   g10072(.A1(new_n8804_), .A2(new_n11080_), .B1(new_n8831_), .B2(new_n8814_), .ZN(new_n11081_));
  NOR3_X1    g10073(.A1(new_n8806_), .A2(new_n11081_), .A3(new_n8802_), .ZN(new_n11082_));
  NOR2_X1    g10074(.A1(new_n11080_), .A2(new_n8804_), .ZN(new_n11083_));
  INV_X1     g10075(.I(new_n11083_), .ZN(new_n11084_));
  INV_X1     g10076(.I(new_n8832_), .ZN(new_n11085_));
  AOI22_X1   g10077(.A1(new_n11084_), .A2(new_n11085_), .B1(new_n8820_), .B2(new_n8822_), .ZN(new_n11086_));
  OAI21_X1   g10078(.A1(new_n11086_), .A2(new_n11082_), .B(new_n11079_), .ZN(new_n11087_));
  NOR2_X1    g10079(.A1(new_n11083_), .A2(new_n8832_), .ZN(new_n11088_));
  NAND3_X1   g10080(.A1(new_n11088_), .A2(new_n8820_), .A3(new_n8822_), .ZN(new_n11089_));
  OAI21_X1   g10081(.A1(new_n8802_), .A2(new_n8806_), .B(new_n11081_), .ZN(new_n11090_));
  NAND3_X1   g10082(.A1(new_n11089_), .A2(new_n11090_), .A3(new_n8830_), .ZN(new_n11091_));
  NAND2_X1   g10083(.A1(new_n11083_), .A2(new_n8832_), .ZN(new_n11092_));
  INV_X1     g10084(.I(new_n11092_), .ZN(new_n11093_));
  NAND3_X1   g10085(.A1(new_n8817_), .A2(new_n8828_), .A3(new_n11081_), .ZN(new_n11094_));
  NAND3_X1   g10086(.A1(new_n11094_), .A2(new_n11087_), .A3(new_n11091_), .ZN(new_n11095_));
  NOR2_X1    g10087(.A1(new_n8725_), .A2(new_n8721_), .ZN(new_n11096_));
  AOI21_X1   g10088(.A1(\A[416] ), .A2(\A[417] ), .B(\A[415] ), .ZN(new_n11097_));
  OAI22_X1   g10089(.A1(new_n8713_), .A2(new_n11097_), .B1(new_n8739_), .B2(new_n8723_), .ZN(new_n11098_));
  NOR3_X1    g10090(.A1(new_n8715_), .A2(new_n11098_), .A3(new_n8711_), .ZN(new_n11099_));
  NOR2_X1    g10091(.A1(new_n11097_), .A2(new_n8713_), .ZN(new_n11100_));
  NOR2_X1    g10092(.A1(new_n11100_), .A2(new_n8740_), .ZN(new_n11101_));
  AOI21_X1   g10093(.A1(new_n8729_), .A2(new_n8731_), .B(new_n11101_), .ZN(new_n11102_));
  OAI21_X1   g10094(.A1(new_n11102_), .A2(new_n11099_), .B(new_n11096_), .ZN(new_n11103_));
  NAND3_X1   g10095(.A1(new_n11101_), .A2(new_n8729_), .A3(new_n8731_), .ZN(new_n11104_));
  OAI21_X1   g10096(.A1(new_n8711_), .A2(new_n8715_), .B(new_n11098_), .ZN(new_n11105_));
  NAND3_X1   g10097(.A1(new_n11104_), .A2(new_n11105_), .A3(new_n8738_), .ZN(new_n11106_));
  NAND2_X1   g10098(.A1(new_n11103_), .A2(new_n11106_), .ZN(new_n11107_));
  NOR3_X1    g10099(.A1(new_n11078_), .A2(new_n11095_), .A3(new_n11107_), .ZN(new_n11108_));
  INV_X1     g10100(.I(new_n8741_), .ZN(new_n11109_));
  NOR2_X1    g10101(.A1(new_n11109_), .A2(new_n11096_), .ZN(new_n11110_));
  AOI22_X1   g10102(.A1(new_n8726_), .A2(new_n8737_), .B1(new_n8817_), .B2(new_n8828_), .ZN(new_n11111_));
  NAND3_X1   g10103(.A1(new_n11111_), .A2(new_n11110_), .A3(new_n8835_), .ZN(new_n11112_));
  AOI21_X1   g10104(.A1(new_n11089_), .A2(new_n11090_), .B(new_n8830_), .ZN(new_n11113_));
  NOR3_X1    g10105(.A1(new_n11086_), .A2(new_n11079_), .A3(new_n11082_), .ZN(new_n11114_));
  NOR3_X1    g10106(.A1(new_n8845_), .A2(new_n8846_), .A3(new_n11088_), .ZN(new_n11115_));
  NOR3_X1    g10107(.A1(new_n11115_), .A2(new_n11114_), .A3(new_n11113_), .ZN(new_n11116_));
  AOI21_X1   g10108(.A1(new_n11104_), .A2(new_n11105_), .B(new_n8738_), .ZN(new_n11117_));
  NOR3_X1    g10109(.A1(new_n11102_), .A2(new_n11096_), .A3(new_n11099_), .ZN(new_n11118_));
  NOR2_X1    g10110(.A1(new_n11118_), .A2(new_n11117_), .ZN(new_n11119_));
  AOI21_X1   g10111(.A1(new_n11112_), .A2(new_n11116_), .B(new_n11119_), .ZN(new_n11120_));
  NOR2_X1    g10112(.A1(new_n11120_), .A2(new_n11108_), .ZN(new_n11121_));
  NAND2_X1   g10113(.A1(new_n11087_), .A2(new_n11091_), .ZN(new_n11122_));
  AOI21_X1   g10114(.A1(new_n8845_), .A2(new_n11092_), .B(new_n11088_), .ZN(new_n11123_));
  NOR3_X1    g10115(.A1(new_n11076_), .A2(new_n11123_), .A3(new_n8847_), .ZN(new_n11124_));
  AOI21_X1   g10116(.A1(new_n11124_), .A2(new_n11122_), .B(new_n11110_), .ZN(new_n11125_));
  OAI21_X1   g10117(.A1(new_n8817_), .A2(new_n11093_), .B(new_n11081_), .ZN(new_n11126_));
  NAND2_X1   g10118(.A1(new_n11126_), .A2(new_n8829_), .ZN(new_n11127_));
  NOR2_X1    g10119(.A1(new_n11116_), .A2(new_n11078_), .ZN(new_n11128_));
  OAI21_X1   g10120(.A1(new_n11125_), .A2(new_n11127_), .B(new_n11128_), .ZN(new_n11129_));
  NOR2_X1    g10121(.A1(new_n8872_), .A2(new_n8867_), .ZN(new_n11130_));
  NOR2_X1    g10122(.A1(new_n8769_), .A2(new_n8743_), .ZN(new_n11131_));
  OAI22_X1   g10123(.A1(new_n8868_), .A2(new_n8869_), .B1(new_n11130_), .B2(new_n11131_), .ZN(new_n11132_));
  NOR4_X1    g10124(.A1(new_n11129_), .A2(new_n11121_), .A3(new_n11132_), .A4(new_n11073_), .ZN(new_n11133_));
  INV_X1     g10125(.I(new_n11073_), .ZN(new_n11134_));
  NAND3_X1   g10126(.A1(new_n11122_), .A2(new_n11111_), .A3(new_n11126_), .ZN(new_n11135_));
  AOI21_X1   g10127(.A1(new_n11135_), .A2(new_n8742_), .B(new_n11127_), .ZN(new_n11136_));
  NOR4_X1    g10128(.A1(new_n11136_), .A2(new_n11078_), .A3(new_n11116_), .A4(new_n11119_), .ZN(new_n11137_));
  NAND2_X1   g10129(.A1(new_n8769_), .A2(new_n8743_), .ZN(new_n11138_));
  NAND2_X1   g10130(.A1(new_n8872_), .A2(new_n8867_), .ZN(new_n11139_));
  AOI22_X1   g10131(.A1(new_n8837_), .A2(new_n8849_), .B1(new_n11139_), .B2(new_n11138_), .ZN(new_n11140_));
  AOI21_X1   g10132(.A1(new_n11137_), .A2(new_n11140_), .B(new_n11134_), .ZN(new_n11141_));
  OAI21_X1   g10133(.A1(new_n11141_), .A2(new_n11133_), .B(new_n11062_), .ZN(new_n11142_));
  OR2_X2     g10134(.A1(new_n11040_), .A2(new_n11037_), .Z(new_n11143_));
  NAND2_X1   g10135(.A1(new_n11063_), .A2(new_n11058_), .ZN(new_n11144_));
  NAND3_X1   g10136(.A1(new_n11049_), .A2(new_n11052_), .A3(new_n11055_), .ZN(new_n11145_));
  AOI21_X1   g10137(.A1(new_n11144_), .A2(new_n11145_), .B(new_n11143_), .ZN(new_n11146_));
  NAND3_X1   g10138(.A1(new_n11137_), .A2(new_n11134_), .A3(new_n11140_), .ZN(new_n11147_));
  NAND3_X1   g10139(.A1(new_n11112_), .A2(new_n11116_), .A3(new_n11119_), .ZN(new_n11148_));
  OAI21_X1   g10140(.A1(new_n11078_), .A2(new_n11095_), .B(new_n11107_), .ZN(new_n11149_));
  NAND2_X1   g10141(.A1(new_n11148_), .A2(new_n11149_), .ZN(new_n11150_));
  NOR2_X1    g10142(.A1(new_n11114_), .A2(new_n11113_), .ZN(new_n11151_));
  NAND2_X1   g10143(.A1(new_n8726_), .A2(new_n8737_), .ZN(new_n11152_));
  NAND3_X1   g10144(.A1(new_n11152_), .A2(new_n11126_), .A3(new_n8829_), .ZN(new_n11153_));
  OAI21_X1   g10145(.A1(new_n11153_), .A2(new_n11151_), .B(new_n8742_), .ZN(new_n11154_));
  INV_X1     g10146(.I(new_n11127_), .ZN(new_n11155_));
  NAND2_X1   g10147(.A1(new_n11154_), .A2(new_n11155_), .ZN(new_n11156_));
  NAND4_X1   g10148(.A1(new_n11150_), .A2(new_n11140_), .A3(new_n11156_), .A4(new_n11128_), .ZN(new_n11157_));
  NAND2_X1   g10149(.A1(new_n11157_), .A2(new_n11073_), .ZN(new_n11158_));
  NAND3_X1   g10150(.A1(new_n11158_), .A2(new_n11147_), .A3(new_n11146_), .ZN(new_n11159_));
  AOI21_X1   g10151(.A1(new_n11159_), .A2(new_n11142_), .B(new_n11033_), .ZN(new_n11160_));
  NOR2_X1    g10152(.A1(new_n11032_), .A2(new_n11160_), .ZN(new_n11161_));
  NOR3_X1    g10153(.A1(new_n8326_), .A2(new_n8354_), .A3(new_n8322_), .ZN(new_n11162_));
  AOI21_X1   g10154(.A1(new_n8340_), .A2(new_n8342_), .B(new_n8370_), .ZN(new_n11163_));
  OAI21_X1   g10155(.A1(new_n11163_), .A2(new_n11162_), .B(new_n8351_), .ZN(new_n11164_));
  NAND3_X1   g10156(.A1(new_n8370_), .A2(new_n8340_), .A3(new_n8342_), .ZN(new_n11165_));
  OAI21_X1   g10157(.A1(new_n8322_), .A2(new_n8326_), .B(new_n8354_), .ZN(new_n11166_));
  NAND3_X1   g10158(.A1(new_n11165_), .A2(new_n11166_), .A3(new_n8367_), .ZN(new_n11167_));
  NAND2_X1   g10159(.A1(new_n11164_), .A2(new_n11167_), .ZN(new_n11168_));
  NOR4_X1    g10160(.A1(new_n8361_), .A2(new_n8349_), .A3(new_n8359_), .A4(new_n8355_), .ZN(new_n11169_));
  NAND2_X1   g10161(.A1(new_n8311_), .A2(new_n8313_), .ZN(new_n11170_));
  NOR2_X1    g10162(.A1(new_n8298_), .A2(new_n8300_), .ZN(new_n11171_));
  NAND3_X1   g10163(.A1(new_n11171_), .A2(new_n8306_), .A3(new_n8308_), .ZN(new_n11172_));
  OAI22_X1   g10164(.A1(new_n8282_), .A2(new_n8299_), .B1(new_n8297_), .B2(new_n8292_), .ZN(new_n11173_));
  OAI21_X1   g10165(.A1(new_n8281_), .A2(new_n8285_), .B(new_n11173_), .ZN(new_n11174_));
  AOI21_X1   g10166(.A1(new_n11172_), .A2(new_n11174_), .B(new_n11170_), .ZN(new_n11175_));
  INV_X1     g10167(.I(new_n11170_), .ZN(new_n11176_));
  NOR3_X1    g10168(.A1(new_n8285_), .A2(new_n11173_), .A3(new_n8281_), .ZN(new_n11177_));
  AOI21_X1   g10169(.A1(new_n8306_), .A2(new_n8308_), .B(new_n11171_), .ZN(new_n11178_));
  NOR3_X1    g10170(.A1(new_n11178_), .A2(new_n11176_), .A3(new_n11177_), .ZN(new_n11179_));
  NOR2_X1    g10171(.A1(new_n11179_), .A2(new_n11175_), .ZN(new_n11180_));
  XOR2_X1    g10172(.A1(new_n11169_), .A2(new_n11180_), .Z(new_n11181_));
  NOR2_X1    g10173(.A1(new_n11181_), .A2(new_n11168_), .ZN(new_n11182_));
  OAI21_X1   g10174(.A1(new_n11178_), .A2(new_n11177_), .B(new_n11176_), .ZN(new_n11183_));
  NAND3_X1   g10175(.A1(new_n11172_), .A2(new_n11174_), .A3(new_n11170_), .ZN(new_n11184_));
  NAND2_X1   g10176(.A1(new_n11183_), .A2(new_n11184_), .ZN(new_n11185_));
  INV_X1     g10177(.I(new_n11168_), .ZN(new_n11186_));
  XNOR2_X1   g10178(.A1(new_n8298_), .A2(new_n8300_), .ZN(new_n11187_));
  NAND2_X1   g10179(.A1(new_n8301_), .A2(new_n11173_), .ZN(new_n11188_));
  NAND2_X1   g10180(.A1(new_n8358_), .A2(new_n11188_), .ZN(new_n11189_));
  OAI21_X1   g10181(.A1(new_n8358_), .A2(new_n11187_), .B(new_n11189_), .ZN(new_n11190_));
  NAND2_X1   g10182(.A1(new_n8314_), .A2(new_n8301_), .ZN(new_n11191_));
  NOR2_X1    g10183(.A1(new_n11191_), .A2(new_n8371_), .ZN(new_n11192_));
  NAND4_X1   g10184(.A1(new_n11190_), .A2(new_n8315_), .A3(new_n8365_), .A4(new_n11192_), .ZN(new_n11193_));
  NOR2_X1    g10185(.A1(new_n11193_), .A2(new_n11186_), .ZN(new_n11194_));
  OAI21_X1   g10186(.A1(new_n11194_), .A2(new_n11185_), .B(new_n11169_), .ZN(new_n11195_));
  NOR4_X1    g10187(.A1(new_n8265_), .A2(new_n8267_), .A3(new_n8272_), .A4(new_n8270_), .ZN(new_n11196_));
  INV_X1     g10188(.I(new_n8261_), .ZN(new_n11197_));
  NAND2_X1   g10189(.A1(new_n11196_), .A2(new_n11197_), .ZN(new_n11198_));
  AOI22_X1   g10190(.A1(new_n8240_), .A2(new_n8245_), .B1(new_n8250_), .B2(new_n8255_), .ZN(new_n11199_));
  NOR2_X1    g10191(.A1(new_n11199_), .A2(new_n11196_), .ZN(new_n11200_));
  NAND4_X1   g10192(.A1(new_n8224_), .A2(new_n8234_), .A3(new_n11200_), .A4(new_n11198_), .ZN(new_n11201_));
  NAND2_X1   g10193(.A1(new_n8250_), .A2(new_n8255_), .ZN(new_n11202_));
  OAI22_X1   g10194(.A1(new_n8242_), .A2(new_n8259_), .B1(new_n8257_), .B2(new_n8252_), .ZN(new_n11203_));
  INV_X1     g10195(.I(new_n11203_), .ZN(new_n11204_));
  NAND3_X1   g10196(.A1(new_n11204_), .A2(new_n8240_), .A3(new_n8245_), .ZN(new_n11205_));
  OAI21_X1   g10197(.A1(new_n8265_), .A2(new_n8267_), .B(new_n11203_), .ZN(new_n11206_));
  AOI21_X1   g10198(.A1(new_n11205_), .A2(new_n11206_), .B(new_n11202_), .ZN(new_n11207_));
  NOR2_X1    g10199(.A1(new_n8272_), .A2(new_n8270_), .ZN(new_n11208_));
  NOR3_X1    g10200(.A1(new_n8267_), .A2(new_n11203_), .A3(new_n8265_), .ZN(new_n11209_));
  NOR2_X1    g10201(.A1(new_n8267_), .A2(new_n8265_), .ZN(new_n11210_));
  NOR2_X1    g10202(.A1(new_n11210_), .A2(new_n11204_), .ZN(new_n11211_));
  NOR3_X1    g10203(.A1(new_n11211_), .A2(new_n11208_), .A3(new_n11209_), .ZN(new_n11212_));
  NOR2_X1    g10204(.A1(new_n11212_), .A2(new_n11207_), .ZN(new_n11213_));
  NOR3_X1    g10205(.A1(new_n8209_), .A2(new_n8388_), .A3(new_n8205_), .ZN(new_n11214_));
  OAI21_X1   g10206(.A1(\A[391] ), .A2(new_n8383_), .B(new_n8208_), .ZN(new_n11215_));
  INV_X1     g10207(.I(new_n8232_), .ZN(new_n11216_));
  AOI22_X1   g10208(.A1(new_n11215_), .A2(new_n11216_), .B1(new_n8382_), .B2(new_n8384_), .ZN(new_n11217_));
  OAI21_X1   g10209(.A1(new_n11217_), .A2(new_n11214_), .B(new_n8221_), .ZN(new_n11218_));
  NAND4_X1   g10210(.A1(new_n8382_), .A2(new_n11215_), .A3(new_n11216_), .A4(new_n8384_), .ZN(new_n11219_));
  OAI21_X1   g10211(.A1(new_n8205_), .A2(new_n8209_), .B(new_n8388_), .ZN(new_n11220_));
  NAND3_X1   g10212(.A1(new_n11219_), .A2(new_n11220_), .A3(new_n8230_), .ZN(new_n11221_));
  NAND2_X1   g10213(.A1(new_n11218_), .A2(new_n11221_), .ZN(new_n11222_));
  XNOR2_X1   g10214(.A1(new_n8258_), .A2(new_n8260_), .ZN(new_n11223_));
  NAND2_X1   g10215(.A1(new_n8261_), .A2(new_n11203_), .ZN(new_n11224_));
  NAND2_X1   g10216(.A1(new_n8256_), .A2(new_n11224_), .ZN(new_n11225_));
  OAI21_X1   g10217(.A1(new_n8256_), .A2(new_n11223_), .B(new_n11225_), .ZN(new_n11226_));
  NAND2_X1   g10218(.A1(new_n11199_), .A2(new_n8261_), .ZN(new_n11227_));
  NOR2_X1    g10219(.A1(new_n11227_), .A2(new_n8234_), .ZN(new_n11228_));
  NAND4_X1   g10220(.A1(new_n11226_), .A2(new_n8224_), .A3(new_n11228_), .A4(new_n11200_), .ZN(new_n11229_));
  NAND4_X1   g10221(.A1(new_n11229_), .A2(new_n11201_), .A3(new_n11213_), .A4(new_n11222_), .ZN(new_n11230_));
  NOR2_X1    g10222(.A1(new_n8372_), .A2(new_n8390_), .ZN(new_n11231_));
  NOR2_X1    g10223(.A1(new_n8235_), .A2(new_n8356_), .ZN(new_n11232_));
  NAND2_X1   g10224(.A1(new_n11200_), .A2(new_n11198_), .ZN(new_n11233_));
  NOR2_X1    g10225(.A1(new_n11233_), .A2(new_n8362_), .ZN(new_n11234_));
  NOR2_X1    g10226(.A1(new_n8316_), .A2(new_n8275_), .ZN(new_n11235_));
  OAI22_X1   g10227(.A1(new_n11232_), .A2(new_n11231_), .B1(new_n11234_), .B2(new_n11235_), .ZN(new_n11236_));
  NOR2_X1    g10228(.A1(new_n11236_), .A2(new_n11230_), .ZN(new_n11237_));
  NAND2_X1   g10229(.A1(new_n11237_), .A2(new_n11195_), .ZN(new_n11238_));
  INV_X1     g10230(.I(new_n11238_), .ZN(new_n11239_));
  NOR2_X1    g10231(.A1(new_n11237_), .A2(new_n11195_), .ZN(new_n11240_));
  OAI21_X1   g10232(.A1(new_n11239_), .A2(new_n11240_), .B(new_n11182_), .ZN(new_n11241_));
  NAND2_X1   g10233(.A1(new_n8467_), .A2(new_n8443_), .ZN(new_n11242_));
  OAI21_X1   g10234(.A1(new_n8464_), .A2(new_n8466_), .B(new_n8442_), .ZN(new_n11243_));
  AOI21_X1   g10235(.A1(new_n11242_), .A2(new_n11243_), .B(new_n8439_), .ZN(new_n11244_));
  NOR2_X1    g10236(.A1(new_n8428_), .A2(new_n8442_), .ZN(new_n11245_));
  INV_X1     g10237(.I(new_n11243_), .ZN(new_n11246_));
  NOR3_X1    g10238(.A1(new_n11246_), .A2(new_n11245_), .A3(new_n8473_), .ZN(new_n11247_));
  NOR2_X1    g10239(.A1(new_n11247_), .A2(new_n11244_), .ZN(new_n11248_));
  NAND2_X1   g10240(.A1(new_n8417_), .A2(new_n8474_), .ZN(new_n11249_));
  NOR3_X1    g10241(.A1(new_n8401_), .A2(new_n8416_), .A3(new_n8397_), .ZN(new_n11250_));
  AOI21_X1   g10242(.A1(new_n8448_), .A2(new_n8450_), .B(new_n8460_), .ZN(new_n11251_));
  OAI21_X1   g10243(.A1(new_n11251_), .A2(new_n11250_), .B(new_n8413_), .ZN(new_n11252_));
  NAND3_X1   g10244(.A1(new_n8460_), .A2(new_n8448_), .A3(new_n8450_), .ZN(new_n11253_));
  OAI21_X1   g10245(.A1(new_n8397_), .A2(new_n8401_), .B(new_n8416_), .ZN(new_n11254_));
  NAND3_X1   g10246(.A1(new_n11253_), .A2(new_n11254_), .A3(new_n8457_), .ZN(new_n11255_));
  NOR2_X1    g10247(.A1(new_n8413_), .A2(new_n8451_), .ZN(new_n11256_));
  NOR2_X1    g10248(.A1(new_n8402_), .A2(new_n8457_), .ZN(new_n11257_));
  OAI21_X1   g10249(.A1(new_n11256_), .A2(new_n11257_), .B(new_n8460_), .ZN(new_n11258_));
  NAND3_X1   g10250(.A1(new_n11258_), .A2(new_n11252_), .A3(new_n11255_), .ZN(new_n11259_));
  XOR2_X1    g10251(.A1(new_n11259_), .A2(new_n11249_), .Z(new_n11260_));
  NAND2_X1   g10252(.A1(new_n11260_), .A2(new_n11248_), .ZN(new_n11261_));
  OAI21_X1   g10253(.A1(new_n11246_), .A2(new_n11245_), .B(new_n8473_), .ZN(new_n11262_));
  NAND3_X1   g10254(.A1(new_n11242_), .A2(new_n8439_), .A3(new_n11243_), .ZN(new_n11263_));
  NAND2_X1   g10255(.A1(new_n11262_), .A2(new_n11263_), .ZN(new_n11264_));
  AOI22_X1   g10256(.A1(new_n8422_), .A2(new_n8427_), .B1(new_n8433_), .B2(new_n8438_), .ZN(new_n11265_));
  NOR4_X1    g10257(.A1(new_n8464_), .A2(new_n8466_), .A3(new_n8472_), .A4(new_n8470_), .ZN(new_n11266_));
  NOR2_X1    g10258(.A1(new_n8441_), .A2(new_n8437_), .ZN(new_n11267_));
  INV_X1     g10259(.I(new_n11267_), .ZN(new_n11268_));
  NAND4_X1   g10260(.A1(new_n11268_), .A2(new_n8423_), .A3(new_n8420_), .A4(new_n8418_), .ZN(new_n11269_));
  OAI22_X1   g10261(.A1(new_n11265_), .A2(new_n11266_), .B1(new_n11269_), .B2(new_n8473_), .ZN(new_n11270_));
  NOR4_X1    g10262(.A1(new_n11270_), .A2(new_n8402_), .A3(new_n8413_), .A4(new_n8416_), .ZN(new_n11271_));
  NAND2_X1   g10263(.A1(new_n11271_), .A2(new_n11264_), .ZN(new_n11272_));
  AOI21_X1   g10264(.A1(new_n11272_), .A2(new_n11259_), .B(new_n11249_), .ZN(new_n11273_));
  NOR4_X1    g10265(.A1(new_n8445_), .A2(new_n8475_), .A3(new_n8529_), .A4(new_n8559_), .ZN(new_n11274_));
  NAND2_X1   g10266(.A1(new_n8501_), .A2(new_n8558_), .ZN(new_n11275_));
  NAND3_X1   g10267(.A1(new_n8544_), .A2(new_n8532_), .A3(new_n8534_), .ZN(new_n11276_));
  OAI21_X1   g10268(.A1(new_n8481_), .A2(new_n8485_), .B(new_n8500_), .ZN(new_n11277_));
  AOI21_X1   g10269(.A1(new_n11276_), .A2(new_n11277_), .B(new_n8541_), .ZN(new_n11278_));
  NOR3_X1    g10270(.A1(new_n8485_), .A2(new_n8500_), .A3(new_n8481_), .ZN(new_n11279_));
  AOI21_X1   g10271(.A1(new_n8532_), .A2(new_n8534_), .B(new_n8544_), .ZN(new_n11280_));
  NOR3_X1    g10272(.A1(new_n11280_), .A2(new_n8497_), .A3(new_n11279_), .ZN(new_n11281_));
  NOR2_X1    g10273(.A1(new_n11281_), .A2(new_n11278_), .ZN(new_n11282_));
  NOR2_X1    g10274(.A1(new_n8497_), .A2(new_n8535_), .ZN(new_n11283_));
  NOR2_X1    g10275(.A1(new_n8486_), .A2(new_n8541_), .ZN(new_n11284_));
  OAI21_X1   g10276(.A1(new_n11283_), .A2(new_n11284_), .B(new_n8544_), .ZN(new_n11285_));
  NAND3_X1   g10277(.A1(new_n11282_), .A2(new_n11275_), .A3(new_n11285_), .ZN(new_n11286_));
  NAND2_X1   g10278(.A1(new_n8551_), .A2(new_n8527_), .ZN(new_n11287_));
  NAND2_X1   g10279(.A1(new_n8512_), .A2(new_n8526_), .ZN(new_n11288_));
  AOI21_X1   g10280(.A1(new_n11287_), .A2(new_n11288_), .B(new_n8523_), .ZN(new_n11289_));
  INV_X1     g10281(.I(new_n11289_), .ZN(new_n11290_));
  NAND3_X1   g10282(.A1(new_n11287_), .A2(new_n11288_), .A3(new_n8523_), .ZN(new_n11291_));
  NAND2_X1   g10283(.A1(new_n11290_), .A2(new_n11291_), .ZN(new_n11292_));
  NAND2_X1   g10284(.A1(new_n8512_), .A2(new_n8523_), .ZN(new_n11293_));
  NOR4_X1    g10285(.A1(new_n8548_), .A2(new_n8550_), .A3(new_n8556_), .A4(new_n8554_), .ZN(new_n11294_));
  INV_X1     g10286(.I(new_n11294_), .ZN(new_n11295_));
  NAND2_X1   g10287(.A1(new_n11295_), .A2(new_n11293_), .ZN(new_n11296_));
  NOR2_X1    g10288(.A1(new_n8525_), .A2(new_n8521_), .ZN(new_n11297_));
  OR4_X2     g10289(.A1(\A[367] ), .A2(new_n11297_), .A3(\A[368] ), .A4(\A[369] ), .Z(new_n11298_));
  NAND4_X1   g10290(.A1(new_n11296_), .A2(new_n8535_), .A3(new_n8541_), .A4(new_n8544_), .ZN(new_n11300_));
  NAND4_X1   g10291(.A1(new_n11274_), .A2(new_n11286_), .A3(new_n11292_), .A4(new_n11300_), .ZN(new_n11301_));
  NOR2_X1    g10292(.A1(new_n11273_), .A2(new_n11301_), .ZN(new_n11302_));
  NAND2_X1   g10293(.A1(new_n11273_), .A2(new_n11301_), .ZN(new_n11303_));
  INV_X1     g10294(.I(new_n11303_), .ZN(new_n11304_));
  OAI21_X1   g10295(.A1(new_n11304_), .A2(new_n11302_), .B(new_n11261_), .ZN(new_n11305_));
  NOR2_X1    g10296(.A1(new_n8461_), .A2(new_n8444_), .ZN(new_n11306_));
  XOR2_X1    g10297(.A1(new_n11259_), .A2(new_n11306_), .Z(new_n11307_));
  NOR2_X1    g10298(.A1(new_n11307_), .A2(new_n11264_), .ZN(new_n11308_));
  INV_X1     g10299(.I(new_n11302_), .ZN(new_n11309_));
  NAND3_X1   g10300(.A1(new_n11309_), .A2(new_n11308_), .A3(new_n11303_), .ZN(new_n11310_));
  NAND2_X1   g10301(.A1(new_n11305_), .A2(new_n11310_), .ZN(new_n11311_));
  NAND3_X1   g10302(.A1(new_n11311_), .A2(new_n8566_), .A3(new_n11241_), .ZN(new_n11312_));
  INV_X1     g10303(.I(new_n11182_), .ZN(new_n11313_));
  INV_X1     g10304(.I(new_n11240_), .ZN(new_n11314_));
  AOI21_X1   g10305(.A1(new_n11314_), .A2(new_n11238_), .B(new_n11313_), .ZN(new_n11315_));
  NAND3_X1   g10306(.A1(new_n11311_), .A2(new_n8566_), .A3(new_n11315_), .ZN(new_n11316_));
  NAND2_X1   g10307(.A1(new_n11316_), .A2(new_n11312_), .ZN(new_n11317_));
  NAND3_X1   g10308(.A1(new_n11317_), .A2(new_n8883_), .A3(new_n8884_), .ZN(new_n11318_));
  NAND2_X1   g10309(.A1(new_n11318_), .A2(new_n11161_), .ZN(new_n11319_));
  NAND2_X1   g10310(.A1(new_n9000_), .A2(new_n8936_), .ZN(new_n11320_));
  INV_X1     g10311(.I(new_n8936_), .ZN(new_n11321_));
  NAND2_X1   g10312(.A1(new_n11321_), .A2(new_n8922_), .ZN(new_n11322_));
  AOI21_X1   g10313(.A1(new_n11322_), .A2(new_n11320_), .B(new_n8933_), .ZN(new_n11323_));
  INV_X1     g10314(.I(new_n8933_), .ZN(new_n11324_));
  NOR2_X1    g10315(.A1(new_n11321_), .A2(new_n8922_), .ZN(new_n11325_));
  NOR2_X1    g10316(.A1(new_n9000_), .A2(new_n8936_), .ZN(new_n11326_));
  NOR3_X1    g10317(.A1(new_n11325_), .A2(new_n11326_), .A3(new_n11324_), .ZN(new_n11327_));
  OR2_X2     g10318(.A1(new_n11327_), .A2(new_n11323_), .Z(new_n11328_));
  NAND2_X1   g10319(.A1(new_n9007_), .A2(new_n8933_), .ZN(new_n11329_));
  NAND3_X1   g10320(.A1(new_n8958_), .A2(new_n8927_), .A3(new_n8932_), .ZN(new_n11330_));
  NAND2_X1   g10321(.A1(new_n9000_), .A2(new_n8947_), .ZN(new_n11331_));
  NAND3_X1   g10322(.A1(new_n8922_), .A2(new_n8942_), .A3(new_n8946_), .ZN(new_n11332_));
  AOI22_X1   g10323(.A1(new_n11329_), .A2(new_n11330_), .B1(new_n11332_), .B2(new_n11331_), .ZN(new_n11333_));
  NAND3_X1   g10324(.A1(new_n8922_), .A2(new_n8933_), .A3(new_n8936_), .ZN(new_n11334_));
  NAND3_X1   g10325(.A1(new_n8958_), .A2(new_n8947_), .A3(new_n8963_), .ZN(new_n11335_));
  NAND2_X1   g10326(.A1(new_n11334_), .A2(new_n11335_), .ZN(new_n11336_));
  INV_X1     g10327(.I(new_n11336_), .ZN(new_n11337_));
  NAND2_X1   g10328(.A1(new_n11337_), .A2(new_n11333_), .ZN(new_n11338_));
  NAND2_X1   g10329(.A1(new_n8940_), .A2(\A[363] ), .ZN(new_n11339_));
  NAND2_X1   g10330(.A1(new_n8938_), .A2(\A[362] ), .ZN(new_n11340_));
  AOI21_X1   g10331(.A1(new_n11339_), .A2(new_n11340_), .B(new_n8943_), .ZN(new_n11341_));
  INV_X1     g10332(.I(new_n8944_), .ZN(new_n11342_));
  NAND2_X1   g10333(.A1(\A[362] ), .A2(\A[363] ), .ZN(new_n11343_));
  AOI21_X1   g10334(.A1(new_n11342_), .A2(new_n11343_), .B(\A[361] ), .ZN(new_n11344_));
  OAI22_X1   g10335(.A1(new_n8944_), .A2(new_n8959_), .B1(new_n8961_), .B2(new_n8956_), .ZN(new_n11345_));
  NOR3_X1    g10336(.A1(new_n11344_), .A2(new_n11345_), .A3(new_n11341_), .ZN(new_n11346_));
  INV_X1     g10337(.I(new_n8960_), .ZN(new_n11347_));
  INV_X1     g10338(.I(new_n8962_), .ZN(new_n11348_));
  AOI22_X1   g10339(.A1(new_n11347_), .A2(new_n11348_), .B1(new_n8942_), .B2(new_n8946_), .ZN(new_n11349_));
  OAI21_X1   g10340(.A1(new_n11349_), .A2(new_n11346_), .B(new_n9007_), .ZN(new_n11350_));
  NAND3_X1   g10341(.A1(new_n8963_), .A2(new_n8942_), .A3(new_n8946_), .ZN(new_n11351_));
  OAI21_X1   g10342(.A1(new_n11341_), .A2(new_n11344_), .B(new_n11345_), .ZN(new_n11352_));
  NAND3_X1   g10343(.A1(new_n11351_), .A2(new_n11352_), .A3(new_n8958_), .ZN(new_n11353_));
  NAND2_X1   g10344(.A1(new_n11350_), .A2(new_n11353_), .ZN(new_n11354_));
  XOR2_X1    g10345(.A1(new_n11338_), .A2(new_n11354_), .Z(new_n11355_));
  NOR2_X1    g10346(.A1(new_n11355_), .A2(new_n11328_), .ZN(new_n11356_));
  INV_X1     g10347(.I(new_n11356_), .ZN(new_n11357_));
  INV_X1     g10348(.I(new_n11338_), .ZN(new_n11358_));
  NOR2_X1    g10349(.A1(new_n11327_), .A2(new_n11323_), .ZN(new_n11359_));
  NAND2_X1   g10350(.A1(new_n8960_), .A2(new_n8962_), .ZN(new_n11360_));
  NAND3_X1   g10351(.A1(new_n8958_), .A2(new_n8947_), .A3(new_n11360_), .ZN(new_n11361_));
  NOR2_X1    g10352(.A1(new_n11334_), .A2(new_n11361_), .ZN(new_n11362_));
  NAND3_X1   g10353(.A1(new_n11333_), .A2(new_n11354_), .A3(new_n11362_), .ZN(new_n11363_));
  NOR2_X1    g10354(.A1(new_n11363_), .A2(new_n11359_), .ZN(new_n11364_));
  OAI21_X1   g10355(.A1(new_n11364_), .A2(new_n11354_), .B(new_n11358_), .ZN(new_n11365_));
  XOR2_X1    g10356(.A1(new_n8911_), .A2(new_n8937_), .Z(new_n11366_));
  NAND3_X1   g10357(.A1(new_n8991_), .A2(new_n9011_), .A3(new_n9013_), .ZN(new_n11367_));
  OAI22_X1   g10358(.A1(new_n8971_), .A2(new_n8987_), .B1(new_n8989_), .B2(new_n8984_), .ZN(new_n11368_));
  OAI21_X1   g10359(.A1(new_n8970_), .A2(new_n8974_), .B(new_n11368_), .ZN(new_n11369_));
  AOI21_X1   g10360(.A1(new_n11367_), .A2(new_n11369_), .B(new_n8986_), .ZN(new_n11370_));
  NAND2_X1   g10361(.A1(new_n8978_), .A2(\A[354] ), .ZN(new_n11371_));
  NAND2_X1   g10362(.A1(new_n8976_), .A2(\A[353] ), .ZN(new_n11372_));
  AOI21_X1   g10363(.A1(new_n11371_), .A2(new_n11372_), .B(new_n8981_), .ZN(new_n11373_));
  INV_X1     g10364(.I(new_n8984_), .ZN(new_n11374_));
  AOI21_X1   g10365(.A1(new_n11374_), .A2(new_n8982_), .B(\A[352] ), .ZN(new_n11375_));
  NOR2_X1    g10366(.A1(new_n11375_), .A2(new_n11373_), .ZN(new_n11376_));
  NOR3_X1    g10367(.A1(new_n8974_), .A2(new_n11368_), .A3(new_n8970_), .ZN(new_n11377_));
  AOI21_X1   g10368(.A1(new_n9011_), .A2(new_n9013_), .B(new_n8991_), .ZN(new_n11378_));
  NOR3_X1    g10369(.A1(new_n11378_), .A2(new_n11376_), .A3(new_n11377_), .ZN(new_n11379_));
  NOR2_X1    g10370(.A1(new_n11379_), .A2(new_n11370_), .ZN(new_n11380_));
  NAND2_X1   g10371(.A1(new_n11376_), .A2(new_n8907_), .ZN(new_n11381_));
  NOR2_X1    g10372(.A1(new_n11376_), .A2(new_n8907_), .ZN(new_n11382_));
  INV_X1     g10373(.I(new_n11382_), .ZN(new_n11383_));
  NAND2_X1   g10374(.A1(new_n8896_), .A2(new_n9014_), .ZN(new_n11384_));
  NOR2_X1    g10375(.A1(new_n8889_), .A2(\A[344] ), .ZN(new_n11385_));
  NOR2_X1    g10376(.A1(new_n8887_), .A2(\A[345] ), .ZN(new_n11386_));
  OAI21_X1   g10377(.A1(new_n11385_), .A2(new_n11386_), .B(\A[343] ), .ZN(new_n11387_));
  INV_X1     g10378(.I(new_n8894_), .ZN(new_n11388_));
  OAI21_X1   g10379(.A1(new_n11388_), .A2(new_n8892_), .B(new_n8886_), .ZN(new_n11389_));
  NAND2_X1   g10380(.A1(new_n11387_), .A2(new_n11389_), .ZN(new_n11390_));
  NAND2_X1   g10381(.A1(new_n8975_), .A2(new_n11390_), .ZN(new_n11391_));
  AOI22_X1   g10382(.A1(new_n11383_), .A2(new_n11381_), .B1(new_n11384_), .B2(new_n11391_), .ZN(new_n11392_));
  NOR4_X1    g10383(.A1(new_n8908_), .A2(\A[346] ), .A3(\A[347] ), .A4(\A[348] ), .ZN(new_n11393_));
  NOR2_X1    g10384(.A1(new_n11376_), .A2(new_n11368_), .ZN(new_n11394_));
  AOI22_X1   g10385(.A1(new_n11394_), .A2(new_n9014_), .B1(new_n11390_), .B2(new_n11393_), .ZN(new_n11395_));
  NAND2_X1   g10386(.A1(new_n11392_), .A2(new_n11395_), .ZN(new_n11396_));
  INV_X1     g10387(.I(new_n8907_), .ZN(new_n11397_));
  NAND2_X1   g10388(.A1(new_n8896_), .A2(new_n8910_), .ZN(new_n11398_));
  INV_X1     g10389(.I(new_n11398_), .ZN(new_n11399_));
  NOR2_X1    g10390(.A1(new_n8896_), .A2(new_n8910_), .ZN(new_n11400_));
  OAI21_X1   g10391(.A1(new_n11399_), .A2(new_n11400_), .B(new_n11397_), .ZN(new_n11401_));
  INV_X1     g10392(.I(new_n11400_), .ZN(new_n11402_));
  NAND3_X1   g10393(.A1(new_n11402_), .A2(new_n11398_), .A3(new_n8907_), .ZN(new_n11403_));
  NAND2_X1   g10394(.A1(new_n11401_), .A2(new_n11403_), .ZN(new_n11404_));
  INV_X1     g10395(.I(new_n11381_), .ZN(new_n11405_));
  NOR2_X1    g10396(.A1(new_n8975_), .A2(new_n11390_), .ZN(new_n11406_));
  NOR2_X1    g10397(.A1(new_n8896_), .A2(new_n9014_), .ZN(new_n11407_));
  OAI22_X1   g10398(.A1(new_n11405_), .A2(new_n11382_), .B1(new_n11406_), .B2(new_n11407_), .ZN(new_n11408_));
  NAND2_X1   g10399(.A1(new_n11390_), .A2(new_n11393_), .ZN(new_n11409_));
  NAND2_X1   g10400(.A1(new_n8988_), .A2(new_n8990_), .ZN(new_n11410_));
  NAND3_X1   g10401(.A1(new_n9014_), .A2(new_n8986_), .A3(new_n11410_), .ZN(new_n11411_));
  OR2_X2     g10402(.A1(new_n11411_), .A2(new_n11409_), .Z(new_n11412_));
  NAND3_X1   g10403(.A1(new_n11396_), .A2(new_n11404_), .A3(new_n11380_), .ZN(new_n11414_));
  NOR3_X1    g10404(.A1(new_n11414_), .A2(new_n11366_), .A3(new_n8993_), .ZN(new_n11415_));
  NAND2_X1   g10405(.A1(new_n11415_), .A2(new_n11365_), .ZN(new_n11416_));
  OR2_X2     g10406(.A1(new_n11415_), .A2(new_n11365_), .Z(new_n11417_));
  AOI21_X1   g10407(.A1(new_n11417_), .A2(new_n11416_), .B(new_n11357_), .ZN(new_n11418_));
  INV_X1     g10408(.I(new_n11418_), .ZN(new_n11419_));
  NAND4_X1   g10409(.A1(new_n9020_), .A2(new_n9024_), .A3(new_n9187_), .A4(new_n9188_), .ZN(new_n11420_));
  NAND2_X1   g10410(.A1(new_n9075_), .A2(new_n9089_), .ZN(new_n11421_));
  INV_X1     g10411(.I(new_n9089_), .ZN(new_n11422_));
  NAND2_X1   g10412(.A1(new_n11422_), .A2(new_n9181_), .ZN(new_n11423_));
  AOI21_X1   g10413(.A1(new_n11423_), .A2(new_n11421_), .B(new_n9086_), .ZN(new_n11424_));
  AND3_X2    g10414(.A1(new_n11423_), .A2(new_n9086_), .A3(new_n11421_), .Z(new_n11425_));
  NOR2_X1    g10415(.A1(new_n11425_), .A2(new_n11424_), .ZN(new_n11426_));
  NAND3_X1   g10416(.A1(new_n9181_), .A2(new_n9086_), .A3(new_n9089_), .ZN(new_n11427_));
  NAND3_X1   g10417(.A1(new_n9101_), .A2(new_n9112_), .A3(new_n9116_), .ZN(new_n11428_));
  NOR2_X1    g10418(.A1(new_n11427_), .A2(new_n11428_), .ZN(new_n11429_));
  NAND2_X1   g10419(.A1(new_n9163_), .A2(new_n9116_), .ZN(new_n11430_));
  OAI21_X1   g10420(.A1(new_n9160_), .A2(new_n9162_), .B(new_n9115_), .ZN(new_n11431_));
  AOI21_X1   g10421(.A1(new_n11430_), .A2(new_n11431_), .B(new_n9112_), .ZN(new_n11432_));
  NAND2_X1   g10422(.A1(new_n9104_), .A2(\A[342] ), .ZN(new_n11433_));
  NAND2_X1   g10423(.A1(new_n9102_), .A2(\A[341] ), .ZN(new_n11434_));
  AOI21_X1   g10424(.A1(new_n11433_), .A2(new_n11434_), .B(new_n9107_), .ZN(new_n11435_));
  INV_X1     g10425(.I(new_n9110_), .ZN(new_n11436_));
  AOI21_X1   g10426(.A1(new_n11436_), .A2(new_n9108_), .B(\A[340] ), .ZN(new_n11437_));
  NOR2_X1    g10427(.A1(new_n11437_), .A2(new_n11435_), .ZN(new_n11438_));
  NOR2_X1    g10428(.A1(new_n9101_), .A2(new_n9115_), .ZN(new_n11439_));
  INV_X1     g10429(.I(new_n11431_), .ZN(new_n11440_));
  NOR3_X1    g10430(.A1(new_n11440_), .A2(new_n11439_), .A3(new_n11438_), .ZN(new_n11441_));
  NOR2_X1    g10431(.A1(new_n11441_), .A2(new_n11432_), .ZN(new_n11442_));
  NOR2_X1    g10432(.A1(new_n11442_), .A2(new_n11429_), .ZN(new_n11443_));
  INV_X1     g10433(.I(new_n11429_), .ZN(new_n11444_));
  OAI21_X1   g10434(.A1(new_n11440_), .A2(new_n11439_), .B(new_n11438_), .ZN(new_n11445_));
  NAND3_X1   g10435(.A1(new_n11430_), .A2(new_n9112_), .A3(new_n11431_), .ZN(new_n11446_));
  NAND2_X1   g10436(.A1(new_n11445_), .A2(new_n11446_), .ZN(new_n11447_));
  NOR2_X1    g10437(.A1(new_n11447_), .A2(new_n11444_), .ZN(new_n11448_));
  OAI21_X1   g10438(.A1(new_n11448_), .A2(new_n11443_), .B(new_n11426_), .ZN(new_n11449_));
  NAND2_X1   g10439(.A1(new_n9078_), .A2(\A[336] ), .ZN(new_n11450_));
  NAND2_X1   g10440(.A1(new_n9076_), .A2(\A[335] ), .ZN(new_n11451_));
  AOI21_X1   g10441(.A1(new_n11450_), .A2(new_n11451_), .B(new_n9081_), .ZN(new_n11452_));
  INV_X1     g10442(.I(new_n9084_), .ZN(new_n11453_));
  AOI21_X1   g10443(.A1(new_n11453_), .A2(new_n9082_), .B(\A[334] ), .ZN(new_n11454_));
  NOR2_X1    g10444(.A1(new_n11454_), .A2(new_n11452_), .ZN(new_n11455_));
  NOR2_X1    g10445(.A1(new_n9075_), .A2(new_n11455_), .ZN(new_n11456_));
  NOR2_X1    g10446(.A1(new_n9181_), .A2(new_n9086_), .ZN(new_n11457_));
  OR4_X2     g10447(.A1(new_n9097_), .A2(new_n9113_), .A3(new_n9114_), .A4(new_n9110_), .Z(new_n11458_));
  NAND3_X1   g10448(.A1(new_n9101_), .A2(new_n9112_), .A3(new_n11458_), .ZN(new_n11459_));
  NOR3_X1    g10449(.A1(new_n11456_), .A2(new_n11459_), .A3(new_n11457_), .ZN(new_n11460_));
  NAND2_X1   g10450(.A1(new_n9181_), .A2(new_n9089_), .ZN(new_n11461_));
  NOR2_X1    g10451(.A1(new_n9163_), .A2(new_n11438_), .ZN(new_n11462_));
  NOR2_X1    g10452(.A1(new_n9101_), .A2(new_n9112_), .ZN(new_n11463_));
  NOR4_X1    g10453(.A1(new_n11462_), .A2(new_n11463_), .A3(new_n11461_), .A4(new_n11455_), .ZN(new_n11464_));
  NAND3_X1   g10454(.A1(new_n11447_), .A2(new_n11460_), .A3(new_n11464_), .ZN(new_n11465_));
  NOR4_X1    g10455(.A1(new_n11427_), .A2(new_n9163_), .A3(new_n11438_), .A4(new_n9115_), .ZN(new_n11467_));
  AOI22_X1   g10456(.A1(new_n9048_), .A2(new_n9050_), .B1(new_n9053_), .B2(new_n9055_), .ZN(new_n11468_));
  NOR4_X1    g10457(.A1(new_n9030_), .A2(new_n9034_), .A3(new_n9044_), .A4(new_n9040_), .ZN(new_n11469_));
  NOR2_X1    g10458(.A1(new_n11468_), .A2(new_n11469_), .ZN(new_n11470_));
  NAND2_X1   g10459(.A1(new_n9053_), .A2(new_n9055_), .ZN(new_n11471_));
  NOR2_X1    g10460(.A1(new_n9061_), .A2(new_n9042_), .ZN(new_n11472_));
  NOR4_X1    g10461(.A1(new_n11472_), .A2(\A[319] ), .A3(\A[320] ), .A4(\A[321] ), .ZN(new_n11473_));
  NAND4_X1   g10462(.A1(new_n11471_), .A2(new_n9151_), .A3(new_n11473_), .A4(new_n9154_), .ZN(new_n11474_));
  NOR3_X1    g10463(.A1(new_n11470_), .A2(new_n9150_), .A3(new_n11474_), .ZN(new_n11475_));
  NOR3_X1    g10464(.A1(new_n9143_), .A2(new_n9171_), .A3(new_n9140_), .ZN(new_n11476_));
  NOR2_X1    g10465(.A1(new_n9170_), .A2(new_n9125_), .ZN(new_n11477_));
  INV_X1     g10466(.I(new_n11477_), .ZN(new_n11478_));
  INV_X1     g10467(.I(new_n9153_), .ZN(new_n11479_));
  AOI22_X1   g10468(.A1(new_n11478_), .A2(new_n11479_), .B1(new_n9122_), .B2(new_n9126_), .ZN(new_n11480_));
  OAI21_X1   g10469(.A1(new_n11480_), .A2(new_n11476_), .B(new_n9169_), .ZN(new_n11481_));
  NOR2_X1    g10470(.A1(new_n11477_), .A2(new_n9153_), .ZN(new_n11482_));
  NAND3_X1   g10471(.A1(new_n11482_), .A2(new_n9122_), .A3(new_n9126_), .ZN(new_n11483_));
  OAI21_X1   g10472(.A1(new_n9140_), .A2(new_n9143_), .B(new_n9171_), .ZN(new_n11484_));
  NAND3_X1   g10473(.A1(new_n11483_), .A2(new_n11484_), .A3(new_n9151_), .ZN(new_n11485_));
  NAND2_X1   g10474(.A1(new_n11477_), .A2(new_n9153_), .ZN(new_n11486_));
  INV_X1     g10475(.I(new_n11486_), .ZN(new_n11487_));
  NAND3_X1   g10476(.A1(new_n9165_), .A2(new_n9166_), .A3(new_n9171_), .ZN(new_n11488_));
  NAND3_X1   g10477(.A1(new_n11488_), .A2(new_n11481_), .A3(new_n11485_), .ZN(new_n11489_));
  NOR3_X1    g10478(.A1(new_n9034_), .A2(new_n9062_), .A3(new_n9030_), .ZN(new_n11490_));
  NOR2_X1    g10479(.A1(new_n9060_), .A2(new_n9032_), .ZN(new_n11491_));
  INV_X1     g10480(.I(new_n11491_), .ZN(new_n11492_));
  INV_X1     g10481(.I(new_n11472_), .ZN(new_n11493_));
  AOI22_X1   g10482(.A1(new_n11492_), .A2(new_n11493_), .B1(new_n9048_), .B2(new_n9050_), .ZN(new_n11494_));
  OAI21_X1   g10483(.A1(new_n11494_), .A2(new_n11490_), .B(new_n9059_), .ZN(new_n11495_));
  NOR2_X1    g10484(.A1(new_n11491_), .A2(new_n11472_), .ZN(new_n11496_));
  NAND3_X1   g10485(.A1(new_n11496_), .A2(new_n9048_), .A3(new_n9050_), .ZN(new_n11497_));
  OAI21_X1   g10486(.A1(new_n9030_), .A2(new_n9034_), .B(new_n9062_), .ZN(new_n11498_));
  NAND3_X1   g10487(.A1(new_n11497_), .A2(new_n11498_), .A3(new_n11471_), .ZN(new_n11499_));
  NAND2_X1   g10488(.A1(new_n11495_), .A2(new_n11499_), .ZN(new_n11500_));
  NOR3_X1    g10489(.A1(new_n11489_), .A2(new_n11475_), .A3(new_n11500_), .ZN(new_n11501_));
  NAND4_X1   g10490(.A1(new_n9057_), .A2(new_n9167_), .A3(new_n9063_), .A4(new_n9172_), .ZN(new_n11502_));
  AOI21_X1   g10491(.A1(new_n11483_), .A2(new_n11484_), .B(new_n9151_), .ZN(new_n11503_));
  NOR3_X1    g10492(.A1(new_n11480_), .A2(new_n11476_), .A3(new_n9169_), .ZN(new_n11504_));
  NOR3_X1    g10493(.A1(new_n9149_), .A2(new_n9137_), .A3(new_n11482_), .ZN(new_n11505_));
  NOR3_X1    g10494(.A1(new_n11505_), .A2(new_n11504_), .A3(new_n11503_), .ZN(new_n11506_));
  AOI21_X1   g10495(.A1(new_n11497_), .A2(new_n11498_), .B(new_n11471_), .ZN(new_n11507_));
  NOR3_X1    g10496(.A1(new_n11494_), .A2(new_n9059_), .A3(new_n11490_), .ZN(new_n11508_));
  NOR2_X1    g10497(.A1(new_n11508_), .A2(new_n11507_), .ZN(new_n11509_));
  AOI21_X1   g10498(.A1(new_n11506_), .A2(new_n11502_), .B(new_n11509_), .ZN(new_n11510_));
  NOR2_X1    g10499(.A1(new_n11510_), .A2(new_n11501_), .ZN(new_n11511_));
  NAND2_X1   g10500(.A1(new_n11481_), .A2(new_n11485_), .ZN(new_n11512_));
  AOI21_X1   g10501(.A1(new_n9137_), .A2(new_n11486_), .B(new_n11482_), .ZN(new_n11513_));
  NOR3_X1    g10502(.A1(new_n11470_), .A2(new_n11513_), .A3(new_n9150_), .ZN(new_n11514_));
  AOI21_X1   g10503(.A1(new_n11514_), .A2(new_n11512_), .B(new_n9063_), .ZN(new_n11515_));
  NOR2_X1    g10504(.A1(new_n11513_), .A2(new_n9150_), .ZN(new_n11516_));
  INV_X1     g10505(.I(new_n11516_), .ZN(new_n11517_));
  NOR2_X1    g10506(.A1(new_n11506_), .A2(new_n11475_), .ZN(new_n11518_));
  OAI21_X1   g10507(.A1(new_n11515_), .A2(new_n11517_), .B(new_n11518_), .ZN(new_n11519_));
  NOR2_X1    g10508(.A1(new_n9064_), .A2(new_n9090_), .ZN(new_n11520_));
  NAND2_X1   g10509(.A1(new_n11471_), .A2(new_n11473_), .ZN(new_n11521_));
  NAND3_X1   g10510(.A1(new_n11521_), .A2(new_n9045_), .A3(new_n9056_), .ZN(new_n11522_));
  NOR2_X1    g10511(.A1(new_n9182_), .A2(new_n11522_), .ZN(new_n11523_));
  OAI22_X1   g10512(.A1(new_n9157_), .A2(new_n9174_), .B1(new_n11520_), .B2(new_n11523_), .ZN(new_n11524_));
  NOR4_X1    g10513(.A1(new_n11519_), .A2(new_n11511_), .A3(new_n11524_), .A4(new_n11467_), .ZN(new_n11525_));
  INV_X1     g10514(.I(new_n11467_), .ZN(new_n11526_));
  AOI22_X1   g10515(.A1(new_n9045_), .A2(new_n9056_), .B1(new_n9165_), .B2(new_n9166_), .ZN(new_n11527_));
  OAI21_X1   g10516(.A1(new_n9165_), .A2(new_n11487_), .B(new_n9171_), .ZN(new_n11528_));
  NAND3_X1   g10517(.A1(new_n11512_), .A2(new_n11527_), .A3(new_n11528_), .ZN(new_n11529_));
  AOI21_X1   g10518(.A1(new_n11529_), .A2(new_n11521_), .B(new_n11517_), .ZN(new_n11530_));
  NOR4_X1    g10519(.A1(new_n11530_), .A2(new_n11475_), .A3(new_n11506_), .A4(new_n11509_), .ZN(new_n11531_));
  NAND2_X1   g10520(.A1(new_n9182_), .A2(new_n11522_), .ZN(new_n11532_));
  NAND2_X1   g10521(.A1(new_n9064_), .A2(new_n9090_), .ZN(new_n11533_));
  AOI22_X1   g10522(.A1(new_n9183_), .A2(new_n9184_), .B1(new_n11533_), .B2(new_n11532_), .ZN(new_n11534_));
  AOI21_X1   g10523(.A1(new_n11531_), .A2(new_n11534_), .B(new_n11526_), .ZN(new_n11535_));
  OAI21_X1   g10524(.A1(new_n11535_), .A2(new_n11525_), .B(new_n11449_), .ZN(new_n11536_));
  INV_X1     g10525(.I(new_n11424_), .ZN(new_n11537_));
  NAND3_X1   g10526(.A1(new_n11423_), .A2(new_n11421_), .A3(new_n9086_), .ZN(new_n11538_));
  NAND2_X1   g10527(.A1(new_n11537_), .A2(new_n11538_), .ZN(new_n11539_));
  NAND2_X1   g10528(.A1(new_n11447_), .A2(new_n11444_), .ZN(new_n11540_));
  NAND2_X1   g10529(.A1(new_n11442_), .A2(new_n11429_), .ZN(new_n11541_));
  AOI21_X1   g10530(.A1(new_n11540_), .A2(new_n11541_), .B(new_n11539_), .ZN(new_n11542_));
  NAND3_X1   g10531(.A1(new_n11531_), .A2(new_n11526_), .A3(new_n11534_), .ZN(new_n11543_));
  NAND3_X1   g10532(.A1(new_n11506_), .A2(new_n11502_), .A3(new_n11509_), .ZN(new_n11544_));
  OAI21_X1   g10533(.A1(new_n11489_), .A2(new_n11475_), .B(new_n11500_), .ZN(new_n11545_));
  NAND2_X1   g10534(.A1(new_n11545_), .A2(new_n11544_), .ZN(new_n11546_));
  NOR2_X1    g10535(.A1(new_n11504_), .A2(new_n11503_), .ZN(new_n11547_));
  NAND3_X1   g10536(.A1(new_n11528_), .A2(new_n9057_), .A3(new_n9167_), .ZN(new_n11548_));
  OAI21_X1   g10537(.A1(new_n11548_), .A2(new_n11547_), .B(new_n11521_), .ZN(new_n11549_));
  NAND2_X1   g10538(.A1(new_n11502_), .A2(new_n11489_), .ZN(new_n11550_));
  AOI21_X1   g10539(.A1(new_n11549_), .A2(new_n11516_), .B(new_n11550_), .ZN(new_n11551_));
  NAND3_X1   g10540(.A1(new_n11551_), .A2(new_n11546_), .A3(new_n11534_), .ZN(new_n11552_));
  NAND2_X1   g10541(.A1(new_n11552_), .A2(new_n11467_), .ZN(new_n11553_));
  NAND3_X1   g10542(.A1(new_n11553_), .A2(new_n11543_), .A3(new_n11542_), .ZN(new_n11554_));
  AOI21_X1   g10543(.A1(new_n11554_), .A2(new_n11536_), .B(new_n11420_), .ZN(new_n11555_));
  NOR2_X1    g10544(.A1(new_n9220_), .A2(new_n9276_), .ZN(new_n11556_));
  INV_X1     g10545(.I(new_n11556_), .ZN(new_n11557_));
  NOR3_X1    g10546(.A1(new_n9252_), .A2(new_n9218_), .A3(new_n9250_), .ZN(new_n11558_));
  OAI21_X1   g10547(.A1(new_n9250_), .A2(new_n9252_), .B(new_n9218_), .ZN(new_n11559_));
  INV_X1     g10548(.I(new_n11559_), .ZN(new_n11560_));
  OAI21_X1   g10549(.A1(new_n11560_), .A2(new_n11558_), .B(new_n9259_), .ZN(new_n11561_));
  INV_X1     g10550(.I(new_n11558_), .ZN(new_n11562_));
  NAND3_X1   g10551(.A1(new_n11562_), .A2(new_n9215_), .A3(new_n11559_), .ZN(new_n11563_));
  NOR2_X1    g10552(.A1(new_n9259_), .A2(new_n9204_), .ZN(new_n11564_));
  NOR2_X1    g10553(.A1(new_n9253_), .A2(new_n9215_), .ZN(new_n11565_));
  OAI21_X1   g10554(.A1(new_n11564_), .A2(new_n11565_), .B(new_n9219_), .ZN(new_n11566_));
  NAND3_X1   g10555(.A1(new_n11566_), .A2(new_n11561_), .A3(new_n11563_), .ZN(new_n11567_));
  NAND2_X1   g10556(.A1(new_n11561_), .A2(new_n11563_), .ZN(new_n11568_));
  AOI22_X1   g10557(.A1(new_n9263_), .A2(new_n9265_), .B1(new_n9269_), .B2(new_n9271_), .ZN(new_n11569_));
  NOR4_X1    g10558(.A1(new_n9226_), .A2(new_n9230_), .A3(new_n9241_), .A4(new_n9237_), .ZN(new_n11570_));
  NOR2_X1    g10559(.A1(new_n11569_), .A2(new_n11570_), .ZN(new_n11571_));
  NOR3_X1    g10560(.A1(new_n9231_), .A2(new_n9242_), .A3(new_n9245_), .ZN(new_n11572_));
  NOR3_X1    g10561(.A1(new_n11571_), .A2(new_n9220_), .A3(new_n11572_), .ZN(new_n11573_));
  NOR3_X1    g10562(.A1(new_n9230_), .A2(new_n9245_), .A3(new_n9226_), .ZN(new_n11574_));
  AOI21_X1   g10563(.A1(new_n9263_), .A2(new_n9265_), .B(new_n9275_), .ZN(new_n11575_));
  OAI21_X1   g10564(.A1(new_n11575_), .A2(new_n11574_), .B(new_n9242_), .ZN(new_n11576_));
  NAND3_X1   g10565(.A1(new_n9275_), .A2(new_n9263_), .A3(new_n9265_), .ZN(new_n11577_));
  OAI21_X1   g10566(.A1(new_n9226_), .A2(new_n9230_), .B(new_n9245_), .ZN(new_n11578_));
  NAND3_X1   g10567(.A1(new_n11577_), .A2(new_n11578_), .A3(new_n9272_), .ZN(new_n11579_));
  NAND2_X1   g10568(.A1(new_n11576_), .A2(new_n11579_), .ZN(new_n11580_));
  NAND4_X1   g10569(.A1(new_n11568_), .A2(new_n11573_), .A3(new_n11580_), .A4(new_n11566_), .ZN(new_n11581_));
  AOI21_X1   g10570(.A1(new_n11581_), .A2(new_n11567_), .B(new_n11557_), .ZN(new_n11582_));
  INV_X1     g10571(.I(new_n11580_), .ZN(new_n11583_));
  NOR2_X1    g10572(.A1(new_n11567_), .A2(new_n11556_), .ZN(new_n11584_));
  AOI21_X1   g10573(.A1(new_n11562_), .A2(new_n11559_), .B(new_n9215_), .ZN(new_n11585_));
  NOR3_X1    g10574(.A1(new_n11560_), .A2(new_n9259_), .A3(new_n11558_), .ZN(new_n11586_));
  NAND2_X1   g10575(.A1(new_n9253_), .A2(new_n9215_), .ZN(new_n11587_));
  NAND2_X1   g10576(.A1(new_n9259_), .A2(new_n9204_), .ZN(new_n11588_));
  AOI21_X1   g10577(.A1(new_n11587_), .A2(new_n11588_), .B(new_n9218_), .ZN(new_n11589_));
  NOR3_X1    g10578(.A1(new_n11589_), .A2(new_n11585_), .A3(new_n11586_), .ZN(new_n11590_));
  NOR2_X1    g10579(.A1(new_n11590_), .A2(new_n11557_), .ZN(new_n11591_));
  OAI21_X1   g10580(.A1(new_n11591_), .A2(new_n11584_), .B(new_n11583_), .ZN(new_n11592_));
  NOR2_X1    g10581(.A1(new_n9305_), .A2(new_n9359_), .ZN(new_n11593_));
  NOR3_X1    g10582(.A1(new_n9337_), .A2(new_n9303_), .A3(new_n9335_), .ZN(new_n11594_));
  NOR2_X1    g10583(.A1(new_n9338_), .A2(new_n9304_), .ZN(new_n11595_));
  OAI21_X1   g10584(.A1(new_n11595_), .A2(new_n11594_), .B(new_n9344_), .ZN(new_n11596_));
  NAND3_X1   g10585(.A1(new_n9304_), .A2(new_n9283_), .A3(new_n9288_), .ZN(new_n11597_));
  OAI21_X1   g10586(.A1(new_n9335_), .A2(new_n9337_), .B(new_n9303_), .ZN(new_n11598_));
  NAND3_X1   g10587(.A1(new_n11597_), .A2(new_n11598_), .A3(new_n9300_), .ZN(new_n11599_));
  NAND2_X1   g10588(.A1(new_n11596_), .A2(new_n11599_), .ZN(new_n11600_));
  NAND2_X1   g10589(.A1(new_n9338_), .A2(new_n9300_), .ZN(new_n11601_));
  NAND2_X1   g10590(.A1(new_n9344_), .A2(new_n9289_), .ZN(new_n11602_));
  AOI21_X1   g10591(.A1(new_n11601_), .A2(new_n11602_), .B(new_n9303_), .ZN(new_n11603_));
  NOR3_X1    g10592(.A1(new_n11600_), .A2(new_n11593_), .A3(new_n11603_), .ZN(new_n11604_));
  NAND2_X1   g10593(.A1(new_n9316_), .A2(new_n9358_), .ZN(new_n11605_));
  NAND2_X1   g10594(.A1(new_n9351_), .A2(new_n9330_), .ZN(new_n11606_));
  AOI21_X1   g10595(.A1(new_n11605_), .A2(new_n11606_), .B(new_n9357_), .ZN(new_n11607_));
  NOR2_X1    g10596(.A1(new_n9351_), .A2(new_n9330_), .ZN(new_n11608_));
  NOR2_X1    g10597(.A1(new_n9316_), .A2(new_n9358_), .ZN(new_n11609_));
  NOR3_X1    g10598(.A1(new_n11609_), .A2(new_n11608_), .A3(new_n9327_), .ZN(new_n11610_));
  NOR2_X1    g10599(.A1(new_n11607_), .A2(new_n11610_), .ZN(new_n11611_));
  OAI22_X1   g10600(.A1(new_n9311_), .A2(new_n9315_), .B1(new_n9326_), .B2(new_n9322_), .ZN(new_n11612_));
  NAND4_X1   g10601(.A1(new_n9348_), .A2(new_n9350_), .A3(new_n9354_), .A4(new_n9356_), .ZN(new_n11613_));
  NAND2_X1   g10602(.A1(new_n11612_), .A2(new_n11613_), .ZN(new_n11614_));
  NOR2_X1    g10603(.A1(new_n9329_), .A2(new_n9324_), .ZN(new_n11615_));
  OR4_X2     g10604(.A1(\A[295] ), .A2(new_n11615_), .A3(\A[296] ), .A4(\A[297] ), .Z(new_n11616_));
  NAND4_X1   g10605(.A1(new_n11614_), .A2(new_n9289_), .A3(new_n9300_), .A4(new_n9304_), .ZN(new_n11618_));
  INV_X1     g10606(.I(new_n11618_), .ZN(new_n11619_));
  NOR4_X1    g10607(.A1(new_n11604_), .A2(new_n9363_), .A3(new_n11611_), .A4(new_n11619_), .ZN(new_n11620_));
  NAND2_X1   g10608(.A1(new_n11592_), .A2(new_n11620_), .ZN(new_n11621_));
  INV_X1     g10609(.I(new_n11621_), .ZN(new_n11622_));
  NOR2_X1    g10610(.A1(new_n11592_), .A2(new_n11620_), .ZN(new_n11623_));
  OAI21_X1   g10611(.A1(new_n11622_), .A2(new_n11623_), .B(new_n11582_), .ZN(new_n11624_));
  NAND3_X1   g10612(.A1(new_n9417_), .A2(new_n9395_), .A3(new_n9400_), .ZN(new_n11625_));
  OAI21_X1   g10613(.A1(new_n9438_), .A2(new_n9440_), .B(new_n9448_), .ZN(new_n11626_));
  AOI21_X1   g10614(.A1(new_n11625_), .A2(new_n11626_), .B(new_n9412_), .ZN(new_n11627_));
  NOR3_X1    g10615(.A1(new_n9440_), .A2(new_n9448_), .A3(new_n9438_), .ZN(new_n11628_));
  AOI21_X1   g10616(.A1(new_n9395_), .A2(new_n9400_), .B(new_n9417_), .ZN(new_n11629_));
  NOR3_X1    g10617(.A1(new_n11629_), .A2(new_n9447_), .A3(new_n11628_), .ZN(new_n11630_));
  NOR2_X1    g10618(.A1(new_n11630_), .A2(new_n11627_), .ZN(new_n11631_));
  NOR2_X1    g10619(.A1(new_n9435_), .A2(new_n9418_), .ZN(new_n11632_));
  INV_X1     g10620(.I(new_n11632_), .ZN(new_n11633_));
  NOR3_X1    g10621(.A1(new_n9374_), .A2(new_n9389_), .A3(new_n9370_), .ZN(new_n11634_));
  INV_X1     g10622(.I(new_n9432_), .ZN(new_n11635_));
  INV_X1     g10623(.I(new_n9433_), .ZN(new_n11636_));
  AOI22_X1   g10624(.A1(new_n11635_), .A2(new_n11636_), .B1(new_n9422_), .B2(new_n9424_), .ZN(new_n11637_));
  OAI21_X1   g10625(.A1(new_n11637_), .A2(new_n11634_), .B(new_n9386_), .ZN(new_n11638_));
  NAND3_X1   g10626(.A1(new_n9434_), .A2(new_n9422_), .A3(new_n9424_), .ZN(new_n11639_));
  OAI21_X1   g10627(.A1(new_n9370_), .A2(new_n9374_), .B(new_n9389_), .ZN(new_n11640_));
  NAND3_X1   g10628(.A1(new_n11639_), .A2(new_n11640_), .A3(new_n9431_), .ZN(new_n11641_));
  NAND2_X1   g10629(.A1(new_n11638_), .A2(new_n11641_), .ZN(new_n11642_));
  NAND2_X1   g10630(.A1(new_n9375_), .A2(new_n9431_), .ZN(new_n11643_));
  NAND2_X1   g10631(.A1(new_n9386_), .A2(new_n9425_), .ZN(new_n11644_));
  AOI21_X1   g10632(.A1(new_n11643_), .A2(new_n11644_), .B(new_n9389_), .ZN(new_n11645_));
  NOR2_X1    g10633(.A1(new_n11642_), .A2(new_n11645_), .ZN(new_n11646_));
  NAND2_X1   g10634(.A1(new_n11646_), .A2(new_n11633_), .ZN(new_n11647_));
  NOR2_X1    g10635(.A1(new_n9386_), .A2(new_n9425_), .ZN(new_n11648_));
  NOR2_X1    g10636(.A1(new_n9375_), .A2(new_n9431_), .ZN(new_n11649_));
  OAI21_X1   g10637(.A1(new_n11648_), .A2(new_n11649_), .B(new_n9434_), .ZN(new_n11650_));
  NAND3_X1   g10638(.A1(new_n11650_), .A2(new_n11638_), .A3(new_n11641_), .ZN(new_n11651_));
  NAND2_X1   g10639(.A1(new_n11651_), .A2(new_n11632_), .ZN(new_n11652_));
  NAND2_X1   g10640(.A1(new_n11647_), .A2(new_n11652_), .ZN(new_n11653_));
  NAND2_X1   g10641(.A1(new_n11653_), .A2(new_n11631_), .ZN(new_n11654_));
  OAI21_X1   g10642(.A1(new_n11629_), .A2(new_n11628_), .B(new_n9447_), .ZN(new_n11655_));
  NAND3_X1   g10643(.A1(new_n11625_), .A2(new_n11626_), .A3(new_n9412_), .ZN(new_n11656_));
  NAND2_X1   g10644(.A1(new_n11655_), .A2(new_n11656_), .ZN(new_n11657_));
  AOI22_X1   g10645(.A1(new_n9395_), .A2(new_n9400_), .B1(new_n9406_), .B2(new_n9411_), .ZN(new_n11658_));
  NOR4_X1    g10646(.A1(new_n9438_), .A2(new_n9440_), .A3(new_n9446_), .A4(new_n9444_), .ZN(new_n11659_));
  NOR2_X1    g10647(.A1(new_n11658_), .A2(new_n11659_), .ZN(new_n11660_));
  NOR3_X1    g10648(.A1(new_n9441_), .A2(new_n9447_), .A3(new_n9448_), .ZN(new_n11661_));
  NOR3_X1    g10649(.A1(new_n11660_), .A2(new_n9435_), .A3(new_n11661_), .ZN(new_n11662_));
  NAND4_X1   g10650(.A1(new_n11662_), .A2(new_n11657_), .A3(new_n11642_), .A4(new_n11650_), .ZN(new_n11663_));
  AOI21_X1   g10651(.A1(new_n11663_), .A2(new_n11651_), .B(new_n11633_), .ZN(new_n11664_));
  NOR4_X1    g10652(.A1(new_n9419_), .A2(new_n9450_), .A3(new_n9504_), .A4(new_n9534_), .ZN(new_n11665_));
  NAND2_X1   g10653(.A1(new_n9476_), .A2(new_n9533_), .ZN(new_n11666_));
  NOR3_X1    g10654(.A1(new_n9460_), .A2(new_n9475_), .A3(new_n9456_), .ZN(new_n11667_));
  AOI21_X1   g10655(.A1(new_n9507_), .A2(new_n9509_), .B(new_n9519_), .ZN(new_n11668_));
  OAI21_X1   g10656(.A1(new_n11668_), .A2(new_n11667_), .B(new_n9472_), .ZN(new_n11669_));
  NAND3_X1   g10657(.A1(new_n9519_), .A2(new_n9507_), .A3(new_n9509_), .ZN(new_n11670_));
  OAI21_X1   g10658(.A1(new_n9456_), .A2(new_n9460_), .B(new_n9475_), .ZN(new_n11671_));
  NAND3_X1   g10659(.A1(new_n11670_), .A2(new_n11671_), .A3(new_n9516_), .ZN(new_n11672_));
  NOR2_X1    g10660(.A1(new_n9472_), .A2(new_n9510_), .ZN(new_n11673_));
  NOR2_X1    g10661(.A1(new_n9461_), .A2(new_n9516_), .ZN(new_n11674_));
  OAI21_X1   g10662(.A1(new_n11673_), .A2(new_n11674_), .B(new_n9519_), .ZN(new_n11675_));
  NAND4_X1   g10663(.A1(new_n11675_), .A2(new_n11666_), .A3(new_n11669_), .A4(new_n11672_), .ZN(new_n11676_));
  NOR2_X1    g10664(.A1(new_n9487_), .A2(new_n9501_), .ZN(new_n11677_));
  OAI21_X1   g10665(.A1(new_n9523_), .A2(new_n9525_), .B(new_n9501_), .ZN(new_n11678_));
  INV_X1     g10666(.I(new_n11678_), .ZN(new_n11679_));
  OAI21_X1   g10667(.A1(new_n11679_), .A2(new_n11677_), .B(new_n9532_), .ZN(new_n11680_));
  NAND2_X1   g10668(.A1(new_n9526_), .A2(new_n9502_), .ZN(new_n11681_));
  NAND3_X1   g10669(.A1(new_n11681_), .A2(new_n9498_), .A3(new_n11678_), .ZN(new_n11682_));
  NAND2_X1   g10670(.A1(new_n11680_), .A2(new_n11682_), .ZN(new_n11683_));
  OAI22_X1   g10671(.A1(new_n9523_), .A2(new_n9525_), .B1(new_n9531_), .B2(new_n9529_), .ZN(new_n11684_));
  NAND4_X1   g10672(.A1(new_n9481_), .A2(new_n9486_), .A3(new_n9492_), .A4(new_n9497_), .ZN(new_n11685_));
  NAND2_X1   g10673(.A1(new_n11684_), .A2(new_n11685_), .ZN(new_n11686_));
  NOR2_X1    g10674(.A1(new_n9500_), .A2(new_n9496_), .ZN(new_n11687_));
  OR4_X2     g10675(.A1(\A[271] ), .A2(new_n11687_), .A3(\A[272] ), .A4(\A[273] ), .Z(new_n11688_));
  NAND4_X1   g10676(.A1(new_n11686_), .A2(new_n9510_), .A3(new_n9516_), .A4(new_n9519_), .ZN(new_n11690_));
  NAND4_X1   g10677(.A1(new_n11665_), .A2(new_n11676_), .A3(new_n11683_), .A4(new_n11690_), .ZN(new_n11691_));
  NOR2_X1    g10678(.A1(new_n11664_), .A2(new_n11691_), .ZN(new_n11692_));
  OAI22_X1   g10679(.A1(new_n9438_), .A2(new_n9440_), .B1(new_n9446_), .B2(new_n9444_), .ZN(new_n11693_));
  NAND4_X1   g10680(.A1(new_n9395_), .A2(new_n9400_), .A3(new_n9406_), .A4(new_n9411_), .ZN(new_n11694_));
  AOI21_X1   g10681(.A1(new_n9395_), .A2(new_n9400_), .B(new_n9448_), .ZN(new_n11695_));
  AOI22_X1   g10682(.A1(new_n11693_), .A2(new_n11694_), .B1(new_n9412_), .B2(new_n11695_), .ZN(new_n11696_));
  NAND4_X1   g10683(.A1(new_n11696_), .A2(new_n9425_), .A3(new_n9431_), .A4(new_n9434_), .ZN(new_n11697_));
  NOR2_X1    g10684(.A1(new_n11697_), .A2(new_n11631_), .ZN(new_n11698_));
  OAI21_X1   g10685(.A1(new_n11698_), .A2(new_n11646_), .B(new_n11632_), .ZN(new_n11699_));
  NOR2_X1    g10686(.A1(new_n9520_), .A2(new_n9503_), .ZN(new_n11700_));
  AOI21_X1   g10687(.A1(new_n11670_), .A2(new_n11671_), .B(new_n9516_), .ZN(new_n11701_));
  NOR3_X1    g10688(.A1(new_n11668_), .A2(new_n9472_), .A3(new_n11667_), .ZN(new_n11702_));
  NAND2_X1   g10689(.A1(new_n9461_), .A2(new_n9516_), .ZN(new_n11703_));
  NAND2_X1   g10690(.A1(new_n9472_), .A2(new_n9510_), .ZN(new_n11704_));
  AOI21_X1   g10691(.A1(new_n11703_), .A2(new_n11704_), .B(new_n9475_), .ZN(new_n11705_));
  NOR4_X1    g10692(.A1(new_n11705_), .A2(new_n11700_), .A3(new_n11701_), .A4(new_n11702_), .ZN(new_n11706_));
  AOI21_X1   g10693(.A1(new_n11681_), .A2(new_n11678_), .B(new_n9498_), .ZN(new_n11707_));
  NOR3_X1    g10694(.A1(new_n11679_), .A2(new_n11677_), .A3(new_n9532_), .ZN(new_n11708_));
  NOR2_X1    g10695(.A1(new_n11708_), .A2(new_n11707_), .ZN(new_n11709_));
  INV_X1     g10696(.I(new_n11690_), .ZN(new_n11710_));
  NOR4_X1    g10697(.A1(new_n9540_), .A2(new_n11706_), .A3(new_n11710_), .A4(new_n11709_), .ZN(new_n11711_));
  NOR2_X1    g10698(.A1(new_n11699_), .A2(new_n11711_), .ZN(new_n11712_));
  OAI21_X1   g10699(.A1(new_n11692_), .A2(new_n11712_), .B(new_n11654_), .ZN(new_n11713_));
  AOI21_X1   g10700(.A1(new_n11647_), .A2(new_n11652_), .B(new_n11657_), .ZN(new_n11714_));
  NAND2_X1   g10701(.A1(new_n11699_), .A2(new_n11711_), .ZN(new_n11715_));
  NAND2_X1   g10702(.A1(new_n11664_), .A2(new_n11691_), .ZN(new_n11716_));
  NAND3_X1   g10703(.A1(new_n11715_), .A2(new_n11716_), .A3(new_n11714_), .ZN(new_n11717_));
  AOI21_X1   g10704(.A1(new_n11713_), .A2(new_n11717_), .B(new_n9544_), .ZN(new_n11718_));
  NAND2_X1   g10705(.A1(new_n11718_), .A2(new_n11624_), .ZN(new_n11719_));
  INV_X1     g10706(.I(new_n11582_), .ZN(new_n11720_));
  INV_X1     g10707(.I(new_n11623_), .ZN(new_n11721_));
  AOI21_X1   g10708(.A1(new_n11721_), .A2(new_n11621_), .B(new_n11720_), .ZN(new_n11722_));
  NAND2_X1   g10709(.A1(new_n11718_), .A2(new_n11722_), .ZN(new_n11723_));
  AOI21_X1   g10710(.A1(new_n11719_), .A2(new_n11723_), .B(new_n9548_), .ZN(new_n11724_));
  OAI21_X1   g10711(.A1(new_n11419_), .A2(new_n11555_), .B(new_n11724_), .ZN(new_n11725_));
  NOR2_X1    g10712(.A1(new_n11419_), .A2(new_n11555_), .ZN(new_n11726_));
  NAND2_X1   g10713(.A1(new_n11724_), .A2(new_n11726_), .ZN(new_n11727_));
  AOI21_X1   g10714(.A1(new_n11725_), .A2(new_n11727_), .B(new_n9550_), .ZN(new_n11728_));
  NOR2_X1    g10715(.A1(new_n11728_), .A2(new_n11319_), .ZN(new_n11729_));
  NAND2_X1   g10716(.A1(new_n9943_), .A2(new_n9957_), .ZN(new_n11730_));
  INV_X1     g10717(.I(new_n9957_), .ZN(new_n11731_));
  NAND2_X1   g10718(.A1(new_n11731_), .A2(new_n10037_), .ZN(new_n11732_));
  AOI21_X1   g10719(.A1(new_n11732_), .A2(new_n11730_), .B(new_n9954_), .ZN(new_n11733_));
  INV_X1     g10720(.I(new_n9954_), .ZN(new_n11734_));
  NOR2_X1    g10721(.A1(new_n11731_), .A2(new_n10037_), .ZN(new_n11735_));
  NOR2_X1    g10722(.A1(new_n9943_), .A2(new_n9957_), .ZN(new_n11736_));
  NOR3_X1    g10723(.A1(new_n11735_), .A2(new_n11736_), .A3(new_n11734_), .ZN(new_n11737_));
  OR2_X2     g10724(.A1(new_n11737_), .A2(new_n11733_), .Z(new_n11738_));
  NAND2_X1   g10725(.A1(new_n9979_), .A2(new_n9954_), .ZN(new_n11739_));
  NAND3_X1   g10726(.A1(new_n10020_), .A2(new_n9948_), .A3(new_n9953_), .ZN(new_n11740_));
  NAND2_X1   g10727(.A1(new_n9943_), .A2(new_n9968_), .ZN(new_n11741_));
  NAND2_X1   g10728(.A1(new_n9961_), .A2(\A[267] ), .ZN(new_n11742_));
  NAND2_X1   g10729(.A1(new_n9959_), .A2(\A[266] ), .ZN(new_n11743_));
  AOI21_X1   g10730(.A1(new_n11742_), .A2(new_n11743_), .B(new_n9964_), .ZN(new_n11744_));
  INV_X1     g10731(.I(new_n9965_), .ZN(new_n11745_));
  NAND2_X1   g10732(.A1(\A[266] ), .A2(\A[267] ), .ZN(new_n11746_));
  AOI21_X1   g10733(.A1(new_n11745_), .A2(new_n11746_), .B(\A[265] ), .ZN(new_n11747_));
  NOR2_X1    g10734(.A1(new_n11747_), .A2(new_n11744_), .ZN(new_n11748_));
  NAND2_X1   g10735(.A1(new_n11748_), .A2(new_n10037_), .ZN(new_n11749_));
  AOI22_X1   g10736(.A1(new_n11739_), .A2(new_n11740_), .B1(new_n11749_), .B2(new_n11741_), .ZN(new_n11750_));
  NAND3_X1   g10737(.A1(new_n10037_), .A2(new_n9954_), .A3(new_n9957_), .ZN(new_n11751_));
  NAND3_X1   g10738(.A1(new_n10020_), .A2(new_n9968_), .A3(new_n9984_), .ZN(new_n11752_));
  NAND2_X1   g10739(.A1(new_n11751_), .A2(new_n11752_), .ZN(new_n11753_));
  INV_X1     g10740(.I(new_n11753_), .ZN(new_n11754_));
  NAND2_X1   g10741(.A1(new_n11754_), .A2(new_n11750_), .ZN(new_n11755_));
  OAI22_X1   g10742(.A1(new_n9965_), .A2(new_n9980_), .B1(new_n9982_), .B2(new_n9976_), .ZN(new_n11756_));
  NOR3_X1    g10743(.A1(new_n11747_), .A2(new_n11756_), .A3(new_n11744_), .ZN(new_n11757_));
  INV_X1     g10744(.I(new_n9981_), .ZN(new_n11758_));
  INV_X1     g10745(.I(new_n9983_), .ZN(new_n11759_));
  AOI22_X1   g10746(.A1(new_n11758_), .A2(new_n11759_), .B1(new_n9963_), .B2(new_n9967_), .ZN(new_n11760_));
  OAI21_X1   g10747(.A1(new_n11760_), .A2(new_n11757_), .B(new_n9979_), .ZN(new_n11761_));
  NAND3_X1   g10748(.A1(new_n9984_), .A2(new_n9963_), .A3(new_n9967_), .ZN(new_n11762_));
  OAI21_X1   g10749(.A1(new_n11744_), .A2(new_n11747_), .B(new_n11756_), .ZN(new_n11763_));
  NAND3_X1   g10750(.A1(new_n11762_), .A2(new_n11763_), .A3(new_n10020_), .ZN(new_n11764_));
  NAND2_X1   g10751(.A1(new_n11761_), .A2(new_n11764_), .ZN(new_n11765_));
  XOR2_X1    g10752(.A1(new_n11755_), .A2(new_n11765_), .Z(new_n11766_));
  NOR2_X1    g10753(.A1(new_n11766_), .A2(new_n11738_), .ZN(new_n11767_));
  INV_X1     g10754(.I(new_n11755_), .ZN(new_n11768_));
  NOR2_X1    g10755(.A1(new_n11737_), .A2(new_n11733_), .ZN(new_n11769_));
  NAND2_X1   g10756(.A1(new_n9981_), .A2(new_n9983_), .ZN(new_n11770_));
  NAND3_X1   g10757(.A1(new_n10020_), .A2(new_n9968_), .A3(new_n11770_), .ZN(new_n11771_));
  NOR2_X1    g10758(.A1(new_n11751_), .A2(new_n11771_), .ZN(new_n11772_));
  NAND3_X1   g10759(.A1(new_n11750_), .A2(new_n11765_), .A3(new_n11772_), .ZN(new_n11773_));
  NOR2_X1    g10760(.A1(new_n11773_), .A2(new_n11769_), .ZN(new_n11774_));
  OAI21_X1   g10761(.A1(new_n11774_), .A2(new_n11765_), .B(new_n11768_), .ZN(new_n11775_));
  XOR2_X1    g10762(.A1(new_n9931_), .A2(new_n10038_), .Z(new_n11776_));
  NAND3_X1   g10763(.A1(new_n10012_), .A2(new_n9990_), .A3(new_n9995_), .ZN(new_n11777_));
  OAI22_X1   g10764(.A1(new_n9992_), .A2(new_n10008_), .B1(new_n10010_), .B2(new_n10005_), .ZN(new_n11778_));
  OAI21_X1   g10765(.A1(new_n10024_), .A2(new_n10026_), .B(new_n11778_), .ZN(new_n11779_));
  AOI21_X1   g10766(.A1(new_n11777_), .A2(new_n11779_), .B(new_n10007_), .ZN(new_n11780_));
  NAND2_X1   g10767(.A1(new_n9999_), .A2(\A[258] ), .ZN(new_n11781_));
  NAND2_X1   g10768(.A1(new_n9997_), .A2(\A[257] ), .ZN(new_n11782_));
  AOI21_X1   g10769(.A1(new_n11781_), .A2(new_n11782_), .B(new_n10002_), .ZN(new_n11783_));
  INV_X1     g10770(.I(new_n10005_), .ZN(new_n11784_));
  AOI21_X1   g10771(.A1(new_n11784_), .A2(new_n10003_), .B(\A[256] ), .ZN(new_n11785_));
  NOR2_X1    g10772(.A1(new_n11785_), .A2(new_n11783_), .ZN(new_n11786_));
  NOR3_X1    g10773(.A1(new_n10026_), .A2(new_n11778_), .A3(new_n10024_), .ZN(new_n11787_));
  INV_X1     g10774(.I(new_n10009_), .ZN(new_n11788_));
  INV_X1     g10775(.I(new_n10011_), .ZN(new_n11789_));
  AOI22_X1   g10776(.A1(new_n11788_), .A2(new_n11789_), .B1(new_n9990_), .B2(new_n9995_), .ZN(new_n11790_));
  NOR3_X1    g10777(.A1(new_n11790_), .A2(new_n11786_), .A3(new_n11787_), .ZN(new_n11791_));
  NOR2_X1    g10778(.A1(new_n11791_), .A2(new_n11780_), .ZN(new_n11792_));
  NAND2_X1   g10779(.A1(new_n11786_), .A2(new_n9927_), .ZN(new_n11793_));
  AND2_X2    g10780(.A1(new_n9921_), .A2(new_n9926_), .Z(new_n11794_));
  NAND2_X1   g10781(.A1(new_n11794_), .A2(new_n10007_), .ZN(new_n11795_));
  NAND2_X1   g10782(.A1(new_n9916_), .A2(new_n9996_), .ZN(new_n11796_));
  NOR2_X1    g10783(.A1(new_n9909_), .A2(\A[248] ), .ZN(new_n11797_));
  NOR2_X1    g10784(.A1(new_n9907_), .A2(\A[249] ), .ZN(new_n11798_));
  OAI21_X1   g10785(.A1(new_n11797_), .A2(new_n11798_), .B(\A[247] ), .ZN(new_n11799_));
  INV_X1     g10786(.I(new_n9914_), .ZN(new_n11800_));
  OAI21_X1   g10787(.A1(new_n11800_), .A2(new_n9912_), .B(new_n9906_), .ZN(new_n11801_));
  NAND2_X1   g10788(.A1(new_n11799_), .A2(new_n11801_), .ZN(new_n11802_));
  NAND2_X1   g10789(.A1(new_n10027_), .A2(new_n11802_), .ZN(new_n11803_));
  AOI22_X1   g10790(.A1(new_n11795_), .A2(new_n11793_), .B1(new_n11796_), .B2(new_n11803_), .ZN(new_n11804_));
  NOR4_X1    g10791(.A1(new_n9928_), .A2(\A[250] ), .A3(\A[251] ), .A4(\A[252] ), .ZN(new_n11805_));
  NOR2_X1    g10792(.A1(new_n11786_), .A2(new_n11778_), .ZN(new_n11806_));
  AOI22_X1   g10793(.A1(new_n11806_), .A2(new_n9996_), .B1(new_n11802_), .B2(new_n11805_), .ZN(new_n11807_));
  NAND2_X1   g10794(.A1(new_n11804_), .A2(new_n11807_), .ZN(new_n11808_));
  INV_X1     g10795(.I(new_n9930_), .ZN(new_n11809_));
  NOR2_X1    g10796(.A1(new_n11809_), .A2(new_n11802_), .ZN(new_n11810_));
  NOR2_X1    g10797(.A1(new_n9916_), .A2(new_n9930_), .ZN(new_n11811_));
  OAI21_X1   g10798(.A1(new_n11810_), .A2(new_n11811_), .B(new_n11794_), .ZN(new_n11812_));
  NAND2_X1   g10799(.A1(new_n9916_), .A2(new_n9930_), .ZN(new_n11813_));
  NAND2_X1   g10800(.A1(new_n11809_), .A2(new_n11802_), .ZN(new_n11814_));
  NAND3_X1   g10801(.A1(new_n11814_), .A2(new_n11813_), .A3(new_n9927_), .ZN(new_n11815_));
  NAND2_X1   g10802(.A1(new_n11812_), .A2(new_n11815_), .ZN(new_n11816_));
  NOR2_X1    g10803(.A1(new_n11794_), .A2(new_n10007_), .ZN(new_n11817_));
  NOR2_X1    g10804(.A1(new_n11786_), .A2(new_n9927_), .ZN(new_n11818_));
  NOR2_X1    g10805(.A1(new_n10027_), .A2(new_n11802_), .ZN(new_n11819_));
  NOR2_X1    g10806(.A1(new_n9916_), .A2(new_n9996_), .ZN(new_n11820_));
  OAI22_X1   g10807(.A1(new_n11817_), .A2(new_n11818_), .B1(new_n11819_), .B2(new_n11820_), .ZN(new_n11821_));
  NAND2_X1   g10808(.A1(new_n11802_), .A2(new_n11805_), .ZN(new_n11822_));
  NAND2_X1   g10809(.A1(new_n10009_), .A2(new_n10011_), .ZN(new_n11823_));
  NAND3_X1   g10810(.A1(new_n9996_), .A2(new_n10007_), .A3(new_n11823_), .ZN(new_n11824_));
  OR2_X2     g10811(.A1(new_n11824_), .A2(new_n11822_), .Z(new_n11825_));
  NAND3_X1   g10812(.A1(new_n11808_), .A2(new_n11792_), .A3(new_n11816_), .ZN(new_n11827_));
  NOR3_X1    g10813(.A1(new_n11776_), .A2(new_n11827_), .A3(new_n10041_), .ZN(new_n11828_));
  NAND2_X1   g10814(.A1(new_n11828_), .A2(new_n11775_), .ZN(new_n11829_));
  OR2_X2     g10815(.A1(new_n11828_), .A2(new_n11775_), .Z(new_n11830_));
  NAND2_X1   g10816(.A1(new_n11830_), .A2(new_n11829_), .ZN(new_n11831_));
  NAND2_X1   g10817(.A1(new_n11831_), .A2(new_n11767_), .ZN(new_n11832_));
  NAND4_X1   g10818(.A1(new_n10223_), .A2(new_n10221_), .A3(new_n10222_), .A4(new_n10218_), .ZN(new_n11833_));
  NAND2_X1   g10819(.A1(new_n10115_), .A2(new_n10125_), .ZN(new_n11834_));
  OR2_X2     g10820(.A1(new_n10123_), .A2(new_n10124_), .Z(new_n11835_));
  NAND2_X1   g10821(.A1(new_n11835_), .A2(new_n10097_), .ZN(new_n11836_));
  AOI21_X1   g10822(.A1(new_n11836_), .A2(new_n11834_), .B(new_n10108_), .ZN(new_n11837_));
  NAND3_X1   g10823(.A1(new_n11836_), .A2(new_n11834_), .A3(new_n10108_), .ZN(new_n11838_));
  INV_X1     g10824(.I(new_n11838_), .ZN(new_n11839_));
  NOR2_X1    g10825(.A1(new_n11839_), .A2(new_n11837_), .ZN(new_n11840_));
  NAND2_X1   g10826(.A1(new_n10141_), .A2(\A[246] ), .ZN(new_n11841_));
  NAND2_X1   g10827(.A1(new_n10139_), .A2(\A[245] ), .ZN(new_n11842_));
  AOI21_X1   g10828(.A1(new_n11841_), .A2(new_n11842_), .B(new_n10144_), .ZN(new_n11843_));
  INV_X1     g10829(.I(new_n10147_), .ZN(new_n11844_));
  AOI21_X1   g10830(.A1(new_n11844_), .A2(new_n10145_), .B(\A[244] ), .ZN(new_n11845_));
  NOR2_X1    g10831(.A1(new_n11845_), .A2(new_n11843_), .ZN(new_n11846_));
  NAND3_X1   g10832(.A1(new_n10097_), .A2(new_n10108_), .A3(new_n10125_), .ZN(new_n11847_));
  NOR4_X1    g10833(.A1(new_n11847_), .A2(new_n10200_), .A3(new_n11846_), .A4(new_n10152_), .ZN(new_n11848_));
  NAND2_X1   g10834(.A1(new_n10200_), .A2(new_n10153_), .ZN(new_n11849_));
  OAI21_X1   g10835(.A1(new_n10197_), .A2(new_n10199_), .B(new_n10152_), .ZN(new_n11850_));
  AOI21_X1   g10836(.A1(new_n11849_), .A2(new_n11850_), .B(new_n10149_), .ZN(new_n11851_));
  NOR2_X1    g10837(.A1(new_n10138_), .A2(new_n10152_), .ZN(new_n11852_));
  INV_X1     g10838(.I(new_n11850_), .ZN(new_n11853_));
  NOR3_X1    g10839(.A1(new_n11853_), .A2(new_n11852_), .A3(new_n11846_), .ZN(new_n11854_));
  NOR2_X1    g10840(.A1(new_n11854_), .A2(new_n11851_), .ZN(new_n11855_));
  NOR2_X1    g10841(.A1(new_n11855_), .A2(new_n11848_), .ZN(new_n11856_));
  NOR3_X1    g10842(.A1(new_n11835_), .A2(new_n10115_), .A3(new_n10121_), .ZN(new_n11857_));
  NAND4_X1   g10843(.A1(new_n11857_), .A2(new_n10138_), .A3(new_n10149_), .A4(new_n10153_), .ZN(new_n11858_));
  OAI21_X1   g10844(.A1(new_n11853_), .A2(new_n11852_), .B(new_n11846_), .ZN(new_n11859_));
  NAND3_X1   g10845(.A1(new_n11849_), .A2(new_n10149_), .A3(new_n11850_), .ZN(new_n11860_));
  NAND2_X1   g10846(.A1(new_n11859_), .A2(new_n11860_), .ZN(new_n11861_));
  NOR2_X1    g10847(.A1(new_n11861_), .A2(new_n11858_), .ZN(new_n11862_));
  OAI21_X1   g10848(.A1(new_n11856_), .A2(new_n11862_), .B(new_n11840_), .ZN(new_n11863_));
  NOR2_X1    g10849(.A1(new_n10115_), .A2(new_n10121_), .ZN(new_n11864_));
  NOR2_X1    g10850(.A1(new_n10097_), .A2(new_n10108_), .ZN(new_n11865_));
  OR4_X2     g10851(.A1(new_n10134_), .A2(new_n10150_), .A3(new_n10151_), .A4(new_n10147_), .Z(new_n11866_));
  NAND3_X1   g10852(.A1(new_n10138_), .A2(new_n10149_), .A3(new_n11866_), .ZN(new_n11867_));
  NOR3_X1    g10853(.A1(new_n11864_), .A2(new_n11867_), .A3(new_n11865_), .ZN(new_n11868_));
  NOR2_X1    g10854(.A1(new_n10200_), .A2(new_n11846_), .ZN(new_n11869_));
  NOR2_X1    g10855(.A1(new_n10138_), .A2(new_n10149_), .ZN(new_n11870_));
  NOR3_X1    g10856(.A1(new_n10126_), .A2(new_n11869_), .A3(new_n11870_), .ZN(new_n11871_));
  NAND3_X1   g10857(.A1(new_n11861_), .A2(new_n11868_), .A3(new_n11871_), .ZN(new_n11872_));
  NOR4_X1    g10858(.A1(new_n11847_), .A2(new_n10200_), .A3(new_n11846_), .A4(new_n10152_), .ZN(new_n11874_));
  AOI22_X1   g10859(.A1(new_n10070_), .A2(new_n10072_), .B1(new_n10075_), .B2(new_n10077_), .ZN(new_n11875_));
  NOR4_X1    g10860(.A1(new_n10052_), .A2(new_n10056_), .A3(new_n10066_), .A4(new_n10062_), .ZN(new_n11876_));
  NOR2_X1    g10861(.A1(new_n11875_), .A2(new_n11876_), .ZN(new_n11877_));
  NAND2_X1   g10862(.A1(new_n10075_), .A2(new_n10077_), .ZN(new_n11878_));
  NOR2_X1    g10863(.A1(new_n10083_), .A2(new_n10064_), .ZN(new_n11879_));
  NOR4_X1    g10864(.A1(new_n11879_), .A2(\A[223] ), .A3(\A[224] ), .A4(\A[225] ), .ZN(new_n11880_));
  NAND4_X1   g10865(.A1(new_n11878_), .A2(new_n10188_), .A3(new_n11880_), .A4(new_n10191_), .ZN(new_n11881_));
  NOR3_X1    g10866(.A1(new_n11877_), .A2(new_n10187_), .A3(new_n11881_), .ZN(new_n11882_));
  NOR3_X1    g10867(.A1(new_n10208_), .A2(new_n10176_), .A3(new_n10179_), .ZN(new_n11883_));
  NOR2_X1    g10868(.A1(new_n10207_), .A2(new_n10162_), .ZN(new_n11884_));
  INV_X1     g10869(.I(new_n11884_), .ZN(new_n11885_));
  INV_X1     g10870(.I(new_n10190_), .ZN(new_n11886_));
  AOI22_X1   g10871(.A1(new_n11885_), .A2(new_n11886_), .B1(new_n10159_), .B2(new_n10163_), .ZN(new_n11887_));
  OAI21_X1   g10872(.A1(new_n11887_), .A2(new_n11883_), .B(new_n10206_), .ZN(new_n11888_));
  NAND4_X1   g10873(.A1(new_n11885_), .A2(new_n11886_), .A3(new_n10159_), .A4(new_n10163_), .ZN(new_n11889_));
  OAI21_X1   g10874(.A1(new_n10176_), .A2(new_n10179_), .B(new_n10208_), .ZN(new_n11890_));
  NAND3_X1   g10875(.A1(new_n11889_), .A2(new_n11890_), .A3(new_n10188_), .ZN(new_n11891_));
  NAND2_X1   g10876(.A1(new_n11884_), .A2(new_n10190_), .ZN(new_n11892_));
  INV_X1     g10877(.I(new_n11892_), .ZN(new_n11893_));
  NAND3_X1   g10878(.A1(new_n10202_), .A2(new_n10203_), .A3(new_n10208_), .ZN(new_n11894_));
  NAND3_X1   g10879(.A1(new_n11888_), .A2(new_n11894_), .A3(new_n11891_), .ZN(new_n11895_));
  NOR3_X1    g10880(.A1(new_n10056_), .A2(new_n10084_), .A3(new_n10052_), .ZN(new_n11896_));
  NOR2_X1    g10881(.A1(new_n10082_), .A2(new_n10054_), .ZN(new_n11897_));
  NOR2_X1    g10882(.A1(new_n11897_), .A2(new_n11879_), .ZN(new_n11898_));
  AOI21_X1   g10883(.A1(new_n10070_), .A2(new_n10072_), .B(new_n11898_), .ZN(new_n11899_));
  OAI21_X1   g10884(.A1(new_n11899_), .A2(new_n11896_), .B(new_n10081_), .ZN(new_n11900_));
  NAND3_X1   g10885(.A1(new_n11898_), .A2(new_n10070_), .A3(new_n10072_), .ZN(new_n11901_));
  OAI21_X1   g10886(.A1(new_n10052_), .A2(new_n10056_), .B(new_n10084_), .ZN(new_n11902_));
  NAND3_X1   g10887(.A1(new_n11901_), .A2(new_n11902_), .A3(new_n11878_), .ZN(new_n11903_));
  NAND2_X1   g10888(.A1(new_n11900_), .A2(new_n11903_), .ZN(new_n11904_));
  NOR3_X1    g10889(.A1(new_n11895_), .A2(new_n11882_), .A3(new_n11904_), .ZN(new_n11905_));
  NAND4_X1   g10890(.A1(new_n10079_), .A2(new_n10204_), .A3(new_n10085_), .A4(new_n10209_), .ZN(new_n11906_));
  AOI21_X1   g10891(.A1(new_n11889_), .A2(new_n11890_), .B(new_n10188_), .ZN(new_n11907_));
  NOR3_X1    g10892(.A1(new_n11887_), .A2(new_n10206_), .A3(new_n11883_), .ZN(new_n11908_));
  INV_X1     g10893(.I(new_n10208_), .ZN(new_n11909_));
  NOR3_X1    g10894(.A1(new_n10173_), .A2(new_n10186_), .A3(new_n11909_), .ZN(new_n11910_));
  NOR3_X1    g10895(.A1(new_n11910_), .A2(new_n11908_), .A3(new_n11907_), .ZN(new_n11911_));
  AOI21_X1   g10896(.A1(new_n11901_), .A2(new_n11902_), .B(new_n11878_), .ZN(new_n11912_));
  NOR3_X1    g10897(.A1(new_n11899_), .A2(new_n10081_), .A3(new_n11896_), .ZN(new_n11913_));
  NOR2_X1    g10898(.A1(new_n11913_), .A2(new_n11912_), .ZN(new_n11914_));
  AOI21_X1   g10899(.A1(new_n11911_), .A2(new_n11906_), .B(new_n11914_), .ZN(new_n11915_));
  NOR2_X1    g10900(.A1(new_n11915_), .A2(new_n11905_), .ZN(new_n11916_));
  NAND2_X1   g10901(.A1(new_n11888_), .A2(new_n11891_), .ZN(new_n11917_));
  AOI21_X1   g10902(.A1(new_n10173_), .A2(new_n11892_), .B(new_n11909_), .ZN(new_n11918_));
  NOR3_X1    g10903(.A1(new_n11877_), .A2(new_n11918_), .A3(new_n10187_), .ZN(new_n11919_));
  AOI21_X1   g10904(.A1(new_n11919_), .A2(new_n11917_), .B(new_n10085_), .ZN(new_n11920_));
  OAI21_X1   g10905(.A1(new_n10202_), .A2(new_n11893_), .B(new_n10208_), .ZN(new_n11921_));
  NAND2_X1   g10906(.A1(new_n11921_), .A2(new_n10204_), .ZN(new_n11922_));
  NOR2_X1    g10907(.A1(new_n11911_), .A2(new_n11882_), .ZN(new_n11923_));
  OAI21_X1   g10908(.A1(new_n11920_), .A2(new_n11922_), .B(new_n11923_), .ZN(new_n11924_));
  NOR2_X1    g10909(.A1(new_n10086_), .A2(new_n10127_), .ZN(new_n11925_));
  NAND2_X1   g10910(.A1(new_n11878_), .A2(new_n11880_), .ZN(new_n11926_));
  NAND3_X1   g10911(.A1(new_n11926_), .A2(new_n10067_), .A3(new_n10078_), .ZN(new_n11927_));
  NOR2_X1    g10912(.A1(new_n10213_), .A2(new_n11927_), .ZN(new_n11928_));
  OAI22_X1   g10913(.A1(new_n10194_), .A2(new_n10211_), .B1(new_n11925_), .B2(new_n11928_), .ZN(new_n11929_));
  NOR4_X1    g10914(.A1(new_n11924_), .A2(new_n11916_), .A3(new_n11929_), .A4(new_n11874_), .ZN(new_n11930_));
  INV_X1     g10915(.I(new_n11874_), .ZN(new_n11931_));
  AOI22_X1   g10916(.A1(new_n10067_), .A2(new_n10078_), .B1(new_n10202_), .B2(new_n10203_), .ZN(new_n11932_));
  NAND3_X1   g10917(.A1(new_n11917_), .A2(new_n11932_), .A3(new_n11921_), .ZN(new_n11933_));
  AOI21_X1   g10918(.A1(new_n11933_), .A2(new_n11926_), .B(new_n11922_), .ZN(new_n11934_));
  NOR4_X1    g10919(.A1(new_n11934_), .A2(new_n11882_), .A3(new_n11911_), .A4(new_n11914_), .ZN(new_n11935_));
  NAND2_X1   g10920(.A1(new_n10213_), .A2(new_n11927_), .ZN(new_n11936_));
  NAND2_X1   g10921(.A1(new_n10086_), .A2(new_n10127_), .ZN(new_n11937_));
  AOI22_X1   g10922(.A1(new_n10214_), .A2(new_n10215_), .B1(new_n11937_), .B2(new_n11936_), .ZN(new_n11938_));
  AOI21_X1   g10923(.A1(new_n11935_), .A2(new_n11938_), .B(new_n11931_), .ZN(new_n11939_));
  OAI21_X1   g10924(.A1(new_n11939_), .A2(new_n11930_), .B(new_n11863_), .ZN(new_n11940_));
  NAND2_X1   g10925(.A1(new_n11836_), .A2(new_n11834_), .ZN(new_n11941_));
  NAND2_X1   g10926(.A1(new_n11941_), .A2(new_n10121_), .ZN(new_n11942_));
  NAND2_X1   g10927(.A1(new_n11942_), .A2(new_n11838_), .ZN(new_n11943_));
  NAND2_X1   g10928(.A1(new_n11861_), .A2(new_n11858_), .ZN(new_n11944_));
  NAND2_X1   g10929(.A1(new_n11855_), .A2(new_n11848_), .ZN(new_n11945_));
  AOI21_X1   g10930(.A1(new_n11945_), .A2(new_n11944_), .B(new_n11943_), .ZN(new_n11946_));
  NAND3_X1   g10931(.A1(new_n11935_), .A2(new_n11931_), .A3(new_n11938_), .ZN(new_n11947_));
  NAND3_X1   g10932(.A1(new_n11911_), .A2(new_n11906_), .A3(new_n11914_), .ZN(new_n11948_));
  OAI21_X1   g10933(.A1(new_n11895_), .A2(new_n11882_), .B(new_n11904_), .ZN(new_n11949_));
  NAND2_X1   g10934(.A1(new_n11948_), .A2(new_n11949_), .ZN(new_n11950_));
  NOR2_X1    g10935(.A1(new_n11908_), .A2(new_n11907_), .ZN(new_n11951_));
  NAND3_X1   g10936(.A1(new_n10079_), .A2(new_n11921_), .A3(new_n10204_), .ZN(new_n11952_));
  OAI21_X1   g10937(.A1(new_n11952_), .A2(new_n11951_), .B(new_n11926_), .ZN(new_n11953_));
  INV_X1     g10938(.I(new_n11922_), .ZN(new_n11954_));
  NAND2_X1   g10939(.A1(new_n11906_), .A2(new_n11895_), .ZN(new_n11955_));
  AOI21_X1   g10940(.A1(new_n11953_), .A2(new_n11954_), .B(new_n11955_), .ZN(new_n11956_));
  NAND3_X1   g10941(.A1(new_n11956_), .A2(new_n11950_), .A3(new_n11938_), .ZN(new_n11957_));
  NAND2_X1   g10942(.A1(new_n11957_), .A2(new_n11874_), .ZN(new_n11958_));
  NAND3_X1   g10943(.A1(new_n11958_), .A2(new_n11947_), .A3(new_n11946_), .ZN(new_n11959_));
  AOI21_X1   g10944(.A1(new_n11959_), .A2(new_n11940_), .B(new_n11833_), .ZN(new_n11960_));
  NOR2_X1    g10945(.A1(new_n11960_), .A2(new_n11832_), .ZN(new_n11961_));
  NOR3_X1    g10946(.A1(new_n9632_), .A2(new_n9647_), .A3(new_n9628_), .ZN(new_n11962_));
  OAI21_X1   g10947(.A1(\A[211] ), .A2(new_n9653_), .B(new_n9630_), .ZN(new_n11963_));
  OAI21_X1   g10948(.A1(\A[214] ), .A2(new_n9658_), .B(new_n9642_), .ZN(new_n11964_));
  AOI22_X1   g10949(.A1(new_n11964_), .A2(new_n11963_), .B1(new_n9652_), .B2(new_n9654_), .ZN(new_n11965_));
  OAI21_X1   g10950(.A1(new_n11965_), .A2(new_n11962_), .B(new_n9644_), .ZN(new_n11966_));
  NAND4_X1   g10951(.A1(new_n11964_), .A2(new_n11963_), .A3(new_n9652_), .A4(new_n9654_), .ZN(new_n11967_));
  OAI21_X1   g10952(.A1(new_n9628_), .A2(new_n9632_), .B(new_n9647_), .ZN(new_n11968_));
  NAND3_X1   g10953(.A1(new_n11967_), .A2(new_n11968_), .A3(new_n9722_), .ZN(new_n11969_));
  NAND2_X1   g10954(.A1(new_n11966_), .A2(new_n11969_), .ZN(new_n11970_));
  NAND4_X1   g10955(.A1(new_n9693_), .A2(new_n9698_), .A3(new_n9695_), .A4(new_n9700_), .ZN(new_n11971_));
  NOR2_X1    g10956(.A1(new_n11971_), .A2(new_n9688_), .ZN(new_n11972_));
  OAI22_X1   g10957(.A1(new_n9668_), .A2(new_n9672_), .B1(new_n9682_), .B2(new_n9678_), .ZN(new_n11973_));
  NAND2_X1   g10958(.A1(new_n11973_), .A2(new_n11971_), .ZN(new_n11974_));
  NOR4_X1    g10959(.A1(new_n9661_), .A2(new_n11974_), .A3(new_n11972_), .A4(new_n9648_), .ZN(new_n11975_));
  NAND2_X1   g10960(.A1(new_n9698_), .A2(new_n9700_), .ZN(new_n11976_));
  NOR2_X1    g10961(.A1(new_n9685_), .A2(new_n9687_), .ZN(new_n11977_));
  NAND3_X1   g10962(.A1(new_n11977_), .A2(new_n9693_), .A3(new_n9695_), .ZN(new_n11978_));
  OAI22_X1   g10963(.A1(new_n9669_), .A2(new_n9686_), .B1(new_n9684_), .B2(new_n9679_), .ZN(new_n11979_));
  OAI21_X1   g10964(.A1(new_n9668_), .A2(new_n9672_), .B(new_n11979_), .ZN(new_n11980_));
  AOI21_X1   g10965(.A1(new_n11978_), .A2(new_n11980_), .B(new_n11976_), .ZN(new_n11981_));
  INV_X1     g10966(.I(new_n11976_), .ZN(new_n11982_));
  NOR3_X1    g10967(.A1(new_n9672_), .A2(new_n11979_), .A3(new_n9668_), .ZN(new_n11983_));
  INV_X1     g10968(.I(new_n9685_), .ZN(new_n11984_));
  INV_X1     g10969(.I(new_n9687_), .ZN(new_n11985_));
  AOI22_X1   g10970(.A1(new_n11984_), .A2(new_n11985_), .B1(new_n9693_), .B2(new_n9695_), .ZN(new_n11986_));
  NOR3_X1    g10971(.A1(new_n11986_), .A2(new_n11982_), .A3(new_n11983_), .ZN(new_n11987_));
  NOR2_X1    g10972(.A1(new_n11987_), .A2(new_n11981_), .ZN(new_n11988_));
  XOR2_X1    g10973(.A1(new_n11975_), .A2(new_n11988_), .Z(new_n11989_));
  NOR2_X1    g10974(.A1(new_n11989_), .A2(new_n11970_), .ZN(new_n11990_));
  INV_X1     g10975(.I(new_n11990_), .ZN(new_n11991_));
  AOI22_X1   g10976(.A1(new_n9657_), .A2(new_n9659_), .B1(new_n9652_), .B2(new_n9654_), .ZN(new_n11992_));
  NOR4_X1    g10977(.A1(new_n9628_), .A2(new_n9632_), .A3(new_n9643_), .A4(new_n9639_), .ZN(new_n11993_));
  NOR2_X1    g10978(.A1(new_n11992_), .A2(new_n11993_), .ZN(new_n11994_));
  NAND4_X1   g10979(.A1(new_n11994_), .A2(new_n9702_), .A3(new_n9690_), .A4(new_n9724_), .ZN(new_n11995_));
  NOR2_X1    g10980(.A1(new_n9661_), .A2(new_n11974_), .ZN(new_n11996_));
  XNOR2_X1   g10981(.A1(new_n9685_), .A2(new_n9687_), .ZN(new_n11997_));
  NAND2_X1   g10982(.A1(new_n9688_), .A2(new_n11979_), .ZN(new_n11998_));
  NAND2_X1   g10983(.A1(new_n11971_), .A2(new_n11998_), .ZN(new_n11999_));
  OAI21_X1   g10984(.A1(new_n11971_), .A2(new_n11997_), .B(new_n11999_), .ZN(new_n12000_));
  NAND2_X1   g10985(.A1(new_n9701_), .A2(new_n9688_), .ZN(new_n12001_));
  NOR2_X1    g10986(.A1(new_n12001_), .A2(new_n9724_), .ZN(new_n12002_));
  NAND4_X1   g10987(.A1(new_n12000_), .A2(new_n11970_), .A3(new_n11996_), .A4(new_n12002_), .ZN(new_n12003_));
  AOI21_X1   g10988(.A1(new_n12003_), .A2(new_n11988_), .B(new_n11995_), .ZN(new_n12004_));
  INV_X1     g10989(.I(new_n12004_), .ZN(new_n12005_));
  NAND4_X1   g10990(.A1(new_n9590_), .A2(new_n9577_), .A3(new_n9718_), .A4(new_n9719_), .ZN(new_n12006_));
  NOR2_X1    g10991(.A1(new_n9616_), .A2(new_n9619_), .ZN(new_n12007_));
  NAND3_X1   g10992(.A1(new_n12007_), .A2(new_n9714_), .A3(new_n9716_), .ZN(new_n12008_));
  OAI22_X1   g10993(.A1(new_n9598_), .A2(new_n9615_), .B1(new_n9618_), .B2(new_n9617_), .ZN(new_n12009_));
  OAI21_X1   g10994(.A1(new_n9608_), .A2(new_n9611_), .B(new_n12009_), .ZN(new_n12010_));
  AOI21_X1   g10995(.A1(new_n12008_), .A2(new_n12010_), .B(new_n9711_), .ZN(new_n12011_));
  NOR3_X1    g10996(.A1(new_n12009_), .A2(new_n9608_), .A3(new_n9611_), .ZN(new_n12012_));
  INV_X1     g10997(.I(new_n9616_), .ZN(new_n12013_));
  INV_X1     g10998(.I(new_n9619_), .ZN(new_n12014_));
  AOI22_X1   g10999(.A1(new_n12013_), .A2(new_n12014_), .B1(new_n9714_), .B2(new_n9716_), .ZN(new_n12015_));
  NOR3_X1    g11000(.A1(new_n12015_), .A2(new_n9602_), .A3(new_n12012_), .ZN(new_n12016_));
  NOR2_X1    g11001(.A1(new_n12016_), .A2(new_n12011_), .ZN(new_n12017_));
  NOR3_X1    g11002(.A1(new_n9584_), .A2(new_n9732_), .A3(new_n9581_), .ZN(new_n12018_));
  AOI22_X1   g11003(.A1(new_n9576_), .A2(new_n9574_), .B1(new_n9556_), .B2(new_n9560_), .ZN(new_n12019_));
  OAI21_X1   g11004(.A1(new_n12019_), .A2(new_n12018_), .B(new_n9730_), .ZN(new_n12020_));
  NAND4_X1   g11005(.A1(new_n9574_), .A2(new_n9576_), .A3(new_n9556_), .A4(new_n9560_), .ZN(new_n12021_));
  OAI21_X1   g11006(.A1(new_n9581_), .A2(new_n9584_), .B(new_n9732_), .ZN(new_n12022_));
  NAND3_X1   g11007(.A1(new_n12021_), .A2(new_n12022_), .A3(new_n9572_), .ZN(new_n12023_));
  NAND2_X1   g11008(.A1(new_n12020_), .A2(new_n12023_), .ZN(new_n12024_));
  NOR3_X1    g11009(.A1(new_n9736_), .A2(new_n9613_), .A3(new_n9614_), .ZN(new_n12025_));
  XOR2_X1    g11010(.A1(new_n9616_), .A2(new_n9619_), .Z(new_n12026_));
  NAND2_X1   g11011(.A1(new_n12026_), .A2(new_n9614_), .ZN(new_n12027_));
  OAI22_X1   g11012(.A1(new_n9621_), .A2(new_n12007_), .B1(new_n9711_), .B2(new_n9717_), .ZN(new_n12028_));
  NAND2_X1   g11013(.A1(new_n12027_), .A2(new_n12028_), .ZN(new_n12029_));
  NOR2_X1    g11014(.A1(new_n9718_), .A2(new_n9621_), .ZN(new_n12030_));
  NAND4_X1   g11015(.A1(new_n12029_), .A2(new_n12025_), .A3(new_n9733_), .A4(new_n12030_), .ZN(new_n12031_));
  NAND4_X1   g11016(.A1(new_n12031_), .A2(new_n12006_), .A3(new_n12017_), .A4(new_n12024_), .ZN(new_n12032_));
  NOR2_X1    g11017(.A1(new_n9737_), .A2(new_n9725_), .ZN(new_n12033_));
  NOR2_X1    g11018(.A1(new_n9662_), .A2(new_n9591_), .ZN(new_n12034_));
  AOI21_X1   g11019(.A1(new_n9690_), .A2(new_n9702_), .B(new_n9720_), .ZN(new_n12035_));
  NOR3_X1    g11020(.A1(new_n9622_), .A2(new_n11972_), .A3(new_n11974_), .ZN(new_n12036_));
  OAI22_X1   g11021(.A1(new_n12034_), .A2(new_n12033_), .B1(new_n12035_), .B2(new_n12036_), .ZN(new_n12037_));
  NOR2_X1    g11022(.A1(new_n12032_), .A2(new_n12037_), .ZN(new_n12038_));
  NAND2_X1   g11023(.A1(new_n12038_), .A2(new_n12005_), .ZN(new_n12039_));
  OAI21_X1   g11024(.A1(new_n12015_), .A2(new_n12012_), .B(new_n9602_), .ZN(new_n12040_));
  NAND3_X1   g11025(.A1(new_n12008_), .A2(new_n12010_), .A3(new_n9711_), .ZN(new_n12041_));
  NAND2_X1   g11026(.A1(new_n12040_), .A2(new_n12041_), .ZN(new_n12042_));
  NAND2_X1   g11027(.A1(new_n12006_), .A2(new_n12042_), .ZN(new_n12043_));
  NOR4_X1    g11028(.A1(new_n9736_), .A2(new_n9733_), .A3(new_n9613_), .A4(new_n9614_), .ZN(new_n12044_));
  NAND3_X1   g11029(.A1(new_n9733_), .A2(new_n9613_), .A3(new_n9620_), .ZN(new_n12045_));
  AOI21_X1   g11030(.A1(new_n12027_), .A2(new_n12028_), .B(new_n12045_), .ZN(new_n12046_));
  AOI21_X1   g11031(.A1(new_n12046_), .A2(new_n12025_), .B(new_n12044_), .ZN(new_n12047_));
  NAND2_X1   g11032(.A1(new_n9662_), .A2(new_n9591_), .ZN(new_n12048_));
  NAND2_X1   g11033(.A1(new_n9737_), .A2(new_n9725_), .ZN(new_n12049_));
  OAI21_X1   g11034(.A1(new_n11972_), .A2(new_n11974_), .B(new_n9622_), .ZN(new_n12050_));
  NAND3_X1   g11035(.A1(new_n9720_), .A2(new_n9690_), .A3(new_n9702_), .ZN(new_n12051_));
  AOI22_X1   g11036(.A1(new_n12048_), .A2(new_n12049_), .B1(new_n12050_), .B2(new_n12051_), .ZN(new_n12052_));
  NAND4_X1   g11037(.A1(new_n12052_), .A2(new_n12047_), .A3(new_n12043_), .A4(new_n12024_), .ZN(new_n12053_));
  NAND2_X1   g11038(.A1(new_n12053_), .A2(new_n12004_), .ZN(new_n12054_));
  AOI21_X1   g11039(.A1(new_n12039_), .A2(new_n12054_), .B(new_n11991_), .ZN(new_n12055_));
  INV_X1     g11040(.I(new_n12055_), .ZN(new_n12056_));
  NAND3_X1   g11041(.A1(new_n9808_), .A2(new_n9798_), .A3(new_n9800_), .ZN(new_n12057_));
  OAI21_X1   g11042(.A1(new_n9773_), .A2(new_n9777_), .B(new_n9792_), .ZN(new_n12058_));
  AOI21_X1   g11043(.A1(new_n12057_), .A2(new_n12058_), .B(new_n9807_), .ZN(new_n12059_));
  NOR3_X1    g11044(.A1(new_n9777_), .A2(new_n9792_), .A3(new_n9773_), .ZN(new_n12060_));
  INV_X1     g11045(.I(new_n12058_), .ZN(new_n12061_));
  NOR3_X1    g11046(.A1(new_n12061_), .A2(new_n9789_), .A3(new_n12060_), .ZN(new_n12062_));
  NOR2_X1    g11047(.A1(new_n12062_), .A2(new_n12059_), .ZN(new_n12063_));
  NOR2_X1    g11048(.A1(new_n9809_), .A2(new_n9767_), .ZN(new_n12064_));
  INV_X1     g11049(.I(new_n12064_), .ZN(new_n12065_));
  NAND2_X1   g11050(.A1(new_n9754_), .A2(\A[198] ), .ZN(new_n12066_));
  NAND2_X1   g11051(.A1(new_n9752_), .A2(\A[197] ), .ZN(new_n12067_));
  AOI21_X1   g11052(.A1(new_n12066_), .A2(new_n12067_), .B(new_n9757_), .ZN(new_n12068_));
  NAND2_X1   g11053(.A1(\A[197] ), .A2(\A[198] ), .ZN(new_n12069_));
  INV_X1     g11054(.I(new_n9759_), .ZN(new_n12070_));
  AOI21_X1   g11055(.A1(new_n12070_), .A2(new_n12069_), .B(\A[196] ), .ZN(new_n12071_));
  NOR2_X1    g11056(.A1(new_n12071_), .A2(new_n12068_), .ZN(new_n12072_));
  NAND2_X1   g11057(.A1(new_n9743_), .A2(\A[195] ), .ZN(new_n12073_));
  NAND2_X1   g11058(.A1(new_n9741_), .A2(\A[194] ), .ZN(new_n12074_));
  AOI21_X1   g11059(.A1(new_n12073_), .A2(new_n12074_), .B(new_n9746_), .ZN(new_n12075_));
  INV_X1     g11060(.I(new_n9749_), .ZN(new_n12076_));
  AOI21_X1   g11061(.A1(new_n12076_), .A2(new_n9747_), .B(\A[193] ), .ZN(new_n12077_));
  OAI22_X1   g11062(.A1(new_n9749_), .A2(new_n9762_), .B1(new_n9764_), .B2(new_n9759_), .ZN(new_n12078_));
  NOR3_X1    g11063(.A1(new_n12077_), .A2(new_n12078_), .A3(new_n12075_), .ZN(new_n12079_));
  AOI21_X1   g11064(.A1(new_n9745_), .A2(new_n9750_), .B(new_n9766_), .ZN(new_n12080_));
  OAI21_X1   g11065(.A1(new_n12080_), .A2(new_n12079_), .B(new_n12072_), .ZN(new_n12081_));
  NAND3_X1   g11066(.A1(new_n9766_), .A2(new_n9745_), .A3(new_n9750_), .ZN(new_n12082_));
  OAI21_X1   g11067(.A1(new_n12075_), .A2(new_n12077_), .B(new_n12078_), .ZN(new_n12083_));
  NAND3_X1   g11068(.A1(new_n12082_), .A2(new_n12083_), .A3(new_n9761_), .ZN(new_n12084_));
  NOR2_X1    g11069(.A1(new_n12072_), .A2(new_n9751_), .ZN(new_n12085_));
  NOR2_X1    g11070(.A1(new_n12077_), .A2(new_n12075_), .ZN(new_n12086_));
  NOR2_X1    g11071(.A1(new_n12086_), .A2(new_n9761_), .ZN(new_n12087_));
  OAI21_X1   g11072(.A1(new_n12085_), .A2(new_n12087_), .B(new_n9766_), .ZN(new_n12088_));
  NAND3_X1   g11073(.A1(new_n12088_), .A2(new_n12081_), .A3(new_n12084_), .ZN(new_n12089_));
  XOR2_X1    g11074(.A1(new_n12089_), .A2(new_n12065_), .Z(new_n12090_));
  NAND2_X1   g11075(.A1(new_n12090_), .A2(new_n12063_), .ZN(new_n12091_));
  OAI21_X1   g11076(.A1(new_n12061_), .A2(new_n12060_), .B(new_n9789_), .ZN(new_n12092_));
  NAND3_X1   g11077(.A1(new_n12057_), .A2(new_n12058_), .A3(new_n9807_), .ZN(new_n12093_));
  NAND2_X1   g11078(.A1(new_n12092_), .A2(new_n12093_), .ZN(new_n12094_));
  AOI22_X1   g11079(.A1(new_n9798_), .A2(new_n9800_), .B1(new_n9804_), .B2(new_n9806_), .ZN(new_n12095_));
  NOR4_X1    g11080(.A1(new_n9773_), .A2(new_n9777_), .A3(new_n9788_), .A4(new_n9784_), .ZN(new_n12096_));
  NOR2_X1    g11081(.A1(new_n9791_), .A2(new_n9786_), .ZN(new_n12097_));
  INV_X1     g11082(.I(new_n12097_), .ZN(new_n12098_));
  NAND4_X1   g11083(.A1(new_n12098_), .A2(new_n9768_), .A3(new_n9769_), .A4(new_n9771_), .ZN(new_n12099_));
  OAI22_X1   g11084(.A1(new_n12095_), .A2(new_n12096_), .B1(new_n12099_), .B2(new_n9789_), .ZN(new_n12100_));
  NOR4_X1    g11085(.A1(new_n12100_), .A2(new_n12086_), .A3(new_n12072_), .A4(new_n12078_), .ZN(new_n12101_));
  NAND2_X1   g11086(.A1(new_n12101_), .A2(new_n12094_), .ZN(new_n12102_));
  AOI21_X1   g11087(.A1(new_n12102_), .A2(new_n12089_), .B(new_n12065_), .ZN(new_n12103_));
  NAND2_X1   g11088(.A1(new_n9879_), .A2(new_n9864_), .ZN(new_n12104_));
  NAND3_X1   g11089(.A1(new_n9837_), .A2(new_n9815_), .A3(new_n9820_), .ZN(new_n12105_));
  OAI21_X1   g11090(.A1(new_n9868_), .A2(new_n9870_), .B(new_n9878_), .ZN(new_n12106_));
  AOI21_X1   g11091(.A1(new_n12105_), .A2(new_n12106_), .B(new_n9832_), .ZN(new_n12107_));
  NOR3_X1    g11092(.A1(new_n9870_), .A2(new_n9878_), .A3(new_n9868_), .ZN(new_n12108_));
  INV_X1     g11093(.I(new_n9834_), .ZN(new_n12109_));
  INV_X1     g11094(.I(new_n9836_), .ZN(new_n12110_));
  AOI22_X1   g11095(.A1(new_n12109_), .A2(new_n12110_), .B1(new_n9815_), .B2(new_n9820_), .ZN(new_n12111_));
  NOR3_X1    g11096(.A1(new_n12111_), .A2(new_n9877_), .A3(new_n12108_), .ZN(new_n12112_));
  NOR2_X1    g11097(.A1(new_n12112_), .A2(new_n12107_), .ZN(new_n12113_));
  NOR2_X1    g11098(.A1(new_n9877_), .A2(new_n9821_), .ZN(new_n12114_));
  NOR2_X1    g11099(.A1(new_n9871_), .A2(new_n9832_), .ZN(new_n12115_));
  OAI21_X1   g11100(.A1(new_n12114_), .A2(new_n12115_), .B(new_n9837_), .ZN(new_n12116_));
  NAND3_X1   g11101(.A1(new_n12113_), .A2(new_n12104_), .A3(new_n12116_), .ZN(new_n12117_));
  NAND2_X1   g11102(.A1(new_n9849_), .A2(new_n9892_), .ZN(new_n12118_));
  OAI21_X1   g11103(.A1(new_n9844_), .A2(new_n9848_), .B(new_n9863_), .ZN(new_n12119_));
  AOI21_X1   g11104(.A1(new_n12118_), .A2(new_n12119_), .B(new_n9891_), .ZN(new_n12120_));
  INV_X1     g11105(.I(new_n12120_), .ZN(new_n12121_));
  NAND3_X1   g11106(.A1(new_n12118_), .A2(new_n9891_), .A3(new_n12119_), .ZN(new_n12122_));
  NAND2_X1   g11107(.A1(new_n12121_), .A2(new_n12122_), .ZN(new_n12123_));
  OAI22_X1   g11108(.A1(new_n9844_), .A2(new_n9848_), .B1(new_n9859_), .B2(new_n9855_), .ZN(new_n12124_));
  NAND4_X1   g11109(.A1(new_n9882_), .A2(new_n9884_), .A3(new_n9888_), .A4(new_n9890_), .ZN(new_n12125_));
  NAND2_X1   g11110(.A1(new_n12124_), .A2(new_n12125_), .ZN(new_n12126_));
  NOR2_X1    g11111(.A1(new_n9862_), .A2(new_n9857_), .ZN(new_n12127_));
  INV_X1     g11112(.I(new_n12127_), .ZN(new_n12128_));
  NAND4_X1   g11113(.A1(new_n12128_), .A2(new_n9839_), .A3(new_n9840_), .A4(new_n9842_), .ZN(new_n12129_));
  NAND4_X1   g11114(.A1(new_n12126_), .A2(new_n9821_), .A3(new_n9832_), .A4(new_n9837_), .ZN(new_n12131_));
  NAND4_X1   g11115(.A1(new_n9900_), .A2(new_n12117_), .A3(new_n12123_), .A4(new_n12131_), .ZN(new_n12132_));
  NOR2_X1    g11116(.A1(new_n12132_), .A2(new_n12103_), .ZN(new_n12133_));
  AOI21_X1   g11117(.A1(new_n12082_), .A2(new_n12083_), .B(new_n9761_), .ZN(new_n12134_));
  NOR3_X1    g11118(.A1(new_n12080_), .A2(new_n12072_), .A3(new_n12079_), .ZN(new_n12135_));
  NAND2_X1   g11119(.A1(new_n12086_), .A2(new_n9761_), .ZN(new_n12136_));
  NAND2_X1   g11120(.A1(new_n12072_), .A2(new_n9751_), .ZN(new_n12137_));
  AOI21_X1   g11121(.A1(new_n12137_), .A2(new_n12136_), .B(new_n12078_), .ZN(new_n12138_));
  NOR3_X1    g11122(.A1(new_n12138_), .A2(new_n12134_), .A3(new_n12135_), .ZN(new_n12139_));
  OAI22_X1   g11123(.A1(new_n9773_), .A2(new_n9777_), .B1(new_n9788_), .B2(new_n9784_), .ZN(new_n12140_));
  NAND4_X1   g11124(.A1(new_n9798_), .A2(new_n9800_), .A3(new_n9804_), .A4(new_n9806_), .ZN(new_n12141_));
  AOI21_X1   g11125(.A1(new_n9798_), .A2(new_n9800_), .B(new_n9792_), .ZN(new_n12142_));
  AOI22_X1   g11126(.A1(new_n12140_), .A2(new_n12141_), .B1(new_n9807_), .B2(new_n12142_), .ZN(new_n12143_));
  NAND4_X1   g11127(.A1(new_n12143_), .A2(new_n9751_), .A3(new_n9761_), .A4(new_n9766_), .ZN(new_n12144_));
  NOR2_X1    g11128(.A1(new_n12144_), .A2(new_n12063_), .ZN(new_n12145_));
  OAI21_X1   g11129(.A1(new_n12145_), .A2(new_n12139_), .B(new_n12064_), .ZN(new_n12146_));
  NAND4_X1   g11130(.A1(new_n9810_), .A2(new_n9865_), .A3(new_n9894_), .A4(new_n9794_), .ZN(new_n12147_));
  NOR2_X1    g11131(.A1(new_n9838_), .A2(new_n9893_), .ZN(new_n12148_));
  OAI21_X1   g11132(.A1(new_n12111_), .A2(new_n12108_), .B(new_n9877_), .ZN(new_n12149_));
  NAND3_X1   g11133(.A1(new_n12105_), .A2(new_n12106_), .A3(new_n9832_), .ZN(new_n12150_));
  NAND2_X1   g11134(.A1(new_n12149_), .A2(new_n12150_), .ZN(new_n12151_));
  NAND2_X1   g11135(.A1(new_n9871_), .A2(new_n9832_), .ZN(new_n12152_));
  NAND2_X1   g11136(.A1(new_n9877_), .A2(new_n9821_), .ZN(new_n12153_));
  AOI21_X1   g11137(.A1(new_n12152_), .A2(new_n12153_), .B(new_n9878_), .ZN(new_n12154_));
  NOR3_X1    g11138(.A1(new_n12151_), .A2(new_n12154_), .A3(new_n12148_), .ZN(new_n12155_));
  NOR2_X1    g11139(.A1(new_n9885_), .A2(new_n9863_), .ZN(new_n12156_));
  INV_X1     g11140(.I(new_n12119_), .ZN(new_n12157_));
  NOR3_X1    g11141(.A1(new_n12157_), .A2(new_n12156_), .A3(new_n9860_), .ZN(new_n12158_));
  NOR2_X1    g11142(.A1(new_n12158_), .A2(new_n12120_), .ZN(new_n12159_));
  INV_X1     g11143(.I(new_n12131_), .ZN(new_n12160_));
  NOR4_X1    g11144(.A1(new_n12147_), .A2(new_n12155_), .A3(new_n12160_), .A4(new_n12159_), .ZN(new_n12161_));
  NOR2_X1    g11145(.A1(new_n12146_), .A2(new_n12161_), .ZN(new_n12162_));
  OAI21_X1   g11146(.A1(new_n12133_), .A2(new_n12162_), .B(new_n12091_), .ZN(new_n12163_));
  XOR2_X1    g11147(.A1(new_n12089_), .A2(new_n12064_), .Z(new_n12164_));
  NOR2_X1    g11148(.A1(new_n12164_), .A2(new_n12094_), .ZN(new_n12165_));
  NAND2_X1   g11149(.A1(new_n12146_), .A2(new_n12161_), .ZN(new_n12166_));
  NAND2_X1   g11150(.A1(new_n12132_), .A2(new_n12103_), .ZN(new_n12167_));
  NAND3_X1   g11151(.A1(new_n12165_), .A2(new_n12167_), .A3(new_n12166_), .ZN(new_n12168_));
  NAND2_X1   g11152(.A1(new_n12163_), .A2(new_n12168_), .ZN(new_n12169_));
  NAND3_X1   g11153(.A1(new_n12056_), .A2(new_n9903_), .A3(new_n12169_), .ZN(new_n12170_));
  NAND3_X1   g11154(.A1(new_n9903_), .A2(new_n12169_), .A3(new_n12055_), .ZN(new_n12171_));
  NAND2_X1   g11155(.A1(new_n12170_), .A2(new_n12171_), .ZN(new_n12172_));
  NAND3_X1   g11156(.A1(new_n12172_), .A2(new_n9905_), .A3(new_n10225_), .ZN(new_n12173_));
  NAND2_X1   g11157(.A1(new_n12173_), .A2(new_n11961_), .ZN(new_n12174_));
  NOR2_X1    g11158(.A1(new_n10380_), .A2(new_n10280_), .ZN(new_n12175_));
  INV_X1     g11159(.I(new_n12175_), .ZN(new_n12176_));
  NOR3_X1    g11160(.A1(new_n10237_), .A2(new_n10252_), .A3(new_n10233_), .ZN(new_n12177_));
  OAI21_X1   g11161(.A1(new_n10233_), .A2(new_n10237_), .B(new_n10252_), .ZN(new_n12178_));
  INV_X1     g11162(.I(new_n12178_), .ZN(new_n12179_));
  OAI21_X1   g11163(.A1(new_n12179_), .A2(new_n12177_), .B(new_n10249_), .ZN(new_n12180_));
  NAND2_X1   g11164(.A1(new_n10238_), .A2(new_n10379_), .ZN(new_n12181_));
  NAND3_X1   g11165(.A1(new_n12181_), .A2(new_n12178_), .A3(new_n10378_), .ZN(new_n12182_));
  NOR2_X1    g11166(.A1(new_n10249_), .A2(new_n10372_), .ZN(new_n12183_));
  NOR2_X1    g11167(.A1(new_n10238_), .A2(new_n10378_), .ZN(new_n12184_));
  OAI21_X1   g11168(.A1(new_n12183_), .A2(new_n12184_), .B(new_n10379_), .ZN(new_n12185_));
  NAND3_X1   g11169(.A1(new_n12185_), .A2(new_n12180_), .A3(new_n12182_), .ZN(new_n12186_));
  NAND2_X1   g11170(.A1(new_n12180_), .A2(new_n12182_), .ZN(new_n12187_));
  AOI22_X1   g11171(.A1(new_n10258_), .A2(new_n10263_), .B1(new_n10269_), .B2(new_n10274_), .ZN(new_n12188_));
  NAND2_X1   g11172(.A1(new_n10256_), .A2(\A[165] ), .ZN(new_n12189_));
  NAND2_X1   g11173(.A1(new_n10254_), .A2(\A[164] ), .ZN(new_n12190_));
  AOI21_X1   g11174(.A1(new_n12189_), .A2(new_n12190_), .B(new_n10259_), .ZN(new_n12191_));
  INV_X1     g11175(.I(new_n10262_), .ZN(new_n12192_));
  AOI21_X1   g11176(.A1(new_n12192_), .A2(new_n10260_), .B(\A[163] ), .ZN(new_n12193_));
  NAND2_X1   g11177(.A1(new_n10267_), .A2(\A[168] ), .ZN(new_n12194_));
  NAND2_X1   g11178(.A1(new_n10265_), .A2(\A[167] ), .ZN(new_n12195_));
  AOI21_X1   g11179(.A1(new_n12194_), .A2(new_n12195_), .B(new_n10270_), .ZN(new_n12196_));
  INV_X1     g11180(.I(new_n10273_), .ZN(new_n12197_));
  AOI21_X1   g11181(.A1(new_n12197_), .A2(new_n10271_), .B(\A[166] ), .ZN(new_n12198_));
  NOR4_X1    g11182(.A1(new_n12191_), .A2(new_n12193_), .A3(new_n12198_), .A4(new_n12196_), .ZN(new_n12199_));
  NOR2_X1    g11183(.A1(new_n12188_), .A2(new_n12199_), .ZN(new_n12200_));
  NOR2_X1    g11184(.A1(new_n12193_), .A2(new_n12191_), .ZN(new_n12201_));
  NOR2_X1    g11185(.A1(new_n12198_), .A2(new_n12196_), .ZN(new_n12202_));
  NOR3_X1    g11186(.A1(new_n12201_), .A2(new_n12202_), .A3(new_n10278_), .ZN(new_n12203_));
  NOR3_X1    g11187(.A1(new_n12200_), .A2(new_n10380_), .A3(new_n12203_), .ZN(new_n12204_));
  NOR3_X1    g11188(.A1(new_n12193_), .A2(new_n10278_), .A3(new_n12191_), .ZN(new_n12205_));
  NOR2_X1    g11189(.A1(new_n10276_), .A2(new_n10262_), .ZN(new_n12206_));
  INV_X1     g11190(.I(new_n12206_), .ZN(new_n12207_));
  NOR2_X1    g11191(.A1(new_n10277_), .A2(new_n10273_), .ZN(new_n12208_));
  INV_X1     g11192(.I(new_n12208_), .ZN(new_n12209_));
  AOI22_X1   g11193(.A1(new_n12207_), .A2(new_n12209_), .B1(new_n10258_), .B2(new_n10263_), .ZN(new_n12210_));
  OAI21_X1   g11194(.A1(new_n12210_), .A2(new_n12205_), .B(new_n12202_), .ZN(new_n12211_));
  NAND3_X1   g11195(.A1(new_n10279_), .A2(new_n10258_), .A3(new_n10263_), .ZN(new_n12212_));
  OAI21_X1   g11196(.A1(new_n12191_), .A2(new_n12193_), .B(new_n10278_), .ZN(new_n12213_));
  NAND3_X1   g11197(.A1(new_n12212_), .A2(new_n12213_), .A3(new_n10275_), .ZN(new_n12214_));
  NAND2_X1   g11198(.A1(new_n12214_), .A2(new_n12211_), .ZN(new_n12215_));
  NAND4_X1   g11199(.A1(new_n12187_), .A2(new_n12204_), .A3(new_n12215_), .A4(new_n12185_), .ZN(new_n12216_));
  AOI21_X1   g11200(.A1(new_n12216_), .A2(new_n12186_), .B(new_n12176_), .ZN(new_n12217_));
  AOI21_X1   g11201(.A1(new_n12181_), .A2(new_n12178_), .B(new_n10378_), .ZN(new_n12218_));
  NOR3_X1    g11202(.A1(new_n12179_), .A2(new_n10249_), .A3(new_n12177_), .ZN(new_n12219_));
  NAND2_X1   g11203(.A1(new_n10238_), .A2(new_n10378_), .ZN(new_n12220_));
  NAND2_X1   g11204(.A1(new_n10249_), .A2(new_n10372_), .ZN(new_n12221_));
  AOI21_X1   g11205(.A1(new_n12220_), .A2(new_n12221_), .B(new_n10252_), .ZN(new_n12222_));
  NOR3_X1    g11206(.A1(new_n12222_), .A2(new_n12219_), .A3(new_n12218_), .ZN(new_n12223_));
  NAND2_X1   g11207(.A1(new_n12223_), .A2(new_n12176_), .ZN(new_n12224_));
  NAND2_X1   g11208(.A1(new_n12186_), .A2(new_n12175_), .ZN(new_n12225_));
  AOI21_X1   g11209(.A1(new_n12224_), .A2(new_n12225_), .B(new_n12215_), .ZN(new_n12226_));
  NOR4_X1    g11210(.A1(new_n10283_), .A2(new_n10337_), .A3(new_n10365_), .A4(new_n10281_), .ZN(new_n12227_));
  NOR2_X1    g11211(.A1(new_n10351_), .A2(new_n10336_), .ZN(new_n12228_));
  INV_X1     g11212(.I(new_n12228_), .ZN(new_n12229_));
  NAND2_X1   g11213(.A1(new_n10294_), .A2(new_n10350_), .ZN(new_n12230_));
  OAI21_X1   g11214(.A1(new_n10289_), .A2(new_n10293_), .B(new_n10308_), .ZN(new_n12231_));
  AOI21_X1   g11215(.A1(new_n12230_), .A2(new_n12231_), .B(new_n10349_), .ZN(new_n12232_));
  NOR2_X1    g11216(.A1(new_n10343_), .A2(new_n10308_), .ZN(new_n12233_));
  INV_X1     g11217(.I(new_n12231_), .ZN(new_n12234_));
  NOR3_X1    g11218(.A1(new_n12234_), .A2(new_n12233_), .A3(new_n10305_), .ZN(new_n12235_));
  NAND2_X1   g11219(.A1(new_n10294_), .A2(new_n10349_), .ZN(new_n12236_));
  NAND2_X1   g11220(.A1(new_n10305_), .A2(new_n10343_), .ZN(new_n12237_));
  AOI21_X1   g11221(.A1(new_n12236_), .A2(new_n12237_), .B(new_n10308_), .ZN(new_n12238_));
  NOR3_X1    g11222(.A1(new_n12238_), .A2(new_n12235_), .A3(new_n12232_), .ZN(new_n12239_));
  NAND2_X1   g11223(.A1(new_n12239_), .A2(new_n12229_), .ZN(new_n12240_));
  NOR2_X1    g11224(.A1(new_n10320_), .A2(new_n10334_), .ZN(new_n12241_));
  NOR2_X1    g11225(.A1(new_n10357_), .A2(new_n10335_), .ZN(new_n12242_));
  OAI21_X1   g11226(.A1(new_n12242_), .A2(new_n12241_), .B(new_n10363_), .ZN(new_n12243_));
  NAND2_X1   g11227(.A1(new_n10357_), .A2(new_n10335_), .ZN(new_n12244_));
  NAND2_X1   g11228(.A1(new_n10320_), .A2(new_n10334_), .ZN(new_n12245_));
  NAND3_X1   g11229(.A1(new_n12244_), .A2(new_n12245_), .A3(new_n10331_), .ZN(new_n12246_));
  NAND2_X1   g11230(.A1(new_n12243_), .A2(new_n12246_), .ZN(new_n12247_));
  OAI22_X1   g11231(.A1(new_n10354_), .A2(new_n10356_), .B1(new_n10362_), .B2(new_n10360_), .ZN(new_n12248_));
  NAND4_X1   g11232(.A1(new_n10314_), .A2(new_n10319_), .A3(new_n10325_), .A4(new_n10330_), .ZN(new_n12249_));
  NAND2_X1   g11233(.A1(new_n12248_), .A2(new_n12249_), .ZN(new_n12250_));
  NOR2_X1    g11234(.A1(new_n10333_), .A2(new_n10329_), .ZN(new_n12251_));
  INV_X1     g11235(.I(new_n12251_), .ZN(new_n12252_));
  NAND4_X1   g11236(.A1(new_n12252_), .A2(new_n10315_), .A3(new_n10312_), .A4(new_n10310_), .ZN(new_n12253_));
  NAND4_X1   g11237(.A1(new_n12250_), .A2(new_n10343_), .A3(new_n10349_), .A4(new_n10350_), .ZN(new_n12255_));
  NAND4_X1   g11238(.A1(new_n12240_), .A2(new_n12227_), .A3(new_n12247_), .A4(new_n12255_), .ZN(new_n12256_));
  NOR2_X1    g11239(.A1(new_n12256_), .A2(new_n12226_), .ZN(new_n12257_));
  NAND2_X1   g11240(.A1(new_n12256_), .A2(new_n12226_), .ZN(new_n12258_));
  INV_X1     g11241(.I(new_n12258_), .ZN(new_n12259_));
  OAI21_X1   g11242(.A1(new_n12259_), .A2(new_n12257_), .B(new_n12217_), .ZN(new_n12260_));
  NAND3_X1   g11243(.A1(new_n10439_), .A2(new_n10417_), .A3(new_n10422_), .ZN(new_n12261_));
  OAI21_X1   g11244(.A1(new_n10460_), .A2(new_n10462_), .B(new_n10470_), .ZN(new_n12262_));
  AOI21_X1   g11245(.A1(new_n12261_), .A2(new_n12262_), .B(new_n10434_), .ZN(new_n12263_));
  NAND3_X1   g11246(.A1(new_n12261_), .A2(new_n12262_), .A3(new_n10434_), .ZN(new_n12264_));
  INV_X1     g11247(.I(new_n12264_), .ZN(new_n12265_));
  NOR2_X1    g11248(.A1(new_n12265_), .A2(new_n12263_), .ZN(new_n12266_));
  NOR2_X1    g11249(.A1(new_n10440_), .A2(new_n10457_), .ZN(new_n12267_));
  NOR3_X1    g11250(.A1(new_n10396_), .A2(new_n10411_), .A3(new_n10392_), .ZN(new_n12268_));
  INV_X1     g11251(.I(new_n10454_), .ZN(new_n12269_));
  INV_X1     g11252(.I(new_n10455_), .ZN(new_n12270_));
  AOI22_X1   g11253(.A1(new_n12269_), .A2(new_n12270_), .B1(new_n10444_), .B2(new_n10446_), .ZN(new_n12271_));
  OAI21_X1   g11254(.A1(new_n12271_), .A2(new_n12268_), .B(new_n10408_), .ZN(new_n12272_));
  NAND3_X1   g11255(.A1(new_n10456_), .A2(new_n10444_), .A3(new_n10446_), .ZN(new_n12273_));
  OAI21_X1   g11256(.A1(new_n10392_), .A2(new_n10396_), .B(new_n10411_), .ZN(new_n12274_));
  NAND3_X1   g11257(.A1(new_n12273_), .A2(new_n12274_), .A3(new_n10453_), .ZN(new_n12275_));
  NOR2_X1    g11258(.A1(new_n10408_), .A2(new_n10447_), .ZN(new_n12276_));
  NOR2_X1    g11259(.A1(new_n10397_), .A2(new_n10453_), .ZN(new_n12277_));
  OAI21_X1   g11260(.A1(new_n12277_), .A2(new_n12276_), .B(new_n10456_), .ZN(new_n12278_));
  NAND3_X1   g11261(.A1(new_n12278_), .A2(new_n12272_), .A3(new_n12275_), .ZN(new_n12279_));
  NOR2_X1    g11262(.A1(new_n12279_), .A2(new_n12267_), .ZN(new_n12280_));
  INV_X1     g11263(.I(new_n12267_), .ZN(new_n12281_));
  NAND2_X1   g11264(.A1(new_n12272_), .A2(new_n12275_), .ZN(new_n12282_));
  NAND2_X1   g11265(.A1(new_n10397_), .A2(new_n10453_), .ZN(new_n12283_));
  NAND2_X1   g11266(.A1(new_n10408_), .A2(new_n10447_), .ZN(new_n12284_));
  AOI21_X1   g11267(.A1(new_n12283_), .A2(new_n12284_), .B(new_n10411_), .ZN(new_n12285_));
  NOR2_X1    g11268(.A1(new_n12282_), .A2(new_n12285_), .ZN(new_n12286_));
  NOR2_X1    g11269(.A1(new_n12286_), .A2(new_n12281_), .ZN(new_n12287_));
  OAI21_X1   g11270(.A1(new_n12287_), .A2(new_n12280_), .B(new_n12266_), .ZN(new_n12288_));
  NOR3_X1    g11271(.A1(new_n10462_), .A2(new_n10470_), .A3(new_n10460_), .ZN(new_n12289_));
  AOI21_X1   g11272(.A1(new_n10417_), .A2(new_n10422_), .B(new_n10439_), .ZN(new_n12290_));
  OAI21_X1   g11273(.A1(new_n12290_), .A2(new_n12289_), .B(new_n10469_), .ZN(new_n12291_));
  NAND2_X1   g11274(.A1(new_n12291_), .A2(new_n12264_), .ZN(new_n12292_));
  AOI22_X1   g11275(.A1(new_n10417_), .A2(new_n10422_), .B1(new_n10428_), .B2(new_n10433_), .ZN(new_n12293_));
  NOR4_X1    g11276(.A1(new_n10460_), .A2(new_n10462_), .A3(new_n10468_), .A4(new_n10466_), .ZN(new_n12294_));
  NOR2_X1    g11277(.A1(new_n12293_), .A2(new_n12294_), .ZN(new_n12295_));
  NOR3_X1    g11278(.A1(new_n10463_), .A2(new_n10469_), .A3(new_n10470_), .ZN(new_n12296_));
  NOR3_X1    g11279(.A1(new_n12295_), .A2(new_n10457_), .A3(new_n12296_), .ZN(new_n12297_));
  NAND4_X1   g11280(.A1(new_n12297_), .A2(new_n12292_), .A3(new_n12282_), .A4(new_n12278_), .ZN(new_n12298_));
  AOI21_X1   g11281(.A1(new_n12298_), .A2(new_n12279_), .B(new_n12281_), .ZN(new_n12299_));
  NOR4_X1    g11282(.A1(new_n10441_), .A2(new_n10472_), .A3(new_n10526_), .A4(new_n10556_), .ZN(new_n12300_));
  NAND2_X1   g11283(.A1(new_n10498_), .A2(new_n10555_), .ZN(new_n12301_));
  NOR3_X1    g11284(.A1(new_n10482_), .A2(new_n10497_), .A3(new_n10478_), .ZN(new_n12302_));
  NOR2_X1    g11285(.A1(new_n10483_), .A2(new_n10541_), .ZN(new_n12303_));
  OAI21_X1   g11286(.A1(new_n12303_), .A2(new_n12302_), .B(new_n10494_), .ZN(new_n12304_));
  NAND3_X1   g11287(.A1(new_n10541_), .A2(new_n10529_), .A3(new_n10531_), .ZN(new_n12305_));
  OAI21_X1   g11288(.A1(new_n10478_), .A2(new_n10482_), .B(new_n10497_), .ZN(new_n12306_));
  NAND3_X1   g11289(.A1(new_n12305_), .A2(new_n12306_), .A3(new_n10538_), .ZN(new_n12307_));
  NOR2_X1    g11290(.A1(new_n10494_), .A2(new_n10532_), .ZN(new_n12308_));
  NOR2_X1    g11291(.A1(new_n10483_), .A2(new_n10538_), .ZN(new_n12309_));
  OAI21_X1   g11292(.A1(new_n12308_), .A2(new_n12309_), .B(new_n10541_), .ZN(new_n12310_));
  NAND4_X1   g11293(.A1(new_n12301_), .A2(new_n12310_), .A3(new_n12304_), .A4(new_n12307_), .ZN(new_n12311_));
  NOR2_X1    g11294(.A1(new_n10509_), .A2(new_n10523_), .ZN(new_n12312_));
  OAI21_X1   g11295(.A1(new_n10545_), .A2(new_n10547_), .B(new_n10523_), .ZN(new_n12313_));
  INV_X1     g11296(.I(new_n12313_), .ZN(new_n12314_));
  OAI21_X1   g11297(.A1(new_n12314_), .A2(new_n12312_), .B(new_n10554_), .ZN(new_n12315_));
  NAND2_X1   g11298(.A1(new_n10548_), .A2(new_n10524_), .ZN(new_n12316_));
  NAND3_X1   g11299(.A1(new_n12316_), .A2(new_n10520_), .A3(new_n12313_), .ZN(new_n12317_));
  NAND2_X1   g11300(.A1(new_n12315_), .A2(new_n12317_), .ZN(new_n12318_));
  OAI22_X1   g11301(.A1(new_n10545_), .A2(new_n10547_), .B1(new_n10553_), .B2(new_n10551_), .ZN(new_n12319_));
  NAND4_X1   g11302(.A1(new_n10503_), .A2(new_n10508_), .A3(new_n10514_), .A4(new_n10519_), .ZN(new_n12320_));
  NAND2_X1   g11303(.A1(new_n12319_), .A2(new_n12320_), .ZN(new_n12321_));
  AOI21_X1   g11304(.A1(new_n10503_), .A2(new_n10508_), .B(new_n10523_), .ZN(new_n12322_));
  NAND4_X1   g11305(.A1(new_n12321_), .A2(new_n10532_), .A3(new_n10538_), .A4(new_n10541_), .ZN(new_n12325_));
  NAND4_X1   g11306(.A1(new_n12300_), .A2(new_n12311_), .A3(new_n12318_), .A4(new_n12325_), .ZN(new_n12326_));
  NOR2_X1    g11307(.A1(new_n12299_), .A2(new_n12326_), .ZN(new_n12327_));
  OAI22_X1   g11308(.A1(new_n10460_), .A2(new_n10462_), .B1(new_n10468_), .B2(new_n10466_), .ZN(new_n12328_));
  NAND4_X1   g11309(.A1(new_n10417_), .A2(new_n10422_), .A3(new_n10428_), .A4(new_n10433_), .ZN(new_n12329_));
  AOI21_X1   g11310(.A1(new_n10417_), .A2(new_n10422_), .B(new_n10470_), .ZN(new_n12330_));
  AOI22_X1   g11311(.A1(new_n12328_), .A2(new_n12329_), .B1(new_n10434_), .B2(new_n12330_), .ZN(new_n12331_));
  NAND4_X1   g11312(.A1(new_n12331_), .A2(new_n10447_), .A3(new_n10453_), .A4(new_n10456_), .ZN(new_n12332_));
  NOR2_X1    g11313(.A1(new_n12332_), .A2(new_n12266_), .ZN(new_n12333_));
  OAI21_X1   g11314(.A1(new_n12333_), .A2(new_n12286_), .B(new_n12267_), .ZN(new_n12334_));
  NOR2_X1    g11315(.A1(new_n10525_), .A2(new_n10542_), .ZN(new_n12335_));
  AOI21_X1   g11316(.A1(new_n12305_), .A2(new_n12306_), .B(new_n10538_), .ZN(new_n12336_));
  NOR3_X1    g11317(.A1(new_n12303_), .A2(new_n10494_), .A3(new_n12302_), .ZN(new_n12337_));
  NAND2_X1   g11318(.A1(new_n10483_), .A2(new_n10538_), .ZN(new_n12338_));
  NAND2_X1   g11319(.A1(new_n10494_), .A2(new_n10532_), .ZN(new_n12339_));
  AOI21_X1   g11320(.A1(new_n12339_), .A2(new_n12338_), .B(new_n10497_), .ZN(new_n12340_));
  NOR4_X1    g11321(.A1(new_n12340_), .A2(new_n12335_), .A3(new_n12337_), .A4(new_n12336_), .ZN(new_n12341_));
  AOI21_X1   g11322(.A1(new_n12316_), .A2(new_n12313_), .B(new_n10520_), .ZN(new_n12342_));
  NOR3_X1    g11323(.A1(new_n12314_), .A2(new_n12312_), .A3(new_n10554_), .ZN(new_n12343_));
  NOR2_X1    g11324(.A1(new_n12343_), .A2(new_n12342_), .ZN(new_n12344_));
  INV_X1     g11325(.I(new_n12325_), .ZN(new_n12345_));
  NOR4_X1    g11326(.A1(new_n10562_), .A2(new_n12341_), .A3(new_n12345_), .A4(new_n12344_), .ZN(new_n12346_));
  NOR2_X1    g11327(.A1(new_n12334_), .A2(new_n12346_), .ZN(new_n12347_));
  OAI21_X1   g11328(.A1(new_n12347_), .A2(new_n12327_), .B(new_n12288_), .ZN(new_n12348_));
  NAND2_X1   g11329(.A1(new_n12286_), .A2(new_n12281_), .ZN(new_n12349_));
  NAND2_X1   g11330(.A1(new_n12279_), .A2(new_n12267_), .ZN(new_n12350_));
  AOI21_X1   g11331(.A1(new_n12349_), .A2(new_n12350_), .B(new_n12292_), .ZN(new_n12351_));
  NAND2_X1   g11332(.A1(new_n12334_), .A2(new_n12346_), .ZN(new_n12352_));
  NAND2_X1   g11333(.A1(new_n12299_), .A2(new_n12326_), .ZN(new_n12353_));
  NAND3_X1   g11334(.A1(new_n12352_), .A2(new_n12353_), .A3(new_n12351_), .ZN(new_n12354_));
  AOI21_X1   g11335(.A1(new_n12348_), .A2(new_n12354_), .B(new_n10566_), .ZN(new_n12355_));
  NOR2_X1    g11336(.A1(new_n12355_), .A2(new_n12260_), .ZN(new_n12356_));
  NOR2_X1    g11337(.A1(new_n10567_), .A2(new_n10921_), .ZN(new_n12357_));
  INV_X1     g11338(.I(new_n12357_), .ZN(new_n12358_));
  NOR2_X1    g11339(.A1(new_n10595_), .A2(new_n10650_), .ZN(new_n12359_));
  INV_X1     g11340(.I(new_n12359_), .ZN(new_n12360_));
  NAND3_X1   g11341(.A1(new_n10594_), .A2(new_n10572_), .A3(new_n10577_), .ZN(new_n12361_));
  OAI21_X1   g11342(.A1(new_n10625_), .A2(new_n10627_), .B(new_n10635_), .ZN(new_n12362_));
  AOI21_X1   g11343(.A1(new_n12361_), .A2(new_n12362_), .B(new_n10589_), .ZN(new_n12363_));
  NOR3_X1    g11344(.A1(new_n10627_), .A2(new_n10635_), .A3(new_n10625_), .ZN(new_n12364_));
  INV_X1     g11345(.I(new_n10591_), .ZN(new_n12365_));
  INV_X1     g11346(.I(new_n10593_), .ZN(new_n12366_));
  AOI22_X1   g11347(.A1(new_n12365_), .A2(new_n12366_), .B1(new_n10572_), .B2(new_n10577_), .ZN(new_n12367_));
  NOR3_X1    g11348(.A1(new_n12367_), .A2(new_n10634_), .A3(new_n12364_), .ZN(new_n12368_));
  NOR2_X1    g11349(.A1(new_n12368_), .A2(new_n12363_), .ZN(new_n12369_));
  NOR2_X1    g11350(.A1(new_n10634_), .A2(new_n10578_), .ZN(new_n12370_));
  NOR2_X1    g11351(.A1(new_n10628_), .A2(new_n10589_), .ZN(new_n12371_));
  OAI21_X1   g11352(.A1(new_n12370_), .A2(new_n12371_), .B(new_n10594_), .ZN(new_n12372_));
  NAND2_X1   g11353(.A1(new_n12369_), .A2(new_n12372_), .ZN(new_n12373_));
  OAI21_X1   g11354(.A1(new_n12367_), .A2(new_n12364_), .B(new_n10634_), .ZN(new_n12374_));
  NAND3_X1   g11355(.A1(new_n12361_), .A2(new_n12362_), .A3(new_n10589_), .ZN(new_n12375_));
  NAND2_X1   g11356(.A1(new_n12374_), .A2(new_n12375_), .ZN(new_n12376_));
  AOI22_X1   g11357(.A1(new_n10645_), .A2(new_n10647_), .B1(new_n10639_), .B2(new_n10641_), .ZN(new_n12377_));
  NOR4_X1    g11358(.A1(new_n10601_), .A2(new_n10615_), .A3(new_n10611_), .A4(new_n10604_), .ZN(new_n12378_));
  NOR2_X1    g11359(.A1(new_n12377_), .A2(new_n12378_), .ZN(new_n12379_));
  NOR3_X1    g11360(.A1(new_n10616_), .A2(new_n10605_), .A3(new_n10620_), .ZN(new_n12380_));
  NOR3_X1    g11361(.A1(new_n12379_), .A2(new_n10595_), .A3(new_n12380_), .ZN(new_n12381_));
  NOR3_X1    g11362(.A1(new_n10620_), .A2(new_n10601_), .A3(new_n10604_), .ZN(new_n12382_));
  NOR2_X1    g11363(.A1(new_n10618_), .A2(new_n10617_), .ZN(new_n12383_));
  INV_X1     g11364(.I(new_n12383_), .ZN(new_n12384_));
  NOR2_X1    g11365(.A1(new_n10619_), .A2(new_n10613_), .ZN(new_n12385_));
  INV_X1     g11366(.I(new_n12385_), .ZN(new_n12386_));
  AOI22_X1   g11367(.A1(new_n12384_), .A2(new_n12386_), .B1(new_n10639_), .B2(new_n10641_), .ZN(new_n12387_));
  OAI21_X1   g11368(.A1(new_n12387_), .A2(new_n12382_), .B(new_n10616_), .ZN(new_n12388_));
  NAND4_X1   g11369(.A1(new_n12384_), .A2(new_n12386_), .A3(new_n10639_), .A4(new_n10641_), .ZN(new_n12389_));
  OAI21_X1   g11370(.A1(new_n10601_), .A2(new_n10604_), .B(new_n10620_), .ZN(new_n12390_));
  NAND3_X1   g11371(.A1(new_n12389_), .A2(new_n12390_), .A3(new_n10648_), .ZN(new_n12391_));
  NAND2_X1   g11372(.A1(new_n12388_), .A2(new_n12391_), .ZN(new_n12392_));
  NAND4_X1   g11373(.A1(new_n12376_), .A2(new_n12381_), .A3(new_n12392_), .A4(new_n12372_), .ZN(new_n12393_));
  AOI21_X1   g11374(.A1(new_n12393_), .A2(new_n12373_), .B(new_n12360_), .ZN(new_n12394_));
  NAND2_X1   g11375(.A1(new_n10628_), .A2(new_n10589_), .ZN(new_n12395_));
  NAND2_X1   g11376(.A1(new_n10634_), .A2(new_n10578_), .ZN(new_n12396_));
  AOI21_X1   g11377(.A1(new_n12395_), .A2(new_n12396_), .B(new_n10635_), .ZN(new_n12397_));
  NOR2_X1    g11378(.A1(new_n12376_), .A2(new_n12397_), .ZN(new_n12398_));
  NAND2_X1   g11379(.A1(new_n12398_), .A2(new_n12360_), .ZN(new_n12399_));
  NAND2_X1   g11380(.A1(new_n12373_), .A2(new_n12359_), .ZN(new_n12400_));
  AOI21_X1   g11381(.A1(new_n12400_), .A2(new_n12399_), .B(new_n12392_), .ZN(new_n12401_));
  NOR2_X1    g11382(.A1(new_n10652_), .A2(new_n10737_), .ZN(new_n12402_));
  NOR2_X1    g11383(.A1(new_n10735_), .A2(new_n10679_), .ZN(new_n12403_));
  NAND3_X1   g11384(.A1(new_n10678_), .A2(new_n10657_), .A3(new_n10662_), .ZN(new_n12404_));
  OAI21_X1   g11385(.A1(new_n10709_), .A2(new_n10711_), .B(new_n10720_), .ZN(new_n12405_));
  AOI21_X1   g11386(.A1(new_n12404_), .A2(new_n12405_), .B(new_n10673_), .ZN(new_n12406_));
  NOR3_X1    g11387(.A1(new_n10711_), .A2(new_n10720_), .A3(new_n10709_), .ZN(new_n12407_));
  INV_X1     g11388(.I(new_n10675_), .ZN(new_n12408_));
  INV_X1     g11389(.I(new_n10677_), .ZN(new_n12409_));
  AOI22_X1   g11390(.A1(new_n12408_), .A2(new_n12409_), .B1(new_n10657_), .B2(new_n10662_), .ZN(new_n12410_));
  NOR3_X1    g11391(.A1(new_n12410_), .A2(new_n10719_), .A3(new_n12407_), .ZN(new_n12411_));
  NAND2_X1   g11392(.A1(new_n10712_), .A2(new_n10673_), .ZN(new_n12412_));
  NAND2_X1   g11393(.A1(new_n10719_), .A2(new_n10663_), .ZN(new_n12413_));
  AOI21_X1   g11394(.A1(new_n12413_), .A2(new_n12412_), .B(new_n10720_), .ZN(new_n12414_));
  NOR4_X1    g11395(.A1(new_n12414_), .A2(new_n12403_), .A3(new_n12406_), .A4(new_n12411_), .ZN(new_n12415_));
  NAND2_X1   g11396(.A1(new_n10690_), .A2(new_n10734_), .ZN(new_n12416_));
  OAI21_X1   g11397(.A1(new_n10685_), .A2(new_n10689_), .B(new_n10704_), .ZN(new_n12417_));
  AOI21_X1   g11398(.A1(new_n12416_), .A2(new_n12417_), .B(new_n10733_), .ZN(new_n12418_));
  NOR3_X1    g11399(.A1(new_n10689_), .A2(new_n10704_), .A3(new_n10685_), .ZN(new_n12419_));
  INV_X1     g11400(.I(new_n12417_), .ZN(new_n12420_));
  NOR3_X1    g11401(.A1(new_n12420_), .A2(new_n10701_), .A3(new_n12419_), .ZN(new_n12421_));
  NOR2_X1    g11402(.A1(new_n12421_), .A2(new_n12418_), .ZN(new_n12422_));
  AOI22_X1   g11403(.A1(new_n10724_), .A2(new_n10726_), .B1(new_n10730_), .B2(new_n10732_), .ZN(new_n12423_));
  NOR4_X1    g11404(.A1(new_n10685_), .A2(new_n10689_), .A3(new_n10700_), .A4(new_n10696_), .ZN(new_n12424_));
  NOR2_X1    g11405(.A1(new_n12423_), .A2(new_n12424_), .ZN(new_n12425_));
  OAI21_X1   g11406(.A1(\A[106] ), .A2(new_n10731_), .B(new_n10699_), .ZN(new_n12426_));
  NAND4_X1   g11407(.A1(new_n12426_), .A2(new_n10680_), .A3(new_n10681_), .A4(new_n10683_), .ZN(new_n12427_));
  NOR4_X1    g11408(.A1(new_n12425_), .A2(new_n10712_), .A3(new_n10719_), .A4(new_n10720_), .ZN(new_n12429_));
  NOR3_X1    g11409(.A1(new_n12415_), .A2(new_n12422_), .A3(new_n12429_), .ZN(new_n12430_));
  NAND2_X1   g11410(.A1(new_n12430_), .A2(new_n12402_), .ZN(new_n12431_));
  NOR2_X1    g11411(.A1(new_n12401_), .A2(new_n12431_), .ZN(new_n12432_));
  NAND2_X1   g11412(.A1(new_n12401_), .A2(new_n12431_), .ZN(new_n12433_));
  INV_X1     g11413(.I(new_n12433_), .ZN(new_n12434_));
  OAI21_X1   g11414(.A1(new_n12434_), .A2(new_n12432_), .B(new_n12394_), .ZN(new_n12435_));
  NAND3_X1   g11415(.A1(new_n10792_), .A2(new_n10771_), .A3(new_n10776_), .ZN(new_n12436_));
  OAI21_X1   g11416(.A1(new_n10813_), .A2(new_n10815_), .B(new_n10824_), .ZN(new_n12437_));
  AOI21_X1   g11417(.A1(new_n12436_), .A2(new_n12437_), .B(new_n10787_), .ZN(new_n12438_));
  NOR3_X1    g11418(.A1(new_n10815_), .A2(new_n10824_), .A3(new_n10813_), .ZN(new_n12439_));
  AOI21_X1   g11419(.A1(new_n10771_), .A2(new_n10776_), .B(new_n10792_), .ZN(new_n12440_));
  NOR3_X1    g11420(.A1(new_n12440_), .A2(new_n10823_), .A3(new_n12439_), .ZN(new_n12441_));
  NOR2_X1    g11421(.A1(new_n12441_), .A2(new_n12438_), .ZN(new_n12442_));
  NOR2_X1    g11422(.A1(new_n10810_), .A2(new_n10793_), .ZN(new_n12443_));
  NAND3_X1   g11423(.A1(new_n10809_), .A2(new_n10797_), .A3(new_n10799_), .ZN(new_n12444_));
  OAI21_X1   g11424(.A1(new_n10746_), .A2(new_n10750_), .B(new_n10765_), .ZN(new_n12445_));
  AOI21_X1   g11425(.A1(new_n12444_), .A2(new_n12445_), .B(new_n10806_), .ZN(new_n12446_));
  NOR3_X1    g11426(.A1(new_n10750_), .A2(new_n10765_), .A3(new_n10746_), .ZN(new_n12447_));
  INV_X1     g11427(.I(new_n10807_), .ZN(new_n12448_));
  INV_X1     g11428(.I(new_n10808_), .ZN(new_n12449_));
  AOI22_X1   g11429(.A1(new_n12448_), .A2(new_n12449_), .B1(new_n10797_), .B2(new_n10799_), .ZN(new_n12450_));
  NOR3_X1    g11430(.A1(new_n12450_), .A2(new_n10762_), .A3(new_n12447_), .ZN(new_n12451_));
  NOR2_X1    g11431(.A1(new_n12451_), .A2(new_n12446_), .ZN(new_n12452_));
  NOR2_X1    g11432(.A1(new_n10762_), .A2(new_n10800_), .ZN(new_n12453_));
  NOR2_X1    g11433(.A1(new_n10751_), .A2(new_n10806_), .ZN(new_n12454_));
  OAI21_X1   g11434(.A1(new_n12453_), .A2(new_n12454_), .B(new_n10809_), .ZN(new_n12455_));
  NAND2_X1   g11435(.A1(new_n12452_), .A2(new_n12455_), .ZN(new_n12456_));
  NOR2_X1    g11436(.A1(new_n12456_), .A2(new_n12443_), .ZN(new_n12457_));
  INV_X1     g11437(.I(new_n12443_), .ZN(new_n12458_));
  OAI21_X1   g11438(.A1(new_n12450_), .A2(new_n12447_), .B(new_n10762_), .ZN(new_n12459_));
  NAND3_X1   g11439(.A1(new_n12444_), .A2(new_n12445_), .A3(new_n10806_), .ZN(new_n12460_));
  NAND2_X1   g11440(.A1(new_n12459_), .A2(new_n12460_), .ZN(new_n12461_));
  NAND2_X1   g11441(.A1(new_n10751_), .A2(new_n10806_), .ZN(new_n12462_));
  NAND2_X1   g11442(.A1(new_n10762_), .A2(new_n10800_), .ZN(new_n12463_));
  AOI21_X1   g11443(.A1(new_n12462_), .A2(new_n12463_), .B(new_n10765_), .ZN(new_n12464_));
  NOR2_X1    g11444(.A1(new_n12461_), .A2(new_n12464_), .ZN(new_n12465_));
  NOR2_X1    g11445(.A1(new_n12465_), .A2(new_n12458_), .ZN(new_n12466_));
  OAI21_X1   g11446(.A1(new_n12457_), .A2(new_n12466_), .B(new_n12442_), .ZN(new_n12467_));
  OAI21_X1   g11447(.A1(new_n12440_), .A2(new_n12439_), .B(new_n10823_), .ZN(new_n12468_));
  NAND3_X1   g11448(.A1(new_n12436_), .A2(new_n12437_), .A3(new_n10787_), .ZN(new_n12469_));
  NAND2_X1   g11449(.A1(new_n12468_), .A2(new_n12469_), .ZN(new_n12470_));
  AOI22_X1   g11450(.A1(new_n10771_), .A2(new_n10776_), .B1(new_n10782_), .B2(new_n10786_), .ZN(new_n12471_));
  NOR4_X1    g11451(.A1(new_n10813_), .A2(new_n10815_), .A3(new_n10822_), .A4(new_n10819_), .ZN(new_n12472_));
  NOR2_X1    g11452(.A1(new_n12472_), .A2(new_n12471_), .ZN(new_n12473_));
  NOR3_X1    g11453(.A1(new_n10816_), .A2(new_n10823_), .A3(new_n10824_), .ZN(new_n12474_));
  NOR3_X1    g11454(.A1(new_n12473_), .A2(new_n10810_), .A3(new_n12474_), .ZN(new_n12475_));
  NAND4_X1   g11455(.A1(new_n12470_), .A2(new_n12475_), .A3(new_n12461_), .A4(new_n12455_), .ZN(new_n12476_));
  AOI21_X1   g11456(.A1(new_n12476_), .A2(new_n12456_), .B(new_n12458_), .ZN(new_n12477_));
  NOR4_X1    g11457(.A1(new_n10794_), .A2(new_n10826_), .A3(new_n10879_), .A4(new_n10910_), .ZN(new_n12478_));
  NAND2_X1   g11458(.A1(new_n10852_), .A2(new_n10909_), .ZN(new_n12479_));
  NOR3_X1    g11459(.A1(new_n10836_), .A2(new_n10851_), .A3(new_n10832_), .ZN(new_n12480_));
  INV_X1     g11460(.I(new_n10892_), .ZN(new_n12481_));
  INV_X1     g11461(.I(new_n10893_), .ZN(new_n12482_));
  AOI22_X1   g11462(.A1(new_n12481_), .A2(new_n12482_), .B1(new_n10882_), .B2(new_n10884_), .ZN(new_n12483_));
  OAI21_X1   g11463(.A1(new_n12483_), .A2(new_n12480_), .B(new_n10848_), .ZN(new_n12484_));
  NAND3_X1   g11464(.A1(new_n10894_), .A2(new_n10882_), .A3(new_n10884_), .ZN(new_n12485_));
  OAI21_X1   g11465(.A1(new_n10832_), .A2(new_n10836_), .B(new_n10851_), .ZN(new_n12486_));
  NAND3_X1   g11466(.A1(new_n12485_), .A2(new_n12486_), .A3(new_n10891_), .ZN(new_n12487_));
  NOR2_X1    g11467(.A1(new_n10848_), .A2(new_n10885_), .ZN(new_n12488_));
  NOR2_X1    g11468(.A1(new_n10837_), .A2(new_n10891_), .ZN(new_n12489_));
  OAI21_X1   g11469(.A1(new_n12488_), .A2(new_n12489_), .B(new_n10894_), .ZN(new_n12490_));
  NAND4_X1   g11470(.A1(new_n12490_), .A2(new_n12479_), .A3(new_n12484_), .A4(new_n12487_), .ZN(new_n12491_));
  NOR2_X1    g11471(.A1(new_n10863_), .A2(new_n10876_), .ZN(new_n12492_));
  OAI21_X1   g11472(.A1(new_n10898_), .A2(new_n10900_), .B(new_n10876_), .ZN(new_n12493_));
  INV_X1     g11473(.I(new_n12493_), .ZN(new_n12494_));
  OAI21_X1   g11474(.A1(new_n12494_), .A2(new_n12492_), .B(new_n10908_), .ZN(new_n12495_));
  NAND2_X1   g11475(.A1(new_n10901_), .A2(new_n10877_), .ZN(new_n12496_));
  NAND3_X1   g11476(.A1(new_n12496_), .A2(new_n10873_), .A3(new_n12493_), .ZN(new_n12497_));
  NAND2_X1   g11477(.A1(new_n12495_), .A2(new_n12497_), .ZN(new_n12498_));
  OAI22_X1   g11478(.A1(new_n10898_), .A2(new_n10900_), .B1(new_n10904_), .B2(new_n10907_), .ZN(new_n12499_));
  NAND4_X1   g11479(.A1(new_n10857_), .A2(new_n10868_), .A3(new_n10862_), .A4(new_n10872_), .ZN(new_n12500_));
  NAND2_X1   g11480(.A1(new_n12499_), .A2(new_n12500_), .ZN(new_n12501_));
  AOI21_X1   g11481(.A1(new_n10857_), .A2(new_n10862_), .B(new_n10876_), .ZN(new_n12502_));
  NAND4_X1   g11482(.A1(new_n12501_), .A2(new_n10885_), .A3(new_n10891_), .A4(new_n10894_), .ZN(new_n12505_));
  NAND4_X1   g11483(.A1(new_n12478_), .A2(new_n12491_), .A3(new_n12498_), .A4(new_n12505_), .ZN(new_n12506_));
  NOR2_X1    g11484(.A1(new_n12477_), .A2(new_n12506_), .ZN(new_n12507_));
  OAI22_X1   g11485(.A1(new_n10813_), .A2(new_n10815_), .B1(new_n10822_), .B2(new_n10819_), .ZN(new_n12508_));
  NAND4_X1   g11486(.A1(new_n10771_), .A2(new_n10782_), .A3(new_n10776_), .A4(new_n10786_), .ZN(new_n12509_));
  AOI21_X1   g11487(.A1(new_n10771_), .A2(new_n10776_), .B(new_n10824_), .ZN(new_n12510_));
  AOI22_X1   g11488(.A1(new_n12508_), .A2(new_n12509_), .B1(new_n12510_), .B2(new_n10787_), .ZN(new_n12511_));
  NAND4_X1   g11489(.A1(new_n12511_), .A2(new_n10800_), .A3(new_n10806_), .A4(new_n10809_), .ZN(new_n12512_));
  NOR2_X1    g11490(.A1(new_n12512_), .A2(new_n12442_), .ZN(new_n12513_));
  OAI21_X1   g11491(.A1(new_n12513_), .A2(new_n12465_), .B(new_n12443_), .ZN(new_n12514_));
  NOR2_X1    g11492(.A1(new_n10878_), .A2(new_n10895_), .ZN(new_n12515_));
  AOI21_X1   g11493(.A1(new_n12485_), .A2(new_n12486_), .B(new_n10891_), .ZN(new_n12516_));
  NOR3_X1    g11494(.A1(new_n12483_), .A2(new_n12480_), .A3(new_n10848_), .ZN(new_n12517_));
  NAND2_X1   g11495(.A1(new_n10837_), .A2(new_n10891_), .ZN(new_n12518_));
  NAND2_X1   g11496(.A1(new_n10848_), .A2(new_n10885_), .ZN(new_n12519_));
  AOI21_X1   g11497(.A1(new_n12518_), .A2(new_n12519_), .B(new_n10851_), .ZN(new_n12520_));
  NOR4_X1    g11498(.A1(new_n12520_), .A2(new_n12515_), .A3(new_n12516_), .A4(new_n12517_), .ZN(new_n12521_));
  AOI21_X1   g11499(.A1(new_n12496_), .A2(new_n12493_), .B(new_n10873_), .ZN(new_n12522_));
  NOR3_X1    g11500(.A1(new_n12494_), .A2(new_n12492_), .A3(new_n10908_), .ZN(new_n12523_));
  NOR2_X1    g11501(.A1(new_n12523_), .A2(new_n12522_), .ZN(new_n12524_));
  INV_X1     g11502(.I(new_n12505_), .ZN(new_n12525_));
  NOR4_X1    g11503(.A1(new_n10916_), .A2(new_n12521_), .A3(new_n12525_), .A4(new_n12524_), .ZN(new_n12526_));
  NOR2_X1    g11504(.A1(new_n12514_), .A2(new_n12526_), .ZN(new_n12527_));
  OAI21_X1   g11505(.A1(new_n12507_), .A2(new_n12527_), .B(new_n12467_), .ZN(new_n12528_));
  NAND2_X1   g11506(.A1(new_n12465_), .A2(new_n12458_), .ZN(new_n12529_));
  NAND2_X1   g11507(.A1(new_n12456_), .A2(new_n12443_), .ZN(new_n12530_));
  AOI21_X1   g11508(.A1(new_n12530_), .A2(new_n12529_), .B(new_n12470_), .ZN(new_n12531_));
  NAND2_X1   g11509(.A1(new_n12514_), .A2(new_n12526_), .ZN(new_n12532_));
  OAI22_X1   g11510(.A1(new_n12512_), .A2(new_n12442_), .B1(new_n12461_), .B2(new_n12464_), .ZN(new_n12533_));
  NAND3_X1   g11511(.A1(new_n12506_), .A2(new_n12443_), .A3(new_n12533_), .ZN(new_n12534_));
  NAND3_X1   g11512(.A1(new_n12532_), .A2(new_n12534_), .A3(new_n12531_), .ZN(new_n12535_));
  AOI21_X1   g11513(.A1(new_n12528_), .A2(new_n12535_), .B(new_n10920_), .ZN(new_n12536_));
  NAND2_X1   g11514(.A1(new_n12536_), .A2(new_n12435_), .ZN(new_n12537_));
  INV_X1     g11515(.I(new_n12394_), .ZN(new_n12538_));
  INV_X1     g11516(.I(new_n12432_), .ZN(new_n12539_));
  AOI21_X1   g11517(.A1(new_n12539_), .A2(new_n12433_), .B(new_n12538_), .ZN(new_n12540_));
  NAND2_X1   g11518(.A1(new_n12536_), .A2(new_n12540_), .ZN(new_n12541_));
  AOI21_X1   g11519(.A1(new_n12537_), .A2(new_n12541_), .B(new_n12358_), .ZN(new_n12542_));
  INV_X1     g11520(.I(new_n12542_), .ZN(new_n12543_));
  NOR2_X1    g11521(.A1(new_n12543_), .A2(new_n12356_), .ZN(new_n12544_));
  NOR3_X1    g11522(.A1(new_n12543_), .A2(new_n12260_), .A3(new_n12355_), .ZN(new_n12545_));
  NOR2_X1    g11523(.A1(new_n12545_), .A2(new_n12544_), .ZN(new_n12546_));
  INV_X1     g11524(.I(new_n12546_), .ZN(new_n12547_));
  NAND3_X1   g11525(.A1(new_n12547_), .A2(new_n10924_), .A3(new_n12174_), .ZN(new_n12548_));
  INV_X1     g11526(.I(new_n12174_), .ZN(new_n12549_));
  NAND3_X1   g11527(.A1(new_n12547_), .A2(new_n10924_), .A3(new_n12549_), .ZN(new_n12550_));
  NAND2_X1   g11528(.A1(new_n12548_), .A2(new_n12550_), .ZN(new_n12551_));
  NAND2_X1   g11529(.A1(new_n12551_), .A2(new_n10926_), .ZN(new_n12552_));
  NAND2_X1   g11530(.A1(new_n12552_), .A2(new_n11729_), .ZN(new_n12553_));
  INV_X1     g11531(.I(new_n12553_), .ZN(new_n12554_));
  NAND2_X1   g11532(.A1(new_n10932_), .A2(new_n8199_), .ZN(new_n12555_));
  AOI21_X1   g11533(.A1(new_n12554_), .A2(new_n12555_), .B(new_n10933_), .ZN(new_n12556_));
  OAI21_X1   g11534(.A1(new_n12551_), .A2(new_n10926_), .B(new_n11729_), .ZN(new_n12557_));
  NAND2_X1   g11535(.A1(new_n12557_), .A2(new_n12552_), .ZN(new_n12558_));
  OAI21_X1   g11536(.A1(new_n12547_), .A2(new_n10924_), .B(new_n12549_), .ZN(new_n12559_));
  INV_X1     g11537(.I(new_n12559_), .ZN(new_n12560_));
  NAND3_X1   g11538(.A1(new_n12358_), .A2(new_n12541_), .A3(new_n12537_), .ZN(new_n12561_));
  NAND2_X1   g11539(.A1(new_n12561_), .A2(new_n12356_), .ZN(new_n12562_));
  NAND2_X1   g11540(.A1(new_n12562_), .A2(new_n12543_), .ZN(new_n12563_));
  AOI21_X1   g11541(.A1(new_n12532_), .A2(new_n12534_), .B(new_n12531_), .ZN(new_n12564_));
  NOR3_X1    g11542(.A1(new_n12507_), .A2(new_n12527_), .A3(new_n12467_), .ZN(new_n12565_));
  OAI21_X1   g11543(.A1(new_n12565_), .A2(new_n12564_), .B(new_n10919_), .ZN(new_n12566_));
  NOR3_X1    g11544(.A1(new_n12565_), .A2(new_n12564_), .A3(new_n10919_), .ZN(new_n12567_));
  OAI21_X1   g11545(.A1(new_n12435_), .A2(new_n12567_), .B(new_n12566_), .ZN(new_n12568_));
  NOR3_X1    g11546(.A1(new_n12521_), .A2(new_n12525_), .A3(new_n12524_), .ZN(new_n12569_));
  NOR2_X1    g11547(.A1(new_n12569_), .A2(new_n12478_), .ZN(new_n12570_));
  NAND4_X1   g11548(.A1(new_n12513_), .A2(new_n12442_), .A3(new_n12443_), .A4(new_n12456_), .ZN(new_n12571_));
  OAI21_X1   g11549(.A1(new_n12570_), .A2(new_n12571_), .B(new_n12506_), .ZN(new_n12572_));
  AOI22_X1   g11550(.A1(new_n12499_), .A2(new_n12500_), .B1(new_n12502_), .B2(new_n10873_), .ZN(new_n12573_));
  NAND4_X1   g11551(.A1(new_n12573_), .A2(new_n10885_), .A3(new_n10891_), .A4(new_n10894_), .ZN(new_n12574_));
  INV_X1     g11552(.I(new_n12574_), .ZN(new_n12575_));
  NAND2_X1   g11553(.A1(new_n10892_), .A2(new_n10893_), .ZN(new_n12576_));
  NAND3_X1   g11554(.A1(new_n10885_), .A2(new_n10891_), .A3(new_n12576_), .ZN(new_n12577_));
  NAND2_X1   g11555(.A1(new_n12577_), .A2(new_n10851_), .ZN(new_n12578_));
  NOR4_X1    g11556(.A1(new_n10874_), .A2(new_n10875_), .A3(new_n10861_), .A4(new_n10871_), .ZN(new_n12579_));
  OAI21_X1   g11557(.A1(new_n12499_), .A2(new_n12579_), .B(new_n10876_), .ZN(new_n12580_));
  XOR2_X1    g11558(.A1(new_n12578_), .A2(new_n12580_), .Z(new_n12581_));
  NAND3_X1   g11559(.A1(new_n12490_), .A2(new_n12484_), .A3(new_n12487_), .ZN(new_n12582_));
  AOI21_X1   g11560(.A1(new_n12582_), .A2(new_n12479_), .B(new_n12524_), .ZN(new_n12583_));
  OAI21_X1   g11561(.A1(new_n12583_), .A2(new_n12575_), .B(new_n12581_), .ZN(new_n12584_));
  NOR2_X1    g11562(.A1(new_n10751_), .A2(new_n10762_), .ZN(new_n12585_));
  NAND2_X1   g11563(.A1(new_n10807_), .A2(new_n10808_), .ZN(new_n12586_));
  AOI21_X1   g11564(.A1(new_n12585_), .A2(new_n12586_), .B(new_n10809_), .ZN(new_n12587_));
  NAND2_X1   g11565(.A1(new_n10789_), .A2(new_n10791_), .ZN(new_n12588_));
  NAND3_X1   g11566(.A1(new_n10777_), .A2(new_n10787_), .A3(new_n12588_), .ZN(new_n12589_));
  NAND2_X1   g11567(.A1(new_n12589_), .A2(new_n10824_), .ZN(new_n12590_));
  XOR2_X1    g11568(.A1(new_n12587_), .A2(new_n12590_), .Z(new_n12591_));
  OAI21_X1   g11569(.A1(new_n12465_), .A2(new_n12443_), .B(new_n12470_), .ZN(new_n12592_));
  AOI21_X1   g11570(.A1(new_n12592_), .A2(new_n12512_), .B(new_n12591_), .ZN(new_n12593_));
  NOR2_X1    g11571(.A1(new_n12593_), .A2(new_n12584_), .ZN(new_n12594_));
  XNOR2_X1   g11572(.A1(new_n12578_), .A2(new_n12580_), .ZN(new_n12595_));
  NOR3_X1    g11573(.A1(new_n12520_), .A2(new_n12516_), .A3(new_n12517_), .ZN(new_n12596_));
  OAI21_X1   g11574(.A1(new_n12596_), .A2(new_n12515_), .B(new_n12498_), .ZN(new_n12597_));
  AOI21_X1   g11575(.A1(new_n12597_), .A2(new_n12574_), .B(new_n12595_), .ZN(new_n12598_));
  INV_X1     g11576(.I(new_n12512_), .ZN(new_n12599_));
  NAND2_X1   g11577(.A1(new_n12587_), .A2(new_n12590_), .ZN(new_n12600_));
  NAND3_X1   g11578(.A1(new_n10800_), .A2(new_n10806_), .A3(new_n12586_), .ZN(new_n12601_));
  NAND2_X1   g11579(.A1(new_n12601_), .A2(new_n10765_), .ZN(new_n12602_));
  NAND3_X1   g11580(.A1(new_n12602_), .A2(new_n10824_), .A3(new_n12589_), .ZN(new_n12603_));
  NAND2_X1   g11581(.A1(new_n12603_), .A2(new_n12600_), .ZN(new_n12604_));
  AOI21_X1   g11582(.A1(new_n12452_), .A2(new_n12455_), .B(new_n12443_), .ZN(new_n12605_));
  NOR2_X1    g11583(.A1(new_n12605_), .A2(new_n12442_), .ZN(new_n12606_));
  OAI21_X1   g11584(.A1(new_n12606_), .A2(new_n12599_), .B(new_n12604_), .ZN(new_n12607_));
  NOR2_X1    g11585(.A1(new_n12607_), .A2(new_n12598_), .ZN(new_n12608_));
  OAI21_X1   g11586(.A1(new_n12608_), .A2(new_n12594_), .B(new_n12572_), .ZN(new_n12609_));
  NAND3_X1   g11587(.A1(new_n12491_), .A2(new_n12498_), .A3(new_n12505_), .ZN(new_n12610_));
  NAND2_X1   g11588(.A1(new_n12610_), .A2(new_n10916_), .ZN(new_n12611_));
  NOR4_X1    g11589(.A1(new_n12476_), .A2(new_n12470_), .A3(new_n12458_), .A4(new_n12465_), .ZN(new_n12612_));
  AOI21_X1   g11590(.A1(new_n12611_), .A2(new_n12612_), .B(new_n12526_), .ZN(new_n12613_));
  NOR2_X1    g11591(.A1(new_n12593_), .A2(new_n12598_), .ZN(new_n12614_));
  NOR2_X1    g11592(.A1(new_n12607_), .A2(new_n12584_), .ZN(new_n12615_));
  OAI21_X1   g11593(.A1(new_n12614_), .A2(new_n12615_), .B(new_n12613_), .ZN(new_n12616_));
  NAND2_X1   g11594(.A1(new_n12609_), .A2(new_n12616_), .ZN(new_n12617_));
  NOR4_X1    g11595(.A1(new_n10739_), .A2(new_n12415_), .A3(new_n12422_), .A4(new_n12429_), .ZN(new_n12618_));
  INV_X1     g11596(.I(new_n12403_), .ZN(new_n12619_));
  OAI21_X1   g11597(.A1(new_n12410_), .A2(new_n12407_), .B(new_n10719_), .ZN(new_n12620_));
  NAND3_X1   g11598(.A1(new_n12404_), .A2(new_n12405_), .A3(new_n10673_), .ZN(new_n12621_));
  NOR2_X1    g11599(.A1(new_n10719_), .A2(new_n10663_), .ZN(new_n12622_));
  NOR2_X1    g11600(.A1(new_n10712_), .A2(new_n10673_), .ZN(new_n12623_));
  OAI21_X1   g11601(.A1(new_n12622_), .A2(new_n12623_), .B(new_n10678_), .ZN(new_n12624_));
  NAND3_X1   g11602(.A1(new_n12624_), .A2(new_n12620_), .A3(new_n12621_), .ZN(new_n12625_));
  OAI21_X1   g11603(.A1(new_n12420_), .A2(new_n12419_), .B(new_n10701_), .ZN(new_n12626_));
  NAND3_X1   g11604(.A1(new_n12416_), .A2(new_n10733_), .A3(new_n12417_), .ZN(new_n12627_));
  NAND2_X1   g11605(.A1(new_n12626_), .A2(new_n12627_), .ZN(new_n12628_));
  OAI22_X1   g11606(.A1(new_n10685_), .A2(new_n10689_), .B1(new_n10700_), .B2(new_n10696_), .ZN(new_n12629_));
  NAND4_X1   g11607(.A1(new_n10724_), .A2(new_n10726_), .A3(new_n10730_), .A4(new_n10732_), .ZN(new_n12630_));
  AOI21_X1   g11608(.A1(new_n10724_), .A2(new_n10726_), .B(new_n10704_), .ZN(new_n12631_));
  AOI22_X1   g11609(.A1(new_n12629_), .A2(new_n12630_), .B1(new_n10733_), .B2(new_n12631_), .ZN(new_n12632_));
  NAND4_X1   g11610(.A1(new_n12632_), .A2(new_n10663_), .A3(new_n10673_), .A4(new_n10678_), .ZN(new_n12633_));
  NAND4_X1   g11611(.A1(new_n12625_), .A2(new_n12633_), .A3(new_n12628_), .A4(new_n12619_), .ZN(new_n12634_));
  NAND2_X1   g11612(.A1(new_n12634_), .A2(new_n10739_), .ZN(new_n12635_));
  NOR4_X1    g11613(.A1(new_n12393_), .A2(new_n12360_), .A3(new_n12398_), .A4(new_n12392_), .ZN(new_n12636_));
  AOI21_X1   g11614(.A1(new_n12635_), .A2(new_n12636_), .B(new_n12618_), .ZN(new_n12637_));
  NAND2_X1   g11615(.A1(new_n10675_), .A2(new_n10677_), .ZN(new_n12638_));
  NAND3_X1   g11616(.A1(new_n10663_), .A2(new_n10673_), .A3(new_n12638_), .ZN(new_n12639_));
  NAND2_X1   g11617(.A1(new_n12639_), .A2(new_n10720_), .ZN(new_n12640_));
  NOR3_X1    g11618(.A1(new_n12426_), .A2(new_n10687_), .A3(new_n10702_), .ZN(new_n12641_));
  OAI21_X1   g11619(.A1(new_n12629_), .A2(new_n12641_), .B(new_n10704_), .ZN(new_n12642_));
  XNOR2_X1   g11620(.A1(new_n12640_), .A2(new_n12642_), .ZN(new_n12643_));
  NOR3_X1    g11621(.A1(new_n12414_), .A2(new_n12406_), .A3(new_n12411_), .ZN(new_n12644_));
  OAI21_X1   g11622(.A1(new_n12644_), .A2(new_n12403_), .B(new_n12628_), .ZN(new_n12645_));
  AOI21_X1   g11623(.A1(new_n12645_), .A2(new_n12633_), .B(new_n12643_), .ZN(new_n12646_));
  OAI22_X1   g11624(.A1(new_n10611_), .A2(new_n10615_), .B1(new_n10601_), .B2(new_n10604_), .ZN(new_n12647_));
  NAND4_X1   g11625(.A1(new_n10639_), .A2(new_n10645_), .A3(new_n10647_), .A4(new_n10641_), .ZN(new_n12648_));
  AOI21_X1   g11626(.A1(new_n10639_), .A2(new_n10641_), .B(new_n10620_), .ZN(new_n12649_));
  AOI22_X1   g11627(.A1(new_n12647_), .A2(new_n12648_), .B1(new_n12649_), .B2(new_n10648_), .ZN(new_n12650_));
  NAND4_X1   g11628(.A1(new_n12650_), .A2(new_n10578_), .A3(new_n10589_), .A4(new_n10594_), .ZN(new_n12651_));
  INV_X1     g11629(.I(new_n12651_), .ZN(new_n12652_));
  NAND2_X1   g11630(.A1(new_n10591_), .A2(new_n10593_), .ZN(new_n12653_));
  NAND3_X1   g11631(.A1(new_n10578_), .A2(new_n10589_), .A3(new_n12653_), .ZN(new_n12654_));
  NAND2_X1   g11632(.A1(new_n12654_), .A2(new_n10635_), .ZN(new_n12655_));
  NOR2_X1    g11633(.A1(new_n12384_), .A2(new_n12386_), .ZN(new_n12656_));
  OAI21_X1   g11634(.A1(new_n12647_), .A2(new_n12656_), .B(new_n10620_), .ZN(new_n12657_));
  XOR2_X1    g11635(.A1(new_n12655_), .A2(new_n12657_), .Z(new_n12658_));
  INV_X1     g11636(.I(new_n12392_), .ZN(new_n12659_));
  AOI21_X1   g11637(.A1(new_n12369_), .A2(new_n12372_), .B(new_n12359_), .ZN(new_n12660_));
  NOR2_X1    g11638(.A1(new_n12660_), .A2(new_n12659_), .ZN(new_n12661_));
  OAI21_X1   g11639(.A1(new_n12661_), .A2(new_n12652_), .B(new_n12658_), .ZN(new_n12662_));
  NAND2_X1   g11640(.A1(new_n12662_), .A2(new_n12646_), .ZN(new_n12663_));
  OAI22_X1   g11641(.A1(new_n12423_), .A2(new_n12424_), .B1(new_n12427_), .B2(new_n10701_), .ZN(new_n12664_));
  NOR4_X1    g11642(.A1(new_n12664_), .A2(new_n10712_), .A3(new_n10719_), .A4(new_n10720_), .ZN(new_n12665_));
  XOR2_X1    g11643(.A1(new_n12640_), .A2(new_n12642_), .Z(new_n12666_));
  AOI21_X1   g11644(.A1(new_n12625_), .A2(new_n12619_), .B(new_n12422_), .ZN(new_n12667_));
  OAI21_X1   g11645(.A1(new_n12667_), .A2(new_n12665_), .B(new_n12666_), .ZN(new_n12668_));
  INV_X1     g11646(.I(new_n12657_), .ZN(new_n12669_));
  NOR2_X1    g11647(.A1(new_n12669_), .A2(new_n12655_), .ZN(new_n12670_));
  NOR2_X1    g11648(.A1(new_n10628_), .A2(new_n10634_), .ZN(new_n12671_));
  AOI21_X1   g11649(.A1(new_n12671_), .A2(new_n12653_), .B(new_n10594_), .ZN(new_n12672_));
  NOR2_X1    g11650(.A1(new_n12672_), .A2(new_n12657_), .ZN(new_n12673_));
  NOR2_X1    g11651(.A1(new_n12670_), .A2(new_n12673_), .ZN(new_n12674_));
  OAI21_X1   g11652(.A1(new_n12398_), .A2(new_n12359_), .B(new_n12392_), .ZN(new_n12675_));
  AOI21_X1   g11653(.A1(new_n12675_), .A2(new_n12651_), .B(new_n12674_), .ZN(new_n12676_));
  NAND2_X1   g11654(.A1(new_n12676_), .A2(new_n12668_), .ZN(new_n12677_));
  AOI21_X1   g11655(.A1(new_n12663_), .A2(new_n12677_), .B(new_n12637_), .ZN(new_n12678_));
  NOR2_X1    g11656(.A1(new_n12430_), .A2(new_n12402_), .ZN(new_n12679_));
  NOR2_X1    g11657(.A1(new_n12659_), .A2(new_n12651_), .ZN(new_n12680_));
  NAND4_X1   g11658(.A1(new_n12680_), .A2(new_n12359_), .A3(new_n12373_), .A4(new_n12659_), .ZN(new_n12681_));
  OAI21_X1   g11659(.A1(new_n12679_), .A2(new_n12681_), .B(new_n12431_), .ZN(new_n12682_));
  NAND2_X1   g11660(.A1(new_n12662_), .A2(new_n12668_), .ZN(new_n12683_));
  NAND2_X1   g11661(.A1(new_n12646_), .A2(new_n12676_), .ZN(new_n12684_));
  AOI21_X1   g11662(.A1(new_n12684_), .A2(new_n12683_), .B(new_n12682_), .ZN(new_n12685_));
  NOR2_X1    g11663(.A1(new_n12685_), .A2(new_n12678_), .ZN(new_n12686_));
  NOR2_X1    g11664(.A1(new_n12686_), .A2(new_n12617_), .ZN(new_n12687_));
  NAND2_X1   g11665(.A1(new_n12607_), .A2(new_n12598_), .ZN(new_n12688_));
  NAND2_X1   g11666(.A1(new_n12593_), .A2(new_n12584_), .ZN(new_n12689_));
  AOI21_X1   g11667(.A1(new_n12688_), .A2(new_n12689_), .B(new_n12613_), .ZN(new_n12690_));
  NAND2_X1   g11668(.A1(new_n12607_), .A2(new_n12584_), .ZN(new_n12691_));
  NAND2_X1   g11669(.A1(new_n12593_), .A2(new_n12598_), .ZN(new_n12692_));
  AOI21_X1   g11670(.A1(new_n12692_), .A2(new_n12691_), .B(new_n12572_), .ZN(new_n12693_));
  NOR2_X1    g11671(.A1(new_n12693_), .A2(new_n12690_), .ZN(new_n12694_));
  NOR2_X1    g11672(.A1(new_n12676_), .A2(new_n12668_), .ZN(new_n12695_));
  NOR2_X1    g11673(.A1(new_n12662_), .A2(new_n12646_), .ZN(new_n12696_));
  OAI21_X1   g11674(.A1(new_n12695_), .A2(new_n12696_), .B(new_n12682_), .ZN(new_n12697_));
  NOR2_X1    g11675(.A1(new_n12646_), .A2(new_n12676_), .ZN(new_n12698_));
  NOR2_X1    g11676(.A1(new_n12662_), .A2(new_n12668_), .ZN(new_n12699_));
  OAI21_X1   g11677(.A1(new_n12698_), .A2(new_n12699_), .B(new_n12637_), .ZN(new_n12700_));
  NAND2_X1   g11678(.A1(new_n12697_), .A2(new_n12700_), .ZN(new_n12701_));
  NOR2_X1    g11679(.A1(new_n12701_), .A2(new_n12694_), .ZN(new_n12702_));
  OAI21_X1   g11680(.A1(new_n12702_), .A2(new_n12687_), .B(new_n12568_), .ZN(new_n12703_));
  NAND3_X1   g11681(.A1(new_n12528_), .A2(new_n12535_), .A3(new_n10920_), .ZN(new_n12704_));
  AOI21_X1   g11682(.A1(new_n12540_), .A2(new_n12704_), .B(new_n12536_), .ZN(new_n12705_));
  AOI22_X1   g11683(.A1(new_n12697_), .A2(new_n12700_), .B1(new_n12609_), .B2(new_n12616_), .ZN(new_n12706_));
  NOR4_X1    g11684(.A1(new_n12685_), .A2(new_n12690_), .A3(new_n12693_), .A4(new_n12678_), .ZN(new_n12707_));
  OAI21_X1   g11685(.A1(new_n12706_), .A2(new_n12707_), .B(new_n12705_), .ZN(new_n12708_));
  NAND2_X1   g11686(.A1(new_n12703_), .A2(new_n12708_), .ZN(new_n12709_));
  INV_X1     g11687(.I(new_n12217_), .ZN(new_n12710_));
  INV_X1     g11688(.I(new_n12257_), .ZN(new_n12711_));
  AOI21_X1   g11689(.A1(new_n12711_), .A2(new_n12258_), .B(new_n12710_), .ZN(new_n12712_));
  NAND3_X1   g11690(.A1(new_n12348_), .A2(new_n12354_), .A3(new_n10566_), .ZN(new_n12713_));
  AOI21_X1   g11691(.A1(new_n12712_), .A2(new_n12713_), .B(new_n12355_), .ZN(new_n12714_));
  NAND3_X1   g11692(.A1(new_n12311_), .A2(new_n12318_), .A3(new_n12325_), .ZN(new_n12715_));
  NAND2_X1   g11693(.A1(new_n12715_), .A2(new_n10562_), .ZN(new_n12716_));
  NOR4_X1    g11694(.A1(new_n12298_), .A2(new_n12292_), .A3(new_n12281_), .A4(new_n12286_), .ZN(new_n12717_));
  AOI21_X1   g11695(.A1(new_n12716_), .A2(new_n12717_), .B(new_n12346_), .ZN(new_n12718_));
  AOI22_X1   g11696(.A1(new_n12319_), .A2(new_n12320_), .B1(new_n12322_), .B2(new_n10520_), .ZN(new_n12719_));
  NAND4_X1   g11697(.A1(new_n12719_), .A2(new_n10532_), .A3(new_n10538_), .A4(new_n10541_), .ZN(new_n12720_));
  NAND2_X1   g11698(.A1(new_n10539_), .A2(new_n10540_), .ZN(new_n12721_));
  NAND3_X1   g11699(.A1(new_n10532_), .A2(new_n10538_), .A3(new_n12721_), .ZN(new_n12722_));
  NAND2_X1   g11700(.A1(new_n12722_), .A2(new_n10497_), .ZN(new_n12723_));
  OR4_X2     g11701(.A1(new_n10507_), .A2(new_n10521_), .A3(new_n10522_), .A4(new_n10518_), .Z(new_n12724_));
  NAND3_X1   g11702(.A1(new_n10509_), .A2(new_n10520_), .A3(new_n12724_), .ZN(new_n12725_));
  NAND2_X1   g11703(.A1(new_n12725_), .A2(new_n10523_), .ZN(new_n12726_));
  XNOR2_X1   g11704(.A1(new_n12726_), .A2(new_n12723_), .ZN(new_n12727_));
  NAND2_X1   g11705(.A1(new_n12304_), .A2(new_n12307_), .ZN(new_n12728_));
  OAI21_X1   g11706(.A1(new_n12728_), .A2(new_n12340_), .B(new_n12301_), .ZN(new_n12729_));
  NAND2_X1   g11707(.A1(new_n12729_), .A2(new_n12318_), .ZN(new_n12730_));
  AOI21_X1   g11708(.A1(new_n12730_), .A2(new_n12720_), .B(new_n12727_), .ZN(new_n12731_));
  INV_X1     g11709(.I(new_n12332_), .ZN(new_n12732_));
  NAND2_X1   g11710(.A1(new_n10454_), .A2(new_n10455_), .ZN(new_n12733_));
  NAND3_X1   g11711(.A1(new_n10453_), .A2(new_n10447_), .A3(new_n12733_), .ZN(new_n12734_));
  NAND2_X1   g11712(.A1(new_n12734_), .A2(new_n10411_), .ZN(new_n12735_));
  NOR4_X1    g11713(.A1(new_n10435_), .A2(new_n10437_), .A3(new_n10421_), .A4(new_n10432_), .ZN(new_n12736_));
  OAI21_X1   g11714(.A1(new_n12328_), .A2(new_n12736_), .B(new_n10470_), .ZN(new_n12737_));
  XOR2_X1    g11715(.A1(new_n12735_), .A2(new_n12737_), .Z(new_n12738_));
  AOI21_X1   g11716(.A1(new_n12279_), .A2(new_n12281_), .B(new_n12266_), .ZN(new_n12739_));
  OAI21_X1   g11717(.A1(new_n12739_), .A2(new_n12732_), .B(new_n12738_), .ZN(new_n12740_));
  NAND2_X1   g11718(.A1(new_n12731_), .A2(new_n12740_), .ZN(new_n12741_));
  INV_X1     g11719(.I(new_n12720_), .ZN(new_n12742_));
  XOR2_X1    g11720(.A1(new_n12726_), .A2(new_n12723_), .Z(new_n12743_));
  NAND3_X1   g11721(.A1(new_n12310_), .A2(new_n12304_), .A3(new_n12307_), .ZN(new_n12744_));
  AOI21_X1   g11722(.A1(new_n12744_), .A2(new_n12301_), .B(new_n12344_), .ZN(new_n12745_));
  OAI21_X1   g11723(.A1(new_n12742_), .A2(new_n12745_), .B(new_n12743_), .ZN(new_n12746_));
  NOR2_X1    g11724(.A1(new_n10397_), .A2(new_n10408_), .ZN(new_n12747_));
  AOI21_X1   g11725(.A1(new_n12747_), .A2(new_n12733_), .B(new_n10456_), .ZN(new_n12748_));
  XOR2_X1    g11726(.A1(new_n12748_), .A2(new_n12737_), .Z(new_n12749_));
  OAI21_X1   g11727(.A1(new_n12286_), .A2(new_n12267_), .B(new_n12292_), .ZN(new_n12750_));
  AOI21_X1   g11728(.A1(new_n12750_), .A2(new_n12332_), .B(new_n12749_), .ZN(new_n12751_));
  NAND2_X1   g11729(.A1(new_n12751_), .A2(new_n12746_), .ZN(new_n12752_));
  AOI21_X1   g11730(.A1(new_n12741_), .A2(new_n12752_), .B(new_n12718_), .ZN(new_n12753_));
  NOR3_X1    g11731(.A1(new_n12341_), .A2(new_n12345_), .A3(new_n12344_), .ZN(new_n12754_));
  NOR2_X1    g11732(.A1(new_n12754_), .A2(new_n12300_), .ZN(new_n12755_));
  NAND4_X1   g11733(.A1(new_n12333_), .A2(new_n12266_), .A3(new_n12267_), .A4(new_n12279_), .ZN(new_n12756_));
  OAI21_X1   g11734(.A1(new_n12755_), .A2(new_n12756_), .B(new_n12326_), .ZN(new_n12757_));
  NAND2_X1   g11735(.A1(new_n12746_), .A2(new_n12740_), .ZN(new_n12758_));
  NAND2_X1   g11736(.A1(new_n12731_), .A2(new_n12751_), .ZN(new_n12759_));
  AOI21_X1   g11737(.A1(new_n12759_), .A2(new_n12758_), .B(new_n12757_), .ZN(new_n12760_));
  NOR2_X1    g11738(.A1(new_n12760_), .A2(new_n12753_), .ZN(new_n12761_));
  NOR4_X1    g11739(.A1(new_n12238_), .A2(new_n12228_), .A3(new_n12235_), .A4(new_n12232_), .ZN(new_n12762_));
  AOI21_X1   g11740(.A1(new_n12244_), .A2(new_n12245_), .B(new_n10331_), .ZN(new_n12763_));
  NOR3_X1    g11741(.A1(new_n12242_), .A2(new_n12241_), .A3(new_n10363_), .ZN(new_n12764_));
  NOR2_X1    g11742(.A1(new_n12763_), .A2(new_n12764_), .ZN(new_n12765_));
  INV_X1     g11743(.I(new_n12255_), .ZN(new_n12766_));
  NOR3_X1    g11744(.A1(new_n12762_), .A2(new_n12766_), .A3(new_n12765_), .ZN(new_n12767_));
  NOR2_X1    g11745(.A1(new_n12767_), .A2(new_n12227_), .ZN(new_n12768_));
  AND2_X2    g11746(.A1(new_n12214_), .A2(new_n12211_), .Z(new_n12769_));
  OAI22_X1   g11747(.A1(new_n12191_), .A2(new_n12193_), .B1(new_n12198_), .B2(new_n12196_), .ZN(new_n12770_));
  NAND4_X1   g11748(.A1(new_n10258_), .A2(new_n10263_), .A3(new_n10269_), .A4(new_n10274_), .ZN(new_n12771_));
  AOI21_X1   g11749(.A1(new_n10258_), .A2(new_n10263_), .B(new_n10278_), .ZN(new_n12772_));
  AOI22_X1   g11750(.A1(new_n12770_), .A2(new_n12771_), .B1(new_n10275_), .B2(new_n12772_), .ZN(new_n12773_));
  NAND4_X1   g11751(.A1(new_n12773_), .A2(new_n10372_), .A3(new_n10378_), .A4(new_n10379_), .ZN(new_n12774_));
  NOR2_X1    g11752(.A1(new_n12769_), .A2(new_n12774_), .ZN(new_n12775_));
  NAND4_X1   g11753(.A1(new_n12775_), .A2(new_n12175_), .A3(new_n12186_), .A4(new_n12769_), .ZN(new_n12776_));
  OAI21_X1   g11754(.A1(new_n12768_), .A2(new_n12776_), .B(new_n12256_), .ZN(new_n12777_));
  AOI22_X1   g11755(.A1(new_n10314_), .A2(new_n10319_), .B1(new_n10325_), .B2(new_n10330_), .ZN(new_n12778_));
  NOR4_X1    g11756(.A1(new_n10354_), .A2(new_n10356_), .A3(new_n10362_), .A4(new_n10360_), .ZN(new_n12779_));
  OAI22_X1   g11757(.A1(new_n12778_), .A2(new_n12779_), .B1(new_n12253_), .B2(new_n10363_), .ZN(new_n12780_));
  NOR4_X1    g11758(.A1(new_n12780_), .A2(new_n10294_), .A3(new_n10305_), .A4(new_n10308_), .ZN(new_n12781_));
  OR4_X2     g11759(.A1(new_n10291_), .A2(new_n10306_), .A3(new_n10307_), .A4(new_n10302_), .Z(new_n12782_));
  NAND3_X1   g11760(.A1(new_n10343_), .A2(new_n10349_), .A3(new_n12782_), .ZN(new_n12783_));
  NAND2_X1   g11761(.A1(new_n12783_), .A2(new_n10308_), .ZN(new_n12784_));
  NOR2_X1    g11762(.A1(new_n10332_), .A2(new_n10318_), .ZN(new_n12785_));
  NAND2_X1   g11763(.A1(new_n12785_), .A2(new_n12251_), .ZN(new_n12786_));
  NAND3_X1   g11764(.A1(new_n10320_), .A2(new_n10331_), .A3(new_n12786_), .ZN(new_n12787_));
  NAND2_X1   g11765(.A1(new_n12787_), .A2(new_n10334_), .ZN(new_n12788_));
  XOR2_X1    g11766(.A1(new_n12784_), .A2(new_n12788_), .Z(new_n12789_));
  OAI21_X1   g11767(.A1(new_n12234_), .A2(new_n12233_), .B(new_n10305_), .ZN(new_n12790_));
  NAND3_X1   g11768(.A1(new_n12230_), .A2(new_n12231_), .A3(new_n10349_), .ZN(new_n12791_));
  NOR2_X1    g11769(.A1(new_n10305_), .A2(new_n10343_), .ZN(new_n12792_));
  NOR2_X1    g11770(.A1(new_n10294_), .A2(new_n10349_), .ZN(new_n12793_));
  OAI21_X1   g11771(.A1(new_n12792_), .A2(new_n12793_), .B(new_n10350_), .ZN(new_n12794_));
  NAND3_X1   g11772(.A1(new_n12794_), .A2(new_n12790_), .A3(new_n12791_), .ZN(new_n12795_));
  AOI21_X1   g11773(.A1(new_n12795_), .A2(new_n12229_), .B(new_n12765_), .ZN(new_n12796_));
  OAI21_X1   g11774(.A1(new_n12796_), .A2(new_n12781_), .B(new_n12789_), .ZN(new_n12797_));
  OR4_X2     g11775(.A1(new_n10235_), .A2(new_n10250_), .A3(new_n10251_), .A4(new_n10246_), .Z(new_n12798_));
  NAND3_X1   g11776(.A1(new_n10372_), .A2(new_n10378_), .A3(new_n12798_), .ZN(new_n12799_));
  NAND2_X1   g11777(.A1(new_n12799_), .A2(new_n10252_), .ZN(new_n12800_));
  NOR2_X1    g11778(.A1(new_n12207_), .A2(new_n12209_), .ZN(new_n12801_));
  OAI21_X1   g11779(.A1(new_n12770_), .A2(new_n12801_), .B(new_n10278_), .ZN(new_n12802_));
  INV_X1     g11780(.I(new_n12802_), .ZN(new_n12803_));
  NOR2_X1    g11781(.A1(new_n12803_), .A2(new_n12800_), .ZN(new_n12804_));
  NOR2_X1    g11782(.A1(new_n10238_), .A2(new_n10249_), .ZN(new_n12805_));
  AOI21_X1   g11783(.A1(new_n12805_), .A2(new_n12798_), .B(new_n10379_), .ZN(new_n12806_));
  NOR2_X1    g11784(.A1(new_n12806_), .A2(new_n12802_), .ZN(new_n12807_));
  NOR2_X1    g11785(.A1(new_n12804_), .A2(new_n12807_), .ZN(new_n12808_));
  OAI21_X1   g11786(.A1(new_n12223_), .A2(new_n12175_), .B(new_n12215_), .ZN(new_n12809_));
  AOI21_X1   g11787(.A1(new_n12809_), .A2(new_n12774_), .B(new_n12808_), .ZN(new_n12810_));
  NOR2_X1    g11788(.A1(new_n12797_), .A2(new_n12810_), .ZN(new_n12811_));
  AOI21_X1   g11789(.A1(new_n10314_), .A2(new_n10319_), .B(new_n10334_), .ZN(new_n12812_));
  AOI22_X1   g11790(.A1(new_n12248_), .A2(new_n12249_), .B1(new_n10331_), .B2(new_n12812_), .ZN(new_n12813_));
  NAND4_X1   g11791(.A1(new_n12813_), .A2(new_n10343_), .A3(new_n10349_), .A4(new_n10350_), .ZN(new_n12814_));
  NOR2_X1    g11792(.A1(new_n10294_), .A2(new_n10305_), .ZN(new_n12815_));
  AOI21_X1   g11793(.A1(new_n12815_), .A2(new_n12782_), .B(new_n10350_), .ZN(new_n12816_));
  XOR2_X1    g11794(.A1(new_n12816_), .A2(new_n12788_), .Z(new_n12817_));
  OAI21_X1   g11795(.A1(new_n12239_), .A2(new_n12228_), .B(new_n12247_), .ZN(new_n12818_));
  AOI21_X1   g11796(.A1(new_n12818_), .A2(new_n12814_), .B(new_n12817_), .ZN(new_n12819_));
  INV_X1     g11797(.I(new_n12774_), .ZN(new_n12820_));
  XOR2_X1    g11798(.A1(new_n12800_), .A2(new_n12802_), .Z(new_n12821_));
  AOI21_X1   g11799(.A1(new_n12186_), .A2(new_n12176_), .B(new_n12769_), .ZN(new_n12822_));
  OAI21_X1   g11800(.A1(new_n12822_), .A2(new_n12820_), .B(new_n12821_), .ZN(new_n12823_));
  NOR2_X1    g11801(.A1(new_n12819_), .A2(new_n12823_), .ZN(new_n12824_));
  OAI21_X1   g11802(.A1(new_n12811_), .A2(new_n12824_), .B(new_n12777_), .ZN(new_n12825_));
  NOR4_X1    g11803(.A1(new_n10385_), .A2(new_n12762_), .A3(new_n12765_), .A4(new_n12766_), .ZN(new_n12826_));
  NAND4_X1   g11804(.A1(new_n12795_), .A2(new_n12814_), .A3(new_n12247_), .A4(new_n12229_), .ZN(new_n12827_));
  NAND2_X1   g11805(.A1(new_n12827_), .A2(new_n10385_), .ZN(new_n12828_));
  NOR4_X1    g11806(.A1(new_n12216_), .A2(new_n12176_), .A3(new_n12223_), .A4(new_n12215_), .ZN(new_n12829_));
  AOI21_X1   g11807(.A1(new_n12829_), .A2(new_n12828_), .B(new_n12826_), .ZN(new_n12830_));
  NOR2_X1    g11808(.A1(new_n12819_), .A2(new_n12810_), .ZN(new_n12831_));
  NOR2_X1    g11809(.A1(new_n12797_), .A2(new_n12823_), .ZN(new_n12832_));
  OAI21_X1   g11810(.A1(new_n12832_), .A2(new_n12831_), .B(new_n12830_), .ZN(new_n12833_));
  NAND2_X1   g11811(.A1(new_n12825_), .A2(new_n12833_), .ZN(new_n12834_));
  NAND2_X1   g11812(.A1(new_n12834_), .A2(new_n12761_), .ZN(new_n12835_));
  NOR2_X1    g11813(.A1(new_n12751_), .A2(new_n12746_), .ZN(new_n12836_));
  NOR2_X1    g11814(.A1(new_n12731_), .A2(new_n12740_), .ZN(new_n12837_));
  OAI21_X1   g11815(.A1(new_n12837_), .A2(new_n12836_), .B(new_n12757_), .ZN(new_n12838_));
  NOR2_X1    g11816(.A1(new_n12731_), .A2(new_n12751_), .ZN(new_n12839_));
  NOR2_X1    g11817(.A1(new_n12746_), .A2(new_n12740_), .ZN(new_n12840_));
  OAI21_X1   g11818(.A1(new_n12839_), .A2(new_n12840_), .B(new_n12718_), .ZN(new_n12841_));
  NAND2_X1   g11819(.A1(new_n12838_), .A2(new_n12841_), .ZN(new_n12842_));
  NAND2_X1   g11820(.A1(new_n12819_), .A2(new_n12823_), .ZN(new_n12843_));
  NAND2_X1   g11821(.A1(new_n12797_), .A2(new_n12810_), .ZN(new_n12844_));
  AOI21_X1   g11822(.A1(new_n12843_), .A2(new_n12844_), .B(new_n12830_), .ZN(new_n12845_));
  NAND2_X1   g11823(.A1(new_n12797_), .A2(new_n12823_), .ZN(new_n12846_));
  NAND2_X1   g11824(.A1(new_n12819_), .A2(new_n12810_), .ZN(new_n12847_));
  AOI21_X1   g11825(.A1(new_n12846_), .A2(new_n12847_), .B(new_n12777_), .ZN(new_n12848_));
  NOR2_X1    g11826(.A1(new_n12848_), .A2(new_n12845_), .ZN(new_n12849_));
  NAND2_X1   g11827(.A1(new_n12849_), .A2(new_n12842_), .ZN(new_n12850_));
  AOI21_X1   g11828(.A1(new_n12835_), .A2(new_n12850_), .B(new_n12714_), .ZN(new_n12851_));
  AOI21_X1   g11829(.A1(new_n12352_), .A2(new_n12353_), .B(new_n12351_), .ZN(new_n12852_));
  NOR3_X1    g11830(.A1(new_n12347_), .A2(new_n12327_), .A3(new_n12288_), .ZN(new_n12853_));
  OAI21_X1   g11831(.A1(new_n12852_), .A2(new_n12853_), .B(new_n10565_), .ZN(new_n12854_));
  NOR3_X1    g11832(.A1(new_n12852_), .A2(new_n12853_), .A3(new_n10565_), .ZN(new_n12855_));
  OAI21_X1   g11833(.A1(new_n12260_), .A2(new_n12855_), .B(new_n12854_), .ZN(new_n12856_));
  OAI22_X1   g11834(.A1(new_n12848_), .A2(new_n12845_), .B1(new_n12760_), .B2(new_n12753_), .ZN(new_n12857_));
  NAND4_X1   g11835(.A1(new_n12838_), .A2(new_n12825_), .A3(new_n12833_), .A4(new_n12841_), .ZN(new_n12858_));
  AOI21_X1   g11836(.A1(new_n12857_), .A2(new_n12858_), .B(new_n12856_), .ZN(new_n12859_));
  NOR2_X1    g11837(.A1(new_n12851_), .A2(new_n12859_), .ZN(new_n12860_));
  NOR2_X1    g11838(.A1(new_n12860_), .A2(new_n12709_), .ZN(new_n12861_));
  NAND2_X1   g11839(.A1(new_n12701_), .A2(new_n12694_), .ZN(new_n12862_));
  NAND2_X1   g11840(.A1(new_n12686_), .A2(new_n12617_), .ZN(new_n12863_));
  AOI21_X1   g11841(.A1(new_n12862_), .A2(new_n12863_), .B(new_n12705_), .ZN(new_n12864_));
  OAI22_X1   g11842(.A1(new_n12685_), .A2(new_n12678_), .B1(new_n12693_), .B2(new_n12690_), .ZN(new_n12865_));
  NAND4_X1   g11843(.A1(new_n12697_), .A2(new_n12609_), .A3(new_n12616_), .A4(new_n12700_), .ZN(new_n12866_));
  AOI21_X1   g11844(.A1(new_n12865_), .A2(new_n12866_), .B(new_n12568_), .ZN(new_n12867_));
  NOR2_X1    g11845(.A1(new_n12864_), .A2(new_n12867_), .ZN(new_n12868_));
  NOR2_X1    g11846(.A1(new_n12849_), .A2(new_n12842_), .ZN(new_n12869_));
  NOR2_X1    g11847(.A1(new_n12834_), .A2(new_n12761_), .ZN(new_n12870_));
  OAI21_X1   g11848(.A1(new_n12870_), .A2(new_n12869_), .B(new_n12856_), .ZN(new_n12871_));
  AOI22_X1   g11849(.A1(new_n12825_), .A2(new_n12833_), .B1(new_n12838_), .B2(new_n12841_), .ZN(new_n12872_));
  NOR4_X1    g11850(.A1(new_n12760_), .A2(new_n12848_), .A3(new_n12845_), .A4(new_n12753_), .ZN(new_n12873_));
  OAI21_X1   g11851(.A1(new_n12872_), .A2(new_n12873_), .B(new_n12714_), .ZN(new_n12874_));
  NAND2_X1   g11852(.A1(new_n12871_), .A2(new_n12874_), .ZN(new_n12875_));
  NOR2_X1    g11853(.A1(new_n12875_), .A2(new_n12868_), .ZN(new_n12876_));
  OAI21_X1   g11854(.A1(new_n12876_), .A2(new_n12861_), .B(new_n12563_), .ZN(new_n12877_));
  AOI21_X1   g11855(.A1(new_n12356_), .A2(new_n12561_), .B(new_n12542_), .ZN(new_n12878_));
  AOI22_X1   g11856(.A1(new_n12871_), .A2(new_n12874_), .B1(new_n12703_), .B2(new_n12708_), .ZN(new_n12879_));
  NOR4_X1    g11857(.A1(new_n12864_), .A2(new_n12851_), .A3(new_n12859_), .A4(new_n12867_), .ZN(new_n12880_));
  OAI21_X1   g11858(.A1(new_n12880_), .A2(new_n12879_), .B(new_n12878_), .ZN(new_n12881_));
  NAND2_X1   g11859(.A1(new_n12877_), .A2(new_n12881_), .ZN(new_n12882_));
  NAND3_X1   g11860(.A1(new_n10226_), .A2(new_n12170_), .A3(new_n12171_), .ZN(new_n12883_));
  NAND2_X1   g11861(.A1(new_n12883_), .A2(new_n11961_), .ZN(new_n12884_));
  NAND2_X1   g11862(.A1(new_n12884_), .A2(new_n12173_), .ZN(new_n12885_));
  AOI21_X1   g11863(.A1(new_n12166_), .A2(new_n12167_), .B(new_n12165_), .ZN(new_n12886_));
  NOR3_X1    g11864(.A1(new_n12091_), .A2(new_n12133_), .A3(new_n12162_), .ZN(new_n12887_));
  NOR2_X1    g11865(.A1(new_n12886_), .A2(new_n12887_), .ZN(new_n12888_));
  AOI21_X1   g11866(.A1(new_n12888_), .A2(new_n9902_), .B(new_n12056_), .ZN(new_n12889_));
  NOR3_X1    g11867(.A1(new_n12155_), .A2(new_n12160_), .A3(new_n12159_), .ZN(new_n12890_));
  NOR2_X1    g11868(.A1(new_n12890_), .A2(new_n9900_), .ZN(new_n12891_));
  NAND4_X1   g11869(.A1(new_n12145_), .A2(new_n12063_), .A3(new_n12064_), .A4(new_n12089_), .ZN(new_n12892_));
  OAI21_X1   g11870(.A1(new_n12891_), .A2(new_n12892_), .B(new_n12132_), .ZN(new_n12893_));
  AOI22_X1   g11871(.A1(new_n9882_), .A2(new_n9884_), .B1(new_n9888_), .B2(new_n9890_), .ZN(new_n12894_));
  NOR4_X1    g11872(.A1(new_n9844_), .A2(new_n9848_), .A3(new_n9859_), .A4(new_n9855_), .ZN(new_n12895_));
  OAI22_X1   g11873(.A1(new_n12894_), .A2(new_n12895_), .B1(new_n12129_), .B2(new_n9860_), .ZN(new_n12896_));
  NOR4_X1    g11874(.A1(new_n12896_), .A2(new_n9871_), .A3(new_n9877_), .A4(new_n9878_), .ZN(new_n12897_));
  NAND2_X1   g11875(.A1(new_n9834_), .A2(new_n9836_), .ZN(new_n12898_));
  NAND3_X1   g11876(.A1(new_n9821_), .A2(new_n9832_), .A3(new_n12898_), .ZN(new_n12899_));
  NAND2_X1   g11877(.A1(new_n12899_), .A2(new_n9878_), .ZN(new_n12900_));
  NOR3_X1    g11878(.A1(new_n12128_), .A2(new_n9846_), .A3(new_n9861_), .ZN(new_n12901_));
  OAI21_X1   g11879(.A1(new_n12124_), .A2(new_n12901_), .B(new_n9863_), .ZN(new_n12902_));
  XOR2_X1    g11880(.A1(new_n12900_), .A2(new_n12902_), .Z(new_n12903_));
  NAND3_X1   g11881(.A1(new_n12116_), .A2(new_n12149_), .A3(new_n12150_), .ZN(new_n12904_));
  AOI21_X1   g11882(.A1(new_n12904_), .A2(new_n12104_), .B(new_n12159_), .ZN(new_n12905_));
  OAI21_X1   g11883(.A1(new_n12905_), .A2(new_n12897_), .B(new_n12903_), .ZN(new_n12906_));
  NOR2_X1    g11884(.A1(new_n12086_), .A2(new_n12072_), .ZN(new_n12907_));
  NAND2_X1   g11885(.A1(new_n9763_), .A2(new_n9765_), .ZN(new_n12908_));
  AOI21_X1   g11886(.A1(new_n12907_), .A2(new_n12908_), .B(new_n9766_), .ZN(new_n12909_));
  NOR2_X1    g11887(.A1(new_n9790_), .A2(new_n9775_), .ZN(new_n12910_));
  NAND2_X1   g11888(.A1(new_n12910_), .A2(new_n12097_), .ZN(new_n12911_));
  NAND3_X1   g11889(.A1(new_n9801_), .A2(new_n9807_), .A3(new_n12911_), .ZN(new_n12912_));
  NAND2_X1   g11890(.A1(new_n12912_), .A2(new_n9792_), .ZN(new_n12913_));
  NAND2_X1   g11891(.A1(new_n12909_), .A2(new_n12913_), .ZN(new_n12914_));
  NAND3_X1   g11892(.A1(new_n9751_), .A2(new_n9761_), .A3(new_n12908_), .ZN(new_n12915_));
  NAND2_X1   g11893(.A1(new_n12915_), .A2(new_n12078_), .ZN(new_n12916_));
  NAND3_X1   g11894(.A1(new_n12916_), .A2(new_n9792_), .A3(new_n12912_), .ZN(new_n12917_));
  OAI21_X1   g11895(.A1(new_n12139_), .A2(new_n12064_), .B(new_n12094_), .ZN(new_n12918_));
  AOI22_X1   g11896(.A1(new_n12918_), .A2(new_n12144_), .B1(new_n12914_), .B2(new_n12917_), .ZN(new_n12919_));
  NOR2_X1    g11897(.A1(new_n12906_), .A2(new_n12919_), .ZN(new_n12920_));
  AOI21_X1   g11898(.A1(new_n9882_), .A2(new_n9884_), .B(new_n9863_), .ZN(new_n12921_));
  AOI22_X1   g11899(.A1(new_n12124_), .A2(new_n12125_), .B1(new_n9891_), .B2(new_n12921_), .ZN(new_n12922_));
  NAND4_X1   g11900(.A1(new_n12922_), .A2(new_n9821_), .A3(new_n9832_), .A4(new_n9837_), .ZN(new_n12923_));
  XNOR2_X1   g11901(.A1(new_n12900_), .A2(new_n12902_), .ZN(new_n12924_));
  NOR2_X1    g11902(.A1(new_n12151_), .A2(new_n12154_), .ZN(new_n12925_));
  OAI21_X1   g11903(.A1(new_n12925_), .A2(new_n12148_), .B(new_n12123_), .ZN(new_n12926_));
  AOI21_X1   g11904(.A1(new_n12926_), .A2(new_n12923_), .B(new_n12924_), .ZN(new_n12927_));
  NAND2_X1   g11905(.A1(new_n12914_), .A2(new_n12917_), .ZN(new_n12928_));
  AOI21_X1   g11906(.A1(new_n12089_), .A2(new_n12065_), .B(new_n12063_), .ZN(new_n12929_));
  OAI21_X1   g11907(.A1(new_n12929_), .A2(new_n12101_), .B(new_n12928_), .ZN(new_n12930_));
  NOR2_X1    g11908(.A1(new_n12927_), .A2(new_n12930_), .ZN(new_n12931_));
  OAI21_X1   g11909(.A1(new_n12931_), .A2(new_n12920_), .B(new_n12893_), .ZN(new_n12932_));
  NAND3_X1   g11910(.A1(new_n12117_), .A2(new_n12123_), .A3(new_n12131_), .ZN(new_n12933_));
  NAND2_X1   g11911(.A1(new_n12933_), .A2(new_n12147_), .ZN(new_n12934_));
  NOR4_X1    g11912(.A1(new_n12102_), .A2(new_n12094_), .A3(new_n12065_), .A4(new_n12139_), .ZN(new_n12935_));
  AOI21_X1   g11913(.A1(new_n12934_), .A2(new_n12935_), .B(new_n12161_), .ZN(new_n12936_));
  NOR2_X1    g11914(.A1(new_n12927_), .A2(new_n12919_), .ZN(new_n12937_));
  NOR2_X1    g11915(.A1(new_n12906_), .A2(new_n12930_), .ZN(new_n12938_));
  OAI21_X1   g11916(.A1(new_n12937_), .A2(new_n12938_), .B(new_n12936_), .ZN(new_n12939_));
  NAND2_X1   g11917(.A1(new_n12939_), .A2(new_n12932_), .ZN(new_n12940_));
  AOI21_X1   g11918(.A1(new_n12021_), .A2(new_n12022_), .B(new_n9572_), .ZN(new_n12941_));
  NOR3_X1    g11919(.A1(new_n12019_), .A2(new_n12018_), .A3(new_n9730_), .ZN(new_n12942_));
  NOR2_X1    g11920(.A1(new_n12942_), .A2(new_n12941_), .ZN(new_n12943_));
  NAND2_X1   g11921(.A1(new_n9719_), .A2(new_n9718_), .ZN(new_n12944_));
  XNOR2_X1   g11922(.A1(new_n9616_), .A2(new_n9619_), .ZN(new_n12945_));
  NOR2_X1    g11923(.A1(new_n9719_), .A2(new_n12945_), .ZN(new_n12946_));
  AOI21_X1   g11924(.A1(new_n9620_), .A2(new_n12009_), .B(new_n9614_), .ZN(new_n12947_));
  NOR2_X1    g11925(.A1(new_n12946_), .A2(new_n12947_), .ZN(new_n12948_));
  NOR4_X1    g11926(.A1(new_n12948_), .A2(new_n9736_), .A3(new_n12944_), .A4(new_n12045_), .ZN(new_n12949_));
  NOR4_X1    g11927(.A1(new_n12949_), .A2(new_n12044_), .A3(new_n12042_), .A4(new_n12943_), .ZN(new_n12950_));
  NOR2_X1    g11928(.A1(new_n12950_), .A2(new_n12052_), .ZN(new_n12951_));
  OAI21_X1   g11929(.A1(new_n11986_), .A2(new_n11983_), .B(new_n11982_), .ZN(new_n12952_));
  NAND3_X1   g11930(.A1(new_n11978_), .A2(new_n11980_), .A3(new_n11976_), .ZN(new_n12953_));
  NAND2_X1   g11931(.A1(new_n12952_), .A2(new_n12953_), .ZN(new_n12954_));
  NOR4_X1    g11932(.A1(new_n12003_), .A2(new_n11970_), .A3(new_n11995_), .A4(new_n12954_), .ZN(new_n12955_));
  INV_X1     g11933(.I(new_n12955_), .ZN(new_n12956_));
  OAI21_X1   g11934(.A1(new_n12951_), .A2(new_n12956_), .B(new_n12053_), .ZN(new_n12957_));
  AOI21_X1   g11935(.A1(new_n12006_), .A2(new_n12017_), .B(new_n12943_), .ZN(new_n12958_));
  OAI21_X1   g11936(.A1(new_n9718_), .A2(new_n9621_), .B(new_n12009_), .ZN(new_n12959_));
  NOR2_X1    g11937(.A1(new_n9576_), .A2(new_n9574_), .ZN(new_n12960_));
  OAI21_X1   g11938(.A1(new_n9734_), .A2(new_n12960_), .B(new_n9732_), .ZN(new_n12961_));
  NAND2_X1   g11939(.A1(new_n12959_), .A2(new_n12961_), .ZN(new_n12962_));
  NOR2_X1    g11940(.A1(new_n12958_), .A2(new_n12962_), .ZN(new_n12963_));
  OAI21_X1   g11941(.A1(new_n12044_), .A2(new_n12042_), .B(new_n12024_), .ZN(new_n12964_));
  INV_X1     g11942(.I(new_n12962_), .ZN(new_n12965_));
  NOR2_X1    g11943(.A1(new_n12964_), .A2(new_n12965_), .ZN(new_n12966_));
  OAI21_X1   g11944(.A1(new_n12963_), .A2(new_n12966_), .B(new_n12031_), .ZN(new_n12967_));
  NAND2_X1   g11945(.A1(new_n12964_), .A2(new_n12965_), .ZN(new_n12968_));
  NAND2_X1   g11946(.A1(new_n12006_), .A2(new_n12017_), .ZN(new_n12969_));
  NAND3_X1   g11947(.A1(new_n12969_), .A2(new_n12024_), .A3(new_n12962_), .ZN(new_n12970_));
  NAND3_X1   g11948(.A1(new_n12968_), .A2(new_n12970_), .A3(new_n12949_), .ZN(new_n12971_));
  NAND2_X1   g11949(.A1(new_n12967_), .A2(new_n12971_), .ZN(new_n12972_));
  NAND2_X1   g11950(.A1(new_n11994_), .A2(new_n9702_), .ZN(new_n12973_));
  NOR2_X1    g11951(.A1(new_n11997_), .A2(new_n11971_), .ZN(new_n12974_));
  AOI21_X1   g11952(.A1(new_n11971_), .A2(new_n11998_), .B(new_n12974_), .ZN(new_n12975_));
  INV_X1     g11953(.I(new_n12002_), .ZN(new_n12976_));
  NOR3_X1    g11954(.A1(new_n12975_), .A2(new_n12976_), .A3(new_n12973_), .ZN(new_n12977_));
  OAI21_X1   g11955(.A1(new_n11975_), .A2(new_n12954_), .B(new_n11970_), .ZN(new_n12978_));
  AOI21_X1   g11956(.A1(new_n9701_), .A2(new_n9688_), .B(new_n11977_), .ZN(new_n12979_));
  OR4_X2     g11957(.A1(new_n9629_), .A2(new_n9645_), .A3(new_n9646_), .A4(new_n9641_), .Z(new_n12980_));
  AOI21_X1   g11958(.A1(new_n11992_), .A2(new_n12980_), .B(new_n9723_), .ZN(new_n12981_));
  NOR2_X1    g11959(.A1(new_n12981_), .A2(new_n12979_), .ZN(new_n12982_));
  NAND2_X1   g11960(.A1(new_n12978_), .A2(new_n12982_), .ZN(new_n12983_));
  NAND2_X1   g11961(.A1(new_n11995_), .A2(new_n11988_), .ZN(new_n12984_));
  INV_X1     g11962(.I(new_n12982_), .ZN(new_n12985_));
  NAND3_X1   g11963(.A1(new_n12984_), .A2(new_n11970_), .A3(new_n12985_), .ZN(new_n12986_));
  AOI21_X1   g11964(.A1(new_n12983_), .A2(new_n12986_), .B(new_n12977_), .ZN(new_n12987_));
  NAND3_X1   g11965(.A1(new_n12000_), .A2(new_n11996_), .A3(new_n12002_), .ZN(new_n12988_));
  AOI21_X1   g11966(.A1(new_n12984_), .A2(new_n11970_), .B(new_n12985_), .ZN(new_n12989_));
  NOR2_X1    g11967(.A1(new_n12978_), .A2(new_n12982_), .ZN(new_n12990_));
  NOR3_X1    g11968(.A1(new_n12990_), .A2(new_n12989_), .A3(new_n12988_), .ZN(new_n12991_));
  NOR2_X1    g11969(.A1(new_n12991_), .A2(new_n12987_), .ZN(new_n12992_));
  NOR2_X1    g11970(.A1(new_n12992_), .A2(new_n12972_), .ZN(new_n12993_));
  AOI21_X1   g11971(.A1(new_n12968_), .A2(new_n12970_), .B(new_n12949_), .ZN(new_n12994_));
  NOR3_X1    g11972(.A1(new_n12963_), .A2(new_n12966_), .A3(new_n12031_), .ZN(new_n12995_));
  NOR2_X1    g11973(.A1(new_n12994_), .A2(new_n12995_), .ZN(new_n12996_));
  OAI21_X1   g11974(.A1(new_n12990_), .A2(new_n12989_), .B(new_n12988_), .ZN(new_n12997_));
  NAND3_X1   g11975(.A1(new_n12983_), .A2(new_n12986_), .A3(new_n12977_), .ZN(new_n12998_));
  NAND2_X1   g11976(.A1(new_n12997_), .A2(new_n12998_), .ZN(new_n12999_));
  NOR2_X1    g11977(.A1(new_n12999_), .A2(new_n12996_), .ZN(new_n13000_));
  OAI21_X1   g11978(.A1(new_n13000_), .A2(new_n12993_), .B(new_n12957_), .ZN(new_n13001_));
  NAND2_X1   g11979(.A1(new_n12032_), .A2(new_n12037_), .ZN(new_n13002_));
  AOI21_X1   g11980(.A1(new_n13002_), .A2(new_n12955_), .B(new_n12038_), .ZN(new_n13003_));
  AOI22_X1   g11981(.A1(new_n12997_), .A2(new_n12998_), .B1(new_n12967_), .B2(new_n12971_), .ZN(new_n13004_));
  NOR4_X1    g11982(.A1(new_n12994_), .A2(new_n12991_), .A3(new_n12987_), .A4(new_n12995_), .ZN(new_n13005_));
  OAI21_X1   g11983(.A1(new_n13005_), .A2(new_n13004_), .B(new_n13003_), .ZN(new_n13006_));
  AOI21_X1   g11984(.A1(new_n13001_), .A2(new_n13006_), .B(new_n12940_), .ZN(new_n13007_));
  NAND2_X1   g11985(.A1(new_n12927_), .A2(new_n12930_), .ZN(new_n13008_));
  NAND2_X1   g11986(.A1(new_n12906_), .A2(new_n12919_), .ZN(new_n13009_));
  AOI21_X1   g11987(.A1(new_n13008_), .A2(new_n13009_), .B(new_n12936_), .ZN(new_n13010_));
  NAND2_X1   g11988(.A1(new_n12906_), .A2(new_n12930_), .ZN(new_n13011_));
  NAND2_X1   g11989(.A1(new_n12927_), .A2(new_n12919_), .ZN(new_n13012_));
  AOI21_X1   g11990(.A1(new_n13012_), .A2(new_n13011_), .B(new_n12893_), .ZN(new_n13013_));
  NOR2_X1    g11991(.A1(new_n13010_), .A2(new_n13013_), .ZN(new_n13014_));
  NAND2_X1   g11992(.A1(new_n12999_), .A2(new_n12996_), .ZN(new_n13015_));
  NAND3_X1   g11993(.A1(new_n12972_), .A2(new_n12997_), .A3(new_n12998_), .ZN(new_n13016_));
  AOI21_X1   g11994(.A1(new_n13015_), .A2(new_n13016_), .B(new_n13003_), .ZN(new_n13017_));
  OAI22_X1   g11995(.A1(new_n12987_), .A2(new_n12991_), .B1(new_n12994_), .B2(new_n12995_), .ZN(new_n13018_));
  NAND4_X1   g11996(.A1(new_n12967_), .A2(new_n12997_), .A3(new_n12998_), .A4(new_n12971_), .ZN(new_n13019_));
  AOI21_X1   g11997(.A1(new_n13018_), .A2(new_n13019_), .B(new_n12957_), .ZN(new_n13020_));
  NOR3_X1    g11998(.A1(new_n13017_), .A2(new_n13014_), .A3(new_n13020_), .ZN(new_n13021_));
  OAI21_X1   g11999(.A1(new_n13007_), .A2(new_n13021_), .B(new_n12889_), .ZN(new_n13022_));
  OAI21_X1   g12000(.A1(new_n9903_), .A2(new_n12169_), .B(new_n12055_), .ZN(new_n13023_));
  AOI21_X1   g12001(.A1(new_n13001_), .A2(new_n13006_), .B(new_n13014_), .ZN(new_n13024_));
  NOR3_X1    g12002(.A1(new_n13017_), .A2(new_n12940_), .A3(new_n13020_), .ZN(new_n13025_));
  OAI21_X1   g12003(.A1(new_n13024_), .A2(new_n13025_), .B(new_n13023_), .ZN(new_n13026_));
  NAND2_X1   g12004(.A1(new_n13022_), .A2(new_n13026_), .ZN(new_n13027_));
  AOI21_X1   g12005(.A1(new_n11958_), .A2(new_n11947_), .B(new_n11946_), .ZN(new_n13028_));
  NOR3_X1    g12006(.A1(new_n11939_), .A2(new_n11863_), .A3(new_n11930_), .ZN(new_n13029_));
  OAI21_X1   g12007(.A1(new_n13028_), .A2(new_n13029_), .B(new_n10220_), .ZN(new_n13030_));
  NOR3_X1    g12008(.A1(new_n13028_), .A2(new_n13029_), .A3(new_n10220_), .ZN(new_n13031_));
  OAI21_X1   g12009(.A1(new_n11832_), .A2(new_n13031_), .B(new_n13030_), .ZN(new_n13032_));
  NOR3_X1    g12010(.A1(new_n11924_), .A2(new_n11916_), .A3(new_n11929_), .ZN(new_n13033_));
  AOI21_X1   g12011(.A1(new_n11956_), .A2(new_n11950_), .B(new_n11938_), .ZN(new_n13034_));
  NAND2_X1   g12012(.A1(new_n11946_), .A2(new_n11874_), .ZN(new_n13035_));
  NOR2_X1    g12013(.A1(new_n13034_), .A2(new_n13035_), .ZN(new_n13036_));
  NAND3_X1   g12014(.A1(new_n10187_), .A2(new_n11888_), .A3(new_n11891_), .ZN(new_n13037_));
  NOR4_X1    g12015(.A1(new_n10082_), .A2(new_n10083_), .A3(new_n10054_), .A4(new_n10064_), .ZN(new_n13038_));
  OAI21_X1   g12016(.A1(new_n10067_), .A2(new_n13038_), .B(new_n10084_), .ZN(new_n13039_));
  INV_X1     g12017(.I(new_n13039_), .ZN(new_n13040_));
  AOI21_X1   g12018(.A1(new_n13037_), .A2(new_n11918_), .B(new_n13040_), .ZN(new_n13041_));
  NOR3_X1    g12019(.A1(new_n11908_), .A2(new_n11907_), .A3(new_n10204_), .ZN(new_n13042_));
  NOR3_X1    g12020(.A1(new_n13042_), .A2(new_n11921_), .A3(new_n13039_), .ZN(new_n13043_));
  AOI21_X1   g12021(.A1(new_n11906_), .A2(new_n11895_), .B(new_n11914_), .ZN(new_n13044_));
  OAI22_X1   g12022(.A1(new_n11934_), .A2(new_n13044_), .B1(new_n13041_), .B2(new_n13043_), .ZN(new_n13045_));
  AOI21_X1   g12023(.A1(new_n11869_), .A2(new_n11866_), .B(new_n10153_), .ZN(new_n13046_));
  NAND2_X1   g12024(.A1(new_n10123_), .A2(new_n10124_), .ZN(new_n13047_));
  NAND3_X1   g12025(.A1(new_n10097_), .A2(new_n10108_), .A3(new_n13047_), .ZN(new_n13048_));
  NAND2_X1   g12026(.A1(new_n13048_), .A2(new_n11835_), .ZN(new_n13049_));
  XOR2_X1    g12027(.A1(new_n13046_), .A2(new_n13049_), .Z(new_n13050_));
  OAI22_X1   g12028(.A1(new_n11861_), .A2(new_n11848_), .B1(new_n11839_), .B2(new_n11837_), .ZN(new_n13051_));
  AOI21_X1   g12029(.A1(new_n11872_), .A2(new_n13051_), .B(new_n13050_), .ZN(new_n13052_));
  NOR2_X1    g12030(.A1(new_n13045_), .A2(new_n13052_), .ZN(new_n13053_));
  NAND2_X1   g12031(.A1(new_n11953_), .A2(new_n11954_), .ZN(new_n13054_));
  INV_X1     g12032(.I(new_n13041_), .ZN(new_n13055_));
  NAND3_X1   g12033(.A1(new_n13037_), .A2(new_n11918_), .A3(new_n13040_), .ZN(new_n13056_));
  OAI21_X1   g12034(.A1(new_n11911_), .A2(new_n11882_), .B(new_n11904_), .ZN(new_n13057_));
  AOI22_X1   g12035(.A1(new_n13054_), .A2(new_n13057_), .B1(new_n13055_), .B2(new_n13056_), .ZN(new_n13058_));
  NAND2_X1   g12036(.A1(new_n11868_), .A2(new_n11871_), .ZN(new_n13059_));
  NOR2_X1    g12037(.A1(new_n13059_), .A2(new_n11855_), .ZN(new_n13060_));
  NAND2_X1   g12038(.A1(new_n11867_), .A2(new_n10152_), .ZN(new_n13061_));
  INV_X1     g12039(.I(new_n13049_), .ZN(new_n13062_));
  NOR2_X1    g12040(.A1(new_n13062_), .A2(new_n13061_), .ZN(new_n13063_));
  NOR2_X1    g12041(.A1(new_n13046_), .A2(new_n13049_), .ZN(new_n13064_));
  AOI22_X1   g12042(.A1(new_n11855_), .A2(new_n11858_), .B1(new_n11942_), .B2(new_n11838_), .ZN(new_n13065_));
  OAI22_X1   g12043(.A1(new_n13060_), .A2(new_n13065_), .B1(new_n13063_), .B2(new_n13064_), .ZN(new_n13066_));
  NOR2_X1    g12044(.A1(new_n13058_), .A2(new_n13066_), .ZN(new_n13067_));
  OAI22_X1   g12045(.A1(new_n13036_), .A2(new_n13033_), .B1(new_n13067_), .B2(new_n13053_), .ZN(new_n13068_));
  OAI21_X1   g12046(.A1(new_n11924_), .A2(new_n11916_), .B(new_n11929_), .ZN(new_n13069_));
  NOR2_X1    g12047(.A1(new_n11863_), .A2(new_n11931_), .ZN(new_n13070_));
  AOI21_X1   g12048(.A1(new_n13069_), .A2(new_n13070_), .B(new_n13033_), .ZN(new_n13071_));
  NAND2_X1   g12049(.A1(new_n13045_), .A2(new_n13066_), .ZN(new_n13072_));
  NAND2_X1   g12050(.A1(new_n13058_), .A2(new_n13052_), .ZN(new_n13073_));
  NAND2_X1   g12051(.A1(new_n13073_), .A2(new_n13072_), .ZN(new_n13074_));
  NAND2_X1   g12052(.A1(new_n13074_), .A2(new_n13071_), .ZN(new_n13075_));
  NAND2_X1   g12053(.A1(new_n13075_), .A2(new_n13068_), .ZN(new_n13076_));
  XOR2_X1    g12054(.A1(new_n9931_), .A2(new_n9958_), .Z(new_n13077_));
  OAI21_X1   g12055(.A1(new_n11790_), .A2(new_n11787_), .B(new_n11786_), .ZN(new_n13078_));
  NAND3_X1   g12056(.A1(new_n11777_), .A2(new_n11779_), .A3(new_n10007_), .ZN(new_n13079_));
  NAND2_X1   g12057(.A1(new_n13078_), .A2(new_n13079_), .ZN(new_n13080_));
  NAND2_X1   g12058(.A1(new_n11806_), .A2(new_n9996_), .ZN(new_n13081_));
  NAND2_X1   g12059(.A1(new_n13081_), .A2(new_n11822_), .ZN(new_n13082_));
  NOR2_X1    g12060(.A1(new_n11821_), .A2(new_n13082_), .ZN(new_n13083_));
  AND2_X2    g12061(.A1(new_n11812_), .A2(new_n11815_), .Z(new_n13084_));
  NOR3_X1    g12062(.A1(new_n13084_), .A2(new_n13083_), .A3(new_n13080_), .ZN(new_n13085_));
  NAND3_X1   g12063(.A1(new_n13085_), .A2(new_n13077_), .A3(new_n10030_), .ZN(new_n13086_));
  AOI21_X1   g12064(.A1(new_n13077_), .A2(new_n10030_), .B(new_n13085_), .ZN(new_n13087_));
  AOI21_X1   g12065(.A1(new_n11762_), .A2(new_n11763_), .B(new_n10020_), .ZN(new_n13088_));
  NOR3_X1    g12066(.A1(new_n11760_), .A2(new_n11757_), .A3(new_n9979_), .ZN(new_n13089_));
  NOR2_X1    g12067(.A1(new_n13089_), .A2(new_n13088_), .ZN(new_n13090_));
  NAND4_X1   g12068(.A1(new_n11774_), .A2(new_n11768_), .A3(new_n11769_), .A4(new_n13090_), .ZN(new_n13091_));
  OAI21_X1   g12069(.A1(new_n13087_), .A2(new_n13091_), .B(new_n13086_), .ZN(new_n13092_));
  NOR3_X1    g12070(.A1(new_n11825_), .A2(new_n11821_), .A3(new_n11792_), .ZN(new_n13093_));
  INV_X1     g12071(.I(new_n13093_), .ZN(new_n13094_));
  OAI21_X1   g12072(.A1(new_n11821_), .A2(new_n13082_), .B(new_n11792_), .ZN(new_n13095_));
  NAND2_X1   g12073(.A1(new_n9928_), .A2(new_n9929_), .ZN(new_n13096_));
  NAND3_X1   g12074(.A1(new_n11802_), .A2(new_n9927_), .A3(new_n13096_), .ZN(new_n13097_));
  AOI22_X1   g12075(.A1(new_n11809_), .A2(new_n13097_), .B1(new_n11824_), .B2(new_n11778_), .ZN(new_n13098_));
  INV_X1     g12076(.I(new_n13098_), .ZN(new_n13099_));
  AOI21_X1   g12077(.A1(new_n13095_), .A2(new_n11816_), .B(new_n13099_), .ZN(new_n13100_));
  AOI21_X1   g12078(.A1(new_n11804_), .A2(new_n11807_), .B(new_n13080_), .ZN(new_n13101_));
  NOR3_X1    g12079(.A1(new_n13101_), .A2(new_n13084_), .A3(new_n13098_), .ZN(new_n13102_));
  OAI21_X1   g12080(.A1(new_n13102_), .A2(new_n13100_), .B(new_n13094_), .ZN(new_n13103_));
  OAI21_X1   g12081(.A1(new_n13101_), .A2(new_n13084_), .B(new_n13098_), .ZN(new_n13104_));
  NAND3_X1   g12082(.A1(new_n13095_), .A2(new_n11816_), .A3(new_n13099_), .ZN(new_n13105_));
  NAND3_X1   g12083(.A1(new_n13104_), .A2(new_n13105_), .A3(new_n13093_), .ZN(new_n13106_));
  NAND2_X1   g12084(.A1(new_n13103_), .A2(new_n13106_), .ZN(new_n13107_));
  NOR2_X1    g12085(.A1(new_n11734_), .A2(new_n10020_), .ZN(new_n13108_));
  NOR2_X1    g12086(.A1(new_n9979_), .A2(new_n9954_), .ZN(new_n13109_));
  NOR2_X1    g12087(.A1(new_n11748_), .A2(new_n10037_), .ZN(new_n13110_));
  NOR2_X1    g12088(.A1(new_n9943_), .A2(new_n9968_), .ZN(new_n13111_));
  OAI22_X1   g12089(.A1(new_n13108_), .A2(new_n13109_), .B1(new_n13110_), .B2(new_n13111_), .ZN(new_n13112_));
  NOR4_X1    g12090(.A1(new_n13112_), .A2(new_n13090_), .A3(new_n11751_), .A4(new_n11771_), .ZN(new_n13113_));
  AOI21_X1   g12091(.A1(new_n11754_), .A2(new_n11750_), .B(new_n11765_), .ZN(new_n13114_));
  NAND2_X1   g12092(.A1(new_n9955_), .A2(new_n9956_), .ZN(new_n13115_));
  NAND3_X1   g12093(.A1(new_n10037_), .A2(new_n9954_), .A3(new_n13115_), .ZN(new_n13116_));
  AOI22_X1   g12094(.A1(new_n13116_), .A2(new_n11731_), .B1(new_n11771_), .B2(new_n11756_), .ZN(new_n13117_));
  OAI21_X1   g12095(.A1(new_n13114_), .A2(new_n11769_), .B(new_n13117_), .ZN(new_n13118_));
  OAI21_X1   g12096(.A1(new_n13112_), .A2(new_n11753_), .B(new_n13090_), .ZN(new_n13119_));
  INV_X1     g12097(.I(new_n13117_), .ZN(new_n13120_));
  NAND3_X1   g12098(.A1(new_n13119_), .A2(new_n11738_), .A3(new_n13120_), .ZN(new_n13121_));
  AOI21_X1   g12099(.A1(new_n13121_), .A2(new_n13118_), .B(new_n13113_), .ZN(new_n13122_));
  AOI21_X1   g12100(.A1(new_n13119_), .A2(new_n11738_), .B(new_n13120_), .ZN(new_n13123_));
  NOR3_X1    g12101(.A1(new_n13114_), .A2(new_n13117_), .A3(new_n11769_), .ZN(new_n13124_));
  NOR3_X1    g12102(.A1(new_n13123_), .A2(new_n13124_), .A3(new_n11773_), .ZN(new_n13125_));
  NOR2_X1    g12103(.A1(new_n13125_), .A2(new_n13122_), .ZN(new_n13126_));
  NOR2_X1    g12104(.A1(new_n13126_), .A2(new_n13107_), .ZN(new_n13127_));
  AOI21_X1   g12105(.A1(new_n13104_), .A2(new_n13105_), .B(new_n13093_), .ZN(new_n13128_));
  NOR3_X1    g12106(.A1(new_n13102_), .A2(new_n13100_), .A3(new_n13094_), .ZN(new_n13129_));
  NOR2_X1    g12107(.A1(new_n13129_), .A2(new_n13128_), .ZN(new_n13130_));
  OAI21_X1   g12108(.A1(new_n13123_), .A2(new_n13124_), .B(new_n11773_), .ZN(new_n13131_));
  NAND3_X1   g12109(.A1(new_n13121_), .A2(new_n13118_), .A3(new_n13113_), .ZN(new_n13132_));
  NAND2_X1   g12110(.A1(new_n13131_), .A2(new_n13132_), .ZN(new_n13133_));
  NOR2_X1    g12111(.A1(new_n13130_), .A2(new_n13133_), .ZN(new_n13134_));
  OAI21_X1   g12112(.A1(new_n13127_), .A2(new_n13134_), .B(new_n13092_), .ZN(new_n13135_));
  OAI21_X1   g12113(.A1(new_n11776_), .A2(new_n10041_), .B(new_n11827_), .ZN(new_n13136_));
  NAND2_X1   g12114(.A1(new_n13113_), .A2(new_n11738_), .ZN(new_n13137_));
  NOR4_X1    g12115(.A1(new_n13137_), .A2(new_n11755_), .A3(new_n11738_), .A4(new_n11765_), .ZN(new_n13138_));
  AOI21_X1   g12116(.A1(new_n13138_), .A2(new_n13136_), .B(new_n11828_), .ZN(new_n13139_));
  AOI22_X1   g12117(.A1(new_n13103_), .A2(new_n13106_), .B1(new_n13131_), .B2(new_n13132_), .ZN(new_n13140_));
  NOR4_X1    g12118(.A1(new_n13128_), .A2(new_n13129_), .A3(new_n13125_), .A4(new_n13122_), .ZN(new_n13141_));
  OAI21_X1   g12119(.A1(new_n13141_), .A2(new_n13140_), .B(new_n13139_), .ZN(new_n13142_));
  AOI21_X1   g12120(.A1(new_n13135_), .A2(new_n13142_), .B(new_n13076_), .ZN(new_n13143_));
  NAND2_X1   g12121(.A1(new_n13069_), .A2(new_n13070_), .ZN(new_n13144_));
  NAND2_X1   g12122(.A1(new_n13058_), .A2(new_n13066_), .ZN(new_n13145_));
  NAND2_X1   g12123(.A1(new_n13045_), .A2(new_n13052_), .ZN(new_n13146_));
  AOI22_X1   g12124(.A1(new_n13144_), .A2(new_n11957_), .B1(new_n13145_), .B2(new_n13146_), .ZN(new_n13147_));
  OAI21_X1   g12125(.A1(new_n13034_), .A2(new_n13035_), .B(new_n11957_), .ZN(new_n13148_));
  NOR2_X1    g12126(.A1(new_n13058_), .A2(new_n13052_), .ZN(new_n13149_));
  NOR2_X1    g12127(.A1(new_n13045_), .A2(new_n13066_), .ZN(new_n13150_));
  NOR2_X1    g12128(.A1(new_n13149_), .A2(new_n13150_), .ZN(new_n13151_));
  NOR2_X1    g12129(.A1(new_n13151_), .A2(new_n13148_), .ZN(new_n13152_));
  NOR2_X1    g12130(.A1(new_n13152_), .A2(new_n13147_), .ZN(new_n13153_));
  NAND2_X1   g12131(.A1(new_n13130_), .A2(new_n13133_), .ZN(new_n13154_));
  NAND2_X1   g12132(.A1(new_n13126_), .A2(new_n13107_), .ZN(new_n13155_));
  AOI21_X1   g12133(.A1(new_n13155_), .A2(new_n13154_), .B(new_n13139_), .ZN(new_n13156_));
  NAND2_X1   g12134(.A1(new_n13107_), .A2(new_n13133_), .ZN(new_n13157_));
  NAND4_X1   g12135(.A1(new_n13103_), .A2(new_n13106_), .A3(new_n13131_), .A4(new_n13132_), .ZN(new_n13158_));
  AOI21_X1   g12136(.A1(new_n13157_), .A2(new_n13158_), .B(new_n13092_), .ZN(new_n13159_));
  NOR3_X1    g12137(.A1(new_n13153_), .A2(new_n13156_), .A3(new_n13159_), .ZN(new_n13160_));
  OAI21_X1   g12138(.A1(new_n13143_), .A2(new_n13160_), .B(new_n13032_), .ZN(new_n13161_));
  INV_X1     g12139(.I(new_n11767_), .ZN(new_n13162_));
  AOI21_X1   g12140(.A1(new_n11830_), .A2(new_n11829_), .B(new_n13162_), .ZN(new_n13163_));
  NAND3_X1   g12141(.A1(new_n11959_), .A2(new_n11940_), .A3(new_n11833_), .ZN(new_n13164_));
  AOI21_X1   g12142(.A1(new_n13163_), .A2(new_n13164_), .B(new_n11960_), .ZN(new_n13165_));
  AOI22_X1   g12143(.A1(new_n13135_), .A2(new_n13142_), .B1(new_n13068_), .B2(new_n13075_), .ZN(new_n13166_));
  NOR3_X1    g12144(.A1(new_n13076_), .A2(new_n13156_), .A3(new_n13159_), .ZN(new_n13167_));
  OAI21_X1   g12145(.A1(new_n13166_), .A2(new_n13167_), .B(new_n13165_), .ZN(new_n13168_));
  AOI21_X1   g12146(.A1(new_n13161_), .A2(new_n13168_), .B(new_n13027_), .ZN(new_n13169_));
  OAI21_X1   g12147(.A1(new_n13017_), .A2(new_n13020_), .B(new_n13014_), .ZN(new_n13170_));
  NAND3_X1   g12148(.A1(new_n13001_), .A2(new_n12940_), .A3(new_n13006_), .ZN(new_n13171_));
  AOI21_X1   g12149(.A1(new_n13170_), .A2(new_n13171_), .B(new_n13023_), .ZN(new_n13172_));
  OAI21_X1   g12150(.A1(new_n13017_), .A2(new_n13020_), .B(new_n12940_), .ZN(new_n13173_));
  NAND3_X1   g12151(.A1(new_n13001_), .A2(new_n13014_), .A3(new_n13006_), .ZN(new_n13174_));
  AOI21_X1   g12152(.A1(new_n13173_), .A2(new_n13174_), .B(new_n12889_), .ZN(new_n13175_));
  NOR2_X1    g12153(.A1(new_n13172_), .A2(new_n13175_), .ZN(new_n13176_));
  OAI21_X1   g12154(.A1(new_n13156_), .A2(new_n13159_), .B(new_n13153_), .ZN(new_n13177_));
  NAND3_X1   g12155(.A1(new_n13076_), .A2(new_n13135_), .A3(new_n13142_), .ZN(new_n13178_));
  AOI21_X1   g12156(.A1(new_n13177_), .A2(new_n13178_), .B(new_n13165_), .ZN(new_n13179_));
  OAI21_X1   g12157(.A1(new_n13156_), .A2(new_n13159_), .B(new_n13076_), .ZN(new_n13180_));
  NAND3_X1   g12158(.A1(new_n13153_), .A2(new_n13135_), .A3(new_n13142_), .ZN(new_n13181_));
  AOI21_X1   g12159(.A1(new_n13180_), .A2(new_n13181_), .B(new_n13032_), .ZN(new_n13182_));
  NOR3_X1    g12160(.A1(new_n13176_), .A2(new_n13179_), .A3(new_n13182_), .ZN(new_n13183_));
  OAI21_X1   g12161(.A1(new_n13169_), .A2(new_n13183_), .B(new_n12885_), .ZN(new_n13184_));
  AOI21_X1   g12162(.A1(new_n12170_), .A2(new_n12171_), .B(new_n10226_), .ZN(new_n13185_));
  AOI21_X1   g12163(.A1(new_n11961_), .A2(new_n12883_), .B(new_n13185_), .ZN(new_n13186_));
  AOI22_X1   g12164(.A1(new_n13161_), .A2(new_n13168_), .B1(new_n13022_), .B2(new_n13026_), .ZN(new_n13187_));
  NOR4_X1    g12165(.A1(new_n13179_), .A2(new_n13182_), .A3(new_n13172_), .A4(new_n13175_), .ZN(new_n13188_));
  OAI21_X1   g12166(.A1(new_n13188_), .A2(new_n13187_), .B(new_n13186_), .ZN(new_n13189_));
  AOI21_X1   g12167(.A1(new_n13184_), .A2(new_n13189_), .B(new_n12882_), .ZN(new_n13190_));
  NAND2_X1   g12168(.A1(new_n12875_), .A2(new_n12868_), .ZN(new_n13191_));
  NAND3_X1   g12169(.A1(new_n12709_), .A2(new_n12871_), .A3(new_n12874_), .ZN(new_n13192_));
  NAND2_X1   g12170(.A1(new_n13191_), .A2(new_n13192_), .ZN(new_n13193_));
  OAI22_X1   g12171(.A1(new_n12851_), .A2(new_n12859_), .B1(new_n12864_), .B2(new_n12867_), .ZN(new_n13194_));
  NAND4_X1   g12172(.A1(new_n12871_), .A2(new_n12703_), .A3(new_n12874_), .A4(new_n12708_), .ZN(new_n13195_));
  AOI21_X1   g12173(.A1(new_n13194_), .A2(new_n13195_), .B(new_n12563_), .ZN(new_n13196_));
  AOI21_X1   g12174(.A1(new_n13193_), .A2(new_n12563_), .B(new_n13196_), .ZN(new_n13197_));
  OAI21_X1   g12175(.A1(new_n13179_), .A2(new_n13182_), .B(new_n13176_), .ZN(new_n13198_));
  NAND3_X1   g12176(.A1(new_n13027_), .A2(new_n13161_), .A3(new_n13168_), .ZN(new_n13199_));
  AOI21_X1   g12177(.A1(new_n13198_), .A2(new_n13199_), .B(new_n13186_), .ZN(new_n13200_));
  OAI22_X1   g12178(.A1(new_n13179_), .A2(new_n13182_), .B1(new_n13172_), .B2(new_n13175_), .ZN(new_n13201_));
  NAND4_X1   g12179(.A1(new_n13161_), .A2(new_n13168_), .A3(new_n13022_), .A4(new_n13026_), .ZN(new_n13202_));
  AOI21_X1   g12180(.A1(new_n13201_), .A2(new_n13202_), .B(new_n12885_), .ZN(new_n13203_));
  NOR3_X1    g12181(.A1(new_n13197_), .A2(new_n13200_), .A3(new_n13203_), .ZN(new_n13204_));
  OAI21_X1   g12182(.A1(new_n13190_), .A2(new_n13204_), .B(new_n12560_), .ZN(new_n13205_));
  AOI22_X1   g12183(.A1(new_n13184_), .A2(new_n13189_), .B1(new_n12877_), .B2(new_n12881_), .ZN(new_n13206_));
  AOI21_X1   g12184(.A1(new_n13191_), .A2(new_n13192_), .B(new_n12878_), .ZN(new_n13207_));
  NOR4_X1    g12185(.A1(new_n13200_), .A2(new_n13207_), .A3(new_n13196_), .A4(new_n13203_), .ZN(new_n13208_));
  OAI21_X1   g12186(.A1(new_n13208_), .A2(new_n13206_), .B(new_n12559_), .ZN(new_n13209_));
  NAND2_X1   g12187(.A1(new_n13205_), .A2(new_n13209_), .ZN(new_n13210_));
  INV_X1     g12188(.I(new_n11319_), .ZN(new_n13211_));
  NAND3_X1   g12189(.A1(new_n11725_), .A2(new_n11727_), .A3(new_n9550_), .ZN(new_n13212_));
  AOI21_X1   g12190(.A1(new_n13211_), .A2(new_n13212_), .B(new_n11728_), .ZN(new_n13213_));
  NAND3_X1   g12191(.A1(new_n9548_), .A2(new_n11719_), .A3(new_n11723_), .ZN(new_n13214_));
  AOI21_X1   g12192(.A1(new_n11726_), .A2(new_n13214_), .B(new_n11724_), .ZN(new_n13215_));
  NAND3_X1   g12193(.A1(new_n11713_), .A2(new_n11717_), .A3(new_n9544_), .ZN(new_n13216_));
  AOI21_X1   g12194(.A1(new_n11722_), .A2(new_n13216_), .B(new_n11718_), .ZN(new_n13217_));
  NAND3_X1   g12195(.A1(new_n11675_), .A2(new_n11669_), .A3(new_n11672_), .ZN(new_n13218_));
  AOI21_X1   g12196(.A1(new_n9481_), .A2(new_n9486_), .B(new_n9501_), .ZN(new_n13219_));
  AOI22_X1   g12197(.A1(new_n11684_), .A2(new_n11685_), .B1(new_n9498_), .B2(new_n13219_), .ZN(new_n13220_));
  NAND4_X1   g12198(.A1(new_n13220_), .A2(new_n9510_), .A3(new_n9516_), .A4(new_n9519_), .ZN(new_n13221_));
  NAND4_X1   g12199(.A1(new_n13218_), .A2(new_n13221_), .A3(new_n11683_), .A4(new_n11666_), .ZN(new_n13222_));
  NAND2_X1   g12200(.A1(new_n13222_), .A2(new_n9540_), .ZN(new_n13223_));
  NOR4_X1    g12201(.A1(new_n11663_), .A2(new_n11657_), .A3(new_n11633_), .A4(new_n11646_), .ZN(new_n13224_));
  AOI21_X1   g12202(.A1(new_n13223_), .A2(new_n13224_), .B(new_n11711_), .ZN(new_n13225_));
  NAND2_X1   g12203(.A1(new_n9517_), .A2(new_n9518_), .ZN(new_n13226_));
  NAND3_X1   g12204(.A1(new_n9510_), .A2(new_n9516_), .A3(new_n13226_), .ZN(new_n13227_));
  NAND2_X1   g12205(.A1(new_n13227_), .A2(new_n9475_), .ZN(new_n13228_));
  NOR2_X1    g12206(.A1(new_n9499_), .A2(new_n9485_), .ZN(new_n13229_));
  NAND2_X1   g12207(.A1(new_n13229_), .A2(new_n11687_), .ZN(new_n13230_));
  NAND3_X1   g12208(.A1(new_n9487_), .A2(new_n9498_), .A3(new_n13230_), .ZN(new_n13231_));
  AOI21_X1   g12209(.A1(new_n9501_), .A2(new_n13231_), .B(new_n13228_), .ZN(new_n13232_));
  NAND2_X1   g12210(.A1(new_n13231_), .A2(new_n9501_), .ZN(new_n13233_));
  AOI21_X1   g12211(.A1(new_n9475_), .A2(new_n13227_), .B(new_n13233_), .ZN(new_n13234_));
  NOR2_X1    g12212(.A1(new_n13232_), .A2(new_n13234_), .ZN(new_n13235_));
  NOR3_X1    g12213(.A1(new_n11705_), .A2(new_n11701_), .A3(new_n11702_), .ZN(new_n13236_));
  OAI21_X1   g12214(.A1(new_n13236_), .A2(new_n11700_), .B(new_n11683_), .ZN(new_n13237_));
  AOI21_X1   g12215(.A1(new_n13237_), .A2(new_n13221_), .B(new_n13235_), .ZN(new_n13238_));
  INV_X1     g12216(.I(new_n11697_), .ZN(new_n13239_));
  NOR2_X1    g12217(.A1(new_n9375_), .A2(new_n9386_), .ZN(new_n13240_));
  NAND2_X1   g12218(.A1(new_n9432_), .A2(new_n9433_), .ZN(new_n13241_));
  AOI21_X1   g12219(.A1(new_n13240_), .A2(new_n13241_), .B(new_n9434_), .ZN(new_n13242_));
  NOR4_X1    g12220(.A1(new_n9413_), .A2(new_n9415_), .A3(new_n9399_), .A4(new_n9410_), .ZN(new_n13243_));
  OAI21_X1   g12221(.A1(new_n11693_), .A2(new_n13243_), .B(new_n9448_), .ZN(new_n13244_));
  NAND2_X1   g12222(.A1(new_n13242_), .A2(new_n13244_), .ZN(new_n13245_));
  NAND3_X1   g12223(.A1(new_n9425_), .A2(new_n9431_), .A3(new_n13241_), .ZN(new_n13246_));
  NAND2_X1   g12224(.A1(new_n13246_), .A2(new_n9389_), .ZN(new_n13247_));
  INV_X1     g12225(.I(new_n13244_), .ZN(new_n13248_));
  NAND2_X1   g12226(.A1(new_n13248_), .A2(new_n13247_), .ZN(new_n13249_));
  NAND2_X1   g12227(.A1(new_n13249_), .A2(new_n13245_), .ZN(new_n13250_));
  AOI21_X1   g12228(.A1(new_n11651_), .A2(new_n11633_), .B(new_n11631_), .ZN(new_n13251_));
  OAI21_X1   g12229(.A1(new_n13251_), .A2(new_n13239_), .B(new_n13250_), .ZN(new_n13252_));
  NAND2_X1   g12230(.A1(new_n13238_), .A2(new_n13252_), .ZN(new_n13253_));
  AOI22_X1   g12231(.A1(new_n9481_), .A2(new_n9486_), .B1(new_n9492_), .B2(new_n9497_), .ZN(new_n13254_));
  NOR4_X1    g12232(.A1(new_n9523_), .A2(new_n9525_), .A3(new_n9531_), .A4(new_n9529_), .ZN(new_n13255_));
  OAI22_X1   g12233(.A1(new_n13254_), .A2(new_n13255_), .B1(new_n11688_), .B2(new_n9532_), .ZN(new_n13256_));
  NOR4_X1    g12234(.A1(new_n13256_), .A2(new_n9461_), .A3(new_n9472_), .A4(new_n9475_), .ZN(new_n13257_));
  AOI21_X1   g12235(.A1(new_n13218_), .A2(new_n11666_), .B(new_n11709_), .ZN(new_n13258_));
  OAI22_X1   g12236(.A1(new_n13258_), .A2(new_n13257_), .B1(new_n13232_), .B2(new_n13234_), .ZN(new_n13259_));
  XOR2_X1    g12237(.A1(new_n13242_), .A2(new_n13244_), .Z(new_n13260_));
  OAI21_X1   g12238(.A1(new_n11646_), .A2(new_n11632_), .B(new_n11657_), .ZN(new_n13261_));
  AOI21_X1   g12239(.A1(new_n13261_), .A2(new_n11697_), .B(new_n13260_), .ZN(new_n13262_));
  NAND2_X1   g12240(.A1(new_n13262_), .A2(new_n13259_), .ZN(new_n13263_));
  AOI21_X1   g12241(.A1(new_n13263_), .A2(new_n13253_), .B(new_n13225_), .ZN(new_n13264_));
  NOR3_X1    g12242(.A1(new_n11706_), .A2(new_n11710_), .A3(new_n11709_), .ZN(new_n13265_));
  NOR2_X1    g12243(.A1(new_n13265_), .A2(new_n11665_), .ZN(new_n13266_));
  NAND4_X1   g12244(.A1(new_n11698_), .A2(new_n11631_), .A3(new_n11632_), .A4(new_n11651_), .ZN(new_n13267_));
  OAI21_X1   g12245(.A1(new_n13266_), .A2(new_n13267_), .B(new_n11691_), .ZN(new_n13268_));
  NAND2_X1   g12246(.A1(new_n13259_), .A2(new_n13252_), .ZN(new_n13269_));
  NAND2_X1   g12247(.A1(new_n13238_), .A2(new_n13262_), .ZN(new_n13270_));
  AOI21_X1   g12248(.A1(new_n13270_), .A2(new_n13269_), .B(new_n13268_), .ZN(new_n13271_));
  NOR2_X1    g12249(.A1(new_n13271_), .A2(new_n13264_), .ZN(new_n13272_));
  NOR2_X1    g12250(.A1(new_n9278_), .A2(new_n9361_), .ZN(new_n13273_));
  NAND2_X1   g12251(.A1(new_n9345_), .A2(new_n9331_), .ZN(new_n13274_));
  AOI21_X1   g12252(.A1(new_n11597_), .A2(new_n11598_), .B(new_n9300_), .ZN(new_n13275_));
  NOR3_X1    g12253(.A1(new_n11595_), .A2(new_n9344_), .A3(new_n11594_), .ZN(new_n13276_));
  NOR2_X1    g12254(.A1(new_n13276_), .A2(new_n13275_), .ZN(new_n13277_));
  NOR2_X1    g12255(.A1(new_n9344_), .A2(new_n9289_), .ZN(new_n13278_));
  NOR2_X1    g12256(.A1(new_n9338_), .A2(new_n9300_), .ZN(new_n13279_));
  OAI21_X1   g12257(.A1(new_n13278_), .A2(new_n13279_), .B(new_n9304_), .ZN(new_n13280_));
  NAND3_X1   g12258(.A1(new_n13277_), .A2(new_n13274_), .A3(new_n13280_), .ZN(new_n13281_));
  OAI21_X1   g12259(.A1(new_n11609_), .A2(new_n11608_), .B(new_n9327_), .ZN(new_n13282_));
  NAND3_X1   g12260(.A1(new_n11605_), .A2(new_n11606_), .A3(new_n9357_), .ZN(new_n13283_));
  NAND2_X1   g12261(.A1(new_n13282_), .A2(new_n13283_), .ZN(new_n13284_));
  NAND4_X1   g12262(.A1(new_n13273_), .A2(new_n13281_), .A3(new_n11618_), .A4(new_n13284_), .ZN(new_n13285_));
  NOR3_X1    g12263(.A1(new_n11603_), .A2(new_n13275_), .A3(new_n13276_), .ZN(new_n13286_));
  AOI22_X1   g12264(.A1(new_n9348_), .A2(new_n9350_), .B1(new_n9354_), .B2(new_n9356_), .ZN(new_n13287_));
  NOR4_X1    g12265(.A1(new_n9311_), .A2(new_n9315_), .A3(new_n9326_), .A4(new_n9322_), .ZN(new_n13288_));
  OAI22_X1   g12266(.A1(new_n13287_), .A2(new_n13288_), .B1(new_n11616_), .B2(new_n9327_), .ZN(new_n13289_));
  NOR4_X1    g12267(.A1(new_n13289_), .A2(new_n9338_), .A3(new_n9344_), .A4(new_n9303_), .ZN(new_n13290_));
  NOR4_X1    g12268(.A1(new_n13286_), .A2(new_n13290_), .A3(new_n11611_), .A4(new_n11593_), .ZN(new_n13291_));
  NOR2_X1    g12269(.A1(new_n13291_), .A2(new_n13273_), .ZN(new_n13292_));
  OAI22_X1   g12270(.A1(new_n9226_), .A2(new_n9230_), .B1(new_n9241_), .B2(new_n9237_), .ZN(new_n13293_));
  NAND4_X1   g12271(.A1(new_n9263_), .A2(new_n9265_), .A3(new_n9269_), .A4(new_n9271_), .ZN(new_n13294_));
  AOI21_X1   g12272(.A1(new_n9263_), .A2(new_n9265_), .B(new_n9245_), .ZN(new_n13295_));
  AOI22_X1   g12273(.A1(new_n13293_), .A2(new_n13294_), .B1(new_n9272_), .B2(new_n13295_), .ZN(new_n13296_));
  NAND4_X1   g12274(.A1(new_n13296_), .A2(new_n9204_), .A3(new_n9215_), .A4(new_n9219_), .ZN(new_n13297_));
  NOR2_X1    g12275(.A1(new_n11583_), .A2(new_n13297_), .ZN(new_n13298_));
  NAND4_X1   g12276(.A1(new_n13298_), .A2(new_n11556_), .A3(new_n11567_), .A4(new_n11583_), .ZN(new_n13299_));
  OAI21_X1   g12277(.A1(new_n13292_), .A2(new_n13299_), .B(new_n13285_), .ZN(new_n13300_));
  OR4_X2     g12278(.A1(new_n9287_), .A2(new_n9301_), .A3(new_n9302_), .A4(new_n9298_), .Z(new_n13301_));
  NAND3_X1   g12279(.A1(new_n9289_), .A2(new_n9300_), .A3(new_n13301_), .ZN(new_n13302_));
  NOR2_X1    g12280(.A1(new_n9328_), .A2(new_n9313_), .ZN(new_n13303_));
  NAND2_X1   g12281(.A1(new_n13303_), .A2(new_n11615_), .ZN(new_n13304_));
  NAND3_X1   g12282(.A1(new_n9351_), .A2(new_n9357_), .A3(new_n13304_), .ZN(new_n13305_));
  NAND2_X1   g12283(.A1(new_n13305_), .A2(new_n9330_), .ZN(new_n13306_));
  NAND3_X1   g12284(.A1(new_n13306_), .A2(new_n9303_), .A3(new_n13302_), .ZN(new_n13307_));
  NAND2_X1   g12285(.A1(new_n13302_), .A2(new_n9303_), .ZN(new_n13308_));
  NAND3_X1   g12286(.A1(new_n13308_), .A2(new_n9330_), .A3(new_n13305_), .ZN(new_n13309_));
  NAND2_X1   g12287(.A1(new_n13307_), .A2(new_n13309_), .ZN(new_n13310_));
  NAND3_X1   g12288(.A1(new_n13280_), .A2(new_n11596_), .A3(new_n11599_), .ZN(new_n13311_));
  AOI21_X1   g12289(.A1(new_n13311_), .A2(new_n13274_), .B(new_n11611_), .ZN(new_n13312_));
  OAI21_X1   g12290(.A1(new_n13312_), .A2(new_n13290_), .B(new_n13310_), .ZN(new_n13313_));
  NOR2_X1    g12291(.A1(new_n9253_), .A2(new_n9259_), .ZN(new_n13314_));
  OR4_X2     g12292(.A1(new_n9202_), .A2(new_n9216_), .A3(new_n9217_), .A4(new_n9213_), .Z(new_n13315_));
  AOI21_X1   g12293(.A1(new_n13314_), .A2(new_n13315_), .B(new_n9219_), .ZN(new_n13316_));
  NAND2_X1   g12294(.A1(new_n9273_), .A2(new_n9274_), .ZN(new_n13317_));
  NAND3_X1   g12295(.A1(new_n9266_), .A2(new_n9272_), .A3(new_n13317_), .ZN(new_n13318_));
  NAND2_X1   g12296(.A1(new_n13318_), .A2(new_n9245_), .ZN(new_n13319_));
  XOR2_X1    g12297(.A1(new_n13316_), .A2(new_n13319_), .Z(new_n13320_));
  OAI21_X1   g12298(.A1(new_n11590_), .A2(new_n11556_), .B(new_n11580_), .ZN(new_n13321_));
  AOI21_X1   g12299(.A1(new_n13297_), .A2(new_n13321_), .B(new_n13320_), .ZN(new_n13322_));
  NOR2_X1    g12300(.A1(new_n13322_), .A2(new_n13313_), .ZN(new_n13323_));
  AOI21_X1   g12301(.A1(new_n9348_), .A2(new_n9350_), .B(new_n9330_), .ZN(new_n13324_));
  AOI22_X1   g12302(.A1(new_n11612_), .A2(new_n11613_), .B1(new_n9357_), .B2(new_n13324_), .ZN(new_n13325_));
  NAND4_X1   g12303(.A1(new_n13325_), .A2(new_n9289_), .A3(new_n9300_), .A4(new_n9304_), .ZN(new_n13326_));
  AND2_X2    g12304(.A1(new_n13307_), .A2(new_n13309_), .Z(new_n13327_));
  OAI21_X1   g12305(.A1(new_n11600_), .A2(new_n11603_), .B(new_n13274_), .ZN(new_n13328_));
  NAND2_X1   g12306(.A1(new_n13328_), .A2(new_n13284_), .ZN(new_n13329_));
  AOI21_X1   g12307(.A1(new_n13329_), .A2(new_n13326_), .B(new_n13327_), .ZN(new_n13330_));
  INV_X1     g12308(.I(new_n13297_), .ZN(new_n13331_));
  NAND3_X1   g12309(.A1(new_n9204_), .A2(new_n9215_), .A3(new_n13315_), .ZN(new_n13332_));
  NAND2_X1   g12310(.A1(new_n13332_), .A2(new_n9218_), .ZN(new_n13333_));
  XOR2_X1    g12311(.A1(new_n13333_), .A2(new_n13319_), .Z(new_n13334_));
  AOI21_X1   g12312(.A1(new_n11567_), .A2(new_n11557_), .B(new_n11583_), .ZN(new_n13335_));
  OAI21_X1   g12313(.A1(new_n13335_), .A2(new_n13331_), .B(new_n13334_), .ZN(new_n13336_));
  NOR2_X1    g12314(.A1(new_n13330_), .A2(new_n13336_), .ZN(new_n13337_));
  OAI21_X1   g12315(.A1(new_n13337_), .A2(new_n13323_), .B(new_n13300_), .ZN(new_n13338_));
  NAND4_X1   g12316(.A1(new_n13311_), .A2(new_n13326_), .A3(new_n13284_), .A4(new_n13274_), .ZN(new_n13339_));
  NAND2_X1   g12317(.A1(new_n13339_), .A2(new_n9363_), .ZN(new_n13340_));
  NOR4_X1    g12318(.A1(new_n11581_), .A2(new_n11557_), .A3(new_n11590_), .A4(new_n11580_), .ZN(new_n13341_));
  AOI21_X1   g12319(.A1(new_n13341_), .A2(new_n13340_), .B(new_n11620_), .ZN(new_n13342_));
  NOR2_X1    g12320(.A1(new_n13330_), .A2(new_n13322_), .ZN(new_n13343_));
  NOR2_X1    g12321(.A1(new_n13336_), .A2(new_n13313_), .ZN(new_n13344_));
  OAI21_X1   g12322(.A1(new_n13343_), .A2(new_n13344_), .B(new_n13342_), .ZN(new_n13345_));
  NAND2_X1   g12323(.A1(new_n13338_), .A2(new_n13345_), .ZN(new_n13346_));
  NAND2_X1   g12324(.A1(new_n13346_), .A2(new_n13272_), .ZN(new_n13347_));
  NOR2_X1    g12325(.A1(new_n13262_), .A2(new_n13259_), .ZN(new_n13348_));
  NOR2_X1    g12326(.A1(new_n13238_), .A2(new_n13252_), .ZN(new_n13349_));
  OAI21_X1   g12327(.A1(new_n13349_), .A2(new_n13348_), .B(new_n13268_), .ZN(new_n13350_));
  NOR2_X1    g12328(.A1(new_n13238_), .A2(new_n13262_), .ZN(new_n13351_));
  NOR2_X1    g12329(.A1(new_n13259_), .A2(new_n13252_), .ZN(new_n13352_));
  OAI21_X1   g12330(.A1(new_n13351_), .A2(new_n13352_), .B(new_n13225_), .ZN(new_n13353_));
  NAND2_X1   g12331(.A1(new_n13350_), .A2(new_n13353_), .ZN(new_n13354_));
  NAND2_X1   g12332(.A1(new_n13330_), .A2(new_n13336_), .ZN(new_n13355_));
  NAND2_X1   g12333(.A1(new_n13322_), .A2(new_n13313_), .ZN(new_n13356_));
  AOI21_X1   g12334(.A1(new_n13355_), .A2(new_n13356_), .B(new_n13342_), .ZN(new_n13357_));
  NAND2_X1   g12335(.A1(new_n13336_), .A2(new_n13313_), .ZN(new_n13358_));
  NAND2_X1   g12336(.A1(new_n13330_), .A2(new_n13322_), .ZN(new_n13359_));
  AOI21_X1   g12337(.A1(new_n13359_), .A2(new_n13358_), .B(new_n13300_), .ZN(new_n13360_));
  NOR2_X1    g12338(.A1(new_n13360_), .A2(new_n13357_), .ZN(new_n13361_));
  NAND2_X1   g12339(.A1(new_n13361_), .A2(new_n13354_), .ZN(new_n13362_));
  AOI21_X1   g12340(.A1(new_n13347_), .A2(new_n13362_), .B(new_n13217_), .ZN(new_n13363_));
  AOI21_X1   g12341(.A1(new_n11715_), .A2(new_n11716_), .B(new_n11714_), .ZN(new_n13364_));
  NOR3_X1    g12342(.A1(new_n11654_), .A2(new_n11712_), .A3(new_n11692_), .ZN(new_n13365_));
  OAI21_X1   g12343(.A1(new_n13365_), .A2(new_n13364_), .B(new_n9543_), .ZN(new_n13366_));
  NOR3_X1    g12344(.A1(new_n13365_), .A2(new_n13364_), .A3(new_n9543_), .ZN(new_n13367_));
  OAI21_X1   g12345(.A1(new_n11624_), .A2(new_n13367_), .B(new_n13366_), .ZN(new_n13368_));
  OAI22_X1   g12346(.A1(new_n13360_), .A2(new_n13357_), .B1(new_n13271_), .B2(new_n13264_), .ZN(new_n13369_));
  NAND4_X1   g12347(.A1(new_n13338_), .A2(new_n13350_), .A3(new_n13345_), .A4(new_n13353_), .ZN(new_n13370_));
  AOI21_X1   g12348(.A1(new_n13369_), .A2(new_n13370_), .B(new_n13368_), .ZN(new_n13371_));
  NOR2_X1    g12349(.A1(new_n13363_), .A2(new_n13371_), .ZN(new_n13372_));
  NAND3_X1   g12350(.A1(new_n11554_), .A2(new_n11536_), .A3(new_n11420_), .ZN(new_n13373_));
  AOI21_X1   g12351(.A1(new_n11418_), .A2(new_n13373_), .B(new_n11555_), .ZN(new_n13374_));
  OAI21_X1   g12352(.A1(new_n11519_), .A2(new_n11511_), .B(new_n11524_), .ZN(new_n13375_));
  NOR2_X1    g12353(.A1(new_n11449_), .A2(new_n11526_), .ZN(new_n13376_));
  NAND2_X1   g12354(.A1(new_n13375_), .A2(new_n13376_), .ZN(new_n13377_));
  NAND2_X1   g12355(.A1(new_n11549_), .A2(new_n11516_), .ZN(new_n13378_));
  NAND3_X1   g12356(.A1(new_n9150_), .A2(new_n11481_), .A3(new_n11485_), .ZN(new_n13379_));
  NAND2_X1   g12357(.A1(new_n11491_), .A2(new_n11472_), .ZN(new_n13380_));
  AOI21_X1   g12358(.A1(new_n11468_), .A2(new_n13380_), .B(new_n11496_), .ZN(new_n13381_));
  AOI21_X1   g12359(.A1(new_n13379_), .A2(new_n11513_), .B(new_n13381_), .ZN(new_n13382_));
  INV_X1     g12360(.I(new_n13382_), .ZN(new_n13383_));
  NAND3_X1   g12361(.A1(new_n13379_), .A2(new_n11513_), .A3(new_n13381_), .ZN(new_n13384_));
  OAI21_X1   g12362(.A1(new_n11506_), .A2(new_n11475_), .B(new_n11500_), .ZN(new_n13385_));
  AOI22_X1   g12363(.A1(new_n13378_), .A2(new_n13385_), .B1(new_n13383_), .B2(new_n13384_), .ZN(new_n13386_));
  NAND2_X1   g12364(.A1(new_n11464_), .A2(new_n11460_), .ZN(new_n13387_));
  NOR2_X1    g12365(.A1(new_n13387_), .A2(new_n11442_), .ZN(new_n13388_));
  NAND2_X1   g12366(.A1(new_n11459_), .A2(new_n9115_), .ZN(new_n13389_));
  NAND2_X1   g12367(.A1(new_n9087_), .A2(new_n9088_), .ZN(new_n13390_));
  NAND3_X1   g12368(.A1(new_n9181_), .A2(new_n9086_), .A3(new_n13390_), .ZN(new_n13391_));
  NAND2_X1   g12369(.A1(new_n13391_), .A2(new_n11422_), .ZN(new_n13392_));
  XOR2_X1    g12370(.A1(new_n13389_), .A2(new_n13392_), .Z(new_n13393_));
  AOI22_X1   g12371(.A1(new_n11442_), .A2(new_n11444_), .B1(new_n11537_), .B2(new_n11538_), .ZN(new_n13394_));
  OAI21_X1   g12372(.A1(new_n13388_), .A2(new_n13394_), .B(new_n13393_), .ZN(new_n13395_));
  NAND2_X1   g12373(.A1(new_n13386_), .A2(new_n13395_), .ZN(new_n13396_));
  NOR3_X1    g12374(.A1(new_n11504_), .A2(new_n11503_), .A3(new_n9167_), .ZN(new_n13397_));
  INV_X1     g12375(.I(new_n13381_), .ZN(new_n13398_));
  NOR3_X1    g12376(.A1(new_n13397_), .A2(new_n11528_), .A3(new_n13398_), .ZN(new_n13399_));
  AOI21_X1   g12377(.A1(new_n11502_), .A2(new_n11489_), .B(new_n11509_), .ZN(new_n13400_));
  OAI22_X1   g12378(.A1(new_n11530_), .A2(new_n13400_), .B1(new_n13382_), .B2(new_n13399_), .ZN(new_n13401_));
  XNOR2_X1   g12379(.A1(new_n13389_), .A2(new_n13392_), .ZN(new_n13402_));
  OAI22_X1   g12380(.A1(new_n11447_), .A2(new_n11429_), .B1(new_n11425_), .B2(new_n11424_), .ZN(new_n13403_));
  AOI21_X1   g12381(.A1(new_n11465_), .A2(new_n13403_), .B(new_n13402_), .ZN(new_n13404_));
  NAND2_X1   g12382(.A1(new_n13401_), .A2(new_n13404_), .ZN(new_n13405_));
  AOI22_X1   g12383(.A1(new_n13377_), .A2(new_n11552_), .B1(new_n13396_), .B2(new_n13405_), .ZN(new_n13406_));
  AOI21_X1   g12384(.A1(new_n11551_), .A2(new_n11546_), .B(new_n11534_), .ZN(new_n13407_));
  NAND2_X1   g12385(.A1(new_n11542_), .A2(new_n11467_), .ZN(new_n13408_));
  OAI21_X1   g12386(.A1(new_n13407_), .A2(new_n13408_), .B(new_n11552_), .ZN(new_n13409_));
  NOR2_X1    g12387(.A1(new_n13386_), .A2(new_n13404_), .ZN(new_n13410_));
  NOR2_X1    g12388(.A1(new_n13401_), .A2(new_n13395_), .ZN(new_n13411_));
  NOR2_X1    g12389(.A1(new_n13410_), .A2(new_n13411_), .ZN(new_n13412_));
  NOR2_X1    g12390(.A1(new_n13412_), .A2(new_n13409_), .ZN(new_n13413_));
  NOR2_X1    g12391(.A1(new_n13413_), .A2(new_n13406_), .ZN(new_n13414_));
  OAI21_X1   g12392(.A1(new_n11366_), .A2(new_n8993_), .B(new_n11414_), .ZN(new_n13415_));
  AOI21_X1   g12393(.A1(new_n11351_), .A2(new_n11352_), .B(new_n8958_), .ZN(new_n13416_));
  NOR3_X1    g12394(.A1(new_n11349_), .A2(new_n11346_), .A3(new_n9007_), .ZN(new_n13417_));
  NOR2_X1    g12395(.A1(new_n13417_), .A2(new_n13416_), .ZN(new_n13418_));
  NAND4_X1   g12396(.A1(new_n11364_), .A2(new_n11358_), .A3(new_n11359_), .A4(new_n13418_), .ZN(new_n13419_));
  INV_X1     g12397(.I(new_n13419_), .ZN(new_n13420_));
  AOI21_X1   g12398(.A1(new_n13420_), .A2(new_n13415_), .B(new_n11415_), .ZN(new_n13421_));
  NOR3_X1    g12399(.A1(new_n11408_), .A2(new_n11412_), .A3(new_n11380_), .ZN(new_n13422_));
  AOI21_X1   g12400(.A1(new_n11402_), .A2(new_n11398_), .B(new_n8907_), .ZN(new_n13423_));
  NOR3_X1    g12401(.A1(new_n11399_), .A2(new_n11400_), .A3(new_n11397_), .ZN(new_n13424_));
  NOR2_X1    g12402(.A1(new_n13423_), .A2(new_n13424_), .ZN(new_n13425_));
  OAI21_X1   g12403(.A1(new_n11378_), .A2(new_n11377_), .B(new_n11376_), .ZN(new_n13426_));
  NAND3_X1   g12404(.A1(new_n11367_), .A2(new_n11369_), .A3(new_n8986_), .ZN(new_n13427_));
  NAND2_X1   g12405(.A1(new_n13426_), .A2(new_n13427_), .ZN(new_n13428_));
  AOI21_X1   g12406(.A1(new_n11392_), .A2(new_n11395_), .B(new_n13428_), .ZN(new_n13429_));
  NAND2_X1   g12407(.A1(new_n11411_), .A2(new_n11368_), .ZN(new_n13430_));
  INV_X1     g12408(.I(new_n8910_), .ZN(new_n13431_));
  NAND2_X1   g12409(.A1(new_n8908_), .A2(new_n8909_), .ZN(new_n13432_));
  NAND3_X1   g12410(.A1(new_n11390_), .A2(new_n8907_), .A3(new_n13432_), .ZN(new_n13433_));
  NAND2_X1   g12411(.A1(new_n13433_), .A2(new_n13431_), .ZN(new_n13434_));
  NAND2_X1   g12412(.A1(new_n13430_), .A2(new_n13434_), .ZN(new_n13435_));
  INV_X1     g12413(.I(new_n13435_), .ZN(new_n13436_));
  OAI21_X1   g12414(.A1(new_n13429_), .A2(new_n13425_), .B(new_n13436_), .ZN(new_n13437_));
  NAND2_X1   g12415(.A1(new_n11394_), .A2(new_n9014_), .ZN(new_n13438_));
  NAND2_X1   g12416(.A1(new_n13438_), .A2(new_n11409_), .ZN(new_n13439_));
  OAI21_X1   g12417(.A1(new_n11408_), .A2(new_n13439_), .B(new_n11380_), .ZN(new_n13440_));
  NAND3_X1   g12418(.A1(new_n13440_), .A2(new_n11404_), .A3(new_n13435_), .ZN(new_n13441_));
  AOI21_X1   g12419(.A1(new_n13437_), .A2(new_n13441_), .B(new_n13422_), .ZN(new_n13442_));
  INV_X1     g12420(.I(new_n13422_), .ZN(new_n13443_));
  AOI21_X1   g12421(.A1(new_n13440_), .A2(new_n11404_), .B(new_n13435_), .ZN(new_n13444_));
  NOR3_X1    g12422(.A1(new_n13429_), .A2(new_n13425_), .A3(new_n13436_), .ZN(new_n13445_));
  NOR3_X1    g12423(.A1(new_n13445_), .A2(new_n13444_), .A3(new_n13443_), .ZN(new_n13446_));
  NOR2_X1    g12424(.A1(new_n13446_), .A2(new_n13442_), .ZN(new_n13447_));
  NAND2_X1   g12425(.A1(new_n11329_), .A2(new_n11330_), .ZN(new_n13448_));
  NAND2_X1   g12426(.A1(new_n11332_), .A2(new_n11331_), .ZN(new_n13449_));
  NAND2_X1   g12427(.A1(new_n13448_), .A2(new_n13449_), .ZN(new_n13450_));
  OAI21_X1   g12428(.A1(new_n13450_), .A2(new_n11336_), .B(new_n13418_), .ZN(new_n13451_));
  NAND2_X1   g12429(.A1(new_n11361_), .A2(new_n11345_), .ZN(new_n13452_));
  NAND2_X1   g12430(.A1(new_n8934_), .A2(new_n8935_), .ZN(new_n13453_));
  NAND3_X1   g12431(.A1(new_n8922_), .A2(new_n8933_), .A3(new_n13453_), .ZN(new_n13454_));
  NAND2_X1   g12432(.A1(new_n13454_), .A2(new_n11321_), .ZN(new_n13455_));
  NAND2_X1   g12433(.A1(new_n13455_), .A2(new_n13452_), .ZN(new_n13456_));
  AOI21_X1   g12434(.A1(new_n13451_), .A2(new_n11328_), .B(new_n13456_), .ZN(new_n13457_));
  AOI21_X1   g12435(.A1(new_n11337_), .A2(new_n11333_), .B(new_n11354_), .ZN(new_n13458_));
  INV_X1     g12436(.I(new_n13456_), .ZN(new_n13459_));
  NOR3_X1    g12437(.A1(new_n13458_), .A2(new_n13459_), .A3(new_n11359_), .ZN(new_n13460_));
  OAI21_X1   g12438(.A1(new_n13457_), .A2(new_n13460_), .B(new_n11363_), .ZN(new_n13461_));
  INV_X1     g12439(.I(new_n11363_), .ZN(new_n13462_));
  OAI21_X1   g12440(.A1(new_n13458_), .A2(new_n11359_), .B(new_n13459_), .ZN(new_n13463_));
  NAND3_X1   g12441(.A1(new_n13451_), .A2(new_n11328_), .A3(new_n13456_), .ZN(new_n13464_));
  NAND3_X1   g12442(.A1(new_n13464_), .A2(new_n13463_), .A3(new_n13462_), .ZN(new_n13465_));
  NAND2_X1   g12443(.A1(new_n13461_), .A2(new_n13465_), .ZN(new_n13466_));
  NAND2_X1   g12444(.A1(new_n13447_), .A2(new_n13466_), .ZN(new_n13467_));
  OAI21_X1   g12445(.A1(new_n13445_), .A2(new_n13444_), .B(new_n13443_), .ZN(new_n13468_));
  NAND3_X1   g12446(.A1(new_n13437_), .A2(new_n13441_), .A3(new_n13422_), .ZN(new_n13469_));
  NAND2_X1   g12447(.A1(new_n13468_), .A2(new_n13469_), .ZN(new_n13470_));
  AOI21_X1   g12448(.A1(new_n13464_), .A2(new_n13463_), .B(new_n13462_), .ZN(new_n13471_));
  NOR3_X1    g12449(.A1(new_n13457_), .A2(new_n13460_), .A3(new_n11363_), .ZN(new_n13472_));
  NOR2_X1    g12450(.A1(new_n13472_), .A2(new_n13471_), .ZN(new_n13473_));
  NAND2_X1   g12451(.A1(new_n13470_), .A2(new_n13473_), .ZN(new_n13474_));
  AOI21_X1   g12452(.A1(new_n13474_), .A2(new_n13467_), .B(new_n13421_), .ZN(new_n13475_));
  XOR2_X1    g12453(.A1(new_n8911_), .A2(new_n9001_), .Z(new_n13476_));
  NOR2_X1    g12454(.A1(new_n11408_), .A2(new_n13439_), .ZN(new_n13477_));
  NOR3_X1    g12455(.A1(new_n13477_), .A2(new_n13425_), .A3(new_n13428_), .ZN(new_n13478_));
  NAND3_X1   g12456(.A1(new_n13478_), .A2(new_n13476_), .A3(new_n9018_), .ZN(new_n13479_));
  AOI21_X1   g12457(.A1(new_n13476_), .A2(new_n9018_), .B(new_n13478_), .ZN(new_n13480_));
  OAI21_X1   g12458(.A1(new_n13480_), .A2(new_n13419_), .B(new_n13479_), .ZN(new_n13481_));
  NAND2_X1   g12459(.A1(new_n13470_), .A2(new_n13466_), .ZN(new_n13482_));
  NAND4_X1   g12460(.A1(new_n13468_), .A2(new_n13469_), .A3(new_n13461_), .A4(new_n13465_), .ZN(new_n13483_));
  AOI21_X1   g12461(.A1(new_n13482_), .A2(new_n13483_), .B(new_n13481_), .ZN(new_n13484_));
  OAI21_X1   g12462(.A1(new_n13475_), .A2(new_n13484_), .B(new_n13414_), .ZN(new_n13485_));
  NOR3_X1    g12463(.A1(new_n11519_), .A2(new_n11511_), .A3(new_n11524_), .ZN(new_n13486_));
  NOR2_X1    g12464(.A1(new_n13407_), .A2(new_n13408_), .ZN(new_n13487_));
  NOR2_X1    g12465(.A1(new_n13401_), .A2(new_n13404_), .ZN(new_n13488_));
  NOR2_X1    g12466(.A1(new_n13386_), .A2(new_n13395_), .ZN(new_n13489_));
  OAI22_X1   g12467(.A1(new_n13487_), .A2(new_n13486_), .B1(new_n13489_), .B2(new_n13488_), .ZN(new_n13490_));
  AOI21_X1   g12468(.A1(new_n13375_), .A2(new_n13376_), .B(new_n13486_), .ZN(new_n13491_));
  NAND2_X1   g12469(.A1(new_n13401_), .A2(new_n13395_), .ZN(new_n13492_));
  NAND2_X1   g12470(.A1(new_n13386_), .A2(new_n13404_), .ZN(new_n13493_));
  NAND2_X1   g12471(.A1(new_n13493_), .A2(new_n13492_), .ZN(new_n13494_));
  NAND2_X1   g12472(.A1(new_n13494_), .A2(new_n13491_), .ZN(new_n13495_));
  NAND2_X1   g12473(.A1(new_n13495_), .A2(new_n13490_), .ZN(new_n13496_));
  NOR2_X1    g12474(.A1(new_n13470_), .A2(new_n13473_), .ZN(new_n13497_));
  NOR2_X1    g12475(.A1(new_n13447_), .A2(new_n13466_), .ZN(new_n13498_));
  OAI21_X1   g12476(.A1(new_n13497_), .A2(new_n13498_), .B(new_n13481_), .ZN(new_n13499_));
  AOI22_X1   g12477(.A1(new_n13468_), .A2(new_n13469_), .B1(new_n13461_), .B2(new_n13465_), .ZN(new_n13500_));
  NOR4_X1    g12478(.A1(new_n13442_), .A2(new_n13446_), .A3(new_n13472_), .A4(new_n13471_), .ZN(new_n13501_));
  OAI21_X1   g12479(.A1(new_n13501_), .A2(new_n13500_), .B(new_n13421_), .ZN(new_n13502_));
  NAND3_X1   g12480(.A1(new_n13496_), .A2(new_n13499_), .A3(new_n13502_), .ZN(new_n13503_));
  AOI21_X1   g12481(.A1(new_n13485_), .A2(new_n13503_), .B(new_n13374_), .ZN(new_n13504_));
  AOI21_X1   g12482(.A1(new_n11553_), .A2(new_n11543_), .B(new_n11542_), .ZN(new_n13505_));
  NOR3_X1    g12483(.A1(new_n11535_), .A2(new_n11449_), .A3(new_n11525_), .ZN(new_n13506_));
  OAI21_X1   g12484(.A1(new_n13505_), .A2(new_n13506_), .B(new_n9193_), .ZN(new_n13507_));
  NOR3_X1    g12485(.A1(new_n13505_), .A2(new_n13506_), .A3(new_n9193_), .ZN(new_n13508_));
  OAI21_X1   g12486(.A1(new_n11419_), .A2(new_n13508_), .B(new_n13507_), .ZN(new_n13509_));
  OAI22_X1   g12487(.A1(new_n13475_), .A2(new_n13484_), .B1(new_n13406_), .B2(new_n13413_), .ZN(new_n13510_));
  NAND3_X1   g12488(.A1(new_n13414_), .A2(new_n13499_), .A3(new_n13502_), .ZN(new_n13511_));
  AOI21_X1   g12489(.A1(new_n13510_), .A2(new_n13511_), .B(new_n13509_), .ZN(new_n13512_));
  OAI21_X1   g12490(.A1(new_n13504_), .A2(new_n13512_), .B(new_n13372_), .ZN(new_n13513_));
  NOR2_X1    g12491(.A1(new_n13361_), .A2(new_n13354_), .ZN(new_n13514_));
  NOR2_X1    g12492(.A1(new_n13346_), .A2(new_n13272_), .ZN(new_n13515_));
  OAI21_X1   g12493(.A1(new_n13515_), .A2(new_n13514_), .B(new_n13368_), .ZN(new_n13516_));
  AOI22_X1   g12494(.A1(new_n13338_), .A2(new_n13345_), .B1(new_n13350_), .B2(new_n13353_), .ZN(new_n13517_));
  NOR4_X1    g12495(.A1(new_n13360_), .A2(new_n13271_), .A3(new_n13357_), .A4(new_n13264_), .ZN(new_n13518_));
  OAI21_X1   g12496(.A1(new_n13517_), .A2(new_n13518_), .B(new_n13217_), .ZN(new_n13519_));
  NAND2_X1   g12497(.A1(new_n13516_), .A2(new_n13519_), .ZN(new_n13520_));
  AOI21_X1   g12498(.A1(new_n13499_), .A2(new_n13502_), .B(new_n13496_), .ZN(new_n13521_));
  NOR3_X1    g12499(.A1(new_n13414_), .A2(new_n13475_), .A3(new_n13484_), .ZN(new_n13522_));
  OAI21_X1   g12500(.A1(new_n13521_), .A2(new_n13522_), .B(new_n13509_), .ZN(new_n13523_));
  AOI22_X1   g12501(.A1(new_n13499_), .A2(new_n13502_), .B1(new_n13490_), .B2(new_n13495_), .ZN(new_n13524_));
  NOR3_X1    g12502(.A1(new_n13496_), .A2(new_n13475_), .A3(new_n13484_), .ZN(new_n13525_));
  OAI21_X1   g12503(.A1(new_n13524_), .A2(new_n13525_), .B(new_n13374_), .ZN(new_n13526_));
  NAND3_X1   g12504(.A1(new_n13520_), .A2(new_n13523_), .A3(new_n13526_), .ZN(new_n13527_));
  AOI21_X1   g12505(.A1(new_n13513_), .A2(new_n13527_), .B(new_n13215_), .ZN(new_n13528_));
  NAND2_X1   g12506(.A1(new_n11719_), .A2(new_n11723_), .ZN(new_n13529_));
  NAND2_X1   g12507(.A1(new_n13529_), .A2(new_n9547_), .ZN(new_n13530_));
  NAND2_X1   g12508(.A1(new_n13214_), .A2(new_n11726_), .ZN(new_n13531_));
  NAND2_X1   g12509(.A1(new_n13531_), .A2(new_n13530_), .ZN(new_n13532_));
  OAI21_X1   g12510(.A1(new_n13504_), .A2(new_n13512_), .B(new_n13520_), .ZN(new_n13533_));
  NAND3_X1   g12511(.A1(new_n13372_), .A2(new_n13523_), .A3(new_n13526_), .ZN(new_n13534_));
  AOI21_X1   g12512(.A1(new_n13533_), .A2(new_n13534_), .B(new_n13532_), .ZN(new_n13535_));
  NOR2_X1    g12513(.A1(new_n13528_), .A2(new_n13535_), .ZN(new_n13536_));
  NAND3_X1   g12514(.A1(new_n8885_), .A2(new_n11312_), .A3(new_n11316_), .ZN(new_n13537_));
  NAND2_X1   g12515(.A1(new_n13537_), .A2(new_n11161_), .ZN(new_n13538_));
  NAND2_X1   g12516(.A1(new_n13538_), .A2(new_n11318_), .ZN(new_n13539_));
  NAND3_X1   g12517(.A1(new_n8378_), .A2(new_n8391_), .A3(new_n8564_), .ZN(new_n13540_));
  AOI21_X1   g12518(.A1(new_n11309_), .A2(new_n11303_), .B(new_n11308_), .ZN(new_n13541_));
  NOR3_X1    g12519(.A1(new_n11304_), .A2(new_n11261_), .A3(new_n11302_), .ZN(new_n13542_));
  NOR2_X1    g12520(.A1(new_n13541_), .A2(new_n13542_), .ZN(new_n13543_));
  AOI21_X1   g12521(.A1(new_n13543_), .A2(new_n13540_), .B(new_n11241_), .ZN(new_n13544_));
  NOR2_X1    g12522(.A1(new_n8545_), .A2(new_n8528_), .ZN(new_n13545_));
  NAND2_X1   g12523(.A1(new_n8486_), .A2(new_n8541_), .ZN(new_n13546_));
  NAND2_X1   g12524(.A1(new_n8497_), .A2(new_n8535_), .ZN(new_n13547_));
  AOI21_X1   g12525(.A1(new_n13546_), .A2(new_n13547_), .B(new_n8500_), .ZN(new_n13548_));
  NOR3_X1    g12526(.A1(new_n13548_), .A2(new_n11278_), .A3(new_n11281_), .ZN(new_n13549_));
  NOR2_X1    g12527(.A1(new_n8512_), .A2(new_n8526_), .ZN(new_n13550_));
  NOR2_X1    g12528(.A1(new_n8551_), .A2(new_n8527_), .ZN(new_n13551_));
  NOR3_X1    g12529(.A1(new_n13551_), .A2(new_n13550_), .A3(new_n8557_), .ZN(new_n13552_));
  NOR2_X1    g12530(.A1(new_n11289_), .A2(new_n13552_), .ZN(new_n13553_));
  AOI22_X1   g12531(.A1(new_n8506_), .A2(new_n8511_), .B1(new_n8517_), .B2(new_n8522_), .ZN(new_n13554_));
  OAI22_X1   g12532(.A1(new_n13554_), .A2(new_n11294_), .B1(new_n11298_), .B2(new_n8557_), .ZN(new_n13555_));
  NOR4_X1    g12533(.A1(new_n13555_), .A2(new_n8486_), .A3(new_n8497_), .A4(new_n8500_), .ZN(new_n13556_));
  NOR4_X1    g12534(.A1(new_n13549_), .A2(new_n13556_), .A3(new_n13553_), .A4(new_n13545_), .ZN(new_n13557_));
  NOR2_X1    g12535(.A1(new_n13557_), .A2(new_n11274_), .ZN(new_n13558_));
  OAI22_X1   g12536(.A1(new_n8464_), .A2(new_n8466_), .B1(new_n8472_), .B2(new_n8470_), .ZN(new_n13559_));
  NAND4_X1   g12537(.A1(new_n8422_), .A2(new_n8427_), .A3(new_n8433_), .A4(new_n8438_), .ZN(new_n13560_));
  AOI21_X1   g12538(.A1(new_n8422_), .A2(new_n8427_), .B(new_n8442_), .ZN(new_n13561_));
  AOI22_X1   g12539(.A1(new_n13559_), .A2(new_n13560_), .B1(new_n8439_), .B2(new_n13561_), .ZN(new_n13562_));
  NAND4_X1   g12540(.A1(new_n13562_), .A2(new_n8451_), .A3(new_n8457_), .A4(new_n8460_), .ZN(new_n13563_));
  NOR2_X1    g12541(.A1(new_n13563_), .A2(new_n11248_), .ZN(new_n13564_));
  NAND4_X1   g12542(.A1(new_n13564_), .A2(new_n11248_), .A3(new_n11306_), .A4(new_n11259_), .ZN(new_n13565_));
  OAI21_X1   g12543(.A1(new_n13558_), .A2(new_n13565_), .B(new_n11301_), .ZN(new_n13566_));
  NAND2_X1   g12544(.A1(new_n8542_), .A2(new_n8543_), .ZN(new_n13567_));
  NAND3_X1   g12545(.A1(new_n8535_), .A2(new_n8541_), .A3(new_n13567_), .ZN(new_n13568_));
  NOR2_X1    g12546(.A1(new_n8524_), .A2(new_n8510_), .ZN(new_n13569_));
  NAND2_X1   g12547(.A1(new_n13569_), .A2(new_n11297_), .ZN(new_n13570_));
  NAND3_X1   g12548(.A1(new_n8512_), .A2(new_n8523_), .A3(new_n13570_), .ZN(new_n13571_));
  NAND2_X1   g12549(.A1(new_n13571_), .A2(new_n8526_), .ZN(new_n13572_));
  NAND3_X1   g12550(.A1(new_n13572_), .A2(new_n8500_), .A3(new_n13568_), .ZN(new_n13573_));
  NAND2_X1   g12551(.A1(new_n13568_), .A2(new_n8500_), .ZN(new_n13574_));
  NAND3_X1   g12552(.A1(new_n13574_), .A2(new_n8526_), .A3(new_n13571_), .ZN(new_n13575_));
  NAND2_X1   g12553(.A1(new_n13573_), .A2(new_n13575_), .ZN(new_n13576_));
  OAI21_X1   g12554(.A1(new_n11280_), .A2(new_n11279_), .B(new_n8497_), .ZN(new_n13577_));
  NAND3_X1   g12555(.A1(new_n11276_), .A2(new_n11277_), .A3(new_n8541_), .ZN(new_n13578_));
  NAND3_X1   g12556(.A1(new_n11285_), .A2(new_n13577_), .A3(new_n13578_), .ZN(new_n13579_));
  AOI21_X1   g12557(.A1(new_n13579_), .A2(new_n11275_), .B(new_n13553_), .ZN(new_n13580_));
  OAI21_X1   g12558(.A1(new_n13580_), .A2(new_n13556_), .B(new_n13576_), .ZN(new_n13581_));
  NAND2_X1   g12559(.A1(new_n8458_), .A2(new_n8459_), .ZN(new_n13582_));
  NAND3_X1   g12560(.A1(new_n8451_), .A2(new_n8457_), .A3(new_n13582_), .ZN(new_n13583_));
  NAND2_X1   g12561(.A1(new_n13583_), .A2(new_n8416_), .ZN(new_n13584_));
  NOR2_X1    g12562(.A1(new_n8440_), .A2(new_n8426_), .ZN(new_n13585_));
  NAND2_X1   g12563(.A1(new_n13585_), .A2(new_n11267_), .ZN(new_n13586_));
  AOI21_X1   g12564(.A1(new_n11265_), .A2(new_n13586_), .B(new_n8443_), .ZN(new_n13587_));
  XOR2_X1    g12565(.A1(new_n13584_), .A2(new_n13587_), .Z(new_n13588_));
  NAND2_X1   g12566(.A1(new_n11252_), .A2(new_n11255_), .ZN(new_n13589_));
  NAND2_X1   g12567(.A1(new_n8402_), .A2(new_n8457_), .ZN(new_n13590_));
  NAND2_X1   g12568(.A1(new_n8413_), .A2(new_n8451_), .ZN(new_n13591_));
  AOI21_X1   g12569(.A1(new_n13590_), .A2(new_n13591_), .B(new_n8416_), .ZN(new_n13592_));
  OAI21_X1   g12570(.A1(new_n13589_), .A2(new_n13592_), .B(new_n11249_), .ZN(new_n13593_));
  NAND2_X1   g12571(.A1(new_n13593_), .A2(new_n11264_), .ZN(new_n13594_));
  AOI21_X1   g12572(.A1(new_n13594_), .A2(new_n13563_), .B(new_n13588_), .ZN(new_n13595_));
  NOR2_X1    g12573(.A1(new_n13595_), .A2(new_n13581_), .ZN(new_n13596_));
  INV_X1     g12574(.I(new_n13555_), .ZN(new_n13597_));
  NAND4_X1   g12575(.A1(new_n13597_), .A2(new_n8535_), .A3(new_n8541_), .A4(new_n8544_), .ZN(new_n13598_));
  XNOR2_X1   g12576(.A1(new_n13574_), .A2(new_n13572_), .ZN(new_n13599_));
  NAND2_X1   g12577(.A1(new_n13577_), .A2(new_n13578_), .ZN(new_n13600_));
  OAI21_X1   g12578(.A1(new_n13600_), .A2(new_n13548_), .B(new_n11275_), .ZN(new_n13601_));
  NAND2_X1   g12579(.A1(new_n13601_), .A2(new_n11292_), .ZN(new_n13602_));
  AOI21_X1   g12580(.A1(new_n13602_), .A2(new_n13598_), .B(new_n13599_), .ZN(new_n13603_));
  NOR2_X1    g12581(.A1(new_n8402_), .A2(new_n8413_), .ZN(new_n13604_));
  AOI21_X1   g12582(.A1(new_n13604_), .A2(new_n13582_), .B(new_n8460_), .ZN(new_n13605_));
  NAND2_X1   g12583(.A1(new_n11265_), .A2(new_n13586_), .ZN(new_n13606_));
  NAND2_X1   g12584(.A1(new_n13606_), .A2(new_n8442_), .ZN(new_n13607_));
  NAND2_X1   g12585(.A1(new_n13607_), .A2(new_n13605_), .ZN(new_n13608_));
  NAND2_X1   g12586(.A1(new_n13584_), .A2(new_n13587_), .ZN(new_n13609_));
  NAND2_X1   g12587(.A1(new_n13608_), .A2(new_n13609_), .ZN(new_n13610_));
  AOI21_X1   g12588(.A1(new_n11259_), .A2(new_n11249_), .B(new_n11248_), .ZN(new_n13611_));
  OAI21_X1   g12589(.A1(new_n13611_), .A2(new_n11271_), .B(new_n13610_), .ZN(new_n13612_));
  NOR2_X1    g12590(.A1(new_n13603_), .A2(new_n13612_), .ZN(new_n13613_));
  OAI21_X1   g12591(.A1(new_n13613_), .A2(new_n13596_), .B(new_n13566_), .ZN(new_n13614_));
  NOR2_X1    g12592(.A1(new_n13579_), .A2(new_n13545_), .ZN(new_n13615_));
  INV_X1     g12593(.I(new_n11300_), .ZN(new_n13616_));
  NOR4_X1    g12594(.A1(new_n8563_), .A2(new_n13615_), .A3(new_n13616_), .A4(new_n13553_), .ZN(new_n13617_));
  NAND3_X1   g12595(.A1(new_n11286_), .A2(new_n11292_), .A3(new_n11300_), .ZN(new_n13618_));
  NAND2_X1   g12596(.A1(new_n13618_), .A2(new_n8563_), .ZN(new_n13619_));
  INV_X1     g12597(.I(new_n11259_), .ZN(new_n13620_));
  NOR4_X1    g12598(.A1(new_n11272_), .A2(new_n13620_), .A3(new_n11264_), .A4(new_n11249_), .ZN(new_n13621_));
  AOI21_X1   g12599(.A1(new_n13619_), .A2(new_n13621_), .B(new_n13617_), .ZN(new_n13622_));
  NAND2_X1   g12600(.A1(new_n13581_), .A2(new_n13612_), .ZN(new_n13623_));
  INV_X1     g12601(.I(new_n13623_), .ZN(new_n13624_));
  NOR2_X1    g12602(.A1(new_n13581_), .A2(new_n13612_), .ZN(new_n13625_));
  OAI21_X1   g12603(.A1(new_n13624_), .A2(new_n13625_), .B(new_n13622_), .ZN(new_n13626_));
  NAND2_X1   g12604(.A1(new_n13626_), .A2(new_n13614_), .ZN(new_n13627_));
  NOR4_X1    g12605(.A1(new_n8386_), .A2(new_n8274_), .A3(new_n8262_), .A4(new_n8389_), .ZN(new_n13628_));
  OAI21_X1   g12606(.A1(new_n11211_), .A2(new_n11209_), .B(new_n11208_), .ZN(new_n13629_));
  NAND3_X1   g12607(.A1(new_n11205_), .A2(new_n11206_), .A3(new_n11202_), .ZN(new_n13630_));
  NAND2_X1   g12608(.A1(new_n13629_), .A2(new_n13630_), .ZN(new_n13631_));
  INV_X1     g12609(.I(new_n11222_), .ZN(new_n13632_));
  NAND2_X1   g12610(.A1(new_n8224_), .A2(new_n11200_), .ZN(new_n13633_));
  NOR2_X1    g12611(.A1(new_n11223_), .A2(new_n8256_), .ZN(new_n13634_));
  AOI21_X1   g12612(.A1(new_n8256_), .A2(new_n11224_), .B(new_n13634_), .ZN(new_n13635_));
  NOR2_X1    g12613(.A1(new_n8273_), .A2(new_n11197_), .ZN(new_n13636_));
  NAND2_X1   g12614(.A1(new_n13636_), .A2(new_n8389_), .ZN(new_n13637_));
  NOR3_X1    g12615(.A1(new_n13635_), .A2(new_n13633_), .A3(new_n13637_), .ZN(new_n13638_));
  NOR4_X1    g12616(.A1(new_n13638_), .A2(new_n13628_), .A3(new_n13631_), .A4(new_n13632_), .ZN(new_n13639_));
  NAND2_X1   g12617(.A1(new_n8235_), .A2(new_n8356_), .ZN(new_n13640_));
  NAND2_X1   g12618(.A1(new_n8372_), .A2(new_n8390_), .ZN(new_n13641_));
  NAND2_X1   g12619(.A1(new_n8316_), .A2(new_n8275_), .ZN(new_n13642_));
  NAND2_X1   g12620(.A1(new_n11233_), .A2(new_n8362_), .ZN(new_n13643_));
  AOI22_X1   g12621(.A1(new_n13640_), .A2(new_n13641_), .B1(new_n13642_), .B2(new_n13643_), .ZN(new_n13644_));
  NAND2_X1   g12622(.A1(new_n13639_), .A2(new_n13644_), .ZN(new_n13645_));
  NOR2_X1    g12623(.A1(new_n13639_), .A2(new_n13644_), .ZN(new_n13646_));
  NAND4_X1   g12624(.A1(new_n11194_), .A2(new_n11186_), .A3(new_n11169_), .A4(new_n11180_), .ZN(new_n13647_));
  OAI21_X1   g12625(.A1(new_n13647_), .A2(new_n13646_), .B(new_n13645_), .ZN(new_n13648_));
  NAND2_X1   g12626(.A1(new_n11201_), .A2(new_n11213_), .ZN(new_n13649_));
  NAND2_X1   g12627(.A1(new_n11227_), .A2(new_n11203_), .ZN(new_n13650_));
  NOR2_X1    g12628(.A1(new_n11215_), .A2(new_n11216_), .ZN(new_n13651_));
  OAI21_X1   g12629(.A1(new_n8379_), .A2(new_n13651_), .B(new_n8388_), .ZN(new_n13652_));
  NAND2_X1   g12630(.A1(new_n13650_), .A2(new_n13652_), .ZN(new_n13653_));
  AOI21_X1   g12631(.A1(new_n13649_), .A2(new_n11222_), .B(new_n13653_), .ZN(new_n13654_));
  OAI21_X1   g12632(.A1(new_n13628_), .A2(new_n13631_), .B(new_n11222_), .ZN(new_n13655_));
  INV_X1     g12633(.I(new_n13653_), .ZN(new_n13656_));
  NOR2_X1    g12634(.A1(new_n13655_), .A2(new_n13656_), .ZN(new_n13657_));
  OAI21_X1   g12635(.A1(new_n13654_), .A2(new_n13657_), .B(new_n11229_), .ZN(new_n13658_));
  NAND2_X1   g12636(.A1(new_n13655_), .A2(new_n13656_), .ZN(new_n13659_));
  NAND3_X1   g12637(.A1(new_n13649_), .A2(new_n11222_), .A3(new_n13653_), .ZN(new_n13660_));
  NAND3_X1   g12638(.A1(new_n13660_), .A2(new_n13659_), .A3(new_n13638_), .ZN(new_n13661_));
  NAND2_X1   g12639(.A1(new_n13658_), .A2(new_n13661_), .ZN(new_n13662_));
  NAND2_X1   g12640(.A1(new_n8315_), .A2(new_n8365_), .ZN(new_n13663_));
  NOR2_X1    g12641(.A1(new_n11187_), .A2(new_n8358_), .ZN(new_n13664_));
  AOI21_X1   g12642(.A1(new_n8358_), .A2(new_n11188_), .B(new_n13664_), .ZN(new_n13665_));
  NOR4_X1    g12643(.A1(new_n13665_), .A2(new_n8371_), .A3(new_n13663_), .A4(new_n11191_), .ZN(new_n13666_));
  OAI21_X1   g12644(.A1(new_n11169_), .A2(new_n11185_), .B(new_n11168_), .ZN(new_n13667_));
  AOI21_X1   g12645(.A1(new_n8314_), .A2(new_n8301_), .B(new_n11171_), .ZN(new_n13668_));
  NAND2_X1   g12646(.A1(new_n8368_), .A2(new_n8369_), .ZN(new_n13669_));
  AOI21_X1   g12647(.A1(new_n8363_), .A2(new_n13669_), .B(new_n8370_), .ZN(new_n13670_));
  NOR2_X1    g12648(.A1(new_n13670_), .A2(new_n13668_), .ZN(new_n13671_));
  NAND2_X1   g12649(.A1(new_n13667_), .A2(new_n13671_), .ZN(new_n13672_));
  NAND4_X1   g12650(.A1(new_n8315_), .A2(new_n8365_), .A3(new_n8303_), .A4(new_n8371_), .ZN(new_n13673_));
  NAND2_X1   g12651(.A1(new_n13673_), .A2(new_n11180_), .ZN(new_n13674_));
  INV_X1     g12652(.I(new_n13671_), .ZN(new_n13675_));
  NAND3_X1   g12653(.A1(new_n13674_), .A2(new_n11168_), .A3(new_n13675_), .ZN(new_n13676_));
  AOI21_X1   g12654(.A1(new_n13672_), .A2(new_n13676_), .B(new_n13666_), .ZN(new_n13677_));
  AOI21_X1   g12655(.A1(new_n13674_), .A2(new_n11168_), .B(new_n13675_), .ZN(new_n13678_));
  NOR2_X1    g12656(.A1(new_n13667_), .A2(new_n13671_), .ZN(new_n13679_));
  NOR3_X1    g12657(.A1(new_n13679_), .A2(new_n13678_), .A3(new_n11193_), .ZN(new_n13680_));
  NOR2_X1    g12658(.A1(new_n13680_), .A2(new_n13677_), .ZN(new_n13681_));
  NOR2_X1    g12659(.A1(new_n13681_), .A2(new_n13662_), .ZN(new_n13682_));
  AOI21_X1   g12660(.A1(new_n13660_), .A2(new_n13659_), .B(new_n13638_), .ZN(new_n13683_));
  NOR3_X1    g12661(.A1(new_n13654_), .A2(new_n13657_), .A3(new_n11229_), .ZN(new_n13684_));
  NOR2_X1    g12662(.A1(new_n13684_), .A2(new_n13683_), .ZN(new_n13685_));
  OAI21_X1   g12663(.A1(new_n13679_), .A2(new_n13678_), .B(new_n11193_), .ZN(new_n13686_));
  NAND3_X1   g12664(.A1(new_n13672_), .A2(new_n13676_), .A3(new_n13666_), .ZN(new_n13687_));
  NAND2_X1   g12665(.A1(new_n13686_), .A2(new_n13687_), .ZN(new_n13688_));
  NOR2_X1    g12666(.A1(new_n13685_), .A2(new_n13688_), .ZN(new_n13689_));
  OAI21_X1   g12667(.A1(new_n13682_), .A2(new_n13689_), .B(new_n13648_), .ZN(new_n13690_));
  NAND2_X1   g12668(.A1(new_n11236_), .A2(new_n11230_), .ZN(new_n13691_));
  NAND2_X1   g12669(.A1(new_n13666_), .A2(new_n11168_), .ZN(new_n13692_));
  NOR4_X1    g12670(.A1(new_n13692_), .A2(new_n11168_), .A3(new_n13673_), .A4(new_n11185_), .ZN(new_n13693_));
  AOI21_X1   g12671(.A1(new_n13693_), .A2(new_n13691_), .B(new_n11237_), .ZN(new_n13694_));
  AOI22_X1   g12672(.A1(new_n13658_), .A2(new_n13661_), .B1(new_n13686_), .B2(new_n13687_), .ZN(new_n13695_));
  NOR4_X1    g12673(.A1(new_n13683_), .A2(new_n13684_), .A3(new_n13680_), .A4(new_n13677_), .ZN(new_n13696_));
  OAI21_X1   g12674(.A1(new_n13696_), .A2(new_n13695_), .B(new_n13694_), .ZN(new_n13697_));
  AOI21_X1   g12675(.A1(new_n13690_), .A2(new_n13697_), .B(new_n13627_), .ZN(new_n13698_));
  NAND2_X1   g12676(.A1(new_n13603_), .A2(new_n13612_), .ZN(new_n13699_));
  NAND2_X1   g12677(.A1(new_n13595_), .A2(new_n13581_), .ZN(new_n13700_));
  AOI21_X1   g12678(.A1(new_n13699_), .A2(new_n13700_), .B(new_n13622_), .ZN(new_n13701_));
  NAND2_X1   g12679(.A1(new_n13603_), .A2(new_n13595_), .ZN(new_n13702_));
  AOI21_X1   g12680(.A1(new_n13702_), .A2(new_n13623_), .B(new_n13566_), .ZN(new_n13703_));
  NOR2_X1    g12681(.A1(new_n13701_), .A2(new_n13703_), .ZN(new_n13704_));
  NAND2_X1   g12682(.A1(new_n13685_), .A2(new_n13688_), .ZN(new_n13705_));
  NAND2_X1   g12683(.A1(new_n13681_), .A2(new_n13662_), .ZN(new_n13706_));
  AOI21_X1   g12684(.A1(new_n13706_), .A2(new_n13705_), .B(new_n13694_), .ZN(new_n13707_));
  NAND2_X1   g12685(.A1(new_n13662_), .A2(new_n13688_), .ZN(new_n13708_));
  NAND4_X1   g12686(.A1(new_n13658_), .A2(new_n13661_), .A3(new_n13686_), .A4(new_n13687_), .ZN(new_n13709_));
  AOI21_X1   g12687(.A1(new_n13708_), .A2(new_n13709_), .B(new_n13648_), .ZN(new_n13710_));
  NOR3_X1    g12688(.A1(new_n13707_), .A2(new_n13710_), .A3(new_n13704_), .ZN(new_n13711_));
  OAI21_X1   g12689(.A1(new_n13711_), .A2(new_n13698_), .B(new_n13544_), .ZN(new_n13712_));
  OAI21_X1   g12690(.A1(new_n11311_), .A2(new_n8566_), .B(new_n11315_), .ZN(new_n13713_));
  AOI21_X1   g12691(.A1(new_n13690_), .A2(new_n13697_), .B(new_n13704_), .ZN(new_n13714_));
  NOR3_X1    g12692(.A1(new_n13707_), .A2(new_n13710_), .A3(new_n13627_), .ZN(new_n13715_));
  OAI21_X1   g12693(.A1(new_n13715_), .A2(new_n13714_), .B(new_n13713_), .ZN(new_n13716_));
  NAND2_X1   g12694(.A1(new_n13712_), .A2(new_n13716_), .ZN(new_n13717_));
  NAND3_X1   g12695(.A1(new_n11159_), .A2(new_n11142_), .A3(new_n11033_), .ZN(new_n13718_));
  AOI21_X1   g12696(.A1(new_n11031_), .A2(new_n13718_), .B(new_n11160_), .ZN(new_n13719_));
  OAI21_X1   g12697(.A1(new_n11129_), .A2(new_n11121_), .B(new_n11132_), .ZN(new_n13720_));
  NOR2_X1    g12698(.A1(new_n11062_), .A2(new_n11134_), .ZN(new_n13721_));
  NAND2_X1   g12699(.A1(new_n13720_), .A2(new_n13721_), .ZN(new_n13722_));
  NAND3_X1   g12700(.A1(new_n11087_), .A2(new_n8847_), .A3(new_n11091_), .ZN(new_n13723_));
  NAND2_X1   g12701(.A1(new_n11100_), .A2(new_n8740_), .ZN(new_n13724_));
  AOI21_X1   g12702(.A1(new_n11074_), .A2(new_n13724_), .B(new_n11101_), .ZN(new_n13725_));
  AOI21_X1   g12703(.A1(new_n13723_), .A2(new_n11123_), .B(new_n13725_), .ZN(new_n13726_));
  INV_X1     g12704(.I(new_n13726_), .ZN(new_n13727_));
  NAND3_X1   g12705(.A1(new_n13723_), .A2(new_n11123_), .A3(new_n13725_), .ZN(new_n13728_));
  OAI21_X1   g12706(.A1(new_n11116_), .A2(new_n11078_), .B(new_n11107_), .ZN(new_n13729_));
  AOI22_X1   g12707(.A1(new_n11156_), .A2(new_n13729_), .B1(new_n13727_), .B2(new_n13728_), .ZN(new_n13730_));
  NOR2_X1    g12708(.A1(new_n11059_), .A2(new_n11060_), .ZN(new_n13731_));
  NAND4_X1   g12709(.A1(new_n8864_), .A2(new_n11068_), .A3(new_n8851_), .A4(new_n11065_), .ZN(new_n13732_));
  INV_X1     g12710(.I(new_n11070_), .ZN(new_n13733_));
  NOR3_X1    g12711(.A1(new_n13731_), .A2(new_n13733_), .A3(new_n13732_), .ZN(new_n13734_));
  NAND2_X1   g12712(.A1(new_n11066_), .A2(new_n8794_), .ZN(new_n13735_));
  NAND2_X1   g12713(.A1(new_n8766_), .A2(new_n8767_), .ZN(new_n13736_));
  NAND3_X1   g12714(.A1(new_n8754_), .A2(new_n8765_), .A3(new_n13736_), .ZN(new_n13737_));
  NAND2_X1   g12715(.A1(new_n13737_), .A2(new_n11035_), .ZN(new_n13738_));
  XOR2_X1    g12716(.A1(new_n13735_), .A2(new_n13738_), .Z(new_n13739_));
  AOI21_X1   g12717(.A1(new_n11058_), .A2(new_n13731_), .B(new_n11041_), .ZN(new_n13740_));
  OAI21_X1   g12718(.A1(new_n13740_), .A2(new_n13734_), .B(new_n13739_), .ZN(new_n13741_));
  NAND2_X1   g12719(.A1(new_n13730_), .A2(new_n13741_), .ZN(new_n13742_));
  NOR3_X1    g12720(.A1(new_n11114_), .A2(new_n8829_), .A3(new_n11113_), .ZN(new_n13743_));
  INV_X1     g12721(.I(new_n13725_), .ZN(new_n13744_));
  NOR3_X1    g12722(.A1(new_n13743_), .A2(new_n11126_), .A3(new_n13744_), .ZN(new_n13745_));
  AOI21_X1   g12723(.A1(new_n11112_), .A2(new_n11095_), .B(new_n11119_), .ZN(new_n13746_));
  OAI22_X1   g12724(.A1(new_n11136_), .A2(new_n13746_), .B1(new_n13726_), .B2(new_n13745_), .ZN(new_n13747_));
  XNOR2_X1   g12725(.A1(new_n13735_), .A2(new_n13738_), .ZN(new_n13748_));
  OAI22_X1   g12726(.A1(new_n11063_), .A2(new_n11049_), .B1(new_n11037_), .B2(new_n11040_), .ZN(new_n13749_));
  AOI21_X1   g12727(.A1(new_n11071_), .A2(new_n13749_), .B(new_n13748_), .ZN(new_n13750_));
  NAND2_X1   g12728(.A1(new_n13747_), .A2(new_n13750_), .ZN(new_n13751_));
  AOI22_X1   g12729(.A1(new_n13722_), .A2(new_n11157_), .B1(new_n13742_), .B2(new_n13751_), .ZN(new_n13752_));
  NAND2_X1   g12730(.A1(new_n11112_), .A2(new_n11095_), .ZN(new_n13753_));
  AOI21_X1   g12731(.A1(new_n11154_), .A2(new_n11155_), .B(new_n13753_), .ZN(new_n13754_));
  AOI21_X1   g12732(.A1(new_n13754_), .A2(new_n11150_), .B(new_n11140_), .ZN(new_n13755_));
  NAND2_X1   g12733(.A1(new_n11146_), .A2(new_n11073_), .ZN(new_n13756_));
  OAI21_X1   g12734(.A1(new_n13755_), .A2(new_n13756_), .B(new_n11157_), .ZN(new_n13757_));
  NOR2_X1    g12735(.A1(new_n13730_), .A2(new_n13750_), .ZN(new_n13758_));
  NOR2_X1    g12736(.A1(new_n13747_), .A2(new_n13741_), .ZN(new_n13759_));
  NOR2_X1    g12737(.A1(new_n13758_), .A2(new_n13759_), .ZN(new_n13760_));
  NOR2_X1    g12738(.A1(new_n13760_), .A2(new_n13757_), .ZN(new_n13761_));
  NOR2_X1    g12739(.A1(new_n13761_), .A2(new_n13752_), .ZN(new_n13762_));
  OAI21_X1   g12740(.A1(new_n8674_), .A2(new_n10984_), .B(new_n11027_), .ZN(new_n13763_));
  INV_X1     g12741(.I(new_n10957_), .ZN(new_n13764_));
  NOR4_X1    g12742(.A1(new_n10953_), .A2(new_n10965_), .A3(new_n10954_), .A4(new_n10979_), .ZN(new_n13765_));
  NAND2_X1   g12743(.A1(new_n13765_), .A2(new_n10942_), .ZN(new_n13766_));
  NOR4_X1    g12744(.A1(new_n13766_), .A2(new_n10942_), .A3(new_n13764_), .A4(new_n10971_), .ZN(new_n13767_));
  AOI21_X1   g12745(.A1(new_n13767_), .A2(new_n13763_), .B(new_n11028_), .ZN(new_n13768_));
  NOR3_X1    g12746(.A1(new_n11022_), .A2(new_n10993_), .A3(new_n11025_), .ZN(new_n13769_));
  AOI21_X1   g12747(.A1(new_n11015_), .A2(new_n11010_), .B(new_n8588_), .ZN(new_n13770_));
  INV_X1     g12748(.I(new_n11016_), .ZN(new_n13771_));
  NOR2_X1    g12749(.A1(new_n13771_), .A2(new_n13770_), .ZN(new_n13772_));
  OAI21_X1   g12750(.A1(new_n10991_), .A2(new_n10990_), .B(new_n10989_), .ZN(new_n13773_));
  NAND3_X1   g12751(.A1(new_n10985_), .A2(new_n10987_), .A3(new_n8667_), .ZN(new_n13774_));
  NAND2_X1   g12752(.A1(new_n13773_), .A2(new_n13774_), .ZN(new_n13775_));
  AOI21_X1   g12753(.A1(new_n11005_), .A2(new_n11008_), .B(new_n13775_), .ZN(new_n13776_));
  NAND3_X1   g12754(.A1(new_n8667_), .A2(new_n8657_), .A3(new_n11023_), .ZN(new_n13777_));
  NAND2_X1   g12755(.A1(new_n13777_), .A2(new_n10986_), .ZN(new_n13778_));
  NAND2_X1   g12756(.A1(new_n8589_), .A2(new_n8590_), .ZN(new_n13779_));
  NAND3_X1   g12757(.A1(new_n11003_), .A2(new_n8588_), .A3(new_n13779_), .ZN(new_n13780_));
  NAND2_X1   g12758(.A1(new_n13780_), .A2(new_n11014_), .ZN(new_n13781_));
  NAND2_X1   g12759(.A1(new_n13778_), .A2(new_n13781_), .ZN(new_n13782_));
  INV_X1     g12760(.I(new_n13782_), .ZN(new_n13783_));
  OAI21_X1   g12761(.A1(new_n13776_), .A2(new_n13772_), .B(new_n13783_), .ZN(new_n13784_));
  INV_X1     g12762(.I(new_n11008_), .ZN(new_n13785_));
  OAI21_X1   g12763(.A1(new_n11022_), .A2(new_n13785_), .B(new_n10993_), .ZN(new_n13786_));
  NAND3_X1   g12764(.A1(new_n13786_), .A2(new_n11017_), .A3(new_n13782_), .ZN(new_n13787_));
  AOI21_X1   g12765(.A1(new_n13784_), .A2(new_n13787_), .B(new_n13769_), .ZN(new_n13788_));
  INV_X1     g12766(.I(new_n13769_), .ZN(new_n13789_));
  AOI21_X1   g12767(.A1(new_n13786_), .A2(new_n11017_), .B(new_n13782_), .ZN(new_n13790_));
  NOR3_X1    g12768(.A1(new_n13776_), .A2(new_n13772_), .A3(new_n13783_), .ZN(new_n13791_));
  NOR3_X1    g12769(.A1(new_n13791_), .A2(new_n13790_), .A3(new_n13789_), .ZN(new_n13792_));
  NOR2_X1    g12770(.A1(new_n13792_), .A2(new_n13788_), .ZN(new_n13793_));
  OAI21_X1   g12771(.A1(new_n10953_), .A2(new_n10956_), .B(new_n10965_), .ZN(new_n13794_));
  NAND2_X1   g12772(.A1(new_n10979_), .A2(new_n10959_), .ZN(new_n13795_));
  NAND2_X1   g12773(.A1(new_n8615_), .A2(new_n8616_), .ZN(new_n13796_));
  NAND3_X1   g12774(.A1(new_n8603_), .A2(new_n8614_), .A3(new_n13796_), .ZN(new_n13797_));
  NAND2_X1   g12775(.A1(new_n13797_), .A2(new_n10935_), .ZN(new_n13798_));
  NAND2_X1   g12776(.A1(new_n13795_), .A2(new_n13798_), .ZN(new_n13799_));
  AOI21_X1   g12777(.A1(new_n13794_), .A2(new_n10942_), .B(new_n13799_), .ZN(new_n13800_));
  INV_X1     g12778(.I(new_n10956_), .ZN(new_n13801_));
  AOI21_X1   g12779(.A1(new_n13801_), .A2(new_n10977_), .B(new_n10971_), .ZN(new_n13802_));
  INV_X1     g12780(.I(new_n13799_), .ZN(new_n13803_));
  NOR3_X1    g12781(.A1(new_n13802_), .A2(new_n13803_), .A3(new_n10972_), .ZN(new_n13804_));
  OAI21_X1   g12782(.A1(new_n13800_), .A2(new_n13804_), .B(new_n10981_), .ZN(new_n13805_));
  OAI21_X1   g12783(.A1(new_n13802_), .A2(new_n10972_), .B(new_n13803_), .ZN(new_n13806_));
  NAND3_X1   g12784(.A1(new_n13794_), .A2(new_n10942_), .A3(new_n13799_), .ZN(new_n13807_));
  NAND3_X1   g12785(.A1(new_n13806_), .A2(new_n13807_), .A3(new_n13765_), .ZN(new_n13808_));
  NAND2_X1   g12786(.A1(new_n13805_), .A2(new_n13808_), .ZN(new_n13809_));
  NAND2_X1   g12787(.A1(new_n13793_), .A2(new_n13809_), .ZN(new_n13810_));
  OAI21_X1   g12788(.A1(new_n13791_), .A2(new_n13790_), .B(new_n13789_), .ZN(new_n13811_));
  NAND3_X1   g12789(.A1(new_n13784_), .A2(new_n13787_), .A3(new_n13769_), .ZN(new_n13812_));
  NAND2_X1   g12790(.A1(new_n13811_), .A2(new_n13812_), .ZN(new_n13813_));
  AOI21_X1   g12791(.A1(new_n13806_), .A2(new_n13807_), .B(new_n13765_), .ZN(new_n13814_));
  NOR3_X1    g12792(.A1(new_n13800_), .A2(new_n13804_), .A3(new_n10981_), .ZN(new_n13815_));
  NOR2_X1    g12793(.A1(new_n13815_), .A2(new_n13814_), .ZN(new_n13816_));
  NAND2_X1   g12794(.A1(new_n13816_), .A2(new_n13813_), .ZN(new_n13817_));
  AOI21_X1   g12795(.A1(new_n13817_), .A2(new_n13810_), .B(new_n13768_), .ZN(new_n13818_));
  XOR2_X1    g12796(.A1(new_n8592_), .A2(new_n8702_), .Z(new_n13819_));
  NOR2_X1    g12797(.A1(new_n11022_), .A2(new_n13785_), .ZN(new_n13820_));
  NOR3_X1    g12798(.A1(new_n13772_), .A2(new_n13820_), .A3(new_n13775_), .ZN(new_n13821_));
  NAND3_X1   g12799(.A1(new_n13821_), .A2(new_n13819_), .A3(new_n8703_), .ZN(new_n13822_));
  AOI21_X1   g12800(.A1(new_n8703_), .A2(new_n13819_), .B(new_n13821_), .ZN(new_n13823_));
  NAND4_X1   g12801(.A1(new_n10982_), .A2(new_n10972_), .A3(new_n10957_), .A4(new_n10965_), .ZN(new_n13824_));
  OAI21_X1   g12802(.A1(new_n13823_), .A2(new_n13824_), .B(new_n13822_), .ZN(new_n13825_));
  NAND2_X1   g12803(.A1(new_n13813_), .A2(new_n13809_), .ZN(new_n13826_));
  NAND4_X1   g12804(.A1(new_n13811_), .A2(new_n13812_), .A3(new_n13805_), .A4(new_n13808_), .ZN(new_n13827_));
  AOI21_X1   g12805(.A1(new_n13826_), .A2(new_n13827_), .B(new_n13825_), .ZN(new_n13828_));
  OAI21_X1   g12806(.A1(new_n13818_), .A2(new_n13828_), .B(new_n13762_), .ZN(new_n13829_));
  NOR3_X1    g12807(.A1(new_n11129_), .A2(new_n11121_), .A3(new_n11132_), .ZN(new_n13830_));
  NAND3_X1   g12808(.A1(new_n11150_), .A2(new_n11156_), .A3(new_n11128_), .ZN(new_n13831_));
  AOI21_X1   g12809(.A1(new_n13831_), .A2(new_n11132_), .B(new_n13756_), .ZN(new_n13832_));
  NOR2_X1    g12810(.A1(new_n13747_), .A2(new_n13750_), .ZN(new_n13833_));
  NOR2_X1    g12811(.A1(new_n13730_), .A2(new_n13741_), .ZN(new_n13834_));
  OAI22_X1   g12812(.A1(new_n13832_), .A2(new_n13830_), .B1(new_n13834_), .B2(new_n13833_), .ZN(new_n13835_));
  AOI21_X1   g12813(.A1(new_n13720_), .A2(new_n13721_), .B(new_n13830_), .ZN(new_n13836_));
  NAND2_X1   g12814(.A1(new_n13747_), .A2(new_n13741_), .ZN(new_n13837_));
  NAND2_X1   g12815(.A1(new_n13730_), .A2(new_n13750_), .ZN(new_n13838_));
  NAND2_X1   g12816(.A1(new_n13838_), .A2(new_n13837_), .ZN(new_n13839_));
  NAND2_X1   g12817(.A1(new_n13839_), .A2(new_n13836_), .ZN(new_n13840_));
  NAND2_X1   g12818(.A1(new_n13840_), .A2(new_n13835_), .ZN(new_n13841_));
  NOR2_X1    g12819(.A1(new_n13816_), .A2(new_n13813_), .ZN(new_n13842_));
  NOR2_X1    g12820(.A1(new_n13793_), .A2(new_n13809_), .ZN(new_n13843_));
  OAI21_X1   g12821(.A1(new_n13842_), .A2(new_n13843_), .B(new_n13825_), .ZN(new_n13844_));
  AOI22_X1   g12822(.A1(new_n13811_), .A2(new_n13812_), .B1(new_n13805_), .B2(new_n13808_), .ZN(new_n13845_));
  NOR4_X1    g12823(.A1(new_n13788_), .A2(new_n13792_), .A3(new_n13815_), .A4(new_n13814_), .ZN(new_n13846_));
  OAI21_X1   g12824(.A1(new_n13846_), .A2(new_n13845_), .B(new_n13768_), .ZN(new_n13847_));
  NAND3_X1   g12825(.A1(new_n13841_), .A2(new_n13844_), .A3(new_n13847_), .ZN(new_n13848_));
  AOI21_X1   g12826(.A1(new_n13829_), .A2(new_n13848_), .B(new_n13719_), .ZN(new_n13849_));
  AOI21_X1   g12827(.A1(new_n11158_), .A2(new_n11147_), .B(new_n11146_), .ZN(new_n13850_));
  NOR3_X1    g12828(.A1(new_n11141_), .A2(new_n11062_), .A3(new_n11133_), .ZN(new_n13851_));
  OAI21_X1   g12829(.A1(new_n13850_), .A2(new_n13851_), .B(new_n8881_), .ZN(new_n13852_));
  NOR3_X1    g12830(.A1(new_n13850_), .A2(new_n13851_), .A3(new_n8881_), .ZN(new_n13853_));
  OAI21_X1   g12831(.A1(new_n11032_), .A2(new_n13853_), .B(new_n13852_), .ZN(new_n13854_));
  OAI21_X1   g12832(.A1(new_n13818_), .A2(new_n13828_), .B(new_n13841_), .ZN(new_n13855_));
  NAND3_X1   g12833(.A1(new_n13762_), .A2(new_n13844_), .A3(new_n13847_), .ZN(new_n13856_));
  AOI21_X1   g12834(.A1(new_n13855_), .A2(new_n13856_), .B(new_n13854_), .ZN(new_n13857_));
  NOR2_X1    g12835(.A1(new_n13849_), .A2(new_n13857_), .ZN(new_n13858_));
  NOR2_X1    g12836(.A1(new_n13858_), .A2(new_n13717_), .ZN(new_n13859_));
  OAI21_X1   g12837(.A1(new_n13707_), .A2(new_n13710_), .B(new_n13704_), .ZN(new_n13860_));
  NAND3_X1   g12838(.A1(new_n13690_), .A2(new_n13627_), .A3(new_n13697_), .ZN(new_n13861_));
  AOI21_X1   g12839(.A1(new_n13860_), .A2(new_n13861_), .B(new_n13713_), .ZN(new_n13862_));
  OAI21_X1   g12840(.A1(new_n13707_), .A2(new_n13710_), .B(new_n13627_), .ZN(new_n13863_));
  NAND3_X1   g12841(.A1(new_n13690_), .A2(new_n13704_), .A3(new_n13697_), .ZN(new_n13864_));
  AOI21_X1   g12842(.A1(new_n13863_), .A2(new_n13864_), .B(new_n13544_), .ZN(new_n13865_));
  NOR2_X1    g12843(.A1(new_n13862_), .A2(new_n13865_), .ZN(new_n13866_));
  NOR3_X1    g12844(.A1(new_n13866_), .A2(new_n13849_), .A3(new_n13857_), .ZN(new_n13867_));
  OAI21_X1   g12845(.A1(new_n13859_), .A2(new_n13867_), .B(new_n13539_), .ZN(new_n13868_));
  AOI21_X1   g12846(.A1(new_n11312_), .A2(new_n11316_), .B(new_n8885_), .ZN(new_n13869_));
  AOI21_X1   g12847(.A1(new_n11161_), .A2(new_n13537_), .B(new_n13869_), .ZN(new_n13870_));
  AOI21_X1   g12848(.A1(new_n13844_), .A2(new_n13847_), .B(new_n13841_), .ZN(new_n13871_));
  NOR3_X1    g12849(.A1(new_n13762_), .A2(new_n13818_), .A3(new_n13828_), .ZN(new_n13872_));
  OAI21_X1   g12850(.A1(new_n13871_), .A2(new_n13872_), .B(new_n13854_), .ZN(new_n13873_));
  AOI22_X1   g12851(.A1(new_n13844_), .A2(new_n13847_), .B1(new_n13835_), .B2(new_n13840_), .ZN(new_n13874_));
  NOR3_X1    g12852(.A1(new_n13841_), .A2(new_n13818_), .A3(new_n13828_), .ZN(new_n13875_));
  OAI21_X1   g12853(.A1(new_n13874_), .A2(new_n13875_), .B(new_n13719_), .ZN(new_n13876_));
  AOI22_X1   g12854(.A1(new_n13873_), .A2(new_n13876_), .B1(new_n13712_), .B2(new_n13716_), .ZN(new_n13877_));
  NOR4_X1    g12855(.A1(new_n13849_), .A2(new_n13857_), .A3(new_n13862_), .A4(new_n13865_), .ZN(new_n13878_));
  OAI21_X1   g12856(.A1(new_n13877_), .A2(new_n13878_), .B(new_n13870_), .ZN(new_n13879_));
  NAND2_X1   g12857(.A1(new_n13868_), .A2(new_n13879_), .ZN(new_n13880_));
  NAND2_X1   g12858(.A1(new_n13880_), .A2(new_n13536_), .ZN(new_n13881_));
  AOI21_X1   g12859(.A1(new_n13523_), .A2(new_n13526_), .B(new_n13520_), .ZN(new_n13882_));
  NOR3_X1    g12860(.A1(new_n13372_), .A2(new_n13504_), .A3(new_n13512_), .ZN(new_n13883_));
  OAI21_X1   g12861(.A1(new_n13882_), .A2(new_n13883_), .B(new_n13532_), .ZN(new_n13884_));
  AOI22_X1   g12862(.A1(new_n13523_), .A2(new_n13526_), .B1(new_n13516_), .B2(new_n13519_), .ZN(new_n13885_));
  NOR3_X1    g12863(.A1(new_n13520_), .A2(new_n13504_), .A3(new_n13512_), .ZN(new_n13886_));
  OAI21_X1   g12864(.A1(new_n13885_), .A2(new_n13886_), .B(new_n13215_), .ZN(new_n13887_));
  NAND2_X1   g12865(.A1(new_n13884_), .A2(new_n13887_), .ZN(new_n13888_));
  NAND3_X1   g12866(.A1(new_n13888_), .A2(new_n13868_), .A3(new_n13879_), .ZN(new_n13889_));
  AOI21_X1   g12867(.A1(new_n13881_), .A2(new_n13889_), .B(new_n13213_), .ZN(new_n13890_));
  INV_X1     g12868(.I(new_n13213_), .ZN(new_n13891_));
  OAI21_X1   g12869(.A1(new_n13849_), .A2(new_n13857_), .B(new_n13866_), .ZN(new_n13892_));
  NAND2_X1   g12870(.A1(new_n13858_), .A2(new_n13717_), .ZN(new_n13893_));
  AOI21_X1   g12871(.A1(new_n13892_), .A2(new_n13893_), .B(new_n13870_), .ZN(new_n13894_));
  OAI22_X1   g12872(.A1(new_n13849_), .A2(new_n13857_), .B1(new_n13862_), .B2(new_n13865_), .ZN(new_n13895_));
  NAND4_X1   g12873(.A1(new_n13873_), .A2(new_n13876_), .A3(new_n13712_), .A4(new_n13716_), .ZN(new_n13896_));
  AOI21_X1   g12874(.A1(new_n13895_), .A2(new_n13896_), .B(new_n13539_), .ZN(new_n13897_));
  OAI22_X1   g12875(.A1(new_n13894_), .A2(new_n13897_), .B1(new_n13528_), .B2(new_n13535_), .ZN(new_n13898_));
  NAND4_X1   g12876(.A1(new_n13868_), .A2(new_n13884_), .A3(new_n13887_), .A4(new_n13879_), .ZN(new_n13899_));
  AOI21_X1   g12877(.A1(new_n13898_), .A2(new_n13899_), .B(new_n13891_), .ZN(new_n13900_));
  NOR2_X1    g12878(.A1(new_n13890_), .A2(new_n13900_), .ZN(new_n13901_));
  NOR2_X1    g12879(.A1(new_n13901_), .A2(new_n13210_), .ZN(new_n13902_));
  OAI21_X1   g12880(.A1(new_n13200_), .A2(new_n13203_), .B(new_n13197_), .ZN(new_n13903_));
  NAND3_X1   g12881(.A1(new_n12882_), .A2(new_n13184_), .A3(new_n13189_), .ZN(new_n13904_));
  AOI21_X1   g12882(.A1(new_n13903_), .A2(new_n13904_), .B(new_n12559_), .ZN(new_n13905_));
  OAI22_X1   g12883(.A1(new_n13200_), .A2(new_n13203_), .B1(new_n13207_), .B2(new_n13196_), .ZN(new_n13906_));
  NAND4_X1   g12884(.A1(new_n13184_), .A2(new_n12877_), .A3(new_n12881_), .A4(new_n13189_), .ZN(new_n13907_));
  AOI21_X1   g12885(.A1(new_n13906_), .A2(new_n13907_), .B(new_n12560_), .ZN(new_n13908_));
  NOR2_X1    g12886(.A1(new_n13905_), .A2(new_n13908_), .ZN(new_n13909_));
  NOR3_X1    g12887(.A1(new_n13909_), .A2(new_n13890_), .A3(new_n13900_), .ZN(new_n13910_));
  OAI21_X1   g12888(.A1(new_n13902_), .A2(new_n13910_), .B(new_n12558_), .ZN(new_n13911_));
  INV_X1     g12889(.I(new_n12558_), .ZN(new_n13912_));
  NOR4_X1    g12890(.A1(new_n13890_), .A2(new_n13905_), .A3(new_n13908_), .A4(new_n13900_), .ZN(new_n13913_));
  AOI21_X1   g12891(.A1(new_n13868_), .A2(new_n13879_), .B(new_n13888_), .ZN(new_n13914_));
  NOR2_X1    g12892(.A1(new_n13880_), .A2(new_n13536_), .ZN(new_n13915_));
  OAI21_X1   g12893(.A1(new_n13914_), .A2(new_n13915_), .B(new_n13891_), .ZN(new_n13916_));
  AOI22_X1   g12894(.A1(new_n13868_), .A2(new_n13879_), .B1(new_n13884_), .B2(new_n13887_), .ZN(new_n13917_));
  NOR4_X1    g12895(.A1(new_n13894_), .A2(new_n13528_), .A3(new_n13535_), .A4(new_n13897_), .ZN(new_n13918_));
  OAI21_X1   g12896(.A1(new_n13918_), .A2(new_n13917_), .B(new_n13213_), .ZN(new_n13919_));
  AOI22_X1   g12897(.A1(new_n13916_), .A2(new_n13919_), .B1(new_n13205_), .B2(new_n13209_), .ZN(new_n13920_));
  OAI21_X1   g12898(.A1(new_n13920_), .A2(new_n13913_), .B(new_n13912_), .ZN(new_n13921_));
  NAND2_X1   g12899(.A1(new_n13911_), .A2(new_n13921_), .ZN(new_n13922_));
  NAND2_X1   g12900(.A1(new_n13922_), .A2(new_n12556_), .ZN(new_n13923_));
  NOR2_X1    g12901(.A1(new_n13922_), .A2(new_n12556_), .ZN(new_n13924_));
  INV_X1     g12902(.I(new_n13924_), .ZN(new_n13925_));
  AOI21_X1   g12903(.A1(new_n13925_), .A2(new_n13923_), .B(new_n8198_), .ZN(new_n13926_));
  AOI21_X1   g12904(.A1(new_n8196_), .A2(new_n8195_), .B(new_n8194_), .ZN(new_n13927_));
  NOR3_X1    g12905(.A1(new_n8182_), .A2(new_n8186_), .A3(new_n6273_), .ZN(new_n13928_));
  NOR2_X1    g12906(.A1(new_n13928_), .A2(new_n13927_), .ZN(new_n13929_));
  INV_X1     g12907(.I(new_n13923_), .ZN(new_n13930_));
  NOR3_X1    g12908(.A1(new_n13930_), .A2(new_n13924_), .A3(new_n13929_), .ZN(new_n13931_));
  OAI21_X1   g12909(.A1(new_n13926_), .A2(new_n13931_), .B(new_n5352_), .ZN(new_n13932_));
  OR3_X2     g12910(.A1(new_n13926_), .A2(new_n13931_), .A3(new_n5352_), .Z(new_n13933_));
  NAND2_X1   g12911(.A1(new_n10927_), .A2(new_n10928_), .ZN(new_n13934_));
  AOI21_X1   g12912(.A1(new_n2688_), .A2(new_n2684_), .B(new_n3597_), .ZN(new_n13935_));
  NOR2_X1    g12913(.A1(new_n3599_), .A2(new_n13935_), .ZN(new_n13936_));
  XOR2_X1    g12914(.A1(new_n13936_), .A2(new_n10931_), .Z(new_n13937_));
  XOR2_X1    g12915(.A1(new_n13937_), .A2(\A[1000] ), .Z(new_n13938_));
  NAND2_X1   g12916(.A1(new_n13938_), .A2(new_n13934_), .ZN(new_n13939_));
  INV_X1     g12917(.I(new_n13939_), .ZN(new_n13940_));
  NAND3_X1   g12918(.A1(new_n13933_), .A2(new_n13932_), .A3(new_n13940_), .ZN(new_n13941_));
  NAND2_X1   g12919(.A1(new_n13933_), .A2(new_n13932_), .ZN(new_n13942_));
  NAND2_X1   g12920(.A1(new_n13942_), .A2(new_n13939_), .ZN(new_n13943_));
  INV_X1     g12921(.I(new_n2686_), .ZN(new_n13944_));
  NAND3_X1   g12922(.A1(new_n4269_), .A2(new_n13944_), .A3(new_n3599_), .ZN(new_n13945_));
  NAND3_X1   g12923(.A1(new_n4269_), .A2(new_n2686_), .A3(new_n3599_), .ZN(new_n13946_));
  NAND2_X1   g12924(.A1(new_n13945_), .A2(new_n13946_), .ZN(new_n13947_));
  INV_X1     g12925(.I(new_n13936_), .ZN(new_n13948_));
  OR2_X2     g12926(.A1(new_n10931_), .A2(new_n13934_), .Z(new_n13949_));
  NAND2_X1   g12927(.A1(new_n10931_), .A2(new_n13934_), .ZN(new_n13950_));
  AOI21_X1   g12928(.A1(new_n13949_), .A2(new_n13950_), .B(new_n13948_), .ZN(new_n13951_));
  NAND2_X1   g12929(.A1(new_n13947_), .A2(new_n13951_), .ZN(new_n13952_));
  NOR2_X1    g12930(.A1(new_n10933_), .A2(new_n12553_), .ZN(new_n13953_));
  AOI21_X1   g12931(.A1(new_n13943_), .A2(new_n13941_), .B(new_n13952_), .ZN(new_n13955_));
  OAI21_X1   g12932(.A1(new_n13890_), .A2(new_n13900_), .B(new_n13909_), .ZN(new_n13956_));
  NAND3_X1   g12933(.A1(new_n13210_), .A2(new_n13916_), .A3(new_n13919_), .ZN(new_n13957_));
  AOI21_X1   g12934(.A1(new_n13956_), .A2(new_n13957_), .B(new_n13912_), .ZN(new_n13958_));
  NAND4_X1   g12935(.A1(new_n13916_), .A2(new_n13205_), .A3(new_n13209_), .A4(new_n13919_), .ZN(new_n13959_));
  OAI22_X1   g12936(.A1(new_n13890_), .A2(new_n13900_), .B1(new_n13905_), .B2(new_n13908_), .ZN(new_n13960_));
  AOI21_X1   g12937(.A1(new_n13959_), .A2(new_n13960_), .B(new_n12558_), .ZN(new_n13961_));
  OAI21_X1   g12938(.A1(new_n13958_), .A2(new_n13961_), .B(new_n13929_), .ZN(new_n13962_));
  NAND3_X1   g12939(.A1(new_n13911_), .A2(new_n8198_), .A3(new_n13921_), .ZN(new_n13963_));
  AOI21_X1   g12940(.A1(new_n13962_), .A2(new_n13963_), .B(new_n12556_), .ZN(new_n13964_));
  INV_X1     g12941(.I(new_n12556_), .ZN(new_n13965_));
  NAND3_X1   g12942(.A1(new_n13911_), .A2(new_n13929_), .A3(new_n13921_), .ZN(new_n13966_));
  OAI21_X1   g12943(.A1(new_n13958_), .A2(new_n13961_), .B(new_n8198_), .ZN(new_n13967_));
  AOI21_X1   g12944(.A1(new_n13967_), .A2(new_n13966_), .B(new_n13965_), .ZN(new_n13968_));
  NOR2_X1    g12945(.A1(new_n13964_), .A2(new_n13968_), .ZN(new_n13969_));
  NOR3_X1    g12946(.A1(new_n5344_), .A2(new_n4780_), .A3(new_n4789_), .ZN(new_n13970_));
  NOR2_X1    g12947(.A1(new_n4790_), .A2(new_n5336_), .ZN(new_n13971_));
  OAI21_X1   g12948(.A1(new_n13971_), .A2(new_n13970_), .B(new_n5347_), .ZN(new_n13972_));
  NOR2_X1    g12949(.A1(new_n4771_), .A2(new_n4778_), .ZN(new_n13973_));
  AOI21_X1   g12950(.A1(new_n4505_), .A2(new_n4508_), .B(new_n4769_), .ZN(new_n13974_));
  OAI21_X1   g12951(.A1(new_n13974_), .A2(new_n13973_), .B(new_n4272_), .ZN(new_n13975_));
  NOR2_X1    g12952(.A1(new_n4771_), .A2(new_n4769_), .ZN(new_n13976_));
  AOI21_X1   g12953(.A1(new_n4505_), .A2(new_n4508_), .B(new_n4778_), .ZN(new_n13977_));
  OAI21_X1   g12954(.A1(new_n13977_), .A2(new_n13976_), .B(new_n4273_), .ZN(new_n13978_));
  AOI22_X1   g12955(.A1(new_n13975_), .A2(new_n13978_), .B1(new_n5331_), .B2(new_n5335_), .ZN(new_n13979_));
  OAI21_X1   g12956(.A1(new_n13979_), .A2(new_n5348_), .B(new_n4270_), .ZN(new_n13980_));
  NAND2_X1   g12957(.A1(new_n13972_), .A2(new_n13980_), .ZN(new_n13981_));
  NAND2_X1   g12958(.A1(new_n13962_), .A2(new_n13963_), .ZN(new_n13982_));
  OAI21_X1   g12959(.A1(new_n13947_), .A2(new_n13951_), .B(new_n13953_), .ZN(new_n13983_));
  AOI21_X1   g12960(.A1(new_n13983_), .A2(new_n13952_), .B(new_n12556_), .ZN(new_n13984_));
  AOI21_X1   g12961(.A1(new_n13982_), .A2(new_n13984_), .B(new_n13981_), .ZN(new_n13985_));
  NOR2_X1    g12962(.A1(new_n13969_), .A2(new_n13985_), .ZN(new_n13986_));
  OAI21_X1   g12963(.A1(new_n5100_), .A2(new_n5103_), .B(new_n5099_), .ZN(new_n13987_));
  OAI21_X1   g12964(.A1(new_n13987_), .A2(new_n5106_), .B(new_n5104_), .ZN(new_n13988_));
  OAI21_X1   g12965(.A1(new_n5115_), .A2(new_n5118_), .B(new_n5130_), .ZN(new_n13989_));
  OAI21_X1   g12966(.A1(new_n13989_), .A2(new_n5127_), .B(new_n5119_), .ZN(new_n13990_));
  XOR2_X1    g12967(.A1(new_n13990_), .A2(new_n13988_), .Z(new_n13991_));
  NOR2_X1    g12968(.A1(new_n5145_), .A2(new_n5098_), .ZN(new_n13992_));
  INV_X1     g12969(.I(new_n5106_), .ZN(new_n13993_));
  INV_X1     g12970(.I(new_n5127_), .ZN(new_n13994_));
  XNOR2_X1   g12971(.A1(new_n5100_), .A2(new_n5103_), .ZN(new_n13995_));
  XNOR2_X1   g12972(.A1(new_n5118_), .A2(new_n5115_), .ZN(new_n13996_));
  NOR4_X1    g12973(.A1(new_n13995_), .A2(new_n13996_), .A3(new_n1576_), .A4(new_n1598_), .ZN(new_n13997_));
  NAND3_X1   g12974(.A1(new_n13997_), .A2(new_n13993_), .A3(new_n13994_), .ZN(new_n13998_));
  OAI22_X1   g12975(.A1(new_n5130_), .A2(new_n13994_), .B1(new_n13993_), .B2(new_n5099_), .ZN(new_n13999_));
  NOR2_X1    g12976(.A1(new_n13998_), .A2(new_n13999_), .ZN(new_n14000_));
  OAI21_X1   g12977(.A1(new_n13992_), .A2(new_n14000_), .B(new_n13991_), .ZN(new_n14001_));
  OAI21_X1   g12978(.A1(new_n5166_), .A2(new_n5164_), .B(new_n5296_), .ZN(new_n14002_));
  AOI21_X1   g12979(.A1(new_n1786_), .A2(new_n5070_), .B(new_n5069_), .ZN(new_n14003_));
  NAND3_X1   g12980(.A1(new_n5078_), .A2(new_n5076_), .A3(new_n5077_), .ZN(new_n14004_));
  NOR4_X1    g12981(.A1(new_n14004_), .A2(new_n1802_), .A3(new_n5073_), .A4(new_n5074_), .ZN(new_n14005_));
  NAND2_X1   g12982(.A1(new_n14005_), .A2(new_n14003_), .ZN(new_n14006_));
  NOR2_X1    g12983(.A1(new_n5055_), .A2(new_n5087_), .ZN(new_n14007_));
  NAND2_X1   g12984(.A1(new_n5068_), .A2(new_n5066_), .ZN(new_n14008_));
  NAND4_X1   g12985(.A1(new_n5067_), .A2(new_n1736_), .A3(new_n1664_), .A4(new_n5065_), .ZN(new_n14009_));
  NAND3_X1   g12986(.A1(new_n5078_), .A2(new_n5076_), .A3(new_n14009_), .ZN(new_n14010_));
  NAND2_X1   g12987(.A1(new_n14010_), .A2(new_n14008_), .ZN(new_n14011_));
  NAND2_X1   g12988(.A1(new_n5060_), .A2(new_n5058_), .ZN(new_n14012_));
  OR2_X2     g12989(.A1(new_n5060_), .A2(new_n5058_), .Z(new_n14013_));
  NAND3_X1   g12990(.A1(new_n5062_), .A2(new_n1781_), .A3(new_n14013_), .ZN(new_n14014_));
  NAND2_X1   g12991(.A1(new_n14014_), .A2(new_n14012_), .ZN(new_n14015_));
  NAND2_X1   g12992(.A1(new_n14011_), .A2(new_n14015_), .ZN(new_n14016_));
  NOR2_X1    g12993(.A1(new_n14007_), .A2(new_n14016_), .ZN(new_n14017_));
  NAND2_X1   g12994(.A1(new_n14007_), .A2(new_n14016_), .ZN(new_n14018_));
  INV_X1     g12995(.I(new_n14018_), .ZN(new_n14019_));
  OAI21_X1   g12996(.A1(new_n14019_), .A2(new_n14017_), .B(new_n14006_), .ZN(new_n14020_));
  INV_X1     g12997(.I(new_n14006_), .ZN(new_n14021_));
  INV_X1     g12998(.I(new_n14017_), .ZN(new_n14022_));
  NAND3_X1   g12999(.A1(new_n14022_), .A2(new_n14021_), .A3(new_n14018_), .ZN(new_n14023_));
  NAND2_X1   g13000(.A1(new_n14020_), .A2(new_n14023_), .ZN(new_n14024_));
  INV_X1     g13001(.I(new_n14024_), .ZN(new_n14025_));
  NOR2_X1    g13002(.A1(new_n14025_), .A2(new_n14002_), .ZN(new_n14026_));
  INV_X1     g13003(.I(new_n14002_), .ZN(new_n14027_));
  NOR2_X1    g13004(.A1(new_n14027_), .A2(new_n14024_), .ZN(new_n14028_));
  OAI21_X1   g13005(.A1(new_n14028_), .A2(new_n14026_), .B(new_n14001_), .ZN(new_n14029_));
  INV_X1     g13006(.I(new_n14001_), .ZN(new_n14030_));
  NAND2_X1   g13007(.A1(new_n14002_), .A2(new_n14024_), .ZN(new_n14031_));
  INV_X1     g13008(.I(new_n14031_), .ZN(new_n14032_));
  NOR2_X1    g13009(.A1(new_n14002_), .A2(new_n14024_), .ZN(new_n14033_));
  OAI21_X1   g13010(.A1(new_n14032_), .A2(new_n14033_), .B(new_n14030_), .ZN(new_n14034_));
  NAND2_X1   g13011(.A1(new_n14029_), .A2(new_n14034_), .ZN(new_n14035_));
  NAND2_X1   g13012(.A1(new_n5312_), .A2(new_n5310_), .ZN(new_n14036_));
  AOI21_X1   g13013(.A1(new_n5172_), .A2(new_n5302_), .B(new_n5289_), .ZN(new_n14037_));
  INV_X1     g13014(.I(new_n14037_), .ZN(new_n14038_));
  OAI21_X1   g13015(.A1(new_n5250_), .A2(new_n5241_), .B(new_n5248_), .ZN(new_n14039_));
  NOR3_X1    g13016(.A1(new_n5257_), .A2(new_n5249_), .A3(new_n5240_), .ZN(new_n14040_));
  NAND4_X1   g13017(.A1(new_n14040_), .A2(new_n5253_), .A3(new_n5254_), .A4(new_n5255_), .ZN(new_n14041_));
  NOR2_X1    g13018(.A1(new_n14041_), .A2(new_n14039_), .ZN(new_n14042_));
  NAND2_X1   g13019(.A1(new_n5264_), .A2(new_n5230_), .ZN(new_n14043_));
  INV_X1     g13020(.I(new_n5247_), .ZN(new_n14044_));
  NAND2_X1   g13021(.A1(new_n14044_), .A2(new_n5243_), .ZN(new_n14045_));
  NAND3_X1   g13022(.A1(new_n5247_), .A2(new_n5242_), .A3(new_n1054_), .ZN(new_n14046_));
  NAND3_X1   g13023(.A1(new_n5250_), .A2(new_n5241_), .A3(new_n14046_), .ZN(new_n14047_));
  NAND2_X1   g13024(.A1(new_n5236_), .A2(new_n5233_), .ZN(new_n14048_));
  OR2_X2     g13025(.A1(new_n5236_), .A2(new_n5233_), .Z(new_n14049_));
  NAND3_X1   g13026(.A1(new_n5255_), .A2(new_n5253_), .A3(new_n14049_), .ZN(new_n14050_));
  AOI22_X1   g13027(.A1(new_n14047_), .A2(new_n14045_), .B1(new_n14048_), .B2(new_n14050_), .ZN(new_n14051_));
  NAND2_X1   g13028(.A1(new_n14043_), .A2(new_n14051_), .ZN(new_n14052_));
  NOR2_X1    g13029(.A1(new_n5262_), .A2(new_n5279_), .ZN(new_n14053_));
  NAND2_X1   g13030(.A1(new_n14047_), .A2(new_n14045_), .ZN(new_n14054_));
  NAND2_X1   g13031(.A1(new_n14050_), .A2(new_n14048_), .ZN(new_n14055_));
  NAND2_X1   g13032(.A1(new_n14054_), .A2(new_n14055_), .ZN(new_n14056_));
  NAND2_X1   g13033(.A1(new_n14053_), .A2(new_n14056_), .ZN(new_n14057_));
  AOI21_X1   g13034(.A1(new_n14057_), .A2(new_n14052_), .B(new_n14042_), .ZN(new_n14058_));
  INV_X1     g13035(.I(new_n14042_), .ZN(new_n14059_));
  NOR2_X1    g13036(.A1(new_n14053_), .A2(new_n14056_), .ZN(new_n14060_));
  NOR2_X1    g13037(.A1(new_n14043_), .A2(new_n14051_), .ZN(new_n14061_));
  NOR3_X1    g13038(.A1(new_n14060_), .A2(new_n14059_), .A3(new_n14061_), .ZN(new_n14062_));
  OR2_X2     g13039(.A1(new_n14062_), .A2(new_n14058_), .Z(new_n14063_));
  OAI21_X1   g13040(.A1(new_n5188_), .A2(new_n5179_), .B(new_n5186_), .ZN(new_n14064_));
  NOR3_X1    g13041(.A1(new_n5200_), .A2(new_n5202_), .A3(new_n5199_), .ZN(new_n14065_));
  NAND4_X1   g13042(.A1(new_n14065_), .A2(new_n1320_), .A3(new_n5204_), .A4(new_n5205_), .ZN(new_n14066_));
  NOR2_X1    g13043(.A1(new_n14066_), .A2(new_n14064_), .ZN(new_n14067_));
  NAND2_X1   g13044(.A1(new_n5272_), .A2(new_n5214_), .ZN(new_n14068_));
  NAND2_X1   g13045(.A1(new_n5194_), .A2(new_n5191_), .ZN(new_n14069_));
  NOR2_X1    g13046(.A1(new_n5194_), .A2(new_n5191_), .ZN(new_n14070_));
  OR3_X2     g13047(.A1(new_n1321_), .A2(new_n5196_), .A3(new_n14070_), .Z(new_n14071_));
  NAND2_X1   g13048(.A1(new_n14071_), .A2(new_n14069_), .ZN(new_n14072_));
  NAND2_X1   g13049(.A1(new_n5185_), .A2(new_n5182_), .ZN(new_n14073_));
  NOR2_X1    g13050(.A1(new_n5185_), .A2(new_n5182_), .ZN(new_n14074_));
  OR3_X2     g13051(.A1(new_n5202_), .A2(new_n5199_), .A3(new_n14074_), .Z(new_n14075_));
  NAND2_X1   g13052(.A1(new_n14075_), .A2(new_n14073_), .ZN(new_n14076_));
  NAND3_X1   g13053(.A1(new_n14068_), .A2(new_n14072_), .A3(new_n14076_), .ZN(new_n14077_));
  NOR2_X1    g13054(.A1(new_n5216_), .A2(new_n5176_), .ZN(new_n14078_));
  INV_X1     g13055(.I(new_n14072_), .ZN(new_n14079_));
  INV_X1     g13056(.I(new_n14076_), .ZN(new_n14080_));
  OAI21_X1   g13057(.A1(new_n14080_), .A2(new_n14079_), .B(new_n14078_), .ZN(new_n14081_));
  AOI21_X1   g13058(.A1(new_n14081_), .A2(new_n14077_), .B(new_n14067_), .ZN(new_n14082_));
  INV_X1     g13059(.I(new_n14067_), .ZN(new_n14083_));
  NOR3_X1    g13060(.A1(new_n14080_), .A2(new_n14078_), .A3(new_n14079_), .ZN(new_n14084_));
  AOI21_X1   g13061(.A1(new_n14072_), .A2(new_n14076_), .B(new_n14068_), .ZN(new_n14085_));
  NOR3_X1    g13062(.A1(new_n14084_), .A2(new_n14085_), .A3(new_n14083_), .ZN(new_n14086_));
  NOR2_X1    g13063(.A1(new_n14086_), .A2(new_n14082_), .ZN(new_n14087_));
  NOR2_X1    g13064(.A1(new_n14063_), .A2(new_n14087_), .ZN(new_n14088_));
  NOR2_X1    g13065(.A1(new_n14062_), .A2(new_n14058_), .ZN(new_n14089_));
  OAI21_X1   g13066(.A1(new_n14084_), .A2(new_n14085_), .B(new_n14083_), .ZN(new_n14090_));
  NAND3_X1   g13067(.A1(new_n14081_), .A2(new_n14067_), .A3(new_n14077_), .ZN(new_n14091_));
  NAND2_X1   g13068(.A1(new_n14090_), .A2(new_n14091_), .ZN(new_n14092_));
  NOR2_X1    g13069(.A1(new_n14092_), .A2(new_n14089_), .ZN(new_n14093_));
  OAI21_X1   g13070(.A1(new_n14088_), .A2(new_n14093_), .B(new_n14038_), .ZN(new_n14094_));
  NOR2_X1    g13071(.A1(new_n14087_), .A2(new_n14089_), .ZN(new_n14095_));
  NOR2_X1    g13072(.A1(new_n14063_), .A2(new_n14092_), .ZN(new_n14096_));
  OAI21_X1   g13073(.A1(new_n14096_), .A2(new_n14095_), .B(new_n14037_), .ZN(new_n14097_));
  NAND2_X1   g13074(.A1(new_n14094_), .A2(new_n14097_), .ZN(new_n14098_));
  NAND3_X1   g13075(.A1(new_n14098_), .A2(new_n14036_), .A3(new_n5311_), .ZN(new_n14099_));
  INV_X1     g13076(.I(new_n14099_), .ZN(new_n14100_));
  AOI21_X1   g13077(.A1(new_n5311_), .A2(new_n14036_), .B(new_n14098_), .ZN(new_n14101_));
  OAI21_X1   g13078(.A1(new_n14100_), .A2(new_n14101_), .B(new_n14035_), .ZN(new_n14102_));
  NAND2_X1   g13079(.A1(new_n14027_), .A2(new_n14024_), .ZN(new_n14103_));
  NAND2_X1   g13080(.A1(new_n14025_), .A2(new_n14002_), .ZN(new_n14104_));
  AOI21_X1   g13081(.A1(new_n14103_), .A2(new_n14104_), .B(new_n14030_), .ZN(new_n14105_));
  NAND2_X1   g13082(.A1(new_n14027_), .A2(new_n14025_), .ZN(new_n14106_));
  AOI21_X1   g13083(.A1(new_n14106_), .A2(new_n14031_), .B(new_n14001_), .ZN(new_n14107_));
  NOR2_X1    g13084(.A1(new_n14107_), .A2(new_n14105_), .ZN(new_n14108_));
  AOI22_X1   g13085(.A1(new_n14036_), .A2(new_n5311_), .B1(new_n14094_), .B2(new_n14097_), .ZN(new_n14109_));
  NAND2_X1   g13086(.A1(new_n14036_), .A2(new_n5311_), .ZN(new_n14110_));
  NOR2_X1    g13087(.A1(new_n14110_), .A2(new_n14098_), .ZN(new_n14111_));
  OAI21_X1   g13088(.A1(new_n14111_), .A2(new_n14109_), .B(new_n14108_), .ZN(new_n14112_));
  NAND2_X1   g13089(.A1(new_n14102_), .A2(new_n14112_), .ZN(new_n14113_));
  NAND2_X1   g13090(.A1(new_n5342_), .A2(new_n4793_), .ZN(new_n14114_));
  NAND2_X1   g13091(.A1(new_n14114_), .A2(new_n5341_), .ZN(new_n14115_));
  AOI21_X1   g13092(.A1(new_n4797_), .A2(new_n5319_), .B(new_n5042_), .ZN(new_n14116_));
  OAI21_X1   g13093(.A1(new_n5034_), .A2(new_n4912_), .B(new_n5021_), .ZN(new_n14117_));
  INV_X1     g13094(.I(new_n14117_), .ZN(new_n14118_));
  AOI21_X1   g13095(.A1(new_n4971_), .A2(new_n4980_), .B(new_n4978_), .ZN(new_n14119_));
  NAND3_X1   g13096(.A1(new_n4989_), .A2(new_n4987_), .A3(new_n4986_), .ZN(new_n14120_));
  NOR4_X1    g13097(.A1(new_n14120_), .A2(new_n4961_), .A3(new_n4983_), .A4(new_n4984_), .ZN(new_n14121_));
  NAND2_X1   g13098(.A1(new_n14121_), .A2(new_n14119_), .ZN(new_n14122_));
  INV_X1     g13099(.I(new_n14122_), .ZN(new_n14123_));
  NAND2_X1   g13100(.A1(new_n5010_), .A2(new_n4994_), .ZN(new_n14124_));
  INV_X1     g13101(.I(new_n4977_), .ZN(new_n14125_));
  NAND2_X1   g13102(.A1(new_n14125_), .A2(new_n4973_), .ZN(new_n14126_));
  NAND3_X1   g13103(.A1(new_n4977_), .A2(new_n1876_), .A3(new_n4972_), .ZN(new_n14127_));
  NAND3_X1   g13104(.A1(new_n4989_), .A2(new_n4986_), .A3(new_n14127_), .ZN(new_n14128_));
  OAI21_X1   g13105(.A1(new_n1961_), .A2(new_n4963_), .B(new_n4967_), .ZN(new_n14129_));
  NAND3_X1   g13106(.A1(new_n4964_), .A2(new_n1935_), .A3(new_n4966_), .ZN(new_n14130_));
  NAND3_X1   g13107(.A1(new_n4969_), .A2(new_n4962_), .A3(new_n14130_), .ZN(new_n14131_));
  AOI22_X1   g13108(.A1(new_n14128_), .A2(new_n14126_), .B1(new_n14131_), .B2(new_n14129_), .ZN(new_n14132_));
  NAND2_X1   g13109(.A1(new_n14124_), .A2(new_n14132_), .ZN(new_n14133_));
  NOR2_X1    g13110(.A1(new_n4996_), .A2(new_n4960_), .ZN(new_n14134_));
  INV_X1     g13111(.I(new_n14132_), .ZN(new_n14135_));
  NAND2_X1   g13112(.A1(new_n14135_), .A2(new_n14134_), .ZN(new_n14136_));
  AOI21_X1   g13113(.A1(new_n14136_), .A2(new_n14133_), .B(new_n14123_), .ZN(new_n14137_));
  NOR2_X1    g13114(.A1(new_n14135_), .A2(new_n14134_), .ZN(new_n14138_));
  NOR2_X1    g13115(.A1(new_n14124_), .A2(new_n14132_), .ZN(new_n14139_));
  NOR3_X1    g13116(.A1(new_n14138_), .A2(new_n14139_), .A3(new_n14122_), .ZN(new_n14140_));
  NOR2_X1    g13117(.A1(new_n14140_), .A2(new_n14137_), .ZN(new_n14141_));
  OAI21_X1   g13118(.A1(new_n4924_), .A2(new_n2198_), .B(new_n4923_), .ZN(new_n14142_));
  NOR3_X1    g13119(.A1(new_n4937_), .A2(new_n4936_), .A3(new_n2199_), .ZN(new_n14143_));
  NAND4_X1   g13120(.A1(new_n14143_), .A2(new_n2091_), .A3(new_n4939_), .A4(new_n4940_), .ZN(new_n14144_));
  NOR2_X1    g13121(.A1(new_n14144_), .A2(new_n14142_), .ZN(new_n14145_));
  INV_X1     g13122(.I(new_n14145_), .ZN(new_n14146_));
  NOR2_X1    g13123(.A1(new_n4916_), .A2(new_n4949_), .ZN(new_n14147_));
  INV_X1     g13124(.I(new_n4928_), .ZN(new_n14148_));
  NAND2_X1   g13125(.A1(new_n14148_), .A2(new_n4931_), .ZN(new_n14149_));
  OAI21_X1   g13126(.A1(new_n14148_), .A2(new_n4931_), .B(new_n2091_), .ZN(new_n14150_));
  OAI21_X1   g13127(.A1(new_n14150_), .A2(new_n4933_), .B(new_n14149_), .ZN(new_n14151_));
  NAND2_X1   g13128(.A1(new_n4919_), .A2(new_n4922_), .ZN(new_n14152_));
  OAI21_X1   g13129(.A1(new_n4919_), .A2(new_n4922_), .B(new_n2198_), .ZN(new_n14153_));
  OAI21_X1   g13130(.A1(new_n4937_), .A2(new_n14153_), .B(new_n14152_), .ZN(new_n14154_));
  NAND2_X1   g13131(.A1(new_n14151_), .A2(new_n14154_), .ZN(new_n14155_));
  NOR2_X1    g13132(.A1(new_n14147_), .A2(new_n14155_), .ZN(new_n14156_));
  NAND2_X1   g13133(.A1(new_n4947_), .A2(new_n5004_), .ZN(new_n14157_));
  AOI21_X1   g13134(.A1(new_n14151_), .A2(new_n14154_), .B(new_n14157_), .ZN(new_n14158_));
  OAI21_X1   g13135(.A1(new_n14158_), .A2(new_n14156_), .B(new_n14146_), .ZN(new_n14159_));
  NAND3_X1   g13136(.A1(new_n14157_), .A2(new_n14151_), .A3(new_n14154_), .ZN(new_n14160_));
  NAND2_X1   g13137(.A1(new_n14147_), .A2(new_n14155_), .ZN(new_n14161_));
  NAND3_X1   g13138(.A1(new_n14160_), .A2(new_n14161_), .A3(new_n14145_), .ZN(new_n14162_));
  NAND2_X1   g13139(.A1(new_n14159_), .A2(new_n14162_), .ZN(new_n14163_));
  NAND2_X1   g13140(.A1(new_n14163_), .A2(new_n14141_), .ZN(new_n14164_));
  OAI21_X1   g13141(.A1(new_n14138_), .A2(new_n14139_), .B(new_n14122_), .ZN(new_n14165_));
  NAND3_X1   g13142(.A1(new_n14136_), .A2(new_n14123_), .A3(new_n14133_), .ZN(new_n14166_));
  NAND2_X1   g13143(.A1(new_n14165_), .A2(new_n14166_), .ZN(new_n14167_));
  NAND3_X1   g13144(.A1(new_n14167_), .A2(new_n14159_), .A3(new_n14162_), .ZN(new_n14168_));
  AOI21_X1   g13145(.A1(new_n14164_), .A2(new_n14168_), .B(new_n14118_), .ZN(new_n14169_));
  NAND2_X1   g13146(.A1(new_n14163_), .A2(new_n14167_), .ZN(new_n14170_));
  NAND3_X1   g13147(.A1(new_n14141_), .A2(new_n14159_), .A3(new_n14162_), .ZN(new_n14171_));
  AOI21_X1   g13148(.A1(new_n14170_), .A2(new_n14171_), .B(new_n14117_), .ZN(new_n14172_));
  NOR2_X1    g13149(.A1(new_n14169_), .A2(new_n14172_), .ZN(new_n14173_));
  AOI21_X1   g13150(.A1(new_n4907_), .A2(new_n4908_), .B(new_n5029_), .ZN(new_n14174_));
  AOI21_X1   g13151(.A1(new_n4872_), .A2(new_n2420_), .B(new_n4871_), .ZN(new_n14175_));
  NOR3_X1    g13152(.A1(new_n4872_), .A2(new_n4871_), .A3(new_n2420_), .ZN(new_n14176_));
  AOI21_X1   g13153(.A1(new_n4868_), .A2(new_n4843_), .B(new_n4862_), .ZN(new_n14177_));
  NOR3_X1    g13154(.A1(new_n4868_), .A2(new_n4862_), .A3(new_n4843_), .ZN(new_n14178_));
  NAND4_X1   g13155(.A1(new_n14178_), .A2(new_n14177_), .A3(new_n14175_), .A4(new_n14176_), .ZN(new_n14179_));
  INV_X1     g13156(.I(new_n14179_), .ZN(new_n14180_));
  NAND2_X1   g13157(.A1(new_n4881_), .A2(new_n4898_), .ZN(new_n14181_));
  NAND2_X1   g13158(.A1(new_n4861_), .A2(new_n4858_), .ZN(new_n14182_));
  NOR2_X1    g13159(.A1(new_n4861_), .A2(new_n4858_), .ZN(new_n14183_));
  NOR2_X1    g13160(.A1(new_n4843_), .A2(new_n14183_), .ZN(new_n14184_));
  NAND2_X1   g13161(.A1(new_n4875_), .A2(new_n14184_), .ZN(new_n14185_));
  NAND2_X1   g13162(.A1(new_n4849_), .A2(new_n4852_), .ZN(new_n14186_));
  NOR2_X1    g13163(.A1(new_n4849_), .A2(new_n4852_), .ZN(new_n14187_));
  NOR2_X1    g13164(.A1(new_n2420_), .A2(new_n14187_), .ZN(new_n14188_));
  NAND2_X1   g13165(.A1(new_n4854_), .A2(new_n14188_), .ZN(new_n14189_));
  AOI22_X1   g13166(.A1(new_n14185_), .A2(new_n14182_), .B1(new_n14186_), .B2(new_n14189_), .ZN(new_n14190_));
  NAND2_X1   g13167(.A1(new_n14181_), .A2(new_n14190_), .ZN(new_n14191_));
  NOR2_X1    g13168(.A1(new_n4846_), .A2(new_n4883_), .ZN(new_n14192_));
  INV_X1     g13169(.I(new_n14190_), .ZN(new_n14193_));
  NAND2_X1   g13170(.A1(new_n14192_), .A2(new_n14193_), .ZN(new_n14194_));
  AOI21_X1   g13171(.A1(new_n14191_), .A2(new_n14194_), .B(new_n14180_), .ZN(new_n14195_));
  NOR2_X1    g13172(.A1(new_n14192_), .A2(new_n14193_), .ZN(new_n14196_));
  NOR2_X1    g13173(.A1(new_n14181_), .A2(new_n14190_), .ZN(new_n14197_));
  NOR3_X1    g13174(.A1(new_n14197_), .A2(new_n14196_), .A3(new_n14179_), .ZN(new_n14198_));
  NOR2_X1    g13175(.A1(new_n14195_), .A2(new_n14198_), .ZN(new_n14199_));
  AOI21_X1   g13176(.A1(new_n4829_), .A2(new_n2641_), .B(new_n4828_), .ZN(new_n14200_));
  NAND3_X1   g13177(.A1(new_n4820_), .A2(new_n4819_), .A3(new_n2522_), .ZN(new_n14201_));
  NOR4_X1    g13178(.A1(new_n14201_), .A2(new_n2648_), .A3(new_n4809_), .A4(new_n4811_), .ZN(new_n14202_));
  NAND2_X1   g13179(.A1(new_n14202_), .A2(new_n14200_), .ZN(new_n14203_));
  NOR2_X1    g13180(.A1(new_n4891_), .A2(new_n4836_), .ZN(new_n14204_));
  NAND2_X1   g13181(.A1(new_n4815_), .A2(new_n4818_), .ZN(new_n14205_));
  OAI21_X1   g13182(.A1(new_n4815_), .A2(new_n4818_), .B(new_n2522_), .ZN(new_n14206_));
  OAI21_X1   g13183(.A1(new_n4829_), .A2(new_n14206_), .B(new_n14205_), .ZN(new_n14207_));
  NAND2_X1   g13184(.A1(new_n4805_), .A2(new_n4808_), .ZN(new_n14208_));
  OAI21_X1   g13185(.A1(new_n4805_), .A2(new_n4808_), .B(new_n4824_), .ZN(new_n14209_));
  OAI21_X1   g13186(.A1(new_n14209_), .A2(new_n4811_), .B(new_n14208_), .ZN(new_n14210_));
  NAND2_X1   g13187(.A1(new_n14210_), .A2(new_n14207_), .ZN(new_n14211_));
  NOR2_X1    g13188(.A1(new_n14204_), .A2(new_n14211_), .ZN(new_n14212_));
  NAND2_X1   g13189(.A1(new_n4838_), .A2(new_n4802_), .ZN(new_n14213_));
  INV_X1     g13190(.I(new_n14211_), .ZN(new_n14214_));
  NOR2_X1    g13191(.A1(new_n14213_), .A2(new_n14214_), .ZN(new_n14215_));
  OAI21_X1   g13192(.A1(new_n14215_), .A2(new_n14212_), .B(new_n14203_), .ZN(new_n14216_));
  NAND2_X1   g13193(.A1(new_n14213_), .A2(new_n14214_), .ZN(new_n14217_));
  NAND2_X1   g13194(.A1(new_n14204_), .A2(new_n14211_), .ZN(new_n14218_));
  NAND4_X1   g13195(.A1(new_n14217_), .A2(new_n14218_), .A3(new_n14200_), .A4(new_n14202_), .ZN(new_n14219_));
  NAND2_X1   g13196(.A1(new_n14219_), .A2(new_n14216_), .ZN(new_n14220_));
  NAND2_X1   g13197(.A1(new_n14199_), .A2(new_n14220_), .ZN(new_n14221_));
  OAI21_X1   g13198(.A1(new_n14197_), .A2(new_n14196_), .B(new_n14179_), .ZN(new_n14222_));
  NAND3_X1   g13199(.A1(new_n14191_), .A2(new_n14194_), .A3(new_n14180_), .ZN(new_n14223_));
  NAND2_X1   g13200(.A1(new_n14222_), .A2(new_n14223_), .ZN(new_n14224_));
  AND2_X2    g13201(.A1(new_n14219_), .A2(new_n14216_), .Z(new_n14225_));
  NAND2_X1   g13202(.A1(new_n14225_), .A2(new_n14224_), .ZN(new_n14226_));
  AOI21_X1   g13203(.A1(new_n14226_), .A2(new_n14221_), .B(new_n14174_), .ZN(new_n14227_));
  OAI21_X1   g13204(.A1(new_n4799_), .A2(new_n5028_), .B(new_n4909_), .ZN(new_n14228_));
  NAND2_X1   g13205(.A1(new_n14224_), .A2(new_n14220_), .ZN(new_n14229_));
  NAND3_X1   g13206(.A1(new_n14199_), .A2(new_n14216_), .A3(new_n14219_), .ZN(new_n14230_));
  AOI21_X1   g13207(.A1(new_n14230_), .A2(new_n14229_), .B(new_n14228_), .ZN(new_n14231_));
  OAI21_X1   g13208(.A1(new_n14227_), .A2(new_n14231_), .B(new_n14173_), .ZN(new_n14232_));
  AOI21_X1   g13209(.A1(new_n14159_), .A2(new_n14162_), .B(new_n14167_), .ZN(new_n14233_));
  NOR2_X1    g13210(.A1(new_n14163_), .A2(new_n14141_), .ZN(new_n14234_));
  OAI21_X1   g13211(.A1(new_n14234_), .A2(new_n14233_), .B(new_n14117_), .ZN(new_n14235_));
  AOI21_X1   g13212(.A1(new_n14159_), .A2(new_n14162_), .B(new_n14141_), .ZN(new_n14236_));
  AOI21_X1   g13213(.A1(new_n14160_), .A2(new_n14161_), .B(new_n14145_), .ZN(new_n14237_));
  NOR3_X1    g13214(.A1(new_n14158_), .A2(new_n14146_), .A3(new_n14156_), .ZN(new_n14238_));
  NOR3_X1    g13215(.A1(new_n14167_), .A2(new_n14238_), .A3(new_n14237_), .ZN(new_n14239_));
  OAI21_X1   g13216(.A1(new_n14236_), .A2(new_n14239_), .B(new_n14118_), .ZN(new_n14240_));
  NAND2_X1   g13217(.A1(new_n14235_), .A2(new_n14240_), .ZN(new_n14241_));
  NOR2_X1    g13218(.A1(new_n14225_), .A2(new_n14224_), .ZN(new_n14242_));
  NOR2_X1    g13219(.A1(new_n14199_), .A2(new_n14220_), .ZN(new_n14243_));
  OAI21_X1   g13220(.A1(new_n14242_), .A2(new_n14243_), .B(new_n14228_), .ZN(new_n14244_));
  NOR2_X1    g13221(.A1(new_n14225_), .A2(new_n14199_), .ZN(new_n14245_));
  NOR2_X1    g13222(.A1(new_n14224_), .A2(new_n14220_), .ZN(new_n14246_));
  OAI21_X1   g13223(.A1(new_n14245_), .A2(new_n14246_), .B(new_n14174_), .ZN(new_n14247_));
  NAND3_X1   g13224(.A1(new_n14241_), .A2(new_n14244_), .A3(new_n14247_), .ZN(new_n14248_));
  AOI21_X1   g13225(.A1(new_n14232_), .A2(new_n14248_), .B(new_n14116_), .ZN(new_n14249_));
  INV_X1     g13226(.I(new_n14116_), .ZN(new_n14250_));
  OAI22_X1   g13227(.A1(new_n14227_), .A2(new_n14231_), .B1(new_n14169_), .B2(new_n14172_), .ZN(new_n14251_));
  NAND4_X1   g13228(.A1(new_n14244_), .A2(new_n14247_), .A3(new_n14235_), .A4(new_n14240_), .ZN(new_n14252_));
  AOI21_X1   g13229(.A1(new_n14252_), .A2(new_n14251_), .B(new_n14250_), .ZN(new_n14253_));
  NOR2_X1    g13230(.A1(new_n14249_), .A2(new_n14253_), .ZN(new_n14254_));
  NOR2_X1    g13231(.A1(new_n14115_), .A2(new_n14254_), .ZN(new_n14255_));
  AOI21_X1   g13232(.A1(new_n14244_), .A2(new_n14247_), .B(new_n14241_), .ZN(new_n14256_));
  NOR3_X1    g13233(.A1(new_n14173_), .A2(new_n14227_), .A3(new_n14231_), .ZN(new_n14257_));
  OAI21_X1   g13234(.A1(new_n14256_), .A2(new_n14257_), .B(new_n14250_), .ZN(new_n14258_));
  AOI22_X1   g13235(.A1(new_n14244_), .A2(new_n14247_), .B1(new_n14235_), .B2(new_n14240_), .ZN(new_n14259_));
  NOR4_X1    g13236(.A1(new_n14227_), .A2(new_n14231_), .A3(new_n14169_), .A4(new_n14172_), .ZN(new_n14260_));
  OAI21_X1   g13237(.A1(new_n14259_), .A2(new_n14260_), .B(new_n14116_), .ZN(new_n14261_));
  NAND2_X1   g13238(.A1(new_n14258_), .A2(new_n14261_), .ZN(new_n14262_));
  AOI21_X1   g13239(.A1(new_n5341_), .A2(new_n14114_), .B(new_n14262_), .ZN(new_n14263_));
  OAI21_X1   g13240(.A1(new_n14263_), .A2(new_n14255_), .B(new_n14113_), .ZN(new_n14264_));
  INV_X1     g13241(.I(new_n14264_), .ZN(new_n14265_));
  NAND2_X1   g13242(.A1(new_n14115_), .A2(new_n14262_), .ZN(new_n14266_));
  NOR2_X1    g13243(.A1(new_n14115_), .A2(new_n14262_), .ZN(new_n14267_));
  INV_X1     g13244(.I(new_n14267_), .ZN(new_n14268_));
  AOI21_X1   g13245(.A1(new_n14268_), .A2(new_n14266_), .B(new_n14113_), .ZN(new_n14269_));
  NOR2_X1    g13246(.A1(new_n14265_), .A2(new_n14269_), .ZN(new_n14270_));
  OAI21_X1   g13247(.A1(new_n13977_), .A2(new_n4273_), .B(new_n4781_), .ZN(new_n14271_));
  NAND2_X1   g13248(.A1(new_n4775_), .A2(new_n4511_), .ZN(new_n14272_));
  NAND2_X1   g13249(.A1(new_n14272_), .A2(new_n4776_), .ZN(new_n14273_));
  OAI21_X1   g13250(.A1(new_n4623_), .A2(new_n4759_), .B(new_n4745_), .ZN(new_n14274_));
  AOI21_X1   g13251(.A1(new_n4712_), .A2(new_n4693_), .B(new_n4711_), .ZN(new_n14275_));
  NAND3_X1   g13252(.A1(new_n4701_), .A2(new_n4694_), .A3(new_n4700_), .ZN(new_n14276_));
  NOR4_X1    g13253(.A1(new_n14276_), .A2(new_n4682_), .A3(new_n4689_), .A4(new_n4691_), .ZN(new_n14277_));
  NAND2_X1   g13254(.A1(new_n14277_), .A2(new_n14275_), .ZN(new_n14278_));
  NOR2_X1    g13255(.A1(new_n4680_), .A2(new_n4720_), .ZN(new_n14279_));
  NOR2_X1    g13256(.A1(new_n4697_), .A2(new_n4699_), .ZN(new_n14280_));
  INV_X1     g13257(.I(new_n14280_), .ZN(new_n14281_));
  NAND2_X1   g13258(.A1(new_n4697_), .A2(new_n4699_), .ZN(new_n14282_));
  NAND3_X1   g13259(.A1(new_n4701_), .A2(new_n4694_), .A3(new_n14282_), .ZN(new_n14283_));
  NAND2_X1   g13260(.A1(new_n4688_), .A2(new_n4685_), .ZN(new_n14284_));
  NOR2_X1    g13261(.A1(new_n4688_), .A2(new_n4685_), .ZN(new_n14285_));
  NOR2_X1    g13262(.A1(new_n4682_), .A2(new_n14285_), .ZN(new_n14286_));
  NAND2_X1   g13263(.A1(new_n4718_), .A2(new_n14286_), .ZN(new_n14287_));
  AOI22_X1   g13264(.A1(new_n14283_), .A2(new_n14281_), .B1(new_n14287_), .B2(new_n14284_), .ZN(new_n14288_));
  INV_X1     g13265(.I(new_n14288_), .ZN(new_n14289_));
  NOR2_X1    g13266(.A1(new_n14279_), .A2(new_n14289_), .ZN(new_n14290_));
  NAND2_X1   g13267(.A1(new_n4710_), .A2(new_n4734_), .ZN(new_n14291_));
  NOR2_X1    g13268(.A1(new_n14291_), .A2(new_n14288_), .ZN(new_n14292_));
  OAI21_X1   g13269(.A1(new_n14290_), .A2(new_n14292_), .B(new_n14278_), .ZN(new_n14293_));
  INV_X1     g13270(.I(new_n14278_), .ZN(new_n14294_));
  NAND2_X1   g13271(.A1(new_n14291_), .A2(new_n14288_), .ZN(new_n14295_));
  NAND2_X1   g13272(.A1(new_n14279_), .A2(new_n14289_), .ZN(new_n14296_));
  NAND3_X1   g13273(.A1(new_n14296_), .A2(new_n14295_), .A3(new_n14294_), .ZN(new_n14297_));
  NAND2_X1   g13274(.A1(new_n14297_), .A2(new_n14293_), .ZN(new_n14298_));
  OAI21_X1   g13275(.A1(new_n4652_), .A2(new_n4644_), .B(new_n4651_), .ZN(new_n14299_));
  NOR3_X1    g13276(.A1(new_n4663_), .A2(new_n4662_), .A3(new_n3754_), .ZN(new_n14300_));
  NAND4_X1   g13277(.A1(new_n14300_), .A2(new_n4655_), .A3(new_n4656_), .A4(new_n4660_), .ZN(new_n14301_));
  NOR2_X1    g13278(.A1(new_n14301_), .A2(new_n14299_), .ZN(new_n14302_));
  NAND2_X1   g13279(.A1(new_n4650_), .A2(new_n4647_), .ZN(new_n14303_));
  NOR2_X1    g13280(.A1(new_n4650_), .A2(new_n4647_), .ZN(new_n14304_));
  NOR2_X1    g13281(.A1(new_n3754_), .A2(new_n14304_), .ZN(new_n14305_));
  NAND2_X1   g13282(.A1(new_n14305_), .A2(new_n4652_), .ZN(new_n14306_));
  NAND2_X1   g13283(.A1(new_n4636_), .A2(new_n4634_), .ZN(new_n14307_));
  NOR2_X1    g13284(.A1(new_n4636_), .A2(new_n4634_), .ZN(new_n14308_));
  NOR2_X1    g13285(.A1(new_n4631_), .A2(new_n14308_), .ZN(new_n14309_));
  NAND2_X1   g13286(.A1(new_n14309_), .A2(new_n4660_), .ZN(new_n14310_));
  AOI22_X1   g13287(.A1(new_n14303_), .A2(new_n14306_), .B1(new_n14310_), .B2(new_n14307_), .ZN(new_n14311_));
  OAI21_X1   g13288(.A1(new_n4672_), .A2(new_n4728_), .B(new_n14311_), .ZN(new_n14312_));
  NOR2_X1    g13289(.A1(new_n4672_), .A2(new_n4728_), .ZN(new_n14313_));
  NAND2_X1   g13290(.A1(new_n14306_), .A2(new_n14303_), .ZN(new_n14314_));
  NAND2_X1   g13291(.A1(new_n14310_), .A2(new_n14307_), .ZN(new_n14315_));
  NAND2_X1   g13292(.A1(new_n14314_), .A2(new_n14315_), .ZN(new_n14316_));
  NAND2_X1   g13293(.A1(new_n14313_), .A2(new_n14316_), .ZN(new_n14317_));
  AOI21_X1   g13294(.A1(new_n14317_), .A2(new_n14312_), .B(new_n14302_), .ZN(new_n14318_));
  INV_X1     g13295(.I(new_n14302_), .ZN(new_n14319_));
  NOR2_X1    g13296(.A1(new_n14313_), .A2(new_n14316_), .ZN(new_n14320_));
  NOR3_X1    g13297(.A1(new_n14311_), .A2(new_n4672_), .A3(new_n4728_), .ZN(new_n14321_));
  NOR3_X1    g13298(.A1(new_n14320_), .A2(new_n14319_), .A3(new_n14321_), .ZN(new_n14322_));
  NOR2_X1    g13299(.A1(new_n14322_), .A2(new_n14318_), .ZN(new_n14323_));
  NOR2_X1    g13300(.A1(new_n14298_), .A2(new_n14323_), .ZN(new_n14324_));
  AOI21_X1   g13301(.A1(new_n14296_), .A2(new_n14295_), .B(new_n14294_), .ZN(new_n14325_));
  NOR3_X1    g13302(.A1(new_n14290_), .A2(new_n14292_), .A3(new_n14278_), .ZN(new_n14326_));
  NOR2_X1    g13303(.A1(new_n14325_), .A2(new_n14326_), .ZN(new_n14327_));
  OAI21_X1   g13304(.A1(new_n14320_), .A2(new_n14321_), .B(new_n14319_), .ZN(new_n14328_));
  NAND3_X1   g13305(.A1(new_n14317_), .A2(new_n14312_), .A3(new_n14302_), .ZN(new_n14329_));
  NAND2_X1   g13306(.A1(new_n14328_), .A2(new_n14329_), .ZN(new_n14330_));
  NOR2_X1    g13307(.A1(new_n14327_), .A2(new_n14330_), .ZN(new_n14331_));
  OAI21_X1   g13308(.A1(new_n14324_), .A2(new_n14331_), .B(new_n14274_), .ZN(new_n14332_));
  AOI21_X1   g13309(.A1(new_n4744_), .A2(new_n4743_), .B(new_n4760_), .ZN(new_n14333_));
  NOR2_X1    g13310(.A1(new_n14327_), .A2(new_n14323_), .ZN(new_n14334_));
  NOR2_X1    g13311(.A1(new_n14298_), .A2(new_n14330_), .ZN(new_n14335_));
  OAI21_X1   g13312(.A1(new_n14334_), .A2(new_n14335_), .B(new_n14333_), .ZN(new_n14336_));
  NAND2_X1   g13313(.A1(new_n14332_), .A2(new_n14336_), .ZN(new_n14337_));
  AOI21_X1   g13314(.A1(new_n4752_), .A2(new_n4516_), .B(new_n4619_), .ZN(new_n14338_));
  AOI21_X1   g13315(.A1(new_n4584_), .A2(new_n4577_), .B(new_n4583_), .ZN(new_n14339_));
  NAND3_X1   g13316(.A1(new_n4593_), .A2(new_n4591_), .A3(new_n4592_), .ZN(new_n14340_));
  NOR4_X1    g13317(.A1(new_n14340_), .A2(new_n3833_), .A3(new_n4587_), .A4(new_n4589_), .ZN(new_n14341_));
  NAND2_X1   g13318(.A1(new_n14341_), .A2(new_n14339_), .ZN(new_n14342_));
  NOR2_X1    g13319(.A1(new_n4566_), .A2(new_n4598_), .ZN(new_n14343_));
  NOR2_X1    g13320(.A1(new_n4580_), .A2(new_n4582_), .ZN(new_n14344_));
  INV_X1     g13321(.I(new_n14344_), .ZN(new_n14345_));
  NAND2_X1   g13322(.A1(new_n4580_), .A2(new_n4582_), .ZN(new_n14346_));
  NAND3_X1   g13323(.A1(new_n4593_), .A2(new_n4591_), .A3(new_n14346_), .ZN(new_n14347_));
  NAND2_X1   g13324(.A1(new_n4573_), .A2(new_n4570_), .ZN(new_n14348_));
  NOR2_X1    g13325(.A1(new_n4573_), .A2(new_n4570_), .ZN(new_n14349_));
  NOR2_X1    g13326(.A1(new_n3833_), .A2(new_n14349_), .ZN(new_n14350_));
  NAND2_X1   g13327(.A1(new_n4575_), .A2(new_n14350_), .ZN(new_n14351_));
  AOI22_X1   g13328(.A1(new_n14347_), .A2(new_n14345_), .B1(new_n14351_), .B2(new_n14348_), .ZN(new_n14352_));
  INV_X1     g13329(.I(new_n14352_), .ZN(new_n14353_));
  NOR2_X1    g13330(.A1(new_n14343_), .A2(new_n14353_), .ZN(new_n14354_));
  NOR3_X1    g13331(.A1(new_n4566_), .A2(new_n14352_), .A3(new_n4598_), .ZN(new_n14355_));
  OAI21_X1   g13332(.A1(new_n14354_), .A2(new_n14355_), .B(new_n14342_), .ZN(new_n14356_));
  INV_X1     g13333(.I(new_n14342_), .ZN(new_n14357_));
  OAI21_X1   g13334(.A1(new_n4566_), .A2(new_n4598_), .B(new_n14352_), .ZN(new_n14358_));
  NAND2_X1   g13335(.A1(new_n14343_), .A2(new_n14353_), .ZN(new_n14359_));
  NAND3_X1   g13336(.A1(new_n14359_), .A2(new_n14357_), .A3(new_n14358_), .ZN(new_n14360_));
  AND2_X2    g13337(.A1(new_n14356_), .A2(new_n14360_), .Z(new_n14361_));
  AOI21_X1   g13338(.A1(new_n4541_), .A2(new_n3916_), .B(new_n4540_), .ZN(new_n14362_));
  NAND3_X1   g13339(.A1(new_n4550_), .A2(new_n4548_), .A3(new_n4549_), .ZN(new_n14363_));
  NOR4_X1    g13340(.A1(new_n14363_), .A2(new_n4522_), .A3(new_n4544_), .A4(new_n4546_), .ZN(new_n14364_));
  NAND2_X1   g13341(.A1(new_n14364_), .A2(new_n14362_), .ZN(new_n14365_));
  NOR2_X1    g13342(.A1(new_n4520_), .A2(new_n4559_), .ZN(new_n14366_));
  NAND2_X1   g13343(.A1(new_n4539_), .A2(new_n4535_), .ZN(new_n14367_));
  NOR2_X1    g13344(.A1(new_n4539_), .A2(new_n4535_), .ZN(new_n14368_));
  NOR2_X1    g13345(.A1(new_n3916_), .A2(new_n14368_), .ZN(new_n14369_));
  NAND2_X1   g13346(.A1(new_n4550_), .A2(new_n14369_), .ZN(new_n14370_));
  NAND2_X1   g13347(.A1(new_n4528_), .A2(new_n4526_), .ZN(new_n14371_));
  NOR2_X1    g13348(.A1(new_n4528_), .A2(new_n4526_), .ZN(new_n14372_));
  NOR2_X1    g13349(.A1(new_n4522_), .A2(new_n14372_), .ZN(new_n14373_));
  NAND2_X1   g13350(.A1(new_n14373_), .A2(new_n4531_), .ZN(new_n14374_));
  AOI22_X1   g13351(.A1(new_n14374_), .A2(new_n14371_), .B1(new_n14370_), .B2(new_n14367_), .ZN(new_n14375_));
  INV_X1     g13352(.I(new_n14375_), .ZN(new_n14376_));
  NOR2_X1    g13353(.A1(new_n14366_), .A2(new_n14376_), .ZN(new_n14377_));
  NAND2_X1   g13354(.A1(new_n4606_), .A2(new_n4557_), .ZN(new_n14378_));
  NOR2_X1    g13355(.A1(new_n14378_), .A2(new_n14375_), .ZN(new_n14379_));
  OAI21_X1   g13356(.A1(new_n14377_), .A2(new_n14379_), .B(new_n14365_), .ZN(new_n14380_));
  INV_X1     g13357(.I(new_n14365_), .ZN(new_n14381_));
  NAND2_X1   g13358(.A1(new_n14378_), .A2(new_n14375_), .ZN(new_n14382_));
  NAND2_X1   g13359(.A1(new_n14366_), .A2(new_n14376_), .ZN(new_n14383_));
  NAND3_X1   g13360(.A1(new_n14383_), .A2(new_n14382_), .A3(new_n14381_), .ZN(new_n14384_));
  NAND2_X1   g13361(.A1(new_n14380_), .A2(new_n14384_), .ZN(new_n14385_));
  NAND2_X1   g13362(.A1(new_n14361_), .A2(new_n14385_), .ZN(new_n14386_));
  NAND2_X1   g13363(.A1(new_n14356_), .A2(new_n14360_), .ZN(new_n14387_));
  AOI21_X1   g13364(.A1(new_n14383_), .A2(new_n14382_), .B(new_n14381_), .ZN(new_n14388_));
  NOR3_X1    g13365(.A1(new_n14377_), .A2(new_n14379_), .A3(new_n14365_), .ZN(new_n14389_));
  NOR2_X1    g13366(.A1(new_n14389_), .A2(new_n14388_), .ZN(new_n14390_));
  NAND2_X1   g13367(.A1(new_n14390_), .A2(new_n14387_), .ZN(new_n14391_));
  AOI21_X1   g13368(.A1(new_n14386_), .A2(new_n14391_), .B(new_n14338_), .ZN(new_n14392_));
  OAI21_X1   g13369(.A1(new_n4617_), .A2(new_n4618_), .B(new_n4753_), .ZN(new_n14393_));
  NAND2_X1   g13370(.A1(new_n14387_), .A2(new_n14385_), .ZN(new_n14394_));
  NAND3_X1   g13371(.A1(new_n14390_), .A2(new_n14356_), .A3(new_n14360_), .ZN(new_n14395_));
  AOI21_X1   g13372(.A1(new_n14395_), .A2(new_n14394_), .B(new_n14393_), .ZN(new_n14396_));
  NOR2_X1    g13373(.A1(new_n14392_), .A2(new_n14396_), .ZN(new_n14397_));
  NOR2_X1    g13374(.A1(new_n14397_), .A2(new_n14337_), .ZN(new_n14398_));
  NAND2_X1   g13375(.A1(new_n14327_), .A2(new_n14330_), .ZN(new_n14399_));
  NAND2_X1   g13376(.A1(new_n14298_), .A2(new_n14323_), .ZN(new_n14400_));
  AOI21_X1   g13377(.A1(new_n14400_), .A2(new_n14399_), .B(new_n14333_), .ZN(new_n14401_));
  NAND2_X1   g13378(.A1(new_n14298_), .A2(new_n14330_), .ZN(new_n14402_));
  NAND2_X1   g13379(.A1(new_n14327_), .A2(new_n14323_), .ZN(new_n14403_));
  AOI21_X1   g13380(.A1(new_n14403_), .A2(new_n14402_), .B(new_n14274_), .ZN(new_n14404_));
  NOR2_X1    g13381(.A1(new_n14401_), .A2(new_n14404_), .ZN(new_n14405_));
  NOR2_X1    g13382(.A1(new_n14390_), .A2(new_n14387_), .ZN(new_n14406_));
  NOR2_X1    g13383(.A1(new_n14361_), .A2(new_n14385_), .ZN(new_n14407_));
  OAI21_X1   g13384(.A1(new_n14407_), .A2(new_n14406_), .B(new_n14393_), .ZN(new_n14408_));
  NOR2_X1    g13385(.A1(new_n14361_), .A2(new_n14390_), .ZN(new_n14409_));
  NOR2_X1    g13386(.A1(new_n14387_), .A2(new_n14385_), .ZN(new_n14410_));
  OAI21_X1   g13387(.A1(new_n14409_), .A2(new_n14410_), .B(new_n14338_), .ZN(new_n14411_));
  NAND2_X1   g13388(.A1(new_n14408_), .A2(new_n14411_), .ZN(new_n14412_));
  NOR2_X1    g13389(.A1(new_n14412_), .A2(new_n14405_), .ZN(new_n14413_));
  OAI21_X1   g13390(.A1(new_n14413_), .A2(new_n14398_), .B(new_n14273_), .ZN(new_n14414_));
  AOI21_X1   g13391(.A1(new_n4511_), .A2(new_n4775_), .B(new_n4767_), .ZN(new_n14415_));
  OAI22_X1   g13392(.A1(new_n14392_), .A2(new_n14396_), .B1(new_n14401_), .B2(new_n14404_), .ZN(new_n14416_));
  NAND4_X1   g13393(.A1(new_n14408_), .A2(new_n14411_), .A3(new_n14332_), .A4(new_n14336_), .ZN(new_n14417_));
  NAND2_X1   g13394(.A1(new_n14417_), .A2(new_n14416_), .ZN(new_n14418_));
  NAND2_X1   g13395(.A1(new_n14418_), .A2(new_n14415_), .ZN(new_n14419_));
  NAND2_X1   g13396(.A1(new_n14419_), .A2(new_n14414_), .ZN(new_n14420_));
  AOI21_X1   g13397(.A1(new_n4785_), .A2(new_n4276_), .B(new_n4507_), .ZN(new_n14421_));
  AOI21_X1   g13398(.A1(new_n4485_), .A2(new_n4484_), .B(new_n4501_), .ZN(new_n14422_));
  AOI21_X1   g13399(.A1(new_n4459_), .A2(new_n4440_), .B(new_n4457_), .ZN(new_n14423_));
  NAND3_X1   g13400(.A1(new_n4448_), .A2(new_n4441_), .A3(new_n4447_), .ZN(new_n14424_));
  NOR4_X1    g13401(.A1(new_n14424_), .A2(new_n3996_), .A3(new_n4437_), .A4(new_n4438_), .ZN(new_n14425_));
  NAND2_X1   g13402(.A1(new_n14425_), .A2(new_n14423_), .ZN(new_n14426_));
  INV_X1     g13403(.I(new_n14426_), .ZN(new_n14427_));
  NAND2_X1   g13404(.A1(new_n4455_), .A2(new_n4475_), .ZN(new_n14428_));
  NAND2_X1   g13405(.A1(new_n4446_), .A2(new_n4444_), .ZN(new_n14429_));
  NAND3_X1   g13406(.A1(new_n4456_), .A2(new_n2960_), .A3(new_n4445_), .ZN(new_n14430_));
  NAND3_X1   g13407(.A1(new_n4448_), .A2(new_n4441_), .A3(new_n14430_), .ZN(new_n14431_));
  NOR2_X1    g13408(.A1(new_n4436_), .A2(new_n4434_), .ZN(new_n14432_));
  NOR2_X1    g13409(.A1(new_n3996_), .A2(new_n14432_), .ZN(new_n14433_));
  AOI22_X1   g13410(.A1(new_n4463_), .A2(new_n14433_), .B1(new_n4434_), .B2(new_n4436_), .ZN(new_n14434_));
  AOI21_X1   g13411(.A1(new_n14429_), .A2(new_n14431_), .B(new_n14434_), .ZN(new_n14435_));
  NAND2_X1   g13412(.A1(new_n14428_), .A2(new_n14435_), .ZN(new_n14436_));
  NOR2_X1    g13413(.A1(new_n4431_), .A2(new_n4465_), .ZN(new_n14437_));
  NAND2_X1   g13414(.A1(new_n14431_), .A2(new_n14429_), .ZN(new_n14438_));
  INV_X1     g13415(.I(new_n14434_), .ZN(new_n14439_));
  NAND2_X1   g13416(.A1(new_n14439_), .A2(new_n14438_), .ZN(new_n14440_));
  NAND2_X1   g13417(.A1(new_n14437_), .A2(new_n14440_), .ZN(new_n14441_));
  AOI21_X1   g13418(.A1(new_n14441_), .A2(new_n14436_), .B(new_n14427_), .ZN(new_n14442_));
  NOR2_X1    g13419(.A1(new_n14437_), .A2(new_n14440_), .ZN(new_n14443_));
  NOR2_X1    g13420(.A1(new_n14428_), .A2(new_n14435_), .ZN(new_n14444_));
  NOR3_X1    g13421(.A1(new_n14443_), .A2(new_n14444_), .A3(new_n14426_), .ZN(new_n14445_));
  NOR2_X1    g13422(.A1(new_n14442_), .A2(new_n14445_), .ZN(new_n14446_));
  OAI21_X1   g13423(.A1(new_n4416_), .A2(new_n4080_), .B(new_n4415_), .ZN(new_n14447_));
  NAND3_X1   g13424(.A1(new_n4416_), .A2(new_n4080_), .A3(new_n4415_), .ZN(new_n14448_));
  INV_X1     g13425(.I(new_n4086_), .ZN(new_n14449_));
  INV_X1     g13426(.I(new_n4410_), .ZN(new_n14450_));
  INV_X1     g13427(.I(new_n4411_), .ZN(new_n14451_));
  OAI21_X1   g13428(.A1(new_n14451_), .A2(new_n14449_), .B(new_n14450_), .ZN(new_n14452_));
  NAND3_X1   g13429(.A1(new_n14451_), .A2(new_n14450_), .A3(new_n14449_), .ZN(new_n14453_));
  NOR4_X1    g13430(.A1(new_n14452_), .A2(new_n14453_), .A3(new_n14447_), .A4(new_n14448_), .ZN(new_n14454_));
  INV_X1     g13431(.I(new_n14454_), .ZN(new_n14455_));
  NAND2_X1   g13432(.A1(new_n4409_), .A2(new_n4407_), .ZN(new_n14456_));
  INV_X1     g13433(.I(new_n14456_), .ZN(new_n14457_));
  NOR2_X1    g13434(.A1(new_n4409_), .A2(new_n4407_), .ZN(new_n14458_));
  OR2_X2     g13435(.A1(new_n4086_), .A2(new_n14458_), .Z(new_n14459_));
  NOR2_X1    g13436(.A1(new_n14459_), .A2(new_n4411_), .ZN(new_n14460_));
  NAND2_X1   g13437(.A1(new_n4401_), .A2(new_n4399_), .ZN(new_n14461_));
  INV_X1     g13438(.I(new_n14461_), .ZN(new_n14462_));
  NOR2_X1    g13439(.A1(new_n4401_), .A2(new_n4399_), .ZN(new_n14463_));
  NOR3_X1    g13440(.A1(new_n4403_), .A2(new_n4093_), .A3(new_n14463_), .ZN(new_n14464_));
  OAI22_X1   g13441(.A1(new_n14464_), .A2(new_n14462_), .B1(new_n14457_), .B2(new_n14460_), .ZN(new_n14465_));
  AOI21_X1   g13442(.A1(new_n4396_), .A2(new_n4424_), .B(new_n14465_), .ZN(new_n14466_));
  NAND3_X1   g13443(.A1(new_n14465_), .A2(new_n4396_), .A3(new_n4424_), .ZN(new_n14467_));
  INV_X1     g13444(.I(new_n14467_), .ZN(new_n14468_));
  OAI21_X1   g13445(.A1(new_n14468_), .A2(new_n14466_), .B(new_n14455_), .ZN(new_n14469_));
  NAND2_X1   g13446(.A1(new_n4396_), .A2(new_n4424_), .ZN(new_n14470_));
  INV_X1     g13447(.I(new_n14465_), .ZN(new_n14471_));
  NAND2_X1   g13448(.A1(new_n14470_), .A2(new_n14471_), .ZN(new_n14472_));
  NAND3_X1   g13449(.A1(new_n14472_), .A2(new_n14467_), .A3(new_n14454_), .ZN(new_n14473_));
  NAND2_X1   g13450(.A1(new_n14469_), .A2(new_n14473_), .ZN(new_n14474_));
  NAND2_X1   g13451(.A1(new_n14446_), .A2(new_n14474_), .ZN(new_n14475_));
  OAI21_X1   g13452(.A1(new_n14443_), .A2(new_n14444_), .B(new_n14426_), .ZN(new_n14476_));
  NAND3_X1   g13453(.A1(new_n14441_), .A2(new_n14436_), .A3(new_n14427_), .ZN(new_n14477_));
  NAND2_X1   g13454(.A1(new_n14476_), .A2(new_n14477_), .ZN(new_n14478_));
  AOI21_X1   g13455(.A1(new_n14472_), .A2(new_n14467_), .B(new_n14454_), .ZN(new_n14479_));
  NOR3_X1    g13456(.A1(new_n14468_), .A2(new_n14455_), .A3(new_n14466_), .ZN(new_n14480_));
  NOR2_X1    g13457(.A1(new_n14480_), .A2(new_n14479_), .ZN(new_n14481_));
  NAND2_X1   g13458(.A1(new_n14478_), .A2(new_n14481_), .ZN(new_n14482_));
  AOI21_X1   g13459(.A1(new_n14482_), .A2(new_n14475_), .B(new_n14422_), .ZN(new_n14483_));
  OAI21_X1   g13460(.A1(new_n4393_), .A2(new_n4500_), .B(new_n4486_), .ZN(new_n14484_));
  NAND2_X1   g13461(.A1(new_n14478_), .A2(new_n14474_), .ZN(new_n14485_));
  NAND2_X1   g13462(.A1(new_n14446_), .A2(new_n14481_), .ZN(new_n14486_));
  AOI21_X1   g13463(.A1(new_n14486_), .A2(new_n14485_), .B(new_n14484_), .ZN(new_n14487_));
  NOR2_X1    g13464(.A1(new_n14483_), .A2(new_n14487_), .ZN(new_n14488_));
  OAI21_X1   g13465(.A1(new_n4387_), .A2(new_n4388_), .B(new_n4494_), .ZN(new_n14489_));
  OAI21_X1   g13466(.A1(new_n4351_), .A2(new_n4344_), .B(new_n4350_), .ZN(new_n14490_));
  NOR3_X1    g13467(.A1(new_n4358_), .A2(new_n4357_), .A3(new_n4343_), .ZN(new_n14491_));
  NAND4_X1   g13468(.A1(new_n14491_), .A2(new_n4172_), .A3(new_n4354_), .A4(new_n4355_), .ZN(new_n14492_));
  NOR2_X1    g13469(.A1(new_n14492_), .A2(new_n14490_), .ZN(new_n14493_));
  INV_X1     g13470(.I(new_n14493_), .ZN(new_n14494_));
  NOR2_X1    g13471(.A1(new_n4365_), .A2(new_n4381_), .ZN(new_n14495_));
  NAND2_X1   g13472(.A1(new_n4349_), .A2(new_n4347_), .ZN(new_n14496_));
  NOR2_X1    g13473(.A1(new_n4349_), .A2(new_n4347_), .ZN(new_n14497_));
  NOR2_X1    g13474(.A1(new_n4343_), .A2(new_n14497_), .ZN(new_n14498_));
  NAND2_X1   g13475(.A1(new_n4351_), .A2(new_n14498_), .ZN(new_n14499_));
  NAND2_X1   g13476(.A1(new_n14499_), .A2(new_n14496_), .ZN(new_n14500_));
  NAND2_X1   g13477(.A1(new_n4338_), .A2(new_n4336_), .ZN(new_n14501_));
  NOR2_X1    g13478(.A1(new_n4338_), .A2(new_n4336_), .ZN(new_n14502_));
  NOR2_X1    g13479(.A1(new_n4160_), .A2(new_n14502_), .ZN(new_n14503_));
  NAND2_X1   g13480(.A1(new_n4355_), .A2(new_n14503_), .ZN(new_n14504_));
  NAND2_X1   g13481(.A1(new_n14504_), .A2(new_n14501_), .ZN(new_n14505_));
  NAND2_X1   g13482(.A1(new_n14500_), .A2(new_n14505_), .ZN(new_n14506_));
  NOR2_X1    g13483(.A1(new_n14495_), .A2(new_n14506_), .ZN(new_n14507_));
  AOI22_X1   g13484(.A1(new_n14501_), .A2(new_n14504_), .B1(new_n14499_), .B2(new_n14496_), .ZN(new_n14508_));
  NOR3_X1    g13485(.A1(new_n14508_), .A2(new_n4365_), .A3(new_n4381_), .ZN(new_n14509_));
  OAI21_X1   g13486(.A1(new_n14507_), .A2(new_n14509_), .B(new_n14494_), .ZN(new_n14510_));
  OAI21_X1   g13487(.A1(new_n4365_), .A2(new_n4381_), .B(new_n14508_), .ZN(new_n14511_));
  NAND3_X1   g13488(.A1(new_n14506_), .A2(new_n4333_), .A3(new_n4367_), .ZN(new_n14512_));
  NAND3_X1   g13489(.A1(new_n14512_), .A2(new_n14511_), .A3(new_n14493_), .ZN(new_n14513_));
  NAND2_X1   g13490(.A1(new_n14510_), .A2(new_n14513_), .ZN(new_n14514_));
  AOI21_X1   g13491(.A1(new_n4318_), .A2(new_n4243_), .B(new_n4317_), .ZN(new_n14515_));
  NAND3_X1   g13492(.A1(new_n4301_), .A2(new_n4300_), .A3(new_n4294_), .ZN(new_n14516_));
  NOR4_X1    g13493(.A1(new_n14516_), .A2(new_n4250_), .A3(new_n4290_), .A4(new_n4292_), .ZN(new_n14517_));
  NAND2_X1   g13494(.A1(new_n14517_), .A2(new_n14515_), .ZN(new_n14518_));
  INV_X1     g13495(.I(new_n14518_), .ZN(new_n14519_));
  NAND2_X1   g13496(.A1(new_n4299_), .A2(new_n4297_), .ZN(new_n14520_));
  NOR2_X1    g13497(.A1(new_n4299_), .A2(new_n4297_), .ZN(new_n14521_));
  NOR2_X1    g13498(.A1(new_n4243_), .A2(new_n14521_), .ZN(new_n14522_));
  NAND2_X1   g13499(.A1(new_n14522_), .A2(new_n4301_), .ZN(new_n14523_));
  NAND2_X1   g13500(.A1(new_n4289_), .A2(new_n4287_), .ZN(new_n14524_));
  NOR2_X1    g13501(.A1(new_n4289_), .A2(new_n4287_), .ZN(new_n14525_));
  NOR2_X1    g13502(.A1(new_n4250_), .A2(new_n14525_), .ZN(new_n14526_));
  NAND2_X1   g13503(.A1(new_n4323_), .A2(new_n14526_), .ZN(new_n14527_));
  AOI22_X1   g13504(.A1(new_n14527_), .A2(new_n14524_), .B1(new_n14523_), .B2(new_n14520_), .ZN(new_n14528_));
  OAI21_X1   g13505(.A1(new_n4284_), .A2(new_n4325_), .B(new_n14528_), .ZN(new_n14529_));
  NOR3_X1    g13506(.A1(new_n4284_), .A2(new_n14528_), .A3(new_n4325_), .ZN(new_n14530_));
  INV_X1     g13507(.I(new_n14530_), .ZN(new_n14531_));
  AOI21_X1   g13508(.A1(new_n14531_), .A2(new_n14529_), .B(new_n14519_), .ZN(new_n14532_));
  INV_X1     g13509(.I(new_n14529_), .ZN(new_n14533_));
  NOR3_X1    g13510(.A1(new_n14533_), .A2(new_n14518_), .A3(new_n14530_), .ZN(new_n14534_));
  NOR2_X1    g13511(.A1(new_n14534_), .A2(new_n14532_), .ZN(new_n14535_));
  NOR2_X1    g13512(.A1(new_n14535_), .A2(new_n14514_), .ZN(new_n14536_));
  AOI21_X1   g13513(.A1(new_n14512_), .A2(new_n14511_), .B(new_n14493_), .ZN(new_n14537_));
  NOR3_X1    g13514(.A1(new_n14507_), .A2(new_n14494_), .A3(new_n14509_), .ZN(new_n14538_));
  NOR2_X1    g13515(.A1(new_n14538_), .A2(new_n14537_), .ZN(new_n14539_));
  OAI21_X1   g13516(.A1(new_n14533_), .A2(new_n14530_), .B(new_n14518_), .ZN(new_n14540_));
  NAND3_X1   g13517(.A1(new_n14531_), .A2(new_n14529_), .A3(new_n14519_), .ZN(new_n14541_));
  NAND2_X1   g13518(.A1(new_n14540_), .A2(new_n14541_), .ZN(new_n14542_));
  NOR2_X1    g13519(.A1(new_n14542_), .A2(new_n14539_), .ZN(new_n14543_));
  OAI21_X1   g13520(.A1(new_n14543_), .A2(new_n14536_), .B(new_n14489_), .ZN(new_n14544_));
  AOI21_X1   g13521(.A1(new_n4281_), .A2(new_n4493_), .B(new_n4389_), .ZN(new_n14545_));
  NOR2_X1    g13522(.A1(new_n14535_), .A2(new_n14539_), .ZN(new_n14546_));
  NOR2_X1    g13523(.A1(new_n14542_), .A2(new_n14514_), .ZN(new_n14547_));
  OAI21_X1   g13524(.A1(new_n14546_), .A2(new_n14547_), .B(new_n14545_), .ZN(new_n14548_));
  NAND2_X1   g13525(.A1(new_n14544_), .A2(new_n14548_), .ZN(new_n14549_));
  NAND2_X1   g13526(.A1(new_n14488_), .A2(new_n14549_), .ZN(new_n14550_));
  NOR2_X1    g13527(.A1(new_n14478_), .A2(new_n14481_), .ZN(new_n14551_));
  NOR2_X1    g13528(.A1(new_n14446_), .A2(new_n14474_), .ZN(new_n14552_));
  OAI21_X1   g13529(.A1(new_n14551_), .A2(new_n14552_), .B(new_n14484_), .ZN(new_n14553_));
  NOR2_X1    g13530(.A1(new_n14446_), .A2(new_n14481_), .ZN(new_n14554_));
  NOR2_X1    g13531(.A1(new_n14478_), .A2(new_n14474_), .ZN(new_n14555_));
  OAI21_X1   g13532(.A1(new_n14554_), .A2(new_n14555_), .B(new_n14422_), .ZN(new_n14556_));
  NAND2_X1   g13533(.A1(new_n14553_), .A2(new_n14556_), .ZN(new_n14557_));
  NAND2_X1   g13534(.A1(new_n14542_), .A2(new_n14539_), .ZN(new_n14558_));
  NAND2_X1   g13535(.A1(new_n14535_), .A2(new_n14514_), .ZN(new_n14559_));
  AOI21_X1   g13536(.A1(new_n14558_), .A2(new_n14559_), .B(new_n14545_), .ZN(new_n14560_));
  NAND2_X1   g13537(.A1(new_n14542_), .A2(new_n14514_), .ZN(new_n14561_));
  NAND2_X1   g13538(.A1(new_n14535_), .A2(new_n14539_), .ZN(new_n14562_));
  AOI21_X1   g13539(.A1(new_n14562_), .A2(new_n14561_), .B(new_n14489_), .ZN(new_n14563_));
  NOR2_X1    g13540(.A1(new_n14560_), .A2(new_n14563_), .ZN(new_n14564_));
  NAND2_X1   g13541(.A1(new_n14557_), .A2(new_n14564_), .ZN(new_n14565_));
  AOI21_X1   g13542(.A1(new_n14565_), .A2(new_n14550_), .B(new_n14421_), .ZN(new_n14566_));
  OAI21_X1   g13543(.A1(new_n4506_), .A2(new_n4275_), .B(new_n4786_), .ZN(new_n14567_));
  OAI22_X1   g13544(.A1(new_n14483_), .A2(new_n14487_), .B1(new_n14560_), .B2(new_n14563_), .ZN(new_n14568_));
  NAND2_X1   g13545(.A1(new_n14488_), .A2(new_n14564_), .ZN(new_n14569_));
  AOI21_X1   g13546(.A1(new_n14569_), .A2(new_n14568_), .B(new_n14567_), .ZN(new_n14570_));
  NOR2_X1    g13547(.A1(new_n14566_), .A2(new_n14570_), .ZN(new_n14571_));
  NOR2_X1    g13548(.A1(new_n14571_), .A2(new_n14420_), .ZN(new_n14572_));
  NAND2_X1   g13549(.A1(new_n14412_), .A2(new_n14405_), .ZN(new_n14573_));
  NAND2_X1   g13550(.A1(new_n14397_), .A2(new_n14337_), .ZN(new_n14574_));
  AOI21_X1   g13551(.A1(new_n14573_), .A2(new_n14574_), .B(new_n14415_), .ZN(new_n14575_));
  AOI21_X1   g13552(.A1(new_n14416_), .A2(new_n14417_), .B(new_n14273_), .ZN(new_n14576_));
  NOR2_X1    g13553(.A1(new_n14575_), .A2(new_n14576_), .ZN(new_n14577_));
  NOR2_X1    g13554(.A1(new_n14557_), .A2(new_n14564_), .ZN(new_n14578_));
  NOR2_X1    g13555(.A1(new_n14488_), .A2(new_n14549_), .ZN(new_n14579_));
  OAI21_X1   g13556(.A1(new_n14578_), .A2(new_n14579_), .B(new_n14567_), .ZN(new_n14580_));
  NOR2_X1    g13557(.A1(new_n14488_), .A2(new_n14564_), .ZN(new_n14581_));
  NOR4_X1    g13558(.A1(new_n14483_), .A2(new_n14487_), .A3(new_n14560_), .A4(new_n14563_), .ZN(new_n14582_));
  OAI21_X1   g13559(.A1(new_n14581_), .A2(new_n14582_), .B(new_n14421_), .ZN(new_n14583_));
  NAND2_X1   g13560(.A1(new_n14580_), .A2(new_n14583_), .ZN(new_n14584_));
  NOR2_X1    g13561(.A1(new_n14584_), .A2(new_n14577_), .ZN(new_n14585_));
  OAI21_X1   g13562(.A1(new_n14572_), .A2(new_n14585_), .B(new_n14271_), .ZN(new_n14586_));
  AOI21_X1   g13563(.A1(new_n4272_), .A2(new_n4788_), .B(new_n13976_), .ZN(new_n14587_));
  NOR2_X1    g13564(.A1(new_n14571_), .A2(new_n14577_), .ZN(new_n14588_));
  NOR4_X1    g13565(.A1(new_n14566_), .A2(new_n14570_), .A3(new_n14575_), .A4(new_n14576_), .ZN(new_n14589_));
  OAI21_X1   g13566(.A1(new_n14588_), .A2(new_n14589_), .B(new_n14587_), .ZN(new_n14590_));
  NAND2_X1   g13567(.A1(new_n14586_), .A2(new_n14590_), .ZN(new_n14591_));
  AOI21_X1   g13568(.A1(new_n5347_), .A2(new_n5350_), .B(new_n5348_), .ZN(new_n14592_));
  NOR2_X1    g13569(.A1(new_n14591_), .A2(new_n14592_), .ZN(new_n14593_));
  INV_X1     g13570(.I(new_n14593_), .ZN(new_n14594_));
  NAND2_X1   g13571(.A1(new_n14591_), .A2(new_n14592_), .ZN(new_n14595_));
  AOI21_X1   g13572(.A1(new_n14594_), .A2(new_n14595_), .B(new_n14270_), .ZN(new_n14596_));
  INV_X1     g13573(.I(new_n14269_), .ZN(new_n14597_));
  NAND2_X1   g13574(.A1(new_n14597_), .A2(new_n14264_), .ZN(new_n14598_));
  INV_X1     g13575(.I(new_n14592_), .ZN(new_n14599_));
  NAND2_X1   g13576(.A1(new_n14599_), .A2(new_n14591_), .ZN(new_n14600_));
  NAND2_X1   g13577(.A1(new_n14584_), .A2(new_n14577_), .ZN(new_n14601_));
  NAND2_X1   g13578(.A1(new_n14571_), .A2(new_n14420_), .ZN(new_n14602_));
  AOI21_X1   g13579(.A1(new_n14602_), .A2(new_n14601_), .B(new_n14587_), .ZN(new_n14603_));
  OAI22_X1   g13580(.A1(new_n14566_), .A2(new_n14570_), .B1(new_n14575_), .B2(new_n14576_), .ZN(new_n14604_));
  NAND3_X1   g13581(.A1(new_n14577_), .A2(new_n14580_), .A3(new_n14583_), .ZN(new_n14605_));
  AOI21_X1   g13582(.A1(new_n14605_), .A2(new_n14604_), .B(new_n14271_), .ZN(new_n14606_));
  NOR2_X1    g13583(.A1(new_n14603_), .A2(new_n14606_), .ZN(new_n14607_));
  NAND2_X1   g13584(.A1(new_n14607_), .A2(new_n14592_), .ZN(new_n14608_));
  AOI21_X1   g13585(.A1(new_n14600_), .A2(new_n14608_), .B(new_n14598_), .ZN(new_n14609_));
  NOR2_X1    g13586(.A1(new_n14596_), .A2(new_n14609_), .ZN(new_n14610_));
  NOR3_X1    g13587(.A1(new_n13958_), .A2(new_n8198_), .A3(new_n13961_), .ZN(new_n14611_));
  AOI21_X1   g13588(.A1(new_n13965_), .A2(new_n13967_), .B(new_n14611_), .ZN(new_n14612_));
  INV_X1     g13589(.I(new_n14612_), .ZN(new_n14613_));
  AOI21_X1   g13590(.A1(new_n12558_), .A2(new_n13960_), .B(new_n13913_), .ZN(new_n14614_));
  OAI21_X1   g13591(.A1(new_n13213_), .A2(new_n13917_), .B(new_n13899_), .ZN(new_n14615_));
  OAI21_X1   g13592(.A1(new_n13877_), .A2(new_n13870_), .B(new_n13896_), .ZN(new_n14616_));
  NAND2_X1   g13593(.A1(new_n13855_), .A2(new_n13854_), .ZN(new_n14617_));
  NOR2_X1    g13594(.A1(new_n13745_), .A2(new_n13726_), .ZN(new_n14618_));
  NAND3_X1   g13595(.A1(new_n13740_), .A2(new_n13739_), .A3(new_n13734_), .ZN(new_n14619_));
  NOR4_X1    g13596(.A1(new_n14619_), .A2(new_n11156_), .A3(new_n14618_), .A4(new_n13729_), .ZN(new_n14620_));
  AOI22_X1   g13597(.A1(new_n11035_), .A2(new_n13737_), .B1(new_n11066_), .B2(new_n8794_), .ZN(new_n14621_));
  NAND4_X1   g13598(.A1(new_n11066_), .A2(new_n13737_), .A3(new_n11035_), .A4(new_n8794_), .ZN(new_n14622_));
  INV_X1     g13599(.I(new_n14622_), .ZN(new_n14623_));
  NOR4_X1    g13600(.A1(new_n14623_), .A2(new_n13731_), .A3(new_n13733_), .A4(new_n13732_), .ZN(new_n14624_));
  AOI21_X1   g13601(.A1(new_n14624_), .A2(new_n13740_), .B(new_n14621_), .ZN(new_n14625_));
  NAND2_X1   g13602(.A1(new_n13723_), .A2(new_n11123_), .ZN(new_n14626_));
  NOR2_X1    g13603(.A1(new_n14626_), .A2(new_n13725_), .ZN(new_n14627_));
  INV_X1     g13604(.I(new_n14627_), .ZN(new_n14628_));
  AOI21_X1   g13605(.A1(new_n13723_), .A2(new_n11123_), .B(new_n13744_), .ZN(new_n14629_));
  INV_X1     g13606(.I(new_n14629_), .ZN(new_n14630_));
  NAND3_X1   g13607(.A1(new_n11136_), .A2(new_n14630_), .A3(new_n13746_), .ZN(new_n14631_));
  AOI21_X1   g13608(.A1(new_n14628_), .A2(new_n14631_), .B(new_n14625_), .ZN(new_n14632_));
  OAI21_X1   g13609(.A1(new_n13757_), .A2(new_n13759_), .B(new_n14632_), .ZN(new_n14633_));
  NOR3_X1    g13610(.A1(new_n13749_), .A2(new_n11071_), .A3(new_n14623_), .ZN(new_n14634_));
  NOR4_X1    g13611(.A1(new_n13729_), .A2(new_n11125_), .A3(new_n14629_), .A4(new_n11127_), .ZN(new_n14635_));
  OAI22_X1   g13612(.A1(new_n14621_), .A2(new_n14634_), .B1(new_n14635_), .B2(new_n14627_), .ZN(new_n14636_));
  NAND4_X1   g13613(.A1(new_n13722_), .A2(new_n13838_), .A3(new_n14636_), .A4(new_n11157_), .ZN(new_n14637_));
  AOI21_X1   g13614(.A1(new_n14633_), .A2(new_n14637_), .B(new_n14620_), .ZN(new_n14638_));
  INV_X1     g13615(.I(new_n14620_), .ZN(new_n14639_));
  AOI21_X1   g13616(.A1(new_n13836_), .A2(new_n13838_), .B(new_n14636_), .ZN(new_n14640_));
  NOR4_X1    g13617(.A1(new_n13832_), .A2(new_n14632_), .A3(new_n13759_), .A4(new_n13830_), .ZN(new_n14641_));
  NOR3_X1    g13618(.A1(new_n14640_), .A2(new_n14641_), .A3(new_n14639_), .ZN(new_n14642_));
  NOR2_X1    g13619(.A1(new_n14642_), .A2(new_n14638_), .ZN(new_n14643_));
  XOR2_X1    g13620(.A1(new_n13795_), .A2(new_n13798_), .Z(new_n14644_));
  XOR2_X1    g13621(.A1(new_n13778_), .A2(new_n13781_), .Z(new_n14645_));
  NAND4_X1   g13622(.A1(new_n14644_), .A2(new_n14645_), .A3(new_n13765_), .A4(new_n13769_), .ZN(new_n14646_));
  NAND2_X1   g13623(.A1(new_n13786_), .A2(new_n11017_), .ZN(new_n14647_));
  INV_X1     g13624(.I(new_n14647_), .ZN(new_n14648_));
  NOR2_X1    g13625(.A1(new_n13802_), .A2(new_n10972_), .ZN(new_n14649_));
  NAND2_X1   g13626(.A1(new_n14648_), .A2(new_n14649_), .ZN(new_n14650_));
  NOR2_X1    g13627(.A1(new_n14648_), .A2(new_n13769_), .ZN(new_n14651_));
  NOR2_X1    g13628(.A1(new_n14649_), .A2(new_n13765_), .ZN(new_n14652_));
  NOR4_X1    g13629(.A1(new_n14651_), .A2(new_n14650_), .A3(new_n14646_), .A4(new_n14652_), .ZN(new_n14653_));
  INV_X1     g13630(.I(new_n14653_), .ZN(new_n14654_));
  NOR2_X1    g13631(.A1(new_n13795_), .A2(new_n13798_), .ZN(new_n14655_));
  NOR2_X1    g13632(.A1(new_n10981_), .A2(new_n14655_), .ZN(new_n14656_));
  AOI21_X1   g13633(.A1(new_n14649_), .A2(new_n14656_), .B(new_n13803_), .ZN(new_n14657_));
  INV_X1     g13634(.I(new_n14657_), .ZN(new_n14658_));
  NOR2_X1    g13635(.A1(new_n13778_), .A2(new_n13781_), .ZN(new_n14659_));
  NOR4_X1    g13636(.A1(new_n14659_), .A2(new_n11022_), .A3(new_n10993_), .A4(new_n11025_), .ZN(new_n14660_));
  INV_X1     g13637(.I(new_n14660_), .ZN(new_n14661_));
  OAI21_X1   g13638(.A1(new_n14661_), .A2(new_n14647_), .B(new_n13782_), .ZN(new_n14662_));
  NAND2_X1   g13639(.A1(new_n14658_), .A2(new_n14662_), .ZN(new_n14663_));
  AOI21_X1   g13640(.A1(new_n13827_), .A2(new_n13768_), .B(new_n14663_), .ZN(new_n14664_));
  AOI21_X1   g13641(.A1(new_n14648_), .A2(new_n14660_), .B(new_n13783_), .ZN(new_n14665_));
  NOR2_X1    g13642(.A1(new_n14665_), .A2(new_n14657_), .ZN(new_n14666_));
  NOR3_X1    g13643(.A1(new_n13846_), .A2(new_n13825_), .A3(new_n14666_), .ZN(new_n14667_));
  OAI21_X1   g13644(.A1(new_n14667_), .A2(new_n14664_), .B(new_n14654_), .ZN(new_n14668_));
  OAI21_X1   g13645(.A1(new_n13846_), .A2(new_n13825_), .B(new_n14666_), .ZN(new_n14669_));
  NAND3_X1   g13646(.A1(new_n13827_), .A2(new_n14663_), .A3(new_n13768_), .ZN(new_n14670_));
  NAND3_X1   g13647(.A1(new_n14669_), .A2(new_n14670_), .A3(new_n14653_), .ZN(new_n14671_));
  NAND2_X1   g13648(.A1(new_n14668_), .A2(new_n14671_), .ZN(new_n14672_));
  NAND2_X1   g13649(.A1(new_n14672_), .A2(new_n14643_), .ZN(new_n14673_));
  OAI21_X1   g13650(.A1(new_n14640_), .A2(new_n14641_), .B(new_n14639_), .ZN(new_n14674_));
  NAND3_X1   g13651(.A1(new_n14633_), .A2(new_n14637_), .A3(new_n14620_), .ZN(new_n14675_));
  NAND2_X1   g13652(.A1(new_n14674_), .A2(new_n14675_), .ZN(new_n14676_));
  NAND3_X1   g13653(.A1(new_n14676_), .A2(new_n14668_), .A3(new_n14671_), .ZN(new_n14677_));
  AOI22_X1   g13654(.A1(new_n14673_), .A2(new_n14677_), .B1(new_n14617_), .B2(new_n13856_), .ZN(new_n14678_));
  OAI21_X1   g13655(.A1(new_n13874_), .A2(new_n13719_), .B(new_n13856_), .ZN(new_n14679_));
  AOI21_X1   g13656(.A1(new_n14669_), .A2(new_n14670_), .B(new_n14653_), .ZN(new_n14680_));
  NOR3_X1    g13657(.A1(new_n14667_), .A2(new_n14664_), .A3(new_n14654_), .ZN(new_n14681_));
  OAI22_X1   g13658(.A1(new_n14681_), .A2(new_n14680_), .B1(new_n14638_), .B2(new_n14642_), .ZN(new_n14682_));
  NAND4_X1   g13659(.A1(new_n14668_), .A2(new_n14671_), .A3(new_n14674_), .A4(new_n14675_), .ZN(new_n14683_));
  AOI21_X1   g13660(.A1(new_n14682_), .A2(new_n14683_), .B(new_n14679_), .ZN(new_n14684_));
  NAND2_X1   g13661(.A1(new_n13863_), .A2(new_n13544_), .ZN(new_n14685_));
  XNOR2_X1   g13662(.A1(new_n13668_), .A2(new_n13670_), .ZN(new_n14686_));
  NOR2_X1    g13663(.A1(new_n13636_), .A2(new_n11204_), .ZN(new_n14687_));
  XOR2_X1    g13664(.A1(new_n14687_), .A2(new_n13652_), .Z(new_n14688_));
  NOR4_X1    g13665(.A1(new_n14688_), .A2(new_n11193_), .A3(new_n14686_), .A4(new_n11229_), .ZN(new_n14689_));
  NOR2_X1    g13666(.A1(new_n13667_), .A2(new_n13655_), .ZN(new_n14690_));
  NAND2_X1   g13667(.A1(new_n13655_), .A2(new_n11229_), .ZN(new_n14691_));
  NAND2_X1   g13668(.A1(new_n13667_), .A2(new_n11193_), .ZN(new_n14692_));
  NAND4_X1   g13669(.A1(new_n14689_), .A2(new_n14690_), .A3(new_n14691_), .A4(new_n14692_), .ZN(new_n14693_));
  NAND2_X1   g13670(.A1(new_n13670_), .A2(new_n13668_), .ZN(new_n14694_));
  NAND2_X1   g13671(.A1(new_n13666_), .A2(new_n14694_), .ZN(new_n14695_));
  OAI21_X1   g13672(.A1(new_n14695_), .A2(new_n13667_), .B(new_n13675_), .ZN(new_n14696_));
  INV_X1     g13673(.I(new_n13652_), .ZN(new_n14697_));
  NAND2_X1   g13674(.A1(new_n14687_), .A2(new_n14697_), .ZN(new_n14698_));
  NAND2_X1   g13675(.A1(new_n13638_), .A2(new_n14698_), .ZN(new_n14699_));
  OAI21_X1   g13676(.A1(new_n14699_), .A2(new_n13655_), .B(new_n13653_), .ZN(new_n14700_));
  NAND2_X1   g13677(.A1(new_n14696_), .A2(new_n14700_), .ZN(new_n14701_));
  AOI21_X1   g13678(.A1(new_n13709_), .A2(new_n13694_), .B(new_n14701_), .ZN(new_n14702_));
  INV_X1     g13679(.I(new_n13667_), .ZN(new_n14703_));
  AOI21_X1   g13680(.A1(new_n13668_), .A2(new_n13670_), .B(new_n11193_), .ZN(new_n14704_));
  AOI21_X1   g13681(.A1(new_n14704_), .A2(new_n14703_), .B(new_n13671_), .ZN(new_n14705_));
  INV_X1     g13682(.I(new_n13655_), .ZN(new_n14706_));
  AOI21_X1   g13683(.A1(new_n14687_), .A2(new_n14697_), .B(new_n11229_), .ZN(new_n14707_));
  AOI21_X1   g13684(.A1(new_n14707_), .A2(new_n14706_), .B(new_n13656_), .ZN(new_n14708_));
  NOR2_X1    g13685(.A1(new_n14705_), .A2(new_n14708_), .ZN(new_n14709_));
  NOR3_X1    g13686(.A1(new_n13696_), .A2(new_n13648_), .A3(new_n14709_), .ZN(new_n14710_));
  OAI21_X1   g13687(.A1(new_n14710_), .A2(new_n14702_), .B(new_n14693_), .ZN(new_n14711_));
  INV_X1     g13688(.I(new_n14693_), .ZN(new_n14712_));
  OAI21_X1   g13689(.A1(new_n13696_), .A2(new_n13648_), .B(new_n14709_), .ZN(new_n14713_));
  NAND3_X1   g13690(.A1(new_n13709_), .A2(new_n13694_), .A3(new_n14701_), .ZN(new_n14714_));
  NAND3_X1   g13691(.A1(new_n14713_), .A2(new_n14714_), .A3(new_n14712_), .ZN(new_n14715_));
  AOI21_X1   g13692(.A1(new_n13602_), .A2(new_n13598_), .B(new_n13599_), .ZN(new_n14716_));
  NOR3_X1    g13693(.A1(new_n13602_), .A2(new_n13599_), .A3(new_n13598_), .ZN(new_n14717_));
  AOI21_X1   g13694(.A1(new_n13594_), .A2(new_n13563_), .B(new_n13588_), .ZN(new_n14718_));
  NOR3_X1    g13695(.A1(new_n13594_), .A2(new_n13563_), .A3(new_n13588_), .ZN(new_n14719_));
  NAND4_X1   g13696(.A1(new_n14716_), .A2(new_n14717_), .A3(new_n14719_), .A4(new_n14718_), .ZN(new_n14720_));
  NOR2_X1    g13697(.A1(new_n13605_), .A2(new_n13587_), .ZN(new_n14721_));
  AOI21_X1   g13698(.A1(new_n11253_), .A2(new_n11254_), .B(new_n8457_), .ZN(new_n14722_));
  NOR3_X1    g13699(.A1(new_n11251_), .A2(new_n8413_), .A3(new_n11250_), .ZN(new_n14723_));
  NOR2_X1    g13700(.A1(new_n14723_), .A2(new_n14722_), .ZN(new_n14724_));
  AOI21_X1   g13701(.A1(new_n14724_), .A2(new_n11258_), .B(new_n11306_), .ZN(new_n14725_));
  NAND2_X1   g13702(.A1(new_n13605_), .A2(new_n13587_), .ZN(new_n14726_));
  NAND2_X1   g13703(.A1(new_n11271_), .A2(new_n14726_), .ZN(new_n14727_));
  NOR3_X1    g13704(.A1(new_n14727_), .A2(new_n11248_), .A3(new_n14725_), .ZN(new_n14728_));
  NAND2_X1   g13705(.A1(new_n13574_), .A2(new_n13572_), .ZN(new_n14729_));
  INV_X1     g13706(.I(new_n14729_), .ZN(new_n14730_));
  AOI21_X1   g13707(.A1(new_n11282_), .A2(new_n11285_), .B(new_n13545_), .ZN(new_n14731_));
  NAND4_X1   g13708(.A1(new_n13568_), .A2(new_n13571_), .A3(new_n8500_), .A4(new_n8526_), .ZN(new_n14732_));
  INV_X1     g13709(.I(new_n14732_), .ZN(new_n14733_));
  NOR4_X1    g13710(.A1(new_n13598_), .A2(new_n14731_), .A3(new_n13553_), .A4(new_n14733_), .ZN(new_n14734_));
  OAI22_X1   g13711(.A1(new_n14730_), .A2(new_n14734_), .B1(new_n14728_), .B2(new_n14721_), .ZN(new_n14735_));
  AOI21_X1   g13712(.A1(new_n13622_), .A2(new_n13702_), .B(new_n14735_), .ZN(new_n14736_));
  INV_X1     g13713(.I(new_n14721_), .ZN(new_n14737_));
  NAND4_X1   g13714(.A1(new_n13593_), .A2(new_n11264_), .A3(new_n11271_), .A4(new_n14726_), .ZN(new_n14738_));
  NAND4_X1   g13715(.A1(new_n13601_), .A2(new_n11292_), .A3(new_n13556_), .A4(new_n14732_), .ZN(new_n14739_));
  AOI22_X1   g13716(.A1(new_n14729_), .A2(new_n14739_), .B1(new_n14738_), .B2(new_n14737_), .ZN(new_n14740_));
  NOR3_X1    g13717(.A1(new_n13566_), .A2(new_n13625_), .A3(new_n14740_), .ZN(new_n14741_));
  OAI21_X1   g13718(.A1(new_n14736_), .A2(new_n14741_), .B(new_n14720_), .ZN(new_n14742_));
  AND4_X2    g13719(.A1(new_n14716_), .A2(new_n14717_), .A3(new_n14719_), .A4(new_n14718_), .Z(new_n14743_));
  OAI21_X1   g13720(.A1(new_n13566_), .A2(new_n13625_), .B(new_n14740_), .ZN(new_n14744_));
  NAND3_X1   g13721(.A1(new_n13622_), .A2(new_n13702_), .A3(new_n14735_), .ZN(new_n14745_));
  NAND3_X1   g13722(.A1(new_n14745_), .A2(new_n14744_), .A3(new_n14743_), .ZN(new_n14746_));
  NAND2_X1   g13723(.A1(new_n14742_), .A2(new_n14746_), .ZN(new_n14747_));
  NAND3_X1   g13724(.A1(new_n14747_), .A2(new_n14711_), .A3(new_n14715_), .ZN(new_n14748_));
  AOI21_X1   g13725(.A1(new_n14713_), .A2(new_n14714_), .B(new_n14712_), .ZN(new_n14749_));
  NOR3_X1    g13726(.A1(new_n14710_), .A2(new_n14702_), .A3(new_n14693_), .ZN(new_n14750_));
  AOI21_X1   g13727(.A1(new_n14745_), .A2(new_n14744_), .B(new_n14743_), .ZN(new_n14751_));
  NOR3_X1    g13728(.A1(new_n14736_), .A2(new_n14741_), .A3(new_n14720_), .ZN(new_n14752_));
  NOR2_X1    g13729(.A1(new_n14752_), .A2(new_n14751_), .ZN(new_n14753_));
  OAI21_X1   g13730(.A1(new_n14749_), .A2(new_n14750_), .B(new_n14753_), .ZN(new_n14754_));
  AOI22_X1   g13731(.A1(new_n14754_), .A2(new_n14748_), .B1(new_n14685_), .B2(new_n13864_), .ZN(new_n14755_));
  OAI21_X1   g13732(.A1(new_n13713_), .A2(new_n13714_), .B(new_n13864_), .ZN(new_n14756_));
  OAI22_X1   g13733(.A1(new_n14750_), .A2(new_n14749_), .B1(new_n14751_), .B2(new_n14752_), .ZN(new_n14757_));
  NAND3_X1   g13734(.A1(new_n14753_), .A2(new_n14711_), .A3(new_n14715_), .ZN(new_n14758_));
  AOI21_X1   g13735(.A1(new_n14757_), .A2(new_n14758_), .B(new_n14756_), .ZN(new_n14759_));
  NOR2_X1    g13736(.A1(new_n14759_), .A2(new_n14755_), .ZN(new_n14760_));
  NOR3_X1    g13737(.A1(new_n14760_), .A2(new_n14678_), .A3(new_n14684_), .ZN(new_n14761_));
  NOR2_X1    g13738(.A1(new_n14684_), .A2(new_n14678_), .ZN(new_n14762_));
  NOR2_X1    g13739(.A1(new_n13714_), .A2(new_n13713_), .ZN(new_n14763_));
  NOR3_X1    g13740(.A1(new_n14753_), .A2(new_n14750_), .A3(new_n14749_), .ZN(new_n14764_));
  AOI21_X1   g13741(.A1(new_n14711_), .A2(new_n14715_), .B(new_n14747_), .ZN(new_n14765_));
  OAI22_X1   g13742(.A1(new_n14764_), .A2(new_n14765_), .B1(new_n14763_), .B2(new_n13715_), .ZN(new_n14766_));
  AOI21_X1   g13743(.A1(new_n13544_), .A2(new_n13863_), .B(new_n13715_), .ZN(new_n14767_));
  NAND2_X1   g13744(.A1(new_n14757_), .A2(new_n14758_), .ZN(new_n14768_));
  NAND2_X1   g13745(.A1(new_n14768_), .A2(new_n14767_), .ZN(new_n14769_));
  NAND2_X1   g13746(.A1(new_n14769_), .A2(new_n14766_), .ZN(new_n14770_));
  NOR2_X1    g13747(.A1(new_n14762_), .A2(new_n14770_), .ZN(new_n14771_));
  OAI21_X1   g13748(.A1(new_n14771_), .A2(new_n14761_), .B(new_n14616_), .ZN(new_n14772_));
  AOI21_X1   g13749(.A1(new_n13539_), .A2(new_n13895_), .B(new_n13878_), .ZN(new_n14773_));
  AOI21_X1   g13750(.A1(new_n14668_), .A2(new_n14671_), .B(new_n14676_), .ZN(new_n14774_));
  NOR2_X1    g13751(.A1(new_n14672_), .A2(new_n14643_), .ZN(new_n14775_));
  OAI21_X1   g13752(.A1(new_n14774_), .A2(new_n14775_), .B(new_n14679_), .ZN(new_n14776_));
  AOI21_X1   g13753(.A1(new_n13855_), .A2(new_n13854_), .B(new_n13875_), .ZN(new_n14777_));
  NAND2_X1   g13754(.A1(new_n14682_), .A2(new_n14683_), .ZN(new_n14778_));
  NAND2_X1   g13755(.A1(new_n14778_), .A2(new_n14777_), .ZN(new_n14779_));
  AOI22_X1   g13756(.A1(new_n14776_), .A2(new_n14779_), .B1(new_n14769_), .B2(new_n14766_), .ZN(new_n14780_));
  NOR4_X1    g13757(.A1(new_n14684_), .A2(new_n14678_), .A3(new_n14755_), .A4(new_n14759_), .ZN(new_n14781_));
  OAI21_X1   g13758(.A1(new_n14780_), .A2(new_n14781_), .B(new_n14773_), .ZN(new_n14782_));
  NAND2_X1   g13759(.A1(new_n14772_), .A2(new_n14782_), .ZN(new_n14783_));
  NOR2_X1    g13760(.A1(new_n13504_), .A2(new_n13512_), .ZN(new_n14784_));
  OAI21_X1   g13761(.A1(new_n14784_), .A2(new_n13372_), .B(new_n13532_), .ZN(new_n14785_));
  OAI21_X1   g13762(.A1(new_n13524_), .A2(new_n13374_), .B(new_n13511_), .ZN(new_n14786_));
  NOR2_X1    g13763(.A1(new_n13382_), .A2(new_n13399_), .ZN(new_n14787_));
  NAND3_X1   g13764(.A1(new_n13393_), .A2(new_n13394_), .A3(new_n13388_), .ZN(new_n14788_));
  NOR4_X1    g13765(.A1(new_n14788_), .A2(new_n13378_), .A3(new_n14787_), .A4(new_n13385_), .ZN(new_n14789_));
  INV_X1     g13766(.I(new_n14789_), .ZN(new_n14790_));
  NAND2_X1   g13767(.A1(new_n13389_), .A2(new_n13392_), .ZN(new_n14791_));
  NAND4_X1   g13768(.A1(new_n11459_), .A2(new_n13391_), .A3(new_n11422_), .A4(new_n9115_), .ZN(new_n14792_));
  NAND4_X1   g13769(.A1(new_n11447_), .A2(new_n11460_), .A3(new_n11464_), .A4(new_n14792_), .ZN(new_n14793_));
  OAI21_X1   g13770(.A1(new_n13403_), .A2(new_n14793_), .B(new_n14791_), .ZN(new_n14794_));
  NOR3_X1    g13771(.A1(new_n13397_), .A2(new_n11528_), .A3(new_n13381_), .ZN(new_n14795_));
  AOI21_X1   g13772(.A1(new_n13379_), .A2(new_n11513_), .B(new_n13398_), .ZN(new_n14796_));
  NOR4_X1    g13773(.A1(new_n13385_), .A2(new_n11515_), .A3(new_n14796_), .A4(new_n11517_), .ZN(new_n14797_));
  OAI21_X1   g13774(.A1(new_n14795_), .A2(new_n14797_), .B(new_n14794_), .ZN(new_n14798_));
  AOI21_X1   g13775(.A1(new_n13491_), .A2(new_n13493_), .B(new_n14798_), .ZN(new_n14799_));
  INV_X1     g13776(.I(new_n14794_), .ZN(new_n14800_));
  NOR2_X1    g13777(.A1(new_n14797_), .A2(new_n14795_), .ZN(new_n14801_));
  NOR2_X1    g13778(.A1(new_n14801_), .A2(new_n14800_), .ZN(new_n14802_));
  NOR4_X1    g13779(.A1(new_n14802_), .A2(new_n13487_), .A3(new_n13486_), .A4(new_n13411_), .ZN(new_n14803_));
  OAI21_X1   g13780(.A1(new_n14799_), .A2(new_n14803_), .B(new_n14790_), .ZN(new_n14804_));
  OAI21_X1   g13781(.A1(new_n13409_), .A2(new_n13411_), .B(new_n14802_), .ZN(new_n14805_));
  NAND4_X1   g13782(.A1(new_n13377_), .A2(new_n13493_), .A3(new_n11552_), .A4(new_n14798_), .ZN(new_n14806_));
  NAND3_X1   g13783(.A1(new_n14805_), .A2(new_n14789_), .A3(new_n14806_), .ZN(new_n14807_));
  NAND2_X1   g13784(.A1(new_n14804_), .A2(new_n14807_), .ZN(new_n14808_));
  XOR2_X1    g13785(.A1(new_n13455_), .A2(new_n13452_), .Z(new_n14809_));
  XOR2_X1    g13786(.A1(new_n13430_), .A2(new_n13434_), .Z(new_n14810_));
  NAND4_X1   g13787(.A1(new_n14810_), .A2(new_n13462_), .A3(new_n14809_), .A4(new_n13422_), .ZN(new_n14811_));
  NOR2_X1    g13788(.A1(new_n13429_), .A2(new_n13425_), .ZN(new_n14812_));
  NOR2_X1    g13789(.A1(new_n13458_), .A2(new_n11359_), .ZN(new_n14813_));
  NAND2_X1   g13790(.A1(new_n14812_), .A2(new_n14813_), .ZN(new_n14814_));
  NOR2_X1    g13791(.A1(new_n14812_), .A2(new_n13422_), .ZN(new_n14815_));
  NOR2_X1    g13792(.A1(new_n14813_), .A2(new_n13462_), .ZN(new_n14816_));
  NOR4_X1    g13793(.A1(new_n14815_), .A2(new_n14814_), .A3(new_n14811_), .A4(new_n14816_), .ZN(new_n14817_));
  NOR2_X1    g13794(.A1(new_n13455_), .A2(new_n13452_), .ZN(new_n14818_));
  NOR2_X1    g13795(.A1(new_n11363_), .A2(new_n14818_), .ZN(new_n14819_));
  AOI21_X1   g13796(.A1(new_n14813_), .A2(new_n14819_), .B(new_n13459_), .ZN(new_n14820_));
  NOR2_X1    g13797(.A1(new_n13430_), .A2(new_n13434_), .ZN(new_n14821_));
  NOR4_X1    g13798(.A1(new_n14821_), .A2(new_n11408_), .A3(new_n11380_), .A4(new_n11412_), .ZN(new_n14822_));
  AOI21_X1   g13799(.A1(new_n14812_), .A2(new_n14822_), .B(new_n13436_), .ZN(new_n14823_));
  NOR2_X1    g13800(.A1(new_n14823_), .A2(new_n14820_), .ZN(new_n14824_));
  OAI21_X1   g13801(.A1(new_n13501_), .A2(new_n13481_), .B(new_n14824_), .ZN(new_n14825_));
  INV_X1     g13802(.I(new_n14820_), .ZN(new_n14826_));
  NAND2_X1   g13803(.A1(new_n13440_), .A2(new_n11404_), .ZN(new_n14827_));
  INV_X1     g13804(.I(new_n14822_), .ZN(new_n14828_));
  OAI21_X1   g13805(.A1(new_n14828_), .A2(new_n14827_), .B(new_n13435_), .ZN(new_n14829_));
  NAND2_X1   g13806(.A1(new_n14826_), .A2(new_n14829_), .ZN(new_n14830_));
  NAND3_X1   g13807(.A1(new_n13483_), .A2(new_n13421_), .A3(new_n14830_), .ZN(new_n14831_));
  AOI21_X1   g13808(.A1(new_n14825_), .A2(new_n14831_), .B(new_n14817_), .ZN(new_n14832_));
  INV_X1     g13809(.I(new_n14817_), .ZN(new_n14833_));
  AOI21_X1   g13810(.A1(new_n13483_), .A2(new_n13421_), .B(new_n14830_), .ZN(new_n14834_));
  NOR3_X1    g13811(.A1(new_n13501_), .A2(new_n13481_), .A3(new_n14824_), .ZN(new_n14835_));
  NOR3_X1    g13812(.A1(new_n14835_), .A2(new_n14834_), .A3(new_n14833_), .ZN(new_n14836_));
  NOR2_X1    g13813(.A1(new_n14836_), .A2(new_n14832_), .ZN(new_n14837_));
  NOR2_X1    g13814(.A1(new_n14837_), .A2(new_n14808_), .ZN(new_n14838_));
  AOI21_X1   g13815(.A1(new_n14805_), .A2(new_n14806_), .B(new_n14789_), .ZN(new_n14839_));
  NOR3_X1    g13816(.A1(new_n14799_), .A2(new_n14803_), .A3(new_n14790_), .ZN(new_n14840_));
  NOR2_X1    g13817(.A1(new_n14840_), .A2(new_n14839_), .ZN(new_n14841_));
  OAI21_X1   g13818(.A1(new_n14835_), .A2(new_n14834_), .B(new_n14833_), .ZN(new_n14842_));
  NAND3_X1   g13819(.A1(new_n14825_), .A2(new_n14831_), .A3(new_n14817_), .ZN(new_n14843_));
  NAND2_X1   g13820(.A1(new_n14842_), .A2(new_n14843_), .ZN(new_n14844_));
  NOR2_X1    g13821(.A1(new_n14844_), .A2(new_n14841_), .ZN(new_n14845_));
  OAI21_X1   g13822(.A1(new_n14838_), .A2(new_n14845_), .B(new_n14786_), .ZN(new_n14846_));
  AOI21_X1   g13823(.A1(new_n13509_), .A2(new_n13510_), .B(new_n13525_), .ZN(new_n14847_));
  OAI22_X1   g13824(.A1(new_n14836_), .A2(new_n14832_), .B1(new_n14840_), .B2(new_n14839_), .ZN(new_n14848_));
  NAND4_X1   g13825(.A1(new_n14842_), .A2(new_n14843_), .A3(new_n14804_), .A4(new_n14807_), .ZN(new_n14849_));
  NAND2_X1   g13826(.A1(new_n14848_), .A2(new_n14849_), .ZN(new_n14850_));
  NAND2_X1   g13827(.A1(new_n14850_), .A2(new_n14847_), .ZN(new_n14851_));
  OAI21_X1   g13828(.A1(new_n13217_), .A2(new_n13517_), .B(new_n13370_), .ZN(new_n14852_));
  AOI21_X1   g13829(.A1(new_n13329_), .A2(new_n13326_), .B(new_n13327_), .ZN(new_n14853_));
  NOR3_X1    g13830(.A1(new_n13329_), .A2(new_n13327_), .A3(new_n13326_), .ZN(new_n14854_));
  AOI21_X1   g13831(.A1(new_n13297_), .A2(new_n13321_), .B(new_n13320_), .ZN(new_n14855_));
  NOR3_X1    g13832(.A1(new_n13321_), .A2(new_n13320_), .A3(new_n13297_), .ZN(new_n14856_));
  NAND4_X1   g13833(.A1(new_n14853_), .A2(new_n14854_), .A3(new_n14855_), .A4(new_n14856_), .ZN(new_n14857_));
  NAND2_X1   g13834(.A1(new_n13333_), .A2(new_n13319_), .ZN(new_n14858_));
  INV_X1     g13835(.I(new_n14858_), .ZN(new_n14859_));
  NOR2_X1    g13836(.A1(new_n13333_), .A2(new_n13319_), .ZN(new_n14860_));
  NOR3_X1    g13837(.A1(new_n13321_), .A2(new_n13297_), .A3(new_n14860_), .ZN(new_n14861_));
  NAND2_X1   g13838(.A1(new_n13308_), .A2(new_n13306_), .ZN(new_n14862_));
  INV_X1     g13839(.I(new_n14862_), .ZN(new_n14863_));
  AOI21_X1   g13840(.A1(new_n13277_), .A2(new_n13280_), .B(new_n11593_), .ZN(new_n14864_));
  NAND4_X1   g13841(.A1(new_n13302_), .A2(new_n13305_), .A3(new_n9303_), .A4(new_n9330_), .ZN(new_n14865_));
  INV_X1     g13842(.I(new_n14865_), .ZN(new_n14866_));
  NOR4_X1    g13843(.A1(new_n14864_), .A2(new_n11611_), .A3(new_n13326_), .A4(new_n14866_), .ZN(new_n14867_));
  OAI22_X1   g13844(.A1(new_n14861_), .A2(new_n14859_), .B1(new_n14867_), .B2(new_n14863_), .ZN(new_n14868_));
  AOI21_X1   g13845(.A1(new_n13359_), .A2(new_n13342_), .B(new_n14868_), .ZN(new_n14869_));
  NAND2_X1   g13846(.A1(new_n11567_), .A2(new_n11557_), .ZN(new_n14870_));
  NOR2_X1    g13847(.A1(new_n13297_), .A2(new_n14860_), .ZN(new_n14871_));
  NAND3_X1   g13848(.A1(new_n14870_), .A2(new_n14871_), .A3(new_n11580_), .ZN(new_n14872_));
  NAND4_X1   g13849(.A1(new_n13328_), .A2(new_n13284_), .A3(new_n13290_), .A4(new_n14865_), .ZN(new_n14873_));
  AOI22_X1   g13850(.A1(new_n14872_), .A2(new_n14858_), .B1(new_n14873_), .B2(new_n14862_), .ZN(new_n14874_));
  NOR3_X1    g13851(.A1(new_n13300_), .A2(new_n13344_), .A3(new_n14874_), .ZN(new_n14875_));
  OAI21_X1   g13852(.A1(new_n14869_), .A2(new_n14875_), .B(new_n14857_), .ZN(new_n14876_));
  INV_X1     g13853(.I(new_n14857_), .ZN(new_n14877_));
  OAI21_X1   g13854(.A1(new_n13300_), .A2(new_n13344_), .B(new_n14874_), .ZN(new_n14878_));
  NAND3_X1   g13855(.A1(new_n13359_), .A2(new_n14868_), .A3(new_n13342_), .ZN(new_n14879_));
  NAND3_X1   g13856(.A1(new_n14879_), .A2(new_n14878_), .A3(new_n14877_), .ZN(new_n14880_));
  NAND2_X1   g13857(.A1(new_n14880_), .A2(new_n14876_), .ZN(new_n14881_));
  AOI21_X1   g13858(.A1(new_n13237_), .A2(new_n13221_), .B(new_n13235_), .ZN(new_n14882_));
  NOR3_X1    g13859(.A1(new_n13237_), .A2(new_n13235_), .A3(new_n13221_), .ZN(new_n14883_));
  AOI21_X1   g13860(.A1(new_n13261_), .A2(new_n11697_), .B(new_n13260_), .ZN(new_n14884_));
  NOR3_X1    g13861(.A1(new_n13261_), .A2(new_n13260_), .A3(new_n11697_), .ZN(new_n14885_));
  AND4_X2    g13862(.A1(new_n14882_), .A2(new_n14884_), .A3(new_n14883_), .A4(new_n14885_), .Z(new_n14886_));
  NOR2_X1    g13863(.A1(new_n13248_), .A2(new_n13242_), .ZN(new_n14887_));
  AOI21_X1   g13864(.A1(new_n11639_), .A2(new_n11640_), .B(new_n9431_), .ZN(new_n14888_));
  NOR3_X1    g13865(.A1(new_n11637_), .A2(new_n9386_), .A3(new_n11634_), .ZN(new_n14889_));
  NOR2_X1    g13866(.A1(new_n14889_), .A2(new_n14888_), .ZN(new_n14890_));
  AOI21_X1   g13867(.A1(new_n14890_), .A2(new_n11650_), .B(new_n11632_), .ZN(new_n14891_));
  NOR2_X1    g13868(.A1(new_n13247_), .A2(new_n13244_), .ZN(new_n14892_));
  NOR4_X1    g13869(.A1(new_n14891_), .A2(new_n11631_), .A3(new_n11697_), .A4(new_n14892_), .ZN(new_n14893_));
  NOR2_X1    g13870(.A1(new_n14893_), .A2(new_n14887_), .ZN(new_n14894_));
  AOI22_X1   g13871(.A1(new_n9475_), .A2(new_n13227_), .B1(new_n13231_), .B2(new_n9501_), .ZN(new_n14895_));
  NOR2_X1    g13872(.A1(new_n13228_), .A2(new_n13233_), .ZN(new_n14896_));
  NOR2_X1    g13873(.A1(new_n13221_), .A2(new_n14896_), .ZN(new_n14897_));
  AOI21_X1   g13874(.A1(new_n13258_), .A2(new_n14897_), .B(new_n14895_), .ZN(new_n14898_));
  NOR2_X1    g13875(.A1(new_n14894_), .A2(new_n14898_), .ZN(new_n14899_));
  OAI21_X1   g13876(.A1(new_n13268_), .A2(new_n13352_), .B(new_n14899_), .ZN(new_n14900_));
  NOR2_X1    g13877(.A1(new_n11702_), .A2(new_n11701_), .ZN(new_n14901_));
  AOI21_X1   g13878(.A1(new_n14901_), .A2(new_n11675_), .B(new_n11700_), .ZN(new_n14902_));
  NOR4_X1    g13879(.A1(new_n14902_), .A2(new_n11709_), .A3(new_n13221_), .A4(new_n14896_), .ZN(new_n14903_));
  OAI22_X1   g13880(.A1(new_n14903_), .A2(new_n14895_), .B1(new_n14893_), .B2(new_n14887_), .ZN(new_n14904_));
  NAND3_X1   g13881(.A1(new_n13270_), .A2(new_n13225_), .A3(new_n14904_), .ZN(new_n14905_));
  AOI21_X1   g13882(.A1(new_n14900_), .A2(new_n14905_), .B(new_n14886_), .ZN(new_n14906_));
  NAND4_X1   g13883(.A1(new_n14882_), .A2(new_n14883_), .A3(new_n14884_), .A4(new_n14885_), .ZN(new_n14907_));
  AOI21_X1   g13884(.A1(new_n13270_), .A2(new_n13225_), .B(new_n14904_), .ZN(new_n14908_));
  NOR3_X1    g13885(.A1(new_n14899_), .A2(new_n13268_), .A3(new_n13352_), .ZN(new_n14909_));
  NOR3_X1    g13886(.A1(new_n14909_), .A2(new_n14908_), .A3(new_n14907_), .ZN(new_n14910_));
  NOR2_X1    g13887(.A1(new_n14906_), .A2(new_n14910_), .ZN(new_n14911_));
  NOR2_X1    g13888(.A1(new_n14881_), .A2(new_n14911_), .ZN(new_n14912_));
  AOI21_X1   g13889(.A1(new_n14879_), .A2(new_n14878_), .B(new_n14877_), .ZN(new_n14913_));
  NOR3_X1    g13890(.A1(new_n14869_), .A2(new_n14875_), .A3(new_n14857_), .ZN(new_n14914_));
  NOR2_X1    g13891(.A1(new_n14913_), .A2(new_n14914_), .ZN(new_n14915_));
  OAI21_X1   g13892(.A1(new_n14909_), .A2(new_n14908_), .B(new_n14907_), .ZN(new_n14916_));
  NAND3_X1   g13893(.A1(new_n14900_), .A2(new_n14905_), .A3(new_n14886_), .ZN(new_n14917_));
  NAND2_X1   g13894(.A1(new_n14916_), .A2(new_n14917_), .ZN(new_n14918_));
  NOR2_X1    g13895(.A1(new_n14915_), .A2(new_n14918_), .ZN(new_n14919_));
  OAI21_X1   g13896(.A1(new_n14912_), .A2(new_n14919_), .B(new_n14852_), .ZN(new_n14920_));
  AOI21_X1   g13897(.A1(new_n13368_), .A2(new_n13369_), .B(new_n13518_), .ZN(new_n14921_));
  NOR2_X1    g13898(.A1(new_n14915_), .A2(new_n14911_), .ZN(new_n14922_));
  NOR4_X1    g13899(.A1(new_n14913_), .A2(new_n14914_), .A3(new_n14906_), .A4(new_n14910_), .ZN(new_n14923_));
  OAI21_X1   g13900(.A1(new_n14922_), .A2(new_n14923_), .B(new_n14921_), .ZN(new_n14924_));
  NAND2_X1   g13901(.A1(new_n14920_), .A2(new_n14924_), .ZN(new_n14925_));
  NAND3_X1   g13902(.A1(new_n14846_), .A2(new_n14925_), .A3(new_n14851_), .ZN(new_n14926_));
  NAND2_X1   g13903(.A1(new_n14844_), .A2(new_n14841_), .ZN(new_n14927_));
  NAND2_X1   g13904(.A1(new_n14837_), .A2(new_n14808_), .ZN(new_n14928_));
  AOI21_X1   g13905(.A1(new_n14927_), .A2(new_n14928_), .B(new_n14847_), .ZN(new_n14929_));
  AOI21_X1   g13906(.A1(new_n14848_), .A2(new_n14849_), .B(new_n14786_), .ZN(new_n14930_));
  NAND2_X1   g13907(.A1(new_n14915_), .A2(new_n14918_), .ZN(new_n14931_));
  NAND2_X1   g13908(.A1(new_n14881_), .A2(new_n14911_), .ZN(new_n14932_));
  AOI21_X1   g13909(.A1(new_n14932_), .A2(new_n14931_), .B(new_n14921_), .ZN(new_n14933_));
  NAND2_X1   g13910(.A1(new_n14881_), .A2(new_n14918_), .ZN(new_n14934_));
  NAND4_X1   g13911(.A1(new_n14876_), .A2(new_n14880_), .A3(new_n14916_), .A4(new_n14917_), .ZN(new_n14935_));
  AOI21_X1   g13912(.A1(new_n14934_), .A2(new_n14935_), .B(new_n14852_), .ZN(new_n14936_));
  NOR2_X1    g13913(.A1(new_n14933_), .A2(new_n14936_), .ZN(new_n14937_));
  OAI21_X1   g13914(.A1(new_n14929_), .A2(new_n14930_), .B(new_n14937_), .ZN(new_n14938_));
  AOI22_X1   g13915(.A1(new_n14938_), .A2(new_n14926_), .B1(new_n13534_), .B2(new_n14785_), .ZN(new_n14939_));
  OAI21_X1   g13916(.A1(new_n13885_), .A2(new_n13215_), .B(new_n13534_), .ZN(new_n14940_));
  OAI21_X1   g13917(.A1(new_n14929_), .A2(new_n14930_), .B(new_n14925_), .ZN(new_n14941_));
  NAND3_X1   g13918(.A1(new_n14846_), .A2(new_n14937_), .A3(new_n14851_), .ZN(new_n14942_));
  AOI21_X1   g13919(.A1(new_n14941_), .A2(new_n14942_), .B(new_n14940_), .ZN(new_n14943_));
  NOR2_X1    g13920(.A1(new_n14943_), .A2(new_n14939_), .ZN(new_n14944_));
  NOR2_X1    g13921(.A1(new_n14783_), .A2(new_n14944_), .ZN(new_n14945_));
  NAND3_X1   g13922(.A1(new_n14770_), .A2(new_n14776_), .A3(new_n14779_), .ZN(new_n14946_));
  NAND2_X1   g13923(.A1(new_n14776_), .A2(new_n14779_), .ZN(new_n14947_));
  NAND2_X1   g13924(.A1(new_n14947_), .A2(new_n14760_), .ZN(new_n14948_));
  AOI21_X1   g13925(.A1(new_n14948_), .A2(new_n14946_), .B(new_n14773_), .ZN(new_n14949_));
  OAI22_X1   g13926(.A1(new_n14684_), .A2(new_n14678_), .B1(new_n14755_), .B2(new_n14759_), .ZN(new_n14950_));
  NAND4_X1   g13927(.A1(new_n14776_), .A2(new_n14779_), .A3(new_n14769_), .A4(new_n14766_), .ZN(new_n14951_));
  AOI21_X1   g13928(.A1(new_n14950_), .A2(new_n14951_), .B(new_n14616_), .ZN(new_n14952_));
  NOR2_X1    g13929(.A1(new_n14949_), .A2(new_n14952_), .ZN(new_n14953_));
  NOR3_X1    g13930(.A1(new_n14929_), .A2(new_n14930_), .A3(new_n14937_), .ZN(new_n14954_));
  AOI21_X1   g13931(.A1(new_n14846_), .A2(new_n14851_), .B(new_n14925_), .ZN(new_n14955_));
  OAI21_X1   g13932(.A1(new_n14954_), .A2(new_n14955_), .B(new_n14940_), .ZN(new_n14956_));
  AOI21_X1   g13933(.A1(new_n13533_), .A2(new_n13532_), .B(new_n13886_), .ZN(new_n14957_));
  AOI21_X1   g13934(.A1(new_n14846_), .A2(new_n14851_), .B(new_n14937_), .ZN(new_n14958_));
  NOR3_X1    g13935(.A1(new_n14929_), .A2(new_n14930_), .A3(new_n14925_), .ZN(new_n14959_));
  OAI21_X1   g13936(.A1(new_n14958_), .A2(new_n14959_), .B(new_n14957_), .ZN(new_n14960_));
  NAND2_X1   g13937(.A1(new_n14960_), .A2(new_n14956_), .ZN(new_n14961_));
  NOR2_X1    g13938(.A1(new_n14953_), .A2(new_n14961_), .ZN(new_n14962_));
  OAI21_X1   g13939(.A1(new_n14945_), .A2(new_n14962_), .B(new_n14615_), .ZN(new_n14963_));
  AOI21_X1   g13940(.A1(new_n13891_), .A2(new_n13898_), .B(new_n13918_), .ZN(new_n14964_));
  AOI22_X1   g13941(.A1(new_n14772_), .A2(new_n14782_), .B1(new_n14960_), .B2(new_n14956_), .ZN(new_n14965_));
  NOR4_X1    g13942(.A1(new_n14949_), .A2(new_n14952_), .A3(new_n14943_), .A4(new_n14939_), .ZN(new_n14966_));
  OAI21_X1   g13943(.A1(new_n14965_), .A2(new_n14966_), .B(new_n14964_), .ZN(new_n14967_));
  OAI21_X1   g13944(.A1(new_n12559_), .A2(new_n13206_), .B(new_n13907_), .ZN(new_n14968_));
  AOI21_X1   g13945(.A1(new_n12885_), .A2(new_n13201_), .B(new_n13188_), .ZN(new_n14969_));
  OAI21_X1   g13946(.A1(new_n13165_), .A2(new_n13166_), .B(new_n13181_), .ZN(new_n14970_));
  NOR2_X1    g13947(.A1(new_n13043_), .A2(new_n13041_), .ZN(new_n14971_));
  OR3_X2     g13948(.A1(new_n13050_), .A2(new_n11872_), .A3(new_n13051_), .Z(new_n14972_));
  NOR4_X1    g13949(.A1(new_n14972_), .A2(new_n13054_), .A3(new_n14971_), .A4(new_n13057_), .ZN(new_n14973_));
  INV_X1     g13950(.I(new_n14973_), .ZN(new_n14974_));
  NAND4_X1   g13951(.A1(new_n11867_), .A2(new_n13048_), .A3(new_n11835_), .A4(new_n10152_), .ZN(new_n14975_));
  NAND4_X1   g13952(.A1(new_n11861_), .A2(new_n11868_), .A3(new_n11871_), .A4(new_n14975_), .ZN(new_n14976_));
  OAI22_X1   g13953(.A1(new_n13051_), .A2(new_n14976_), .B1(new_n13046_), .B2(new_n13062_), .ZN(new_n14977_));
  NOR3_X1    g13954(.A1(new_n13042_), .A2(new_n11921_), .A3(new_n13040_), .ZN(new_n14978_));
  AOI21_X1   g13955(.A1(new_n13037_), .A2(new_n11918_), .B(new_n13039_), .ZN(new_n14979_));
  NOR4_X1    g13956(.A1(new_n13057_), .A2(new_n11920_), .A3(new_n14979_), .A4(new_n11922_), .ZN(new_n14980_));
  OAI21_X1   g13957(.A1(new_n14978_), .A2(new_n14980_), .B(new_n14977_), .ZN(new_n14981_));
  AOI21_X1   g13958(.A1(new_n13071_), .A2(new_n13073_), .B(new_n14981_), .ZN(new_n14982_));
  INV_X1     g13959(.I(new_n14975_), .ZN(new_n14983_));
  NOR3_X1    g13960(.A1(new_n13059_), .A2(new_n11855_), .A3(new_n14983_), .ZN(new_n14984_));
  AOI22_X1   g13961(.A1(new_n14984_), .A2(new_n13065_), .B1(new_n13061_), .B2(new_n13049_), .ZN(new_n14985_));
  NOR2_X1    g13962(.A1(new_n14980_), .A2(new_n14978_), .ZN(new_n14986_));
  NOR2_X1    g13963(.A1(new_n14986_), .A2(new_n14985_), .ZN(new_n14987_));
  NOR4_X1    g13964(.A1(new_n13036_), .A2(new_n14987_), .A3(new_n13150_), .A4(new_n13033_), .ZN(new_n14988_));
  OAI21_X1   g13965(.A1(new_n14982_), .A2(new_n14988_), .B(new_n14974_), .ZN(new_n14989_));
  OAI21_X1   g13966(.A1(new_n13148_), .A2(new_n13150_), .B(new_n14987_), .ZN(new_n14990_));
  NAND4_X1   g13967(.A1(new_n13144_), .A2(new_n13073_), .A3(new_n14981_), .A4(new_n11957_), .ZN(new_n14991_));
  NAND3_X1   g13968(.A1(new_n14990_), .A2(new_n14991_), .A3(new_n14973_), .ZN(new_n14992_));
  NAND2_X1   g13969(.A1(new_n14989_), .A2(new_n14992_), .ZN(new_n14993_));
  NAND2_X1   g13970(.A1(new_n11771_), .A2(new_n11756_), .ZN(new_n14994_));
  NAND2_X1   g13971(.A1(new_n13116_), .A2(new_n11731_), .ZN(new_n14995_));
  XOR2_X1    g13972(.A1(new_n14995_), .A2(new_n14994_), .Z(new_n14996_));
  NAND2_X1   g13973(.A1(new_n11824_), .A2(new_n11778_), .ZN(new_n14997_));
  NAND2_X1   g13974(.A1(new_n13097_), .A2(new_n11809_), .ZN(new_n14998_));
  XOR2_X1    g13975(.A1(new_n14997_), .A2(new_n14998_), .Z(new_n14999_));
  NAND4_X1   g13976(.A1(new_n14999_), .A2(new_n14996_), .A3(new_n13113_), .A4(new_n13093_), .ZN(new_n15000_));
  NOR2_X1    g13977(.A1(new_n13101_), .A2(new_n13084_), .ZN(new_n15001_));
  NOR2_X1    g13978(.A1(new_n13114_), .A2(new_n11769_), .ZN(new_n15002_));
  NAND2_X1   g13979(.A1(new_n15001_), .A2(new_n15002_), .ZN(new_n15003_));
  NOR2_X1    g13980(.A1(new_n15001_), .A2(new_n13093_), .ZN(new_n15004_));
  NOR2_X1    g13981(.A1(new_n15002_), .A2(new_n13113_), .ZN(new_n15005_));
  NOR4_X1    g13982(.A1(new_n15003_), .A2(new_n15004_), .A3(new_n15005_), .A4(new_n15000_), .ZN(new_n15006_));
  NOR2_X1    g13983(.A1(new_n14995_), .A2(new_n14994_), .ZN(new_n15007_));
  NOR2_X1    g13984(.A1(new_n11773_), .A2(new_n15007_), .ZN(new_n15008_));
  AOI21_X1   g13985(.A1(new_n15002_), .A2(new_n15008_), .B(new_n13117_), .ZN(new_n15009_));
  NOR2_X1    g13986(.A1(new_n14997_), .A2(new_n14998_), .ZN(new_n15010_));
  NOR4_X1    g13987(.A1(new_n15010_), .A2(new_n11792_), .A3(new_n11821_), .A4(new_n11825_), .ZN(new_n15011_));
  AOI21_X1   g13988(.A1(new_n15001_), .A2(new_n15011_), .B(new_n13098_), .ZN(new_n15012_));
  NOR2_X1    g13989(.A1(new_n15012_), .A2(new_n15009_), .ZN(new_n15013_));
  OAI21_X1   g13990(.A1(new_n13141_), .A2(new_n13092_), .B(new_n15013_), .ZN(new_n15014_));
  INV_X1     g13991(.I(new_n15009_), .ZN(new_n15015_));
  NAND2_X1   g13992(.A1(new_n13095_), .A2(new_n11816_), .ZN(new_n15016_));
  INV_X1     g13993(.I(new_n15011_), .ZN(new_n15017_));
  OAI21_X1   g13994(.A1(new_n15017_), .A2(new_n15016_), .B(new_n13099_), .ZN(new_n15018_));
  NAND2_X1   g13995(.A1(new_n15015_), .A2(new_n15018_), .ZN(new_n15019_));
  NAND3_X1   g13996(.A1(new_n13158_), .A2(new_n15019_), .A3(new_n13139_), .ZN(new_n15020_));
  AOI21_X1   g13997(.A1(new_n15014_), .A2(new_n15020_), .B(new_n15006_), .ZN(new_n15021_));
  INV_X1     g13998(.I(new_n15006_), .ZN(new_n15022_));
  AOI21_X1   g13999(.A1(new_n13158_), .A2(new_n13139_), .B(new_n15019_), .ZN(new_n15023_));
  NOR3_X1    g14000(.A1(new_n13141_), .A2(new_n13092_), .A3(new_n15013_), .ZN(new_n15024_));
  NOR3_X1    g14001(.A1(new_n15024_), .A2(new_n15023_), .A3(new_n15022_), .ZN(new_n15025_));
  NOR2_X1    g14002(.A1(new_n15025_), .A2(new_n15021_), .ZN(new_n15026_));
  NOR2_X1    g14003(.A1(new_n15026_), .A2(new_n14993_), .ZN(new_n15027_));
  AOI21_X1   g14004(.A1(new_n14990_), .A2(new_n14991_), .B(new_n14973_), .ZN(new_n15028_));
  NOR3_X1    g14005(.A1(new_n14982_), .A2(new_n14988_), .A3(new_n14974_), .ZN(new_n15029_));
  NOR2_X1    g14006(.A1(new_n15029_), .A2(new_n15028_), .ZN(new_n15030_));
  OAI21_X1   g14007(.A1(new_n15024_), .A2(new_n15023_), .B(new_n15022_), .ZN(new_n15031_));
  NAND3_X1   g14008(.A1(new_n15014_), .A2(new_n15020_), .A3(new_n15006_), .ZN(new_n15032_));
  NAND2_X1   g14009(.A1(new_n15031_), .A2(new_n15032_), .ZN(new_n15033_));
  NOR2_X1    g14010(.A1(new_n15033_), .A2(new_n15030_), .ZN(new_n15034_));
  OAI21_X1   g14011(.A1(new_n15027_), .A2(new_n15034_), .B(new_n14970_), .ZN(new_n15035_));
  AOI21_X1   g14012(.A1(new_n13180_), .A2(new_n13032_), .B(new_n13167_), .ZN(new_n15036_));
  OAI22_X1   g14013(.A1(new_n15025_), .A2(new_n15021_), .B1(new_n15029_), .B2(new_n15028_), .ZN(new_n15037_));
  NAND4_X1   g14014(.A1(new_n15031_), .A2(new_n15032_), .A3(new_n14989_), .A4(new_n14992_), .ZN(new_n15038_));
  NAND2_X1   g14015(.A1(new_n15037_), .A2(new_n15038_), .ZN(new_n15039_));
  NAND2_X1   g14016(.A1(new_n15039_), .A2(new_n15036_), .ZN(new_n15040_));
  NAND2_X1   g14017(.A1(new_n13001_), .A2(new_n13006_), .ZN(new_n15041_));
  AOI21_X1   g14018(.A1(new_n15041_), .A2(new_n12940_), .B(new_n13023_), .ZN(new_n15042_));
  XNOR2_X1   g14019(.A1(new_n12981_), .A2(new_n12979_), .ZN(new_n15043_));
  XNOR2_X1   g14020(.A1(new_n12959_), .A2(new_n12961_), .ZN(new_n15044_));
  NOR4_X1    g14021(.A1(new_n15044_), .A2(new_n12988_), .A3(new_n15043_), .A4(new_n12031_), .ZN(new_n15045_));
  NOR2_X1    g14022(.A1(new_n12978_), .A2(new_n12964_), .ZN(new_n15046_));
  AOI22_X1   g14023(.A1(new_n12988_), .A2(new_n12978_), .B1(new_n12031_), .B2(new_n12964_), .ZN(new_n15047_));
  NAND3_X1   g14024(.A1(new_n15045_), .A2(new_n15047_), .A3(new_n15046_), .ZN(new_n15048_));
  INV_X1     g14025(.I(new_n15048_), .ZN(new_n15049_));
  INV_X1     g14026(.I(new_n12978_), .ZN(new_n15050_));
  AOI21_X1   g14027(.A1(new_n12979_), .A2(new_n12981_), .B(new_n12988_), .ZN(new_n15051_));
  AOI21_X1   g14028(.A1(new_n15051_), .A2(new_n15050_), .B(new_n12982_), .ZN(new_n15052_));
  NOR2_X1    g14029(.A1(new_n12959_), .A2(new_n12961_), .ZN(new_n15053_));
  NOR2_X1    g14030(.A1(new_n12031_), .A2(new_n15053_), .ZN(new_n15054_));
  AOI21_X1   g14031(.A1(new_n15054_), .A2(new_n12958_), .B(new_n12965_), .ZN(new_n15055_));
  NOR2_X1    g14032(.A1(new_n15052_), .A2(new_n15055_), .ZN(new_n15056_));
  OAI21_X1   g14033(.A1(new_n13005_), .A2(new_n12957_), .B(new_n15056_), .ZN(new_n15057_));
  NAND2_X1   g14034(.A1(new_n12981_), .A2(new_n12979_), .ZN(new_n15058_));
  NAND2_X1   g14035(.A1(new_n12977_), .A2(new_n15058_), .ZN(new_n15059_));
  OAI21_X1   g14036(.A1(new_n15059_), .A2(new_n12978_), .B(new_n12985_), .ZN(new_n15060_));
  INV_X1     g14037(.I(new_n15053_), .ZN(new_n15061_));
  NAND3_X1   g14038(.A1(new_n12949_), .A2(new_n12958_), .A3(new_n15061_), .ZN(new_n15062_));
  NAND2_X1   g14039(.A1(new_n15062_), .A2(new_n12962_), .ZN(new_n15063_));
  NAND2_X1   g14040(.A1(new_n15060_), .A2(new_n15063_), .ZN(new_n15064_));
  NAND3_X1   g14041(.A1(new_n13019_), .A2(new_n13003_), .A3(new_n15064_), .ZN(new_n15065_));
  AOI21_X1   g14042(.A1(new_n15057_), .A2(new_n15065_), .B(new_n15049_), .ZN(new_n15066_));
  AOI21_X1   g14043(.A1(new_n13019_), .A2(new_n13003_), .B(new_n15064_), .ZN(new_n15067_));
  NOR3_X1    g14044(.A1(new_n13005_), .A2(new_n12957_), .A3(new_n15056_), .ZN(new_n15068_));
  NOR3_X1    g14045(.A1(new_n15068_), .A2(new_n15067_), .A3(new_n15048_), .ZN(new_n15069_));
  OAI21_X1   g14046(.A1(new_n12905_), .A2(new_n12897_), .B(new_n12903_), .ZN(new_n15070_));
  NAND3_X1   g14047(.A1(new_n12905_), .A2(new_n12903_), .A3(new_n12897_), .ZN(new_n15071_));
  OAI21_X1   g14048(.A1(new_n12929_), .A2(new_n12101_), .B(new_n12928_), .ZN(new_n15072_));
  NAND3_X1   g14049(.A1(new_n12929_), .A2(new_n12928_), .A3(new_n12101_), .ZN(new_n15073_));
  NOR4_X1    g14050(.A1(new_n15070_), .A2(new_n15071_), .A3(new_n15072_), .A4(new_n15073_), .ZN(new_n15074_));
  AOI21_X1   g14051(.A1(new_n9792_), .A2(new_n12912_), .B(new_n12909_), .ZN(new_n15075_));
  NOR2_X1    g14052(.A1(new_n12913_), .A2(new_n12916_), .ZN(new_n15076_));
  NOR2_X1    g14053(.A1(new_n12144_), .A2(new_n15076_), .ZN(new_n15077_));
  AOI21_X1   g14054(.A1(new_n12929_), .A2(new_n15077_), .B(new_n15075_), .ZN(new_n15078_));
  AND2_X2    g14055(.A1(new_n12900_), .A2(new_n12902_), .Z(new_n15079_));
  NOR2_X1    g14056(.A1(new_n12900_), .A2(new_n12902_), .ZN(new_n15080_));
  NOR2_X1    g14057(.A1(new_n12923_), .A2(new_n15080_), .ZN(new_n15081_));
  AOI21_X1   g14058(.A1(new_n12905_), .A2(new_n15081_), .B(new_n15079_), .ZN(new_n15082_));
  NOR2_X1    g14059(.A1(new_n15082_), .A2(new_n15078_), .ZN(new_n15083_));
  OAI21_X1   g14060(.A1(new_n12893_), .A2(new_n12938_), .B(new_n15083_), .ZN(new_n15084_));
  NOR2_X1    g14061(.A1(new_n12135_), .A2(new_n12134_), .ZN(new_n15085_));
  AOI21_X1   g14062(.A1(new_n15085_), .A2(new_n12088_), .B(new_n12064_), .ZN(new_n15086_));
  NOR4_X1    g14063(.A1(new_n15086_), .A2(new_n12063_), .A3(new_n12144_), .A4(new_n15076_), .ZN(new_n15087_));
  AOI21_X1   g14064(.A1(new_n12113_), .A2(new_n12116_), .B(new_n12148_), .ZN(new_n15088_));
  NOR4_X1    g14065(.A1(new_n15088_), .A2(new_n12159_), .A3(new_n12923_), .A4(new_n15080_), .ZN(new_n15089_));
  OAI22_X1   g14066(.A1(new_n15087_), .A2(new_n15075_), .B1(new_n15089_), .B2(new_n15079_), .ZN(new_n15090_));
  NAND3_X1   g14067(.A1(new_n13012_), .A2(new_n12936_), .A3(new_n15090_), .ZN(new_n15091_));
  AOI21_X1   g14068(.A1(new_n15091_), .A2(new_n15084_), .B(new_n15074_), .ZN(new_n15092_));
  INV_X1     g14069(.I(new_n15074_), .ZN(new_n15093_));
  AOI21_X1   g14070(.A1(new_n13012_), .A2(new_n12936_), .B(new_n15090_), .ZN(new_n15094_));
  NOR3_X1    g14071(.A1(new_n12893_), .A2(new_n12938_), .A3(new_n15083_), .ZN(new_n15095_));
  NOR3_X1    g14072(.A1(new_n15094_), .A2(new_n15095_), .A3(new_n15093_), .ZN(new_n15096_));
  NOR2_X1    g14073(.A1(new_n15096_), .A2(new_n15092_), .ZN(new_n15097_));
  NOR3_X1    g14074(.A1(new_n15097_), .A2(new_n15066_), .A3(new_n15069_), .ZN(new_n15098_));
  OAI21_X1   g14075(.A1(new_n15068_), .A2(new_n15067_), .B(new_n15048_), .ZN(new_n15099_));
  NAND3_X1   g14076(.A1(new_n15057_), .A2(new_n15065_), .A3(new_n15049_), .ZN(new_n15100_));
  OAI21_X1   g14077(.A1(new_n15094_), .A2(new_n15095_), .B(new_n15093_), .ZN(new_n15101_));
  NAND3_X1   g14078(.A1(new_n15091_), .A2(new_n15084_), .A3(new_n15074_), .ZN(new_n15102_));
  NAND2_X1   g14079(.A1(new_n15101_), .A2(new_n15102_), .ZN(new_n15103_));
  AOI21_X1   g14080(.A1(new_n15099_), .A2(new_n15100_), .B(new_n15103_), .ZN(new_n15104_));
  OAI22_X1   g14081(.A1(new_n15104_), .A2(new_n15098_), .B1(new_n15042_), .B2(new_n13025_), .ZN(new_n15105_));
  AOI21_X1   g14082(.A1(new_n12889_), .A2(new_n13173_), .B(new_n13025_), .ZN(new_n15106_));
  OAI22_X1   g14083(.A1(new_n15069_), .A2(new_n15066_), .B1(new_n15092_), .B2(new_n15096_), .ZN(new_n15107_));
  NAND4_X1   g14084(.A1(new_n15099_), .A2(new_n15100_), .A3(new_n15101_), .A4(new_n15102_), .ZN(new_n15108_));
  NAND2_X1   g14085(.A1(new_n15107_), .A2(new_n15108_), .ZN(new_n15109_));
  NAND2_X1   g14086(.A1(new_n15109_), .A2(new_n15106_), .ZN(new_n15110_));
  NAND2_X1   g14087(.A1(new_n15110_), .A2(new_n15105_), .ZN(new_n15111_));
  NAND3_X1   g14088(.A1(new_n15111_), .A2(new_n15035_), .A3(new_n15040_), .ZN(new_n15112_));
  NAND2_X1   g14089(.A1(new_n15033_), .A2(new_n15030_), .ZN(new_n15113_));
  NAND2_X1   g14090(.A1(new_n15026_), .A2(new_n14993_), .ZN(new_n15114_));
  AOI21_X1   g14091(.A1(new_n15113_), .A2(new_n15114_), .B(new_n15036_), .ZN(new_n15115_));
  AOI21_X1   g14092(.A1(new_n15037_), .A2(new_n15038_), .B(new_n14970_), .ZN(new_n15116_));
  NAND2_X1   g14093(.A1(new_n13173_), .A2(new_n12889_), .ZN(new_n15117_));
  NAND3_X1   g14094(.A1(new_n15103_), .A2(new_n15099_), .A3(new_n15100_), .ZN(new_n15118_));
  OAI21_X1   g14095(.A1(new_n15066_), .A2(new_n15069_), .B(new_n15097_), .ZN(new_n15119_));
  AOI22_X1   g14096(.A1(new_n15119_), .A2(new_n15118_), .B1(new_n15117_), .B2(new_n13174_), .ZN(new_n15120_));
  OAI21_X1   g14097(.A1(new_n13024_), .A2(new_n13023_), .B(new_n13174_), .ZN(new_n15121_));
  AOI21_X1   g14098(.A1(new_n15107_), .A2(new_n15108_), .B(new_n15121_), .ZN(new_n15122_));
  NOR2_X1    g14099(.A1(new_n15122_), .A2(new_n15120_), .ZN(new_n15123_));
  OAI21_X1   g14100(.A1(new_n15115_), .A2(new_n15116_), .B(new_n15123_), .ZN(new_n15124_));
  AOI21_X1   g14101(.A1(new_n15124_), .A2(new_n15112_), .B(new_n14969_), .ZN(new_n15125_));
  OAI21_X1   g14102(.A1(new_n13187_), .A2(new_n13186_), .B(new_n13202_), .ZN(new_n15126_));
  OAI22_X1   g14103(.A1(new_n15116_), .A2(new_n15115_), .B1(new_n15120_), .B2(new_n15122_), .ZN(new_n15127_));
  NAND4_X1   g14104(.A1(new_n15035_), .A2(new_n15040_), .A3(new_n15105_), .A4(new_n15110_), .ZN(new_n15128_));
  AOI21_X1   g14105(.A1(new_n15127_), .A2(new_n15128_), .B(new_n15126_), .ZN(new_n15129_));
  AOI21_X1   g14106(.A1(new_n12563_), .A2(new_n13194_), .B(new_n12880_), .ZN(new_n15130_));
  AOI21_X1   g14107(.A1(new_n12856_), .A2(new_n12857_), .B(new_n12873_), .ZN(new_n15131_));
  AOI21_X1   g14108(.A1(new_n12809_), .A2(new_n12774_), .B(new_n12808_), .ZN(new_n15132_));
  INV_X1     g14109(.I(new_n15132_), .ZN(new_n15133_));
  NOR3_X1    g14110(.A1(new_n12809_), .A2(new_n12774_), .A3(new_n12808_), .ZN(new_n15134_));
  NAND4_X1   g14111(.A1(new_n15134_), .A2(new_n12781_), .A3(new_n12789_), .A4(new_n12796_), .ZN(new_n15135_));
  NOR2_X1    g14112(.A1(new_n15135_), .A2(new_n15133_), .ZN(new_n15136_));
  NOR2_X1    g14113(.A1(new_n12803_), .A2(new_n12806_), .ZN(new_n15137_));
  NOR2_X1    g14114(.A1(new_n12800_), .A2(new_n12802_), .ZN(new_n15138_));
  NOR2_X1    g14115(.A1(new_n12774_), .A2(new_n15138_), .ZN(new_n15139_));
  AOI21_X1   g14116(.A1(new_n12822_), .A2(new_n15139_), .B(new_n15137_), .ZN(new_n15140_));
  AOI21_X1   g14117(.A1(new_n10334_), .A2(new_n12787_), .B(new_n12816_), .ZN(new_n15141_));
  NOR2_X1    g14118(.A1(new_n12784_), .A2(new_n12788_), .ZN(new_n15142_));
  NOR2_X1    g14119(.A1(new_n12814_), .A2(new_n15142_), .ZN(new_n15143_));
  AOI21_X1   g14120(.A1(new_n12796_), .A2(new_n15143_), .B(new_n15141_), .ZN(new_n15144_));
  NOR2_X1    g14121(.A1(new_n15140_), .A2(new_n15144_), .ZN(new_n15145_));
  OAI21_X1   g14122(.A1(new_n12777_), .A2(new_n12832_), .B(new_n15145_), .ZN(new_n15146_));
  NOR3_X1    g14123(.A1(new_n12809_), .A2(new_n12774_), .A3(new_n15138_), .ZN(new_n15147_));
  NOR2_X1    g14124(.A1(new_n12235_), .A2(new_n12232_), .ZN(new_n15148_));
  AOI21_X1   g14125(.A1(new_n15148_), .A2(new_n12794_), .B(new_n12228_), .ZN(new_n15149_));
  NOR4_X1    g14126(.A1(new_n15149_), .A2(new_n12765_), .A3(new_n12814_), .A4(new_n15142_), .ZN(new_n15150_));
  OAI22_X1   g14127(.A1(new_n15147_), .A2(new_n15137_), .B1(new_n15150_), .B2(new_n15141_), .ZN(new_n15151_));
  NAND3_X1   g14128(.A1(new_n15151_), .A2(new_n12847_), .A3(new_n12830_), .ZN(new_n15152_));
  AOI21_X1   g14129(.A1(new_n15146_), .A2(new_n15152_), .B(new_n15136_), .ZN(new_n15153_));
  NAND3_X1   g14130(.A1(new_n12822_), .A2(new_n12820_), .A3(new_n12821_), .ZN(new_n15154_));
  NOR4_X1    g14131(.A1(new_n15154_), .A2(new_n12814_), .A3(new_n12817_), .A4(new_n12818_), .ZN(new_n15155_));
  NAND2_X1   g14132(.A1(new_n15155_), .A2(new_n15132_), .ZN(new_n15156_));
  AOI21_X1   g14133(.A1(new_n12830_), .A2(new_n12847_), .B(new_n15151_), .ZN(new_n15157_));
  NOR3_X1    g14134(.A1(new_n12777_), .A2(new_n12832_), .A3(new_n15145_), .ZN(new_n15158_));
  NOR3_X1    g14135(.A1(new_n15157_), .A2(new_n15158_), .A3(new_n15156_), .ZN(new_n15159_));
  NOR2_X1    g14136(.A1(new_n15159_), .A2(new_n15153_), .ZN(new_n15160_));
  AOI21_X1   g14137(.A1(new_n12750_), .A2(new_n12332_), .B(new_n12749_), .ZN(new_n15161_));
  NAND3_X1   g14138(.A1(new_n12739_), .A2(new_n12738_), .A3(new_n12732_), .ZN(new_n15162_));
  NOR4_X1    g14139(.A1(new_n15162_), .A2(new_n12720_), .A3(new_n12727_), .A4(new_n12730_), .ZN(new_n15163_));
  NAND2_X1   g14140(.A1(new_n15163_), .A2(new_n15161_), .ZN(new_n15164_));
  NAND2_X1   g14141(.A1(new_n12735_), .A2(new_n12737_), .ZN(new_n15165_));
  INV_X1     g14142(.I(new_n15165_), .ZN(new_n15166_));
  AOI21_X1   g14143(.A1(new_n12273_), .A2(new_n12274_), .B(new_n10453_), .ZN(new_n15167_));
  NOR3_X1    g14144(.A1(new_n12271_), .A2(new_n12268_), .A3(new_n10408_), .ZN(new_n15168_));
  NOR2_X1    g14145(.A1(new_n15168_), .A2(new_n15167_), .ZN(new_n15169_));
  AOI21_X1   g14146(.A1(new_n15169_), .A2(new_n12278_), .B(new_n12267_), .ZN(new_n15170_));
  NOR2_X1    g14147(.A1(new_n12735_), .A2(new_n12737_), .ZN(new_n15171_));
  NOR4_X1    g14148(.A1(new_n15170_), .A2(new_n12266_), .A3(new_n12332_), .A4(new_n15171_), .ZN(new_n15172_));
  NAND2_X1   g14149(.A1(new_n12726_), .A2(new_n12723_), .ZN(new_n15173_));
  INV_X1     g14150(.I(new_n15173_), .ZN(new_n15174_));
  NOR2_X1    g14151(.A1(new_n12337_), .A2(new_n12336_), .ZN(new_n15175_));
  AOI21_X1   g14152(.A1(new_n15175_), .A2(new_n12310_), .B(new_n12335_), .ZN(new_n15176_));
  NOR2_X1    g14153(.A1(new_n12726_), .A2(new_n12723_), .ZN(new_n15177_));
  NOR4_X1    g14154(.A1(new_n15176_), .A2(new_n12344_), .A3(new_n12720_), .A4(new_n15177_), .ZN(new_n15178_));
  OAI22_X1   g14155(.A1(new_n15178_), .A2(new_n15174_), .B1(new_n15172_), .B2(new_n15166_), .ZN(new_n15179_));
  AOI21_X1   g14156(.A1(new_n12759_), .A2(new_n12718_), .B(new_n15179_), .ZN(new_n15180_));
  NOR2_X1    g14157(.A1(new_n12332_), .A2(new_n15171_), .ZN(new_n15181_));
  NAND2_X1   g14158(.A1(new_n12739_), .A2(new_n15181_), .ZN(new_n15182_));
  NOR2_X1    g14159(.A1(new_n12720_), .A2(new_n15177_), .ZN(new_n15183_));
  NAND2_X1   g14160(.A1(new_n12745_), .A2(new_n15183_), .ZN(new_n15184_));
  AOI22_X1   g14161(.A1(new_n15165_), .A2(new_n15182_), .B1(new_n15184_), .B2(new_n15173_), .ZN(new_n15185_));
  NOR3_X1    g14162(.A1(new_n15185_), .A2(new_n12757_), .A3(new_n12840_), .ZN(new_n15186_));
  OAI21_X1   g14163(.A1(new_n15186_), .A2(new_n15180_), .B(new_n15164_), .ZN(new_n15187_));
  INV_X1     g14164(.I(new_n15161_), .ZN(new_n15188_));
  NOR3_X1    g14165(.A1(new_n12750_), .A2(new_n12749_), .A3(new_n12332_), .ZN(new_n15189_));
  NAND4_X1   g14166(.A1(new_n15189_), .A2(new_n12742_), .A3(new_n12743_), .A4(new_n12745_), .ZN(new_n15190_));
  NOR2_X1    g14167(.A1(new_n15190_), .A2(new_n15188_), .ZN(new_n15191_));
  OAI21_X1   g14168(.A1(new_n12757_), .A2(new_n12840_), .B(new_n15185_), .ZN(new_n15192_));
  NAND3_X1   g14169(.A1(new_n12759_), .A2(new_n12718_), .A3(new_n15179_), .ZN(new_n15193_));
  NAND3_X1   g14170(.A1(new_n15192_), .A2(new_n15193_), .A3(new_n15191_), .ZN(new_n15194_));
  NAND2_X1   g14171(.A1(new_n15194_), .A2(new_n15187_), .ZN(new_n15195_));
  NAND2_X1   g14172(.A1(new_n15160_), .A2(new_n15195_), .ZN(new_n15196_));
  OAI21_X1   g14173(.A1(new_n15157_), .A2(new_n15158_), .B(new_n15156_), .ZN(new_n15197_));
  NAND3_X1   g14174(.A1(new_n15146_), .A2(new_n15152_), .A3(new_n15136_), .ZN(new_n15198_));
  NAND2_X1   g14175(.A1(new_n15197_), .A2(new_n15198_), .ZN(new_n15199_));
  AOI21_X1   g14176(.A1(new_n15192_), .A2(new_n15193_), .B(new_n15191_), .ZN(new_n15200_));
  NOR3_X1    g14177(.A1(new_n15186_), .A2(new_n15180_), .A3(new_n15164_), .ZN(new_n15201_));
  NOR2_X1    g14178(.A1(new_n15200_), .A2(new_n15201_), .ZN(new_n15202_));
  NAND2_X1   g14179(.A1(new_n15199_), .A2(new_n15202_), .ZN(new_n15203_));
  AOI21_X1   g14180(.A1(new_n15203_), .A2(new_n15196_), .B(new_n15131_), .ZN(new_n15204_));
  OAI21_X1   g14181(.A1(new_n12714_), .A2(new_n12872_), .B(new_n12858_), .ZN(new_n15205_));
  NAND2_X1   g14182(.A1(new_n15199_), .A2(new_n15195_), .ZN(new_n15206_));
  NAND4_X1   g14183(.A1(new_n15197_), .A2(new_n15198_), .A3(new_n15194_), .A4(new_n15187_), .ZN(new_n15207_));
  AOI21_X1   g14184(.A1(new_n15206_), .A2(new_n15207_), .B(new_n15205_), .ZN(new_n15208_));
  NOR2_X1    g14185(.A1(new_n15204_), .A2(new_n15208_), .ZN(new_n15209_));
  OAI21_X1   g14186(.A1(new_n12705_), .A2(new_n12706_), .B(new_n12866_), .ZN(new_n15210_));
  OAI21_X1   g14187(.A1(new_n12667_), .A2(new_n12665_), .B(new_n12666_), .ZN(new_n15211_));
  NAND3_X1   g14188(.A1(new_n12667_), .A2(new_n12666_), .A3(new_n12665_), .ZN(new_n15212_));
  OAI21_X1   g14189(.A1(new_n12661_), .A2(new_n12652_), .B(new_n12658_), .ZN(new_n15213_));
  NAND3_X1   g14190(.A1(new_n12661_), .A2(new_n12652_), .A3(new_n12658_), .ZN(new_n15214_));
  OR4_X2     g14191(.A1(new_n15211_), .A2(new_n15213_), .A3(new_n15214_), .A4(new_n15212_), .Z(new_n15215_));
  NOR2_X1    g14192(.A1(new_n12669_), .A2(new_n12672_), .ZN(new_n15216_));
  NOR2_X1    g14193(.A1(new_n12655_), .A2(new_n12657_), .ZN(new_n15217_));
  NOR4_X1    g14194(.A1(new_n12660_), .A2(new_n12651_), .A3(new_n12659_), .A4(new_n15217_), .ZN(new_n15218_));
  AND2_X2    g14195(.A1(new_n12640_), .A2(new_n12642_), .Z(new_n15219_));
  NOR2_X1    g14196(.A1(new_n12411_), .A2(new_n12406_), .ZN(new_n15220_));
  AOI21_X1   g14197(.A1(new_n15220_), .A2(new_n12624_), .B(new_n12403_), .ZN(new_n15221_));
  NOR2_X1    g14198(.A1(new_n12640_), .A2(new_n12642_), .ZN(new_n15222_));
  NOR4_X1    g14199(.A1(new_n15221_), .A2(new_n12422_), .A3(new_n12633_), .A4(new_n15222_), .ZN(new_n15223_));
  OAI22_X1   g14200(.A1(new_n15219_), .A2(new_n15223_), .B1(new_n15218_), .B2(new_n15216_), .ZN(new_n15224_));
  AOI21_X1   g14201(.A1(new_n12684_), .A2(new_n12637_), .B(new_n15224_), .ZN(new_n15225_));
  NOR2_X1    g14202(.A1(new_n12651_), .A2(new_n15217_), .ZN(new_n15226_));
  AOI21_X1   g14203(.A1(new_n12661_), .A2(new_n15226_), .B(new_n15216_), .ZN(new_n15227_));
  NOR2_X1    g14204(.A1(new_n12633_), .A2(new_n15222_), .ZN(new_n15228_));
  AOI21_X1   g14205(.A1(new_n12667_), .A2(new_n15228_), .B(new_n15219_), .ZN(new_n15229_));
  NOR2_X1    g14206(.A1(new_n15227_), .A2(new_n15229_), .ZN(new_n15230_));
  NOR3_X1    g14207(.A1(new_n12682_), .A2(new_n15230_), .A3(new_n12699_), .ZN(new_n15231_));
  OAI21_X1   g14208(.A1(new_n15231_), .A2(new_n15225_), .B(new_n15215_), .ZN(new_n15232_));
  NOR4_X1    g14209(.A1(new_n15213_), .A2(new_n15214_), .A3(new_n15211_), .A4(new_n15212_), .ZN(new_n15233_));
  OAI21_X1   g14210(.A1(new_n12682_), .A2(new_n12699_), .B(new_n15230_), .ZN(new_n15234_));
  NAND3_X1   g14211(.A1(new_n12684_), .A2(new_n15224_), .A3(new_n12637_), .ZN(new_n15235_));
  NAND3_X1   g14212(.A1(new_n15234_), .A2(new_n15235_), .A3(new_n15233_), .ZN(new_n15236_));
  NAND2_X1   g14213(.A1(new_n15232_), .A2(new_n15236_), .ZN(new_n15237_));
  AOI21_X1   g14214(.A1(new_n12592_), .A2(new_n12512_), .B(new_n12591_), .ZN(new_n15238_));
  INV_X1     g14215(.I(new_n15238_), .ZN(new_n15239_));
  NOR3_X1    g14216(.A1(new_n12592_), .A2(new_n12591_), .A3(new_n12512_), .ZN(new_n15240_));
  NAND4_X1   g14217(.A1(new_n15240_), .A2(new_n12575_), .A3(new_n12581_), .A4(new_n12583_), .ZN(new_n15241_));
  NOR2_X1    g14218(.A1(new_n15241_), .A2(new_n15239_), .ZN(new_n15242_));
  AOI21_X1   g14219(.A1(new_n10824_), .A2(new_n12589_), .B(new_n12587_), .ZN(new_n15243_));
  NOR2_X1    g14220(.A1(new_n12602_), .A2(new_n12590_), .ZN(new_n15244_));
  NOR2_X1    g14221(.A1(new_n12512_), .A2(new_n15244_), .ZN(new_n15245_));
  AOI21_X1   g14222(.A1(new_n12606_), .A2(new_n15245_), .B(new_n15243_), .ZN(new_n15246_));
  AND2_X2    g14223(.A1(new_n12578_), .A2(new_n12580_), .Z(new_n15247_));
  NOR2_X1    g14224(.A1(new_n12578_), .A2(new_n12580_), .ZN(new_n15248_));
  NOR2_X1    g14225(.A1(new_n12574_), .A2(new_n15248_), .ZN(new_n15249_));
  AOI21_X1   g14226(.A1(new_n12583_), .A2(new_n15249_), .B(new_n15247_), .ZN(new_n15250_));
  NOR2_X1    g14227(.A1(new_n15246_), .A2(new_n15250_), .ZN(new_n15251_));
  OAI21_X1   g14228(.A1(new_n12572_), .A2(new_n12615_), .B(new_n15251_), .ZN(new_n15252_));
  NOR4_X1    g14229(.A1(new_n12605_), .A2(new_n12442_), .A3(new_n12512_), .A4(new_n15244_), .ZN(new_n15253_));
  NOR2_X1    g14230(.A1(new_n12517_), .A2(new_n12516_), .ZN(new_n15254_));
  AOI21_X1   g14231(.A1(new_n15254_), .A2(new_n12490_), .B(new_n12515_), .ZN(new_n15255_));
  NOR4_X1    g14232(.A1(new_n15255_), .A2(new_n12524_), .A3(new_n12574_), .A4(new_n15248_), .ZN(new_n15256_));
  OAI22_X1   g14233(.A1(new_n15243_), .A2(new_n15253_), .B1(new_n15256_), .B2(new_n15247_), .ZN(new_n15257_));
  NAND3_X1   g14234(.A1(new_n12692_), .A2(new_n12613_), .A3(new_n15257_), .ZN(new_n15258_));
  AOI21_X1   g14235(.A1(new_n15252_), .A2(new_n15258_), .B(new_n15242_), .ZN(new_n15259_));
  NAND3_X1   g14236(.A1(new_n12606_), .A2(new_n12599_), .A3(new_n12604_), .ZN(new_n15260_));
  NOR4_X1    g14237(.A1(new_n15260_), .A2(new_n12574_), .A3(new_n12595_), .A4(new_n12597_), .ZN(new_n15261_));
  NAND2_X1   g14238(.A1(new_n15261_), .A2(new_n15238_), .ZN(new_n15262_));
  AOI21_X1   g14239(.A1(new_n12692_), .A2(new_n12613_), .B(new_n15257_), .ZN(new_n15263_));
  NOR3_X1    g14240(.A1(new_n12615_), .A2(new_n15251_), .A3(new_n12572_), .ZN(new_n15264_));
  NOR3_X1    g14241(.A1(new_n15264_), .A2(new_n15263_), .A3(new_n15262_), .ZN(new_n15265_));
  NOR2_X1    g14242(.A1(new_n15265_), .A2(new_n15259_), .ZN(new_n15266_));
  NOR2_X1    g14243(.A1(new_n15266_), .A2(new_n15237_), .ZN(new_n15267_));
  AOI21_X1   g14244(.A1(new_n15234_), .A2(new_n15235_), .B(new_n15233_), .ZN(new_n15268_));
  NOR3_X1    g14245(.A1(new_n15231_), .A2(new_n15225_), .A3(new_n15215_), .ZN(new_n15269_));
  NOR2_X1    g14246(.A1(new_n15269_), .A2(new_n15268_), .ZN(new_n15270_));
  OAI21_X1   g14247(.A1(new_n15264_), .A2(new_n15263_), .B(new_n15262_), .ZN(new_n15271_));
  NAND3_X1   g14248(.A1(new_n15252_), .A2(new_n15258_), .A3(new_n15242_), .ZN(new_n15272_));
  NAND2_X1   g14249(.A1(new_n15271_), .A2(new_n15272_), .ZN(new_n15273_));
  NOR2_X1    g14250(.A1(new_n15273_), .A2(new_n15270_), .ZN(new_n15274_));
  OAI21_X1   g14251(.A1(new_n15274_), .A2(new_n15267_), .B(new_n15210_), .ZN(new_n15275_));
  AOI21_X1   g14252(.A1(new_n12568_), .A2(new_n12865_), .B(new_n12707_), .ZN(new_n15276_));
  NOR2_X1    g14253(.A1(new_n15266_), .A2(new_n15270_), .ZN(new_n15277_));
  NOR4_X1    g14254(.A1(new_n15269_), .A2(new_n15259_), .A3(new_n15265_), .A4(new_n15268_), .ZN(new_n15278_));
  OAI21_X1   g14255(.A1(new_n15277_), .A2(new_n15278_), .B(new_n15276_), .ZN(new_n15279_));
  NAND2_X1   g14256(.A1(new_n15275_), .A2(new_n15279_), .ZN(new_n15280_));
  NAND2_X1   g14257(.A1(new_n15209_), .A2(new_n15280_), .ZN(new_n15281_));
  NOR2_X1    g14258(.A1(new_n15199_), .A2(new_n15202_), .ZN(new_n15282_));
  NOR2_X1    g14259(.A1(new_n15160_), .A2(new_n15195_), .ZN(new_n15283_));
  OAI21_X1   g14260(.A1(new_n15282_), .A2(new_n15283_), .B(new_n15205_), .ZN(new_n15284_));
  NOR2_X1    g14261(.A1(new_n15160_), .A2(new_n15202_), .ZN(new_n15285_));
  NOR4_X1    g14262(.A1(new_n15153_), .A2(new_n15159_), .A3(new_n15200_), .A4(new_n15201_), .ZN(new_n15286_));
  OAI21_X1   g14263(.A1(new_n15285_), .A2(new_n15286_), .B(new_n15131_), .ZN(new_n15287_));
  NAND2_X1   g14264(.A1(new_n15284_), .A2(new_n15287_), .ZN(new_n15288_));
  NAND2_X1   g14265(.A1(new_n15273_), .A2(new_n15270_), .ZN(new_n15289_));
  NAND2_X1   g14266(.A1(new_n15266_), .A2(new_n15237_), .ZN(new_n15290_));
  AOI21_X1   g14267(.A1(new_n15289_), .A2(new_n15290_), .B(new_n15276_), .ZN(new_n15291_));
  NAND2_X1   g14268(.A1(new_n15273_), .A2(new_n15237_), .ZN(new_n15292_));
  NAND4_X1   g14269(.A1(new_n15232_), .A2(new_n15271_), .A3(new_n15272_), .A4(new_n15236_), .ZN(new_n15293_));
  AOI21_X1   g14270(.A1(new_n15292_), .A2(new_n15293_), .B(new_n15210_), .ZN(new_n15294_));
  NOR2_X1    g14271(.A1(new_n15291_), .A2(new_n15294_), .ZN(new_n15295_));
  NAND2_X1   g14272(.A1(new_n15288_), .A2(new_n15295_), .ZN(new_n15296_));
  AOI21_X1   g14273(.A1(new_n15281_), .A2(new_n15296_), .B(new_n15130_), .ZN(new_n15297_));
  OAI21_X1   g14274(.A1(new_n12879_), .A2(new_n12878_), .B(new_n13195_), .ZN(new_n15298_));
  OAI22_X1   g14275(.A1(new_n15204_), .A2(new_n15208_), .B1(new_n15291_), .B2(new_n15294_), .ZN(new_n15299_));
  NAND4_X1   g14276(.A1(new_n15284_), .A2(new_n15287_), .A3(new_n15275_), .A4(new_n15279_), .ZN(new_n15300_));
  AOI21_X1   g14277(.A1(new_n15299_), .A2(new_n15300_), .B(new_n15298_), .ZN(new_n15301_));
  NOR2_X1    g14278(.A1(new_n15297_), .A2(new_n15301_), .ZN(new_n15302_));
  NOR3_X1    g14279(.A1(new_n15302_), .A2(new_n15125_), .A3(new_n15129_), .ZN(new_n15303_));
  NOR3_X1    g14280(.A1(new_n15123_), .A2(new_n15115_), .A3(new_n15116_), .ZN(new_n15304_));
  AOI21_X1   g14281(.A1(new_n15035_), .A2(new_n15040_), .B(new_n15111_), .ZN(new_n15305_));
  OAI21_X1   g14282(.A1(new_n15305_), .A2(new_n15304_), .B(new_n15126_), .ZN(new_n15306_));
  AOI22_X1   g14283(.A1(new_n15035_), .A2(new_n15040_), .B1(new_n15105_), .B2(new_n15110_), .ZN(new_n15307_));
  NOR4_X1    g14284(.A1(new_n15116_), .A2(new_n15115_), .A3(new_n15120_), .A4(new_n15122_), .ZN(new_n15308_));
  OAI21_X1   g14285(.A1(new_n15307_), .A2(new_n15308_), .B(new_n14969_), .ZN(new_n15309_));
  NOR2_X1    g14286(.A1(new_n15288_), .A2(new_n15295_), .ZN(new_n15310_));
  NOR2_X1    g14287(.A1(new_n15209_), .A2(new_n15280_), .ZN(new_n15311_));
  OAI21_X1   g14288(.A1(new_n15311_), .A2(new_n15310_), .B(new_n15298_), .ZN(new_n15312_));
  AOI22_X1   g14289(.A1(new_n15284_), .A2(new_n15287_), .B1(new_n15275_), .B2(new_n15279_), .ZN(new_n15313_));
  NOR4_X1    g14290(.A1(new_n15204_), .A2(new_n15208_), .A3(new_n15291_), .A4(new_n15294_), .ZN(new_n15314_));
  OAI21_X1   g14291(.A1(new_n15313_), .A2(new_n15314_), .B(new_n15130_), .ZN(new_n15315_));
  NAND2_X1   g14292(.A1(new_n15312_), .A2(new_n15315_), .ZN(new_n15316_));
  AOI21_X1   g14293(.A1(new_n15306_), .A2(new_n15309_), .B(new_n15316_), .ZN(new_n15317_));
  OAI21_X1   g14294(.A1(new_n15317_), .A2(new_n15303_), .B(new_n14968_), .ZN(new_n15318_));
  AOI21_X1   g14295(.A1(new_n12560_), .A2(new_n13906_), .B(new_n13208_), .ZN(new_n15319_));
  AOI22_X1   g14296(.A1(new_n15306_), .A2(new_n15309_), .B1(new_n15312_), .B2(new_n15315_), .ZN(new_n15320_));
  NOR3_X1    g14297(.A1(new_n15316_), .A2(new_n15125_), .A3(new_n15129_), .ZN(new_n15321_));
  OAI21_X1   g14298(.A1(new_n15320_), .A2(new_n15321_), .B(new_n15319_), .ZN(new_n15322_));
  NAND2_X1   g14299(.A1(new_n15322_), .A2(new_n15318_), .ZN(new_n15323_));
  NAND3_X1   g14300(.A1(new_n15323_), .A2(new_n14963_), .A3(new_n14967_), .ZN(new_n15324_));
  NAND2_X1   g14301(.A1(new_n14963_), .A2(new_n14967_), .ZN(new_n15325_));
  NAND3_X1   g14302(.A1(new_n15316_), .A2(new_n15306_), .A3(new_n15309_), .ZN(new_n15326_));
  OAI21_X1   g14303(.A1(new_n15125_), .A2(new_n15129_), .B(new_n15302_), .ZN(new_n15327_));
  AOI21_X1   g14304(.A1(new_n15327_), .A2(new_n15326_), .B(new_n15319_), .ZN(new_n15328_));
  OAI22_X1   g14305(.A1(new_n15125_), .A2(new_n15129_), .B1(new_n15297_), .B2(new_n15301_), .ZN(new_n15329_));
  NAND4_X1   g14306(.A1(new_n15306_), .A2(new_n15309_), .A3(new_n15312_), .A4(new_n15315_), .ZN(new_n15330_));
  AOI21_X1   g14307(.A1(new_n15329_), .A2(new_n15330_), .B(new_n14968_), .ZN(new_n15331_));
  NOR2_X1    g14308(.A1(new_n15328_), .A2(new_n15331_), .ZN(new_n15332_));
  NAND2_X1   g14309(.A1(new_n15325_), .A2(new_n15332_), .ZN(new_n15333_));
  AOI21_X1   g14310(.A1(new_n15333_), .A2(new_n15324_), .B(new_n14614_), .ZN(new_n15334_));
  OAI21_X1   g14311(.A1(new_n13912_), .A2(new_n13920_), .B(new_n13959_), .ZN(new_n15335_));
  NAND4_X1   g14312(.A1(new_n14963_), .A2(new_n14967_), .A3(new_n15318_), .A4(new_n15322_), .ZN(new_n15336_));
  NAND3_X1   g14313(.A1(new_n14961_), .A2(new_n14772_), .A3(new_n14782_), .ZN(new_n15337_));
  NAND2_X1   g14314(.A1(new_n14783_), .A2(new_n14944_), .ZN(new_n15338_));
  AOI21_X1   g14315(.A1(new_n15338_), .A2(new_n15337_), .B(new_n14964_), .ZN(new_n15339_));
  OAI22_X1   g14316(.A1(new_n14949_), .A2(new_n14952_), .B1(new_n14943_), .B2(new_n14939_), .ZN(new_n15340_));
  NAND4_X1   g14317(.A1(new_n14772_), .A2(new_n14782_), .A3(new_n14960_), .A4(new_n14956_), .ZN(new_n15341_));
  AOI21_X1   g14318(.A1(new_n15340_), .A2(new_n15341_), .B(new_n14615_), .ZN(new_n15342_));
  OAI22_X1   g14319(.A1(new_n15339_), .A2(new_n15342_), .B1(new_n15328_), .B2(new_n15331_), .ZN(new_n15343_));
  AOI21_X1   g14320(.A1(new_n15336_), .A2(new_n15343_), .B(new_n15335_), .ZN(new_n15344_));
  NOR2_X1    g14321(.A1(new_n15334_), .A2(new_n15344_), .ZN(new_n15345_));
  AOI21_X1   g14322(.A1(new_n6017_), .A2(new_n6270_), .B(new_n8192_), .ZN(new_n15346_));
  AOI21_X1   g14323(.A1(new_n6264_), .A2(new_n6130_), .B(new_n6251_), .ZN(new_n15347_));
  AOI21_X1   g14324(.A1(new_n6214_), .A2(new_n5924_), .B(new_n6205_), .ZN(new_n15348_));
  INV_X1     g14325(.I(new_n15348_), .ZN(new_n15349_));
  NOR3_X1    g14326(.A1(new_n6214_), .A2(new_n5924_), .A3(new_n6205_), .ZN(new_n15350_));
  NAND4_X1   g14327(.A1(new_n15350_), .A2(new_n6210_), .A3(new_n6211_), .A4(new_n6212_), .ZN(new_n15351_));
  NOR2_X1    g14328(.A1(new_n15351_), .A2(new_n15349_), .ZN(new_n15352_));
  NAND2_X1   g14329(.A1(new_n6204_), .A2(new_n6201_), .ZN(new_n15353_));
  NOR2_X1    g14330(.A1(new_n6204_), .A2(new_n6201_), .ZN(new_n15354_));
  NOR2_X1    g14331(.A1(new_n5924_), .A2(new_n15354_), .ZN(new_n15355_));
  NAND2_X1   g14332(.A1(new_n6207_), .A2(new_n15355_), .ZN(new_n15356_));
  NAND2_X1   g14333(.A1(new_n6193_), .A2(new_n6190_), .ZN(new_n15357_));
  OR2_X2     g14334(.A1(new_n6193_), .A2(new_n6190_), .Z(new_n15358_));
  NAND4_X1   g14335(.A1(new_n6195_), .A2(new_n6182_), .A3(new_n6210_), .A4(new_n15358_), .ZN(new_n15359_));
  AOI22_X1   g14336(.A1(new_n15356_), .A2(new_n15353_), .B1(new_n15357_), .B2(new_n15359_), .ZN(new_n15360_));
  OAI21_X1   g14337(.A1(new_n6224_), .A2(new_n6241_), .B(new_n15360_), .ZN(new_n15361_));
  INV_X1     g14338(.I(new_n15355_), .ZN(new_n15362_));
  OAI21_X1   g14339(.A1(new_n6214_), .A2(new_n15362_), .B(new_n15353_), .ZN(new_n15363_));
  NAND2_X1   g14340(.A1(new_n15359_), .A2(new_n15357_), .ZN(new_n15364_));
  NAND2_X1   g14341(.A1(new_n15363_), .A2(new_n15364_), .ZN(new_n15365_));
  NAND3_X1   g14342(.A1(new_n6187_), .A2(new_n15365_), .A3(new_n6226_), .ZN(new_n15366_));
  AOI21_X1   g14343(.A1(new_n15361_), .A2(new_n15366_), .B(new_n15352_), .ZN(new_n15367_));
  NAND3_X1   g14344(.A1(new_n6207_), .A2(new_n6198_), .A3(new_n6206_), .ZN(new_n15368_));
  NOR4_X1    g14345(.A1(new_n15368_), .A2(new_n5951_), .A3(new_n6194_), .A4(new_n6196_), .ZN(new_n15369_));
  NAND2_X1   g14346(.A1(new_n15369_), .A2(new_n15348_), .ZN(new_n15370_));
  AOI21_X1   g14347(.A1(new_n6187_), .A2(new_n6226_), .B(new_n15365_), .ZN(new_n15371_));
  NOR3_X1    g14348(.A1(new_n6224_), .A2(new_n15360_), .A3(new_n6241_), .ZN(new_n15372_));
  NOR3_X1    g14349(.A1(new_n15371_), .A2(new_n15372_), .A3(new_n15370_), .ZN(new_n15373_));
  NOR2_X1    g14350(.A1(new_n15373_), .A2(new_n15367_), .ZN(new_n15374_));
  AOI21_X1   g14351(.A1(new_n6157_), .A2(new_n5976_), .B(new_n6155_), .ZN(new_n15375_));
  NAND3_X1   g14352(.A1(new_n6167_), .A2(new_n6165_), .A3(new_n6166_), .ZN(new_n15376_));
  NOR4_X1    g14353(.A1(new_n15376_), .A2(new_n5994_), .A3(new_n6143_), .A4(new_n6163_), .ZN(new_n15377_));
  NAND2_X1   g14354(.A1(new_n15377_), .A2(new_n15375_), .ZN(new_n15378_));
  NAND2_X1   g14355(.A1(new_n6154_), .A2(new_n6151_), .ZN(new_n15379_));
  INV_X1     g14356(.I(new_n15379_), .ZN(new_n15380_));
  OR2_X2     g14357(.A1(new_n6154_), .A2(new_n6151_), .Z(new_n15381_));
  NAND2_X1   g14358(.A1(new_n6165_), .A2(new_n15381_), .ZN(new_n15382_));
  NOR2_X1    g14359(.A1(new_n6157_), .A2(new_n15382_), .ZN(new_n15383_));
  NAND2_X1   g14360(.A1(new_n6142_), .A2(new_n6139_), .ZN(new_n15384_));
  INV_X1     g14361(.I(new_n15384_), .ZN(new_n15385_));
  OR2_X2     g14362(.A1(new_n6142_), .A2(new_n6139_), .Z(new_n15386_));
  INV_X1     g14363(.I(new_n15386_), .ZN(new_n15387_));
  NOR4_X1    g14364(.A1(new_n6146_), .A2(new_n15387_), .A3(new_n5989_), .A4(new_n5994_), .ZN(new_n15388_));
  OAI22_X1   g14365(.A1(new_n15383_), .A2(new_n15380_), .B1(new_n15388_), .B2(new_n15385_), .ZN(new_n15389_));
  AOI21_X1   g14366(.A1(new_n6234_), .A2(new_n6174_), .B(new_n15389_), .ZN(new_n15390_));
  NAND4_X1   g14367(.A1(new_n6156_), .A2(new_n6001_), .A3(new_n6165_), .A4(new_n15381_), .ZN(new_n15391_));
  NAND3_X1   g14368(.A1(new_n6147_), .A2(new_n6136_), .A3(new_n15386_), .ZN(new_n15392_));
  AOI22_X1   g14369(.A1(new_n15392_), .A2(new_n15384_), .B1(new_n15391_), .B2(new_n15379_), .ZN(new_n15393_));
  NOR3_X1    g14370(.A1(new_n15393_), .A2(new_n6176_), .A3(new_n6135_), .ZN(new_n15394_));
  OAI21_X1   g14371(.A1(new_n15390_), .A2(new_n15394_), .B(new_n15378_), .ZN(new_n15395_));
  INV_X1     g14372(.I(new_n15375_), .ZN(new_n15396_));
  NOR3_X1    g14373(.A1(new_n6157_), .A2(new_n5976_), .A3(new_n6155_), .ZN(new_n15397_));
  NAND4_X1   g14374(.A1(new_n15397_), .A2(new_n6136_), .A3(new_n6144_), .A4(new_n6147_), .ZN(new_n15398_));
  NOR2_X1    g14375(.A1(new_n15398_), .A2(new_n15396_), .ZN(new_n15399_));
  OAI21_X1   g14376(.A1(new_n6176_), .A2(new_n6135_), .B(new_n15393_), .ZN(new_n15400_));
  NAND3_X1   g14377(.A1(new_n6234_), .A2(new_n15389_), .A3(new_n6174_), .ZN(new_n15401_));
  NAND3_X1   g14378(.A1(new_n15400_), .A2(new_n15401_), .A3(new_n15399_), .ZN(new_n15402_));
  NAND2_X1   g14379(.A1(new_n15395_), .A2(new_n15402_), .ZN(new_n15403_));
  NAND2_X1   g14380(.A1(new_n15374_), .A2(new_n15403_), .ZN(new_n15404_));
  OAI21_X1   g14381(.A1(new_n15371_), .A2(new_n15372_), .B(new_n15370_), .ZN(new_n15405_));
  NAND3_X1   g14382(.A1(new_n15361_), .A2(new_n15366_), .A3(new_n15352_), .ZN(new_n15406_));
  NAND2_X1   g14383(.A1(new_n15405_), .A2(new_n15406_), .ZN(new_n15407_));
  AOI21_X1   g14384(.A1(new_n15400_), .A2(new_n15401_), .B(new_n15399_), .ZN(new_n15408_));
  NOR3_X1    g14385(.A1(new_n15390_), .A2(new_n15394_), .A3(new_n15378_), .ZN(new_n15409_));
  NOR2_X1    g14386(.A1(new_n15409_), .A2(new_n15408_), .ZN(new_n15410_));
  NAND2_X1   g14387(.A1(new_n15407_), .A2(new_n15410_), .ZN(new_n15411_));
  AOI21_X1   g14388(.A1(new_n15411_), .A2(new_n15404_), .B(new_n15347_), .ZN(new_n15412_));
  OAI21_X1   g14389(.A1(new_n6249_), .A2(new_n6250_), .B(new_n6265_), .ZN(new_n15413_));
  NAND2_X1   g14390(.A1(new_n15407_), .A2(new_n15403_), .ZN(new_n15414_));
  NAND2_X1   g14391(.A1(new_n15374_), .A2(new_n15410_), .ZN(new_n15415_));
  AOI21_X1   g14392(.A1(new_n15415_), .A2(new_n15414_), .B(new_n15413_), .ZN(new_n15416_));
  NOR2_X1    g14393(.A1(new_n15412_), .A2(new_n15416_), .ZN(new_n15417_));
  OAI21_X1   g14394(.A1(new_n6020_), .A2(new_n6121_), .B(new_n6123_), .ZN(new_n15418_));
  AOI21_X1   g14395(.A1(new_n6082_), .A2(new_n5811_), .B(new_n6081_), .ZN(new_n15419_));
  NAND3_X1   g14396(.A1(new_n6095_), .A2(new_n6093_), .A3(new_n6094_), .ZN(new_n15420_));
  NOR4_X1    g14397(.A1(new_n15420_), .A2(new_n5845_), .A3(new_n6085_), .A4(new_n6091_), .ZN(new_n15421_));
  NAND2_X1   g14398(.A1(new_n15421_), .A2(new_n15419_), .ZN(new_n15422_));
  NAND2_X1   g14399(.A1(new_n6092_), .A2(new_n6083_), .ZN(new_n15423_));
  NAND2_X1   g14400(.A1(new_n6080_), .A2(new_n6077_), .ZN(new_n15424_));
  INV_X1     g14401(.I(new_n15424_), .ZN(new_n15425_));
  NAND4_X1   g14402(.A1(new_n6079_), .A2(new_n5599_), .A3(new_n5626_), .A4(new_n6076_), .ZN(new_n15426_));
  NAND3_X1   g14403(.A1(new_n6095_), .A2(new_n6093_), .A3(new_n15426_), .ZN(new_n15427_));
  INV_X1     g14404(.I(new_n15427_), .ZN(new_n15428_));
  NAND2_X1   g14405(.A1(new_n6070_), .A2(new_n6067_), .ZN(new_n15429_));
  NOR2_X1    g14406(.A1(new_n6070_), .A2(new_n6067_), .ZN(new_n15430_));
  NOR2_X1    g14407(.A1(new_n5845_), .A2(new_n15430_), .ZN(new_n15431_));
  NAND2_X1   g14408(.A1(new_n6073_), .A2(new_n15431_), .ZN(new_n15432_));
  NAND2_X1   g14409(.A1(new_n15432_), .A2(new_n15429_), .ZN(new_n15433_));
  OAI21_X1   g14410(.A1(new_n15425_), .A2(new_n15428_), .B(new_n15433_), .ZN(new_n15434_));
  AOI21_X1   g14411(.A1(new_n6100_), .A2(new_n15423_), .B(new_n15434_), .ZN(new_n15435_));
  NAND2_X1   g14412(.A1(new_n6100_), .A2(new_n15423_), .ZN(new_n15436_));
  AOI22_X1   g14413(.A1(new_n6073_), .A2(new_n15431_), .B1(new_n6067_), .B2(new_n6070_), .ZN(new_n15437_));
  AOI21_X1   g14414(.A1(new_n15424_), .A2(new_n15427_), .B(new_n15437_), .ZN(new_n15438_));
  NOR2_X1    g14415(.A1(new_n15436_), .A2(new_n15438_), .ZN(new_n15439_));
  OAI21_X1   g14416(.A1(new_n15439_), .A2(new_n15435_), .B(new_n15422_), .ZN(new_n15440_));
  INV_X1     g14417(.I(new_n15422_), .ZN(new_n15441_));
  NAND2_X1   g14418(.A1(new_n15436_), .A2(new_n15438_), .ZN(new_n15442_));
  NAND3_X1   g14419(.A1(new_n15434_), .A2(new_n6100_), .A3(new_n15423_), .ZN(new_n15443_));
  NAND3_X1   g14420(.A1(new_n15442_), .A2(new_n15441_), .A3(new_n15443_), .ZN(new_n15444_));
  NAND2_X1   g14421(.A1(new_n15440_), .A2(new_n15444_), .ZN(new_n15445_));
  OAI21_X1   g14422(.A1(new_n6052_), .A2(new_n6051_), .B(new_n6042_), .ZN(new_n15446_));
  NOR3_X1    g14423(.A1(new_n6044_), .A2(new_n6043_), .A3(new_n5875_), .ZN(new_n15447_));
  NAND4_X1   g14424(.A1(new_n15447_), .A2(new_n6026_), .A3(new_n6033_), .A4(new_n6034_), .ZN(new_n15448_));
  NOR2_X1    g14425(.A1(new_n15448_), .A2(new_n15446_), .ZN(new_n15449_));
  NAND2_X1   g14426(.A1(new_n6045_), .A2(new_n6050_), .ZN(new_n15450_));
  NAND2_X1   g14427(.A1(new_n6109_), .A2(new_n15450_), .ZN(new_n15451_));
  NOR2_X1    g14428(.A1(new_n6041_), .A2(new_n6038_), .ZN(new_n15452_));
  NOR2_X1    g14429(.A1(new_n5875_), .A2(new_n15452_), .ZN(new_n15453_));
  AOI22_X1   g14430(.A1(new_n6052_), .A2(new_n15453_), .B1(new_n6038_), .B2(new_n6041_), .ZN(new_n15454_));
  NAND2_X1   g14431(.A1(new_n6032_), .A2(new_n6029_), .ZN(new_n15455_));
  INV_X1     g14432(.I(new_n15455_), .ZN(new_n15456_));
  NOR2_X1    g14433(.A1(new_n6032_), .A2(new_n6029_), .ZN(new_n15457_));
  NOR3_X1    g14434(.A1(new_n6049_), .A2(new_n5893_), .A3(new_n15457_), .ZN(new_n15458_));
  NOR2_X1    g14435(.A1(new_n15458_), .A2(new_n15456_), .ZN(new_n15459_));
  NOR2_X1    g14436(.A1(new_n15459_), .A2(new_n15454_), .ZN(new_n15460_));
  NAND2_X1   g14437(.A1(new_n15451_), .A2(new_n15460_), .ZN(new_n15461_));
  NAND2_X1   g14438(.A1(new_n6041_), .A2(new_n6038_), .ZN(new_n15462_));
  NAND2_X1   g14439(.A1(new_n6052_), .A2(new_n15453_), .ZN(new_n15463_));
  NAND2_X1   g14440(.A1(new_n15463_), .A2(new_n15462_), .ZN(new_n15464_));
  OAI21_X1   g14441(.A1(new_n15456_), .A2(new_n15458_), .B(new_n15464_), .ZN(new_n15465_));
  NAND3_X1   g14442(.A1(new_n15465_), .A2(new_n6109_), .A3(new_n15450_), .ZN(new_n15466_));
  AOI21_X1   g14443(.A1(new_n15461_), .A2(new_n15466_), .B(new_n15449_), .ZN(new_n15467_));
  INV_X1     g14444(.I(new_n15449_), .ZN(new_n15468_));
  AOI21_X1   g14445(.A1(new_n6109_), .A2(new_n15450_), .B(new_n15465_), .ZN(new_n15469_));
  NOR2_X1    g14446(.A1(new_n15451_), .A2(new_n15460_), .ZN(new_n15470_));
  NOR3_X1    g14447(.A1(new_n15469_), .A2(new_n15470_), .A3(new_n15468_), .ZN(new_n15471_));
  NOR2_X1    g14448(.A1(new_n15471_), .A2(new_n15467_), .ZN(new_n15472_));
  NOR2_X1    g14449(.A1(new_n15472_), .A2(new_n15445_), .ZN(new_n15473_));
  AOI21_X1   g14450(.A1(new_n15442_), .A2(new_n15443_), .B(new_n15441_), .ZN(new_n15474_));
  NOR3_X1    g14451(.A1(new_n15439_), .A2(new_n15435_), .A3(new_n15422_), .ZN(new_n15475_));
  NOR2_X1    g14452(.A1(new_n15475_), .A2(new_n15474_), .ZN(new_n15476_));
  OAI21_X1   g14453(.A1(new_n15469_), .A2(new_n15470_), .B(new_n15468_), .ZN(new_n15477_));
  NAND3_X1   g14454(.A1(new_n15461_), .A2(new_n15466_), .A3(new_n15449_), .ZN(new_n15478_));
  NAND2_X1   g14455(.A1(new_n15477_), .A2(new_n15478_), .ZN(new_n15479_));
  NOR2_X1    g14456(.A1(new_n15479_), .A2(new_n15476_), .ZN(new_n15480_));
  OAI21_X1   g14457(.A1(new_n15473_), .A2(new_n15480_), .B(new_n15418_), .ZN(new_n15481_));
  AOI21_X1   g14458(.A1(new_n6122_), .A2(new_n6120_), .B(new_n6258_), .ZN(new_n15482_));
  NOR2_X1    g14459(.A1(new_n15472_), .A2(new_n15476_), .ZN(new_n15483_));
  NOR2_X1    g14460(.A1(new_n15479_), .A2(new_n15445_), .ZN(new_n15484_));
  OAI21_X1   g14461(.A1(new_n15483_), .A2(new_n15484_), .B(new_n15482_), .ZN(new_n15485_));
  NAND2_X1   g14462(.A1(new_n15481_), .A2(new_n15485_), .ZN(new_n15486_));
  NAND2_X1   g14463(.A1(new_n15486_), .A2(new_n15417_), .ZN(new_n15487_));
  NOR2_X1    g14464(.A1(new_n15407_), .A2(new_n15410_), .ZN(new_n15488_));
  NOR2_X1    g14465(.A1(new_n15374_), .A2(new_n15403_), .ZN(new_n15489_));
  OAI21_X1   g14466(.A1(new_n15488_), .A2(new_n15489_), .B(new_n15413_), .ZN(new_n15490_));
  NOR2_X1    g14467(.A1(new_n15374_), .A2(new_n15410_), .ZN(new_n15491_));
  NOR2_X1    g14468(.A1(new_n15407_), .A2(new_n15403_), .ZN(new_n15492_));
  OAI21_X1   g14469(.A1(new_n15491_), .A2(new_n15492_), .B(new_n15347_), .ZN(new_n15493_));
  NAND2_X1   g14470(.A1(new_n15490_), .A2(new_n15493_), .ZN(new_n15494_));
  NAND2_X1   g14471(.A1(new_n15479_), .A2(new_n15476_), .ZN(new_n15495_));
  NAND2_X1   g14472(.A1(new_n15472_), .A2(new_n15445_), .ZN(new_n15496_));
  AOI21_X1   g14473(.A1(new_n15495_), .A2(new_n15496_), .B(new_n15482_), .ZN(new_n15497_));
  NAND2_X1   g14474(.A1(new_n15479_), .A2(new_n15445_), .ZN(new_n15498_));
  NAND2_X1   g14475(.A1(new_n15472_), .A2(new_n15476_), .ZN(new_n15499_));
  AOI21_X1   g14476(.A1(new_n15498_), .A2(new_n15499_), .B(new_n15418_), .ZN(new_n15500_));
  NOR2_X1    g14477(.A1(new_n15500_), .A2(new_n15497_), .ZN(new_n15501_));
  NAND2_X1   g14478(.A1(new_n15501_), .A2(new_n15494_), .ZN(new_n15502_));
  AOI21_X1   g14479(.A1(new_n15487_), .A2(new_n15502_), .B(new_n15346_), .ZN(new_n15503_));
  OAI21_X1   g14480(.A1(new_n8191_), .A2(new_n6018_), .B(new_n6271_), .ZN(new_n15504_));
  NAND2_X1   g14481(.A1(new_n15486_), .A2(new_n15494_), .ZN(new_n15505_));
  NAND2_X1   g14482(.A1(new_n15501_), .A2(new_n15417_), .ZN(new_n15506_));
  AOI21_X1   g14483(.A1(new_n15506_), .A2(new_n15505_), .B(new_n15504_), .ZN(new_n15507_));
  NOR2_X1    g14484(.A1(new_n15503_), .A2(new_n15507_), .ZN(new_n15508_));
  NAND2_X1   g14485(.A1(new_n8119_), .A2(new_n7860_), .ZN(new_n15509_));
  NOR2_X1    g14486(.A1(new_n7941_), .A2(new_n7589_), .ZN(new_n15510_));
  NOR2_X1    g14487(.A1(new_n7968_), .A2(new_n7495_), .ZN(new_n15511_));
  NAND2_X1   g14488(.A1(new_n7536_), .A2(new_n7160_), .ZN(new_n15512_));
  NAND2_X1   g14489(.A1(new_n7958_), .A2(new_n7488_), .ZN(new_n15513_));
  XNOR2_X1   g14490(.A1(new_n15513_), .A2(new_n15512_), .ZN(new_n15514_));
  NAND2_X1   g14491(.A1(new_n7591_), .A2(new_n7186_), .ZN(new_n15515_));
  NAND2_X1   g14492(.A1(new_n7943_), .A2(new_n7583_), .ZN(new_n15516_));
  XNOR2_X1   g14493(.A1(new_n15516_), .A2(new_n15515_), .ZN(new_n15517_));
  NOR4_X1    g14494(.A1(new_n7955_), .A2(new_n7950_), .A3(new_n15514_), .A4(new_n15517_), .ZN(new_n15518_));
  INV_X1     g14495(.I(new_n15510_), .ZN(new_n15519_));
  INV_X1     g14496(.I(new_n15511_), .ZN(new_n15520_));
  AOI22_X1   g14497(.A1(new_n7955_), .A2(new_n15520_), .B1(new_n15519_), .B2(new_n7950_), .ZN(new_n15521_));
  NAND4_X1   g14498(.A1(new_n15521_), .A2(new_n15510_), .A3(new_n15518_), .A4(new_n15511_), .ZN(new_n15522_));
  INV_X1     g14499(.I(new_n15522_), .ZN(new_n15523_));
  NOR2_X1    g14500(.A1(new_n15513_), .A2(new_n15512_), .ZN(new_n15524_));
  NOR2_X1    g14501(.A1(new_n7955_), .A2(new_n15524_), .ZN(new_n15525_));
  NAND2_X1   g14502(.A1(new_n15525_), .A2(new_n15511_), .ZN(new_n15526_));
  NAND4_X1   g14503(.A1(new_n7943_), .A2(new_n7591_), .A3(new_n7583_), .A4(new_n7186_), .ZN(new_n15527_));
  NAND4_X1   g14504(.A1(new_n15510_), .A2(new_n7564_), .A3(new_n7593_), .A4(new_n15527_), .ZN(new_n15528_));
  AOI22_X1   g14505(.A1(new_n15526_), .A2(new_n7960_), .B1(new_n7947_), .B2(new_n15528_), .ZN(new_n15529_));
  OAI21_X1   g14506(.A1(new_n7997_), .A2(new_n7985_), .B(new_n15529_), .ZN(new_n15530_));
  OAI21_X1   g14507(.A1(new_n15512_), .A2(new_n15513_), .B(new_n7538_), .ZN(new_n15531_));
  OAI21_X1   g14508(.A1(new_n15520_), .A2(new_n15531_), .B(new_n7960_), .ZN(new_n15532_));
  NAND2_X1   g14509(.A1(new_n15528_), .A2(new_n7947_), .ZN(new_n15533_));
  NAND2_X1   g14510(.A1(new_n15533_), .A2(new_n15532_), .ZN(new_n15534_));
  NAND3_X1   g14511(.A1(new_n15534_), .A2(new_n7987_), .A3(new_n7939_), .ZN(new_n15535_));
  AOI21_X1   g14512(.A1(new_n15530_), .A2(new_n15535_), .B(new_n15523_), .ZN(new_n15536_));
  AOI21_X1   g14513(.A1(new_n7987_), .A2(new_n7939_), .B(new_n15534_), .ZN(new_n15537_));
  NOR3_X1    g14514(.A1(new_n7997_), .A2(new_n15529_), .A3(new_n7985_), .ZN(new_n15538_));
  NOR3_X1    g14515(.A1(new_n15537_), .A2(new_n15538_), .A3(new_n15522_), .ZN(new_n15539_));
  NOR2_X1    g14516(.A1(new_n15536_), .A2(new_n15539_), .ZN(new_n15540_));
  NOR2_X1    g14517(.A1(new_n7849_), .A2(new_n7640_), .ZN(new_n15541_));
  XOR2_X1    g14518(.A1(new_n7891_), .A2(new_n7888_), .Z(new_n15542_));
  NAND3_X1   g14519(.A1(new_n7845_), .A2(new_n15542_), .A3(new_n7869_), .ZN(new_n15543_));
  NOR2_X1    g14520(.A1(new_n15543_), .A2(new_n7868_), .ZN(new_n15544_));
  INV_X1     g14521(.I(new_n15541_), .ZN(new_n15545_));
  NAND2_X1   g14522(.A1(new_n15545_), .A2(new_n7691_), .ZN(new_n15546_));
  NAND2_X1   g14523(.A1(new_n7870_), .A2(new_n7789_), .ZN(new_n15547_));
  NAND2_X1   g14524(.A1(new_n15547_), .A2(new_n7873_), .ZN(new_n15548_));
  NAND3_X1   g14525(.A1(new_n7879_), .A2(new_n7870_), .A3(new_n7789_), .ZN(new_n15549_));
  AOI22_X1   g14526(.A1(new_n7868_), .A2(new_n7877_), .B1(new_n15549_), .B2(new_n15548_), .ZN(new_n15550_));
  NAND4_X1   g14527(.A1(new_n15546_), .A2(new_n15544_), .A3(new_n15550_), .A4(new_n15541_), .ZN(new_n15551_));
  AOI22_X1   g14528(.A1(new_n7864_), .A2(new_n7865_), .B1(new_n7882_), .B2(new_n7886_), .ZN(new_n15552_));
  AOI21_X1   g14529(.A1(new_n7896_), .A2(new_n7899_), .B(new_n7867_), .ZN(new_n15553_));
  NOR2_X1    g14530(.A1(new_n7891_), .A2(new_n7888_), .ZN(new_n15554_));
  NOR2_X1    g14531(.A1(new_n7691_), .A2(new_n15554_), .ZN(new_n15555_));
  NAND2_X1   g14532(.A1(new_n15541_), .A2(new_n15555_), .ZN(new_n15556_));
  NAND2_X1   g14533(.A1(new_n15556_), .A2(new_n7892_), .ZN(new_n15557_));
  NAND2_X1   g14534(.A1(new_n15547_), .A2(new_n7879_), .ZN(new_n15558_));
  NAND3_X1   g14535(.A1(new_n7883_), .A2(new_n15558_), .A3(new_n7869_), .ZN(new_n15559_));
  NAND2_X1   g14536(.A1(new_n15559_), .A2(new_n7874_), .ZN(new_n15560_));
  NAND2_X1   g14537(.A1(new_n15557_), .A2(new_n15560_), .ZN(new_n15561_));
  NOR3_X1    g14538(.A1(new_n15552_), .A2(new_n15553_), .A3(new_n15561_), .ZN(new_n15562_));
  OAI22_X1   g14539(.A1(new_n7913_), .A2(new_n7914_), .B1(new_n7903_), .B2(new_n7904_), .ZN(new_n15563_));
  OAI21_X1   g14540(.A1(new_n7906_), .A2(new_n7907_), .B(new_n7902_), .ZN(new_n15564_));
  AOI22_X1   g14541(.A1(new_n15556_), .A2(new_n7892_), .B1(new_n15559_), .B2(new_n7874_), .ZN(new_n15565_));
  AOI21_X1   g14542(.A1(new_n15563_), .A2(new_n15564_), .B(new_n15565_), .ZN(new_n15566_));
  OAI21_X1   g14543(.A1(new_n15566_), .A2(new_n15562_), .B(new_n15551_), .ZN(new_n15567_));
  INV_X1     g14544(.I(new_n15551_), .ZN(new_n15568_));
  NAND3_X1   g14545(.A1(new_n15563_), .A2(new_n15564_), .A3(new_n15565_), .ZN(new_n15569_));
  OAI21_X1   g14546(.A1(new_n15552_), .A2(new_n15553_), .B(new_n15561_), .ZN(new_n15570_));
  NAND3_X1   g14547(.A1(new_n15569_), .A2(new_n15570_), .A3(new_n15568_), .ZN(new_n15571_));
  NAND2_X1   g14548(.A1(new_n15567_), .A2(new_n15571_), .ZN(new_n15572_));
  NAND2_X1   g14549(.A1(new_n15572_), .A2(new_n15540_), .ZN(new_n15573_));
  OAI21_X1   g14550(.A1(new_n15537_), .A2(new_n15538_), .B(new_n15522_), .ZN(new_n15574_));
  NAND3_X1   g14551(.A1(new_n15530_), .A2(new_n15523_), .A3(new_n15535_), .ZN(new_n15575_));
  NAND2_X1   g14552(.A1(new_n15574_), .A2(new_n15575_), .ZN(new_n15576_));
  AOI21_X1   g14553(.A1(new_n15569_), .A2(new_n15570_), .B(new_n15568_), .ZN(new_n15577_));
  NOR3_X1    g14554(.A1(new_n15566_), .A2(new_n15562_), .A3(new_n15551_), .ZN(new_n15578_));
  NOR2_X1    g14555(.A1(new_n15577_), .A2(new_n15578_), .ZN(new_n15579_));
  NAND2_X1   g14556(.A1(new_n15579_), .A2(new_n15576_), .ZN(new_n15580_));
  AOI22_X1   g14557(.A1(new_n15580_), .A2(new_n15573_), .B1(new_n15509_), .B2(new_n8120_), .ZN(new_n15581_));
  OAI21_X1   g14558(.A1(new_n8007_), .A2(new_n8006_), .B(new_n8120_), .ZN(new_n15582_));
  OAI22_X1   g14559(.A1(new_n15577_), .A2(new_n15578_), .B1(new_n15536_), .B2(new_n15539_), .ZN(new_n15583_));
  NAND4_X1   g14560(.A1(new_n15567_), .A2(new_n15571_), .A3(new_n15574_), .A4(new_n15575_), .ZN(new_n15584_));
  AOI21_X1   g14561(.A1(new_n15583_), .A2(new_n15584_), .B(new_n15582_), .ZN(new_n15585_));
  NAND2_X1   g14562(.A1(new_n8090_), .A2(new_n8036_), .ZN(new_n15586_));
  NOR2_X1    g14563(.A1(new_n8090_), .A2(new_n8036_), .ZN(new_n15587_));
  NOR3_X1    g14564(.A1(new_n8092_), .A2(new_n8091_), .A3(new_n8012_), .ZN(new_n15588_));
  AOI21_X1   g14565(.A1(new_n8082_), .A2(new_n8087_), .B(new_n8103_), .ZN(new_n15589_));
  NOR2_X1    g14566(.A1(new_n15589_), .A2(new_n15588_), .ZN(new_n15590_));
  OAI21_X1   g14567(.A1(new_n15590_), .A2(new_n15587_), .B(new_n15586_), .ZN(new_n15591_));
  NOR3_X1    g14568(.A1(new_n7073_), .A2(new_n7067_), .A3(new_n7022_), .ZN(new_n15592_));
  OAI21_X1   g14569(.A1(new_n7431_), .A2(new_n7466_), .B(new_n15592_), .ZN(new_n15593_));
  NOR2_X1    g14570(.A1(new_n7078_), .A2(new_n7430_), .ZN(new_n15594_));
  OAI21_X1   g14571(.A1(new_n15594_), .A2(new_n7464_), .B(new_n7469_), .ZN(new_n15595_));
  NAND2_X1   g14572(.A1(new_n15595_), .A2(new_n15593_), .ZN(new_n15596_));
  AOI21_X1   g14573(.A1(new_n7432_), .A2(new_n8037_), .B(new_n7078_), .ZN(new_n15597_));
  NOR3_X1    g14574(.A1(new_n15597_), .A2(new_n8026_), .A3(new_n8018_), .ZN(new_n15598_));
  AOI21_X1   g14575(.A1(new_n7464_), .A2(new_n7465_), .B(new_n8021_), .ZN(new_n15599_));
  INV_X1     g14576(.I(new_n15599_), .ZN(new_n15600_));
  OAI21_X1   g14577(.A1(new_n15598_), .A2(new_n15595_), .B(new_n15600_), .ZN(new_n15601_));
  NAND3_X1   g14578(.A1(new_n15601_), .A2(new_n8026_), .A3(new_n15596_), .ZN(new_n15602_));
  NAND2_X1   g14579(.A1(new_n15592_), .A2(new_n7465_), .ZN(new_n15603_));
  AOI21_X1   g14580(.A1(new_n15603_), .A2(new_n7428_), .B(new_n7457_), .ZN(new_n15604_));
  NOR2_X1    g14581(.A1(new_n15604_), .A2(new_n15597_), .ZN(new_n15605_));
  NAND3_X1   g14582(.A1(new_n15593_), .A2(new_n8032_), .A3(new_n8017_), .ZN(new_n15606_));
  AOI21_X1   g14583(.A1(new_n15606_), .A2(new_n15604_), .B(new_n15599_), .ZN(new_n15607_));
  OAI21_X1   g14584(.A1(new_n15607_), .A2(new_n8032_), .B(new_n15605_), .ZN(new_n15608_));
  NAND2_X1   g14585(.A1(new_n15608_), .A2(new_n15602_), .ZN(new_n15609_));
  XOR2_X1    g14586(.A1(new_n8075_), .A2(new_n8074_), .Z(new_n15610_));
  XOR2_X1    g14587(.A1(new_n8052_), .A2(new_n8055_), .Z(new_n15611_));
  NAND4_X1   g14588(.A1(new_n15610_), .A2(new_n8067_), .A3(new_n8044_), .A4(new_n15611_), .ZN(new_n15612_));
  NOR2_X1    g14589(.A1(new_n8050_), .A2(new_n8045_), .ZN(new_n15613_));
  NOR2_X1    g14590(.A1(new_n8068_), .A2(new_n7269_), .ZN(new_n15614_));
  NAND2_X1   g14591(.A1(new_n15613_), .A2(new_n15614_), .ZN(new_n15615_));
  NOR2_X1    g14592(.A1(new_n15613_), .A2(new_n8044_), .ZN(new_n15616_));
  NOR2_X1    g14593(.A1(new_n15614_), .A2(new_n8067_), .ZN(new_n15617_));
  NOR4_X1    g14594(.A1(new_n15612_), .A2(new_n15615_), .A3(new_n15616_), .A4(new_n15617_), .ZN(new_n15618_));
  INV_X1     g14595(.I(new_n15618_), .ZN(new_n15619_));
  NOR2_X1    g14596(.A1(new_n8075_), .A2(new_n8074_), .ZN(new_n15620_));
  NOR2_X1    g14597(.A1(new_n8066_), .A2(new_n15620_), .ZN(new_n15621_));
  NAND2_X1   g14598(.A1(new_n15614_), .A2(new_n15621_), .ZN(new_n15622_));
  NAND2_X1   g14599(.A1(new_n15622_), .A2(new_n8076_), .ZN(new_n15623_));
  NAND2_X1   g14600(.A1(new_n8059_), .A2(new_n7370_), .ZN(new_n15624_));
  OAI21_X1   g14601(.A1(new_n8052_), .A2(new_n8055_), .B(new_n8044_), .ZN(new_n15625_));
  OAI21_X1   g14602(.A1(new_n15625_), .A2(new_n15624_), .B(new_n8056_), .ZN(new_n15626_));
  NAND2_X1   g14603(.A1(new_n15623_), .A2(new_n15626_), .ZN(new_n15627_));
  AOI21_X1   g14604(.A1(new_n8087_), .A2(new_n8012_), .B(new_n15627_), .ZN(new_n15628_));
  NOR2_X1    g14605(.A1(new_n8052_), .A2(new_n8055_), .ZN(new_n15629_));
  NOR2_X1    g14606(.A1(new_n8062_), .A2(new_n15629_), .ZN(new_n15630_));
  NAND2_X1   g14607(.A1(new_n15630_), .A2(new_n15613_), .ZN(new_n15631_));
  AOI22_X1   g14608(.A1(new_n15631_), .A2(new_n8056_), .B1(new_n8076_), .B2(new_n15622_), .ZN(new_n15632_));
  NOR3_X1    g14609(.A1(new_n8092_), .A2(new_n8103_), .A3(new_n15632_), .ZN(new_n15633_));
  OAI21_X1   g14610(.A1(new_n15633_), .A2(new_n15628_), .B(new_n15619_), .ZN(new_n15634_));
  OAI21_X1   g14611(.A1(new_n8092_), .A2(new_n8103_), .B(new_n15632_), .ZN(new_n15635_));
  NAND3_X1   g14612(.A1(new_n8087_), .A2(new_n15627_), .A3(new_n8012_), .ZN(new_n15636_));
  NAND3_X1   g14613(.A1(new_n15635_), .A2(new_n15636_), .A3(new_n15618_), .ZN(new_n15637_));
  AOI21_X1   g14614(.A1(new_n15634_), .A2(new_n15637_), .B(new_n15609_), .ZN(new_n15638_));
  NOR3_X1    g14615(.A1(new_n15607_), .A2(new_n8032_), .A3(new_n15605_), .ZN(new_n15639_));
  AOI21_X1   g14616(.A1(new_n15601_), .A2(new_n8026_), .B(new_n15596_), .ZN(new_n15640_));
  NOR2_X1    g14617(.A1(new_n15640_), .A2(new_n15639_), .ZN(new_n15641_));
  AOI21_X1   g14618(.A1(new_n15635_), .A2(new_n15636_), .B(new_n15618_), .ZN(new_n15642_));
  NOR3_X1    g14619(.A1(new_n15633_), .A2(new_n15628_), .A3(new_n15619_), .ZN(new_n15643_));
  NOR3_X1    g14620(.A1(new_n15643_), .A2(new_n15642_), .A3(new_n15641_), .ZN(new_n15644_));
  OAI21_X1   g14621(.A1(new_n15644_), .A2(new_n15638_), .B(new_n15591_), .ZN(new_n15645_));
  NOR2_X1    g14622(.A1(new_n8043_), .A2(new_n8098_), .ZN(new_n15646_));
  NAND2_X1   g14623(.A1(new_n8043_), .A2(new_n8098_), .ZN(new_n15647_));
  NAND3_X1   g14624(.A1(new_n8103_), .A2(new_n8082_), .A3(new_n8087_), .ZN(new_n15648_));
  OAI21_X1   g14625(.A1(new_n8092_), .A2(new_n8091_), .B(new_n8012_), .ZN(new_n15649_));
  NAND2_X1   g14626(.A1(new_n15648_), .A2(new_n15649_), .ZN(new_n15650_));
  AOI21_X1   g14627(.A1(new_n15650_), .A2(new_n15647_), .B(new_n15646_), .ZN(new_n15651_));
  AOI21_X1   g14628(.A1(new_n15634_), .A2(new_n15637_), .B(new_n15641_), .ZN(new_n15652_));
  NOR3_X1    g14629(.A1(new_n15643_), .A2(new_n15642_), .A3(new_n15609_), .ZN(new_n15653_));
  OAI21_X1   g14630(.A1(new_n15653_), .A2(new_n15652_), .B(new_n15651_), .ZN(new_n15654_));
  NAND2_X1   g14631(.A1(new_n15645_), .A2(new_n15654_), .ZN(new_n15655_));
  OAI21_X1   g14632(.A1(new_n15581_), .A2(new_n15585_), .B(new_n15655_), .ZN(new_n15656_));
  NOR2_X1    g14633(.A1(new_n15579_), .A2(new_n15576_), .ZN(new_n15657_));
  NOR2_X1    g14634(.A1(new_n15572_), .A2(new_n15540_), .ZN(new_n15658_));
  OAI21_X1   g14635(.A1(new_n15657_), .A2(new_n15658_), .B(new_n15582_), .ZN(new_n15659_));
  AOI21_X1   g14636(.A1(new_n7860_), .A2(new_n8119_), .B(new_n8008_), .ZN(new_n15660_));
  NAND2_X1   g14637(.A1(new_n15583_), .A2(new_n15584_), .ZN(new_n15661_));
  NAND2_X1   g14638(.A1(new_n15661_), .A2(new_n15660_), .ZN(new_n15662_));
  OAI21_X1   g14639(.A1(new_n15643_), .A2(new_n15642_), .B(new_n15641_), .ZN(new_n15663_));
  NAND3_X1   g14640(.A1(new_n15634_), .A2(new_n15637_), .A3(new_n15609_), .ZN(new_n15664_));
  AOI21_X1   g14641(.A1(new_n15663_), .A2(new_n15664_), .B(new_n15651_), .ZN(new_n15665_));
  OAI21_X1   g14642(.A1(new_n15643_), .A2(new_n15642_), .B(new_n15609_), .ZN(new_n15666_));
  NAND3_X1   g14643(.A1(new_n15634_), .A2(new_n15637_), .A3(new_n15641_), .ZN(new_n15667_));
  AOI21_X1   g14644(.A1(new_n15666_), .A2(new_n15667_), .B(new_n15591_), .ZN(new_n15668_));
  NOR2_X1    g14645(.A1(new_n15668_), .A2(new_n15665_), .ZN(new_n15669_));
  NAND3_X1   g14646(.A1(new_n15662_), .A2(new_n15659_), .A3(new_n15669_), .ZN(new_n15670_));
  NAND2_X1   g14647(.A1(new_n15656_), .A2(new_n15670_), .ZN(new_n15671_));
  OAI21_X1   g14648(.A1(new_n8115_), .A2(new_n8129_), .B(new_n8123_), .ZN(new_n15672_));
  INV_X1     g14649(.I(new_n6788_), .ZN(new_n15673_));
  NOR3_X1    g14650(.A1(new_n6834_), .A2(new_n6882_), .A3(new_n6887_), .ZN(new_n15674_));
  AOI21_X1   g14651(.A1(new_n6890_), .A2(new_n15673_), .B(new_n15674_), .ZN(new_n15675_));
  XOR2_X1    g14652(.A1(new_n6860_), .A2(new_n6862_), .Z(new_n15676_));
  XOR2_X1    g14653(.A1(new_n6845_), .A2(new_n6847_), .Z(new_n15677_));
  NAND4_X1   g14654(.A1(new_n6869_), .A2(new_n6839_), .A3(new_n15676_), .A4(new_n15677_), .ZN(new_n15678_));
  INV_X1     g14655(.I(new_n6844_), .ZN(new_n15679_));
  AOI21_X1   g14656(.A1(new_n6836_), .A2(new_n6629_), .B(new_n6611_), .ZN(new_n15680_));
  NAND2_X1   g14657(.A1(new_n15679_), .A2(new_n15680_), .ZN(new_n15681_));
  NOR2_X1    g14658(.A1(new_n15679_), .A2(new_n6839_), .ZN(new_n15682_));
  NOR2_X1    g14659(.A1(new_n15680_), .A2(new_n6869_), .ZN(new_n15683_));
  NOR4_X1    g14660(.A1(new_n15678_), .A2(new_n15682_), .A3(new_n15681_), .A4(new_n15683_), .ZN(new_n15684_));
  AND2_X2    g14661(.A1(new_n6860_), .A2(new_n6862_), .Z(new_n15685_));
  NOR2_X1    g14662(.A1(new_n6858_), .A2(new_n15685_), .ZN(new_n15686_));
  AOI21_X1   g14663(.A1(new_n15686_), .A2(new_n15680_), .B(new_n6863_), .ZN(new_n15687_));
  AOI21_X1   g14664(.A1(new_n6845_), .A2(new_n6847_), .B(new_n6673_), .ZN(new_n15688_));
  AOI21_X1   g14665(.A1(new_n15688_), .A2(new_n15679_), .B(new_n6848_), .ZN(new_n15689_));
  NOR2_X1    g14666(.A1(new_n15689_), .A2(new_n15687_), .ZN(new_n15690_));
  OAI21_X1   g14667(.A1(new_n6884_), .A2(new_n6897_), .B(new_n15690_), .ZN(new_n15691_));
  INV_X1     g14668(.I(new_n15687_), .ZN(new_n15692_));
  NAND2_X1   g14669(.A1(new_n6845_), .A2(new_n6847_), .ZN(new_n15693_));
  NAND2_X1   g14670(.A1(new_n6839_), .A2(new_n15693_), .ZN(new_n15694_));
  OAI21_X1   g14671(.A1(new_n15694_), .A2(new_n6844_), .B(new_n6851_), .ZN(new_n15695_));
  NAND2_X1   g14672(.A1(new_n15692_), .A2(new_n15695_), .ZN(new_n15696_));
  NAND3_X1   g14673(.A1(new_n6886_), .A2(new_n15696_), .A3(new_n6838_), .ZN(new_n15697_));
  AOI21_X1   g14674(.A1(new_n15691_), .A2(new_n15697_), .B(new_n15684_), .ZN(new_n15698_));
  INV_X1     g14675(.I(new_n15684_), .ZN(new_n15699_));
  AOI21_X1   g14676(.A1(new_n6886_), .A2(new_n6838_), .B(new_n15696_), .ZN(new_n15700_));
  NOR3_X1    g14677(.A1(new_n6884_), .A2(new_n6897_), .A3(new_n15690_), .ZN(new_n15701_));
  NOR3_X1    g14678(.A1(new_n15701_), .A2(new_n15700_), .A3(new_n15699_), .ZN(new_n15702_));
  AOI21_X1   g14679(.A1(new_n6829_), .A2(new_n6727_), .B(new_n6828_), .ZN(new_n15703_));
  INV_X1     g14680(.I(new_n15703_), .ZN(new_n15704_));
  NOR3_X1    g14681(.A1(new_n6829_), .A2(new_n6727_), .A3(new_n6828_), .ZN(new_n15705_));
  NAND4_X1   g14682(.A1(new_n15705_), .A2(new_n6795_), .A3(new_n6802_), .A4(new_n6804_), .ZN(new_n15706_));
  NOR2_X1    g14683(.A1(new_n15706_), .A2(new_n15704_), .ZN(new_n15707_));
  NOR2_X1    g14684(.A1(new_n6805_), .A2(new_n6814_), .ZN(new_n15708_));
  INV_X1     g14685(.I(new_n6810_), .ZN(new_n15709_));
  NAND2_X1   g14686(.A1(new_n15709_), .A2(new_n6808_), .ZN(new_n15710_));
  NOR2_X1    g14687(.A1(new_n15709_), .A2(new_n6808_), .ZN(new_n15711_));
  NOR2_X1    g14688(.A1(new_n6727_), .A2(new_n15711_), .ZN(new_n15712_));
  NAND2_X1   g14689(.A1(new_n15712_), .A2(new_n6813_), .ZN(new_n15713_));
  INV_X1     g14690(.I(new_n6801_), .ZN(new_n15714_));
  NAND2_X1   g14691(.A1(new_n15714_), .A2(new_n6798_), .ZN(new_n15715_));
  NAND3_X1   g14692(.A1(new_n6801_), .A2(new_n6732_), .A3(new_n6797_), .ZN(new_n15716_));
  NAND4_X1   g14693(.A1(new_n6825_), .A2(new_n6781_), .A3(new_n6795_), .A4(new_n15716_), .ZN(new_n15717_));
  AOI22_X1   g14694(.A1(new_n15713_), .A2(new_n15710_), .B1(new_n15717_), .B2(new_n15715_), .ZN(new_n15718_));
  OAI21_X1   g14695(.A1(new_n6792_), .A2(new_n15708_), .B(new_n15718_), .ZN(new_n15719_));
  INV_X1     g14696(.I(new_n15710_), .ZN(new_n15720_));
  NOR2_X1    g14697(.A1(new_n6721_), .A2(new_n6694_), .ZN(new_n15721_));
  NOR4_X1    g14698(.A1(new_n15721_), .A2(new_n6722_), .A3(new_n6727_), .A4(new_n15711_), .ZN(new_n15722_));
  INV_X1     g14699(.I(new_n15715_), .ZN(new_n15723_));
  INV_X1     g14700(.I(new_n15716_), .ZN(new_n15724_));
  NOR4_X1    g14701(.A1(new_n6803_), .A2(new_n6757_), .A3(new_n6823_), .A4(new_n15724_), .ZN(new_n15725_));
  OAI22_X1   g14702(.A1(new_n15722_), .A2(new_n15720_), .B1(new_n15725_), .B2(new_n15723_), .ZN(new_n15726_));
  NAND3_X1   g14703(.A1(new_n6820_), .A2(new_n6831_), .A3(new_n15726_), .ZN(new_n15727_));
  AOI21_X1   g14704(.A1(new_n15719_), .A2(new_n15727_), .B(new_n15707_), .ZN(new_n15728_));
  NAND3_X1   g14705(.A1(new_n6813_), .A2(new_n6811_), .A3(new_n6770_), .ZN(new_n15729_));
  NOR4_X1    g14706(.A1(new_n15729_), .A2(new_n6823_), .A3(new_n6824_), .A4(new_n6826_), .ZN(new_n15730_));
  NAND2_X1   g14707(.A1(new_n15730_), .A2(new_n15703_), .ZN(new_n15731_));
  AOI21_X1   g14708(.A1(new_n6820_), .A2(new_n6831_), .B(new_n15726_), .ZN(new_n15732_));
  NOR3_X1    g14709(.A1(new_n6792_), .A2(new_n15718_), .A3(new_n15708_), .ZN(new_n15733_));
  NOR3_X1    g14710(.A1(new_n15732_), .A2(new_n15733_), .A3(new_n15731_), .ZN(new_n15734_));
  NOR2_X1    g14711(.A1(new_n15728_), .A2(new_n15734_), .ZN(new_n15735_));
  NOR3_X1    g14712(.A1(new_n15735_), .A2(new_n15702_), .A3(new_n15698_), .ZN(new_n15736_));
  OAI21_X1   g14713(.A1(new_n15701_), .A2(new_n15700_), .B(new_n15699_), .ZN(new_n15737_));
  NAND3_X1   g14714(.A1(new_n15691_), .A2(new_n15697_), .A3(new_n15684_), .ZN(new_n15738_));
  OAI21_X1   g14715(.A1(new_n15732_), .A2(new_n15733_), .B(new_n15731_), .ZN(new_n15739_));
  NAND3_X1   g14716(.A1(new_n15719_), .A2(new_n15727_), .A3(new_n15707_), .ZN(new_n15740_));
  NAND2_X1   g14717(.A1(new_n15739_), .A2(new_n15740_), .ZN(new_n15741_));
  AOI21_X1   g14718(.A1(new_n15737_), .A2(new_n15738_), .B(new_n15741_), .ZN(new_n15742_));
  NOR2_X1    g14719(.A1(new_n15742_), .A2(new_n15736_), .ZN(new_n15743_));
  NOR2_X1    g14720(.A1(new_n15743_), .A2(new_n15675_), .ZN(new_n15744_));
  NOR2_X1    g14721(.A1(new_n6888_), .A2(new_n6892_), .ZN(new_n15745_));
  OAI21_X1   g14722(.A1(new_n15745_), .A2(new_n6788_), .B(new_n6899_), .ZN(new_n15746_));
  OAI21_X1   g14723(.A1(new_n15698_), .A2(new_n15702_), .B(new_n15741_), .ZN(new_n15747_));
  NAND3_X1   g14724(.A1(new_n15735_), .A2(new_n15737_), .A3(new_n15738_), .ZN(new_n15748_));
  AOI21_X1   g14725(.A1(new_n15747_), .A2(new_n15748_), .B(new_n15746_), .ZN(new_n15749_));
  NOR2_X1    g14726(.A1(new_n15749_), .A2(new_n15744_), .ZN(new_n15750_));
  NOR2_X1    g14727(.A1(new_n15672_), .A2(new_n15750_), .ZN(new_n15751_));
  NOR2_X1    g14728(.A1(new_n8118_), .A2(new_n8121_), .ZN(new_n15752_));
  OAI21_X1   g14729(.A1(new_n15752_), .A2(new_n8112_), .B(new_n7857_), .ZN(new_n15753_));
  NAND2_X1   g14730(.A1(new_n6895_), .A2(new_n6898_), .ZN(new_n15754_));
  AOI21_X1   g14731(.A1(new_n15754_), .A2(new_n6834_), .B(new_n6788_), .ZN(new_n15755_));
  OAI22_X1   g14732(.A1(new_n15674_), .A2(new_n15755_), .B1(new_n15742_), .B2(new_n15736_), .ZN(new_n15756_));
  NAND2_X1   g14733(.A1(new_n15747_), .A2(new_n15748_), .ZN(new_n15757_));
  NAND2_X1   g14734(.A1(new_n15757_), .A2(new_n15675_), .ZN(new_n15758_));
  NAND2_X1   g14735(.A1(new_n15758_), .A2(new_n15756_), .ZN(new_n15759_));
  AOI21_X1   g14736(.A1(new_n8123_), .A2(new_n15753_), .B(new_n15759_), .ZN(new_n15760_));
  OAI21_X1   g14737(.A1(new_n15751_), .A2(new_n15760_), .B(new_n15671_), .ZN(new_n15761_));
  AOI21_X1   g14738(.A1(new_n15662_), .A2(new_n15659_), .B(new_n15669_), .ZN(new_n15762_));
  NOR3_X1    g14739(.A1(new_n15581_), .A2(new_n15585_), .A3(new_n15655_), .ZN(new_n15763_));
  NOR2_X1    g14740(.A1(new_n15763_), .A2(new_n15762_), .ZN(new_n15764_));
  AOI21_X1   g14741(.A1(new_n7857_), .A2(new_n8122_), .B(new_n8130_), .ZN(new_n15765_));
  NOR2_X1    g14742(.A1(new_n15765_), .A2(new_n15750_), .ZN(new_n15766_));
  NOR2_X1    g14743(.A1(new_n15672_), .A2(new_n15759_), .ZN(new_n15767_));
  OAI21_X1   g14744(.A1(new_n15766_), .A2(new_n15767_), .B(new_n15764_), .ZN(new_n15768_));
  NAND2_X1   g14745(.A1(new_n15768_), .A2(new_n15761_), .ZN(new_n15769_));
  NAND2_X1   g14746(.A1(new_n8178_), .A2(new_n8175_), .ZN(new_n15770_));
  NAND2_X1   g14747(.A1(new_n8194_), .A2(new_n15770_), .ZN(new_n15771_));
  NOR2_X1    g14748(.A1(new_n8170_), .A2(new_n8154_), .ZN(new_n15772_));
  NAND3_X1   g14749(.A1(new_n8190_), .A2(new_n8193_), .A3(new_n15772_), .ZN(new_n15773_));
  AOI21_X1   g14750(.A1(new_n8125_), .A2(new_n8132_), .B(new_n8179_), .ZN(new_n15774_));
  AOI21_X1   g14751(.A1(new_n8128_), .A2(new_n8131_), .B(new_n6902_), .ZN(new_n15775_));
  NOR3_X1    g14752(.A1(new_n8114_), .A2(new_n6903_), .A3(new_n8124_), .ZN(new_n15776_));
  NOR3_X1    g14753(.A1(new_n15776_), .A2(new_n15775_), .A3(new_n8173_), .ZN(new_n15777_));
  OAI21_X1   g14754(.A1(new_n15777_), .A2(new_n15774_), .B(new_n15773_), .ZN(new_n15778_));
  NAND2_X1   g14755(.A1(new_n8114_), .A2(new_n8179_), .ZN(new_n15779_));
  NOR2_X1    g14756(.A1(new_n8114_), .A2(new_n8179_), .ZN(new_n15780_));
  NAND2_X1   g14757(.A1(new_n8124_), .A2(new_n6902_), .ZN(new_n15781_));
  OAI21_X1   g14758(.A1(new_n15780_), .A2(new_n15781_), .B(new_n15779_), .ZN(new_n15782_));
  NAND3_X1   g14759(.A1(new_n15778_), .A2(new_n15771_), .A3(new_n15782_), .ZN(new_n15783_));
  NOR2_X1    g14760(.A1(new_n6273_), .A2(new_n15772_), .ZN(new_n15784_));
  NOR3_X1    g14761(.A1(new_n6269_), .A2(new_n6272_), .A3(new_n15770_), .ZN(new_n15785_));
  OAI21_X1   g14762(.A1(new_n15776_), .A2(new_n15775_), .B(new_n8173_), .ZN(new_n15786_));
  NAND3_X1   g14763(.A1(new_n8125_), .A2(new_n8132_), .A3(new_n8179_), .ZN(new_n15787_));
  AOI21_X1   g14764(.A1(new_n15786_), .A2(new_n15787_), .B(new_n15785_), .ZN(new_n15788_));
  NOR2_X1    g14765(.A1(new_n8128_), .A2(new_n8173_), .ZN(new_n15789_));
  NAND2_X1   g14766(.A1(new_n8128_), .A2(new_n8173_), .ZN(new_n15790_));
  NOR2_X1    g14767(.A1(new_n6903_), .A2(new_n8131_), .ZN(new_n15791_));
  AOI21_X1   g14768(.A1(new_n15790_), .A2(new_n15791_), .B(new_n15789_), .ZN(new_n15792_));
  OAI21_X1   g14769(.A1(new_n15788_), .A2(new_n15784_), .B(new_n15792_), .ZN(new_n15793_));
  AOI21_X1   g14770(.A1(new_n15783_), .A2(new_n15793_), .B(new_n15769_), .ZN(new_n15794_));
  INV_X1     g14771(.I(new_n15769_), .ZN(new_n15795_));
  NOR3_X1    g14772(.A1(new_n15788_), .A2(new_n15784_), .A3(new_n15792_), .ZN(new_n15796_));
  AOI21_X1   g14773(.A1(new_n15778_), .A2(new_n15771_), .B(new_n15782_), .ZN(new_n15797_));
  NOR3_X1    g14774(.A1(new_n15797_), .A2(new_n15796_), .A3(new_n15795_), .ZN(new_n15798_));
  OAI21_X1   g14775(.A1(new_n15794_), .A2(new_n15798_), .B(new_n15508_), .ZN(new_n15799_));
  INV_X1     g14776(.I(new_n15508_), .ZN(new_n15800_));
  OAI21_X1   g14777(.A1(new_n15797_), .A2(new_n15796_), .B(new_n15795_), .ZN(new_n15801_));
  NAND3_X1   g14778(.A1(new_n15783_), .A2(new_n15793_), .A3(new_n15769_), .ZN(new_n15802_));
  NAND3_X1   g14779(.A1(new_n15801_), .A2(new_n15802_), .A3(new_n15800_), .ZN(new_n15803_));
  NAND2_X1   g14780(.A1(new_n15799_), .A2(new_n15803_), .ZN(new_n15804_));
  NAND2_X1   g14781(.A1(new_n15804_), .A2(new_n15345_), .ZN(new_n15805_));
  NOR3_X1    g14782(.A1(new_n15332_), .A2(new_n15339_), .A3(new_n15342_), .ZN(new_n15806_));
  NOR2_X1    g14783(.A1(new_n15339_), .A2(new_n15342_), .ZN(new_n15807_));
  NOR2_X1    g14784(.A1(new_n15807_), .A2(new_n15323_), .ZN(new_n15808_));
  OAI21_X1   g14785(.A1(new_n15808_), .A2(new_n15806_), .B(new_n15335_), .ZN(new_n15809_));
  NOR4_X1    g14786(.A1(new_n15339_), .A2(new_n15342_), .A3(new_n15328_), .A4(new_n15331_), .ZN(new_n15810_));
  AOI22_X1   g14787(.A1(new_n14963_), .A2(new_n14967_), .B1(new_n15318_), .B2(new_n15322_), .ZN(new_n15811_));
  OAI21_X1   g14788(.A1(new_n15811_), .A2(new_n15810_), .B(new_n14614_), .ZN(new_n15812_));
  NAND2_X1   g14789(.A1(new_n15809_), .A2(new_n15812_), .ZN(new_n15813_));
  NAND3_X1   g14790(.A1(new_n15813_), .A2(new_n15799_), .A3(new_n15803_), .ZN(new_n15814_));
  AOI21_X1   g14791(.A1(new_n15805_), .A2(new_n15814_), .B(new_n14613_), .ZN(new_n15815_));
  NAND3_X1   g14792(.A1(new_n15345_), .A2(new_n15799_), .A3(new_n15803_), .ZN(new_n15816_));
  NAND2_X1   g14793(.A1(new_n15804_), .A2(new_n15813_), .ZN(new_n15817_));
  AOI21_X1   g14794(.A1(new_n15817_), .A2(new_n15816_), .B(new_n14612_), .ZN(new_n15818_));
  OAI21_X1   g14795(.A1(new_n15818_), .A2(new_n15815_), .B(new_n14610_), .ZN(new_n15819_));
  NOR2_X1    g14796(.A1(new_n14599_), .A2(new_n14607_), .ZN(new_n15820_));
  OAI21_X1   g14797(.A1(new_n15820_), .A2(new_n14593_), .B(new_n14598_), .ZN(new_n15821_));
  NOR2_X1    g14798(.A1(new_n14607_), .A2(new_n14592_), .ZN(new_n15822_));
  NOR2_X1    g14799(.A1(new_n14599_), .A2(new_n14591_), .ZN(new_n15823_));
  OAI21_X1   g14800(.A1(new_n15823_), .A2(new_n15822_), .B(new_n14270_), .ZN(new_n15824_));
  NAND2_X1   g14801(.A1(new_n15821_), .A2(new_n15824_), .ZN(new_n15825_));
  AOI21_X1   g14802(.A1(new_n15799_), .A2(new_n15803_), .B(new_n15813_), .ZN(new_n15826_));
  AOI21_X1   g14803(.A1(new_n15801_), .A2(new_n15802_), .B(new_n15800_), .ZN(new_n15827_));
  NOR3_X1    g14804(.A1(new_n15794_), .A2(new_n15798_), .A3(new_n15508_), .ZN(new_n15828_));
  NOR3_X1    g14805(.A1(new_n15345_), .A2(new_n15827_), .A3(new_n15828_), .ZN(new_n15829_));
  OAI21_X1   g14806(.A1(new_n15826_), .A2(new_n15829_), .B(new_n14612_), .ZN(new_n15830_));
  NOR3_X1    g14807(.A1(new_n15813_), .A2(new_n15827_), .A3(new_n15828_), .ZN(new_n15831_));
  AOI22_X1   g14808(.A1(new_n15799_), .A2(new_n15803_), .B1(new_n15809_), .B2(new_n15812_), .ZN(new_n15832_));
  OAI21_X1   g14809(.A1(new_n15831_), .A2(new_n15832_), .B(new_n14613_), .ZN(new_n15833_));
  NAND3_X1   g14810(.A1(new_n15830_), .A2(new_n15833_), .A3(new_n15825_), .ZN(new_n15834_));
  NAND3_X1   g14811(.A1(new_n15819_), .A2(new_n15834_), .A3(new_n13986_), .ZN(new_n15835_));
  AOI21_X1   g14812(.A1(new_n13911_), .A2(new_n13921_), .B(new_n8198_), .ZN(new_n15836_));
  NOR3_X1    g14813(.A1(new_n13958_), .A2(new_n13929_), .A3(new_n13961_), .ZN(new_n15837_));
  OAI21_X1   g14814(.A1(new_n15837_), .A2(new_n15836_), .B(new_n13965_), .ZN(new_n15838_));
  AOI21_X1   g14815(.A1(new_n13911_), .A2(new_n13921_), .B(new_n13929_), .ZN(new_n15839_));
  OAI21_X1   g14816(.A1(new_n15839_), .A2(new_n14611_), .B(new_n12556_), .ZN(new_n15840_));
  NAND2_X1   g14817(.A1(new_n15840_), .A2(new_n15838_), .ZN(new_n15841_));
  NOR2_X1    g14818(.A1(new_n15837_), .A2(new_n15836_), .ZN(new_n15842_));
  INV_X1     g14819(.I(new_n13984_), .ZN(new_n15843_));
  OAI21_X1   g14820(.A1(new_n15842_), .A2(new_n15843_), .B(new_n5352_), .ZN(new_n15844_));
  NAND2_X1   g14821(.A1(new_n15844_), .A2(new_n15841_), .ZN(new_n15845_));
  NAND2_X1   g14822(.A1(new_n15819_), .A2(new_n15834_), .ZN(new_n15846_));
  NAND2_X1   g14823(.A1(new_n15846_), .A2(new_n15845_), .ZN(new_n15847_));
  NAND2_X1   g14824(.A1(new_n15847_), .A2(new_n15835_), .ZN(new_n15848_));
  NAND2_X1   g14825(.A1(new_n15848_), .A2(new_n13955_), .ZN(new_n15849_));
  NAND2_X1   g14826(.A1(new_n15805_), .A2(new_n15814_), .ZN(new_n15850_));
  NAND3_X1   g14827(.A1(new_n15850_), .A2(new_n13986_), .A3(new_n14612_), .ZN(new_n15851_));
  NOR2_X1    g14828(.A1(new_n15815_), .A2(new_n13986_), .ZN(new_n15852_));
  NAND2_X1   g14829(.A1(new_n15818_), .A2(new_n15825_), .ZN(new_n15853_));
  OAI21_X1   g14830(.A1(new_n15852_), .A2(new_n15853_), .B(new_n15851_), .ZN(new_n15854_));
  NAND2_X1   g14831(.A1(new_n15505_), .A2(new_n15504_), .ZN(new_n15855_));
  NAND2_X1   g14832(.A1(new_n15855_), .A2(new_n15506_), .ZN(new_n15856_));
  INV_X1     g14833(.I(new_n15436_), .ZN(new_n15857_));
  XOR2_X1    g14834(.A1(new_n15459_), .A2(new_n15464_), .Z(new_n15858_));
  NOR2_X1    g14835(.A1(new_n15428_), .A2(new_n15425_), .ZN(new_n15859_));
  XOR2_X1    g14836(.A1(new_n15859_), .A2(new_n15433_), .Z(new_n15860_));
  NOR2_X1    g14837(.A1(new_n15860_), .A2(new_n15858_), .ZN(new_n15861_));
  NAND4_X1   g14838(.A1(new_n15861_), .A2(new_n15441_), .A3(new_n15857_), .A4(new_n15449_), .ZN(new_n15862_));
  AOI21_X1   g14839(.A1(new_n6109_), .A2(new_n15450_), .B(new_n15449_), .ZN(new_n15863_));
  INV_X1     g14840(.I(new_n15863_), .ZN(new_n15864_));
  OAI21_X1   g14841(.A1(new_n15441_), .A2(new_n15857_), .B(new_n15864_), .ZN(new_n15865_));
  NOR3_X1    g14842(.A1(new_n15862_), .A2(new_n15865_), .A3(new_n15451_), .ZN(new_n15866_));
  INV_X1     g14843(.I(new_n15866_), .ZN(new_n15867_));
  NOR2_X1    g14844(.A1(new_n15484_), .A2(new_n15418_), .ZN(new_n15868_));
  NOR2_X1    g14845(.A1(new_n15857_), .A2(new_n15441_), .ZN(new_n15869_));
  NAND2_X1   g14846(.A1(new_n15859_), .A2(new_n15437_), .ZN(new_n15870_));
  NAND2_X1   g14847(.A1(new_n15869_), .A2(new_n15870_), .ZN(new_n15871_));
  NAND2_X1   g14848(.A1(new_n15459_), .A2(new_n15454_), .ZN(new_n15872_));
  NAND2_X1   g14849(.A1(new_n15863_), .A2(new_n15872_), .ZN(new_n15873_));
  AOI22_X1   g14850(.A1(new_n15871_), .A2(new_n15434_), .B1(new_n15873_), .B2(new_n15465_), .ZN(new_n15874_));
  INV_X1     g14851(.I(new_n15874_), .ZN(new_n15875_));
  NOR2_X1    g14852(.A1(new_n15868_), .A2(new_n15875_), .ZN(new_n15876_));
  NAND2_X1   g14853(.A1(new_n15499_), .A2(new_n15482_), .ZN(new_n15877_));
  NOR2_X1    g14854(.A1(new_n15877_), .A2(new_n15874_), .ZN(new_n15878_));
  OAI21_X1   g14855(.A1(new_n15876_), .A2(new_n15878_), .B(new_n15867_), .ZN(new_n15879_));
  NAND2_X1   g14856(.A1(new_n15877_), .A2(new_n15874_), .ZN(new_n15880_));
  NAND2_X1   g14857(.A1(new_n15868_), .A2(new_n15875_), .ZN(new_n15881_));
  NAND3_X1   g14858(.A1(new_n15881_), .A2(new_n15880_), .A3(new_n15866_), .ZN(new_n15882_));
  NAND2_X1   g14859(.A1(new_n15879_), .A2(new_n15882_), .ZN(new_n15883_));
  NOR2_X1    g14860(.A1(new_n6176_), .A2(new_n6135_), .ZN(new_n15884_));
  INV_X1     g14861(.I(new_n15884_), .ZN(new_n15885_));
  NOR2_X1    g14862(.A1(new_n6224_), .A2(new_n6241_), .ZN(new_n15886_));
  NAND2_X1   g14863(.A1(new_n15391_), .A2(new_n15379_), .ZN(new_n15887_));
  NOR2_X1    g14864(.A1(new_n15388_), .A2(new_n15385_), .ZN(new_n15888_));
  XOR2_X1    g14865(.A1(new_n15887_), .A2(new_n15888_), .Z(new_n15889_));
  XNOR2_X1   g14866(.A1(new_n15363_), .A2(new_n15364_), .ZN(new_n15890_));
  NOR2_X1    g14867(.A1(new_n15890_), .A2(new_n15889_), .ZN(new_n15891_));
  NAND4_X1   g14868(.A1(new_n15891_), .A2(new_n15352_), .A3(new_n15886_), .A4(new_n15399_), .ZN(new_n15892_));
  OAI21_X1   g14869(.A1(new_n6224_), .A2(new_n6241_), .B(new_n15370_), .ZN(new_n15893_));
  OAI21_X1   g14870(.A1(new_n15399_), .A2(new_n15884_), .B(new_n15893_), .ZN(new_n15894_));
  NOR3_X1    g14871(.A1(new_n15892_), .A2(new_n15894_), .A3(new_n15885_), .ZN(new_n15895_));
  INV_X1     g14872(.I(new_n15895_), .ZN(new_n15896_));
  NOR2_X1    g14873(.A1(new_n15492_), .A2(new_n15413_), .ZN(new_n15897_));
  NOR2_X1    g14874(.A1(new_n15363_), .A2(new_n15364_), .ZN(new_n15898_));
  OAI21_X1   g14875(.A1(new_n15893_), .A2(new_n15898_), .B(new_n15365_), .ZN(new_n15899_));
  NOR2_X1    g14876(.A1(new_n15399_), .A2(new_n15884_), .ZN(new_n15900_));
  INV_X1     g14877(.I(new_n15900_), .ZN(new_n15901_));
  INV_X1     g14878(.I(new_n15888_), .ZN(new_n15902_));
  NOR2_X1    g14879(.A1(new_n15902_), .A2(new_n15887_), .ZN(new_n15903_));
  OAI21_X1   g14880(.A1(new_n15901_), .A2(new_n15903_), .B(new_n15389_), .ZN(new_n15904_));
  NAND2_X1   g14881(.A1(new_n15904_), .A2(new_n15899_), .ZN(new_n15905_));
  NOR2_X1    g14882(.A1(new_n15897_), .A2(new_n15905_), .ZN(new_n15906_));
  NAND2_X1   g14883(.A1(new_n15415_), .A2(new_n15347_), .ZN(new_n15907_));
  AOI21_X1   g14884(.A1(new_n15899_), .A2(new_n15904_), .B(new_n15907_), .ZN(new_n15908_));
  OAI21_X1   g14885(.A1(new_n15908_), .A2(new_n15906_), .B(new_n15896_), .ZN(new_n15909_));
  NAND3_X1   g14886(.A1(new_n15907_), .A2(new_n15899_), .A3(new_n15904_), .ZN(new_n15910_));
  NAND2_X1   g14887(.A1(new_n15897_), .A2(new_n15905_), .ZN(new_n15911_));
  NAND3_X1   g14888(.A1(new_n15910_), .A2(new_n15911_), .A3(new_n15895_), .ZN(new_n15912_));
  AOI21_X1   g14889(.A1(new_n15909_), .A2(new_n15912_), .B(new_n15883_), .ZN(new_n15913_));
  NAND2_X1   g14890(.A1(new_n15909_), .A2(new_n15912_), .ZN(new_n15914_));
  AOI21_X1   g14891(.A1(new_n15879_), .A2(new_n15882_), .B(new_n15914_), .ZN(new_n15915_));
  OAI21_X1   g14892(.A1(new_n15915_), .A2(new_n15913_), .B(new_n15856_), .ZN(new_n15916_));
  XOR2_X1    g14893(.A1(new_n15914_), .A2(new_n15883_), .Z(new_n15917_));
  OAI21_X1   g14894(.A1(new_n15917_), .A2(new_n15856_), .B(new_n15916_), .ZN(new_n15918_));
  INV_X1     g14895(.I(new_n15918_), .ZN(new_n15919_));
  NOR2_X1    g14896(.A1(new_n6884_), .A2(new_n6897_), .ZN(new_n15920_));
  INV_X1     g14897(.I(new_n15920_), .ZN(new_n15921_));
  NOR2_X1    g14898(.A1(new_n6792_), .A2(new_n15708_), .ZN(new_n15922_));
  NOR2_X1    g14899(.A1(new_n15707_), .A2(new_n15922_), .ZN(new_n15923_));
  NOR2_X1    g14900(.A1(new_n15722_), .A2(new_n15720_), .ZN(new_n15924_));
  NOR2_X1    g14901(.A1(new_n15725_), .A2(new_n15723_), .ZN(new_n15925_));
  XNOR2_X1   g14902(.A1(new_n15924_), .A2(new_n15925_), .ZN(new_n15926_));
  XNOR2_X1   g14903(.A1(new_n15689_), .A2(new_n15687_), .ZN(new_n15927_));
  NOR4_X1    g14904(.A1(new_n15926_), .A2(new_n15927_), .A3(new_n15699_), .A4(new_n15731_), .ZN(new_n15928_));
  INV_X1     g14905(.I(new_n15928_), .ZN(new_n15929_));
  OAI21_X1   g14906(.A1(new_n15920_), .A2(new_n15684_), .B(new_n15922_), .ZN(new_n15930_));
  NOR4_X1    g14907(.A1(new_n15929_), .A2(new_n15921_), .A3(new_n15923_), .A4(new_n15930_), .ZN(new_n15931_));
  INV_X1     g14908(.I(new_n15748_), .ZN(new_n15932_));
  NOR2_X1    g14909(.A1(new_n15746_), .A2(new_n15932_), .ZN(new_n15933_));
  NOR2_X1    g14910(.A1(new_n15692_), .A2(new_n15695_), .ZN(new_n15934_));
  AOI21_X1   g14911(.A1(new_n15684_), .A2(new_n15692_), .B(new_n15934_), .ZN(new_n15935_));
  OAI21_X1   g14912(.A1(new_n15921_), .A2(new_n15689_), .B(new_n15935_), .ZN(new_n15936_));
  INV_X1     g14913(.I(new_n15923_), .ZN(new_n15937_));
  NOR4_X1    g14914(.A1(new_n15722_), .A2(new_n15725_), .A3(new_n15720_), .A4(new_n15723_), .ZN(new_n15938_));
  OAI21_X1   g14915(.A1(new_n15937_), .A2(new_n15938_), .B(new_n15726_), .ZN(new_n15939_));
  INV_X1     g14916(.I(new_n15939_), .ZN(new_n15940_));
  NOR2_X1    g14917(.A1(new_n15940_), .A2(new_n15936_), .ZN(new_n15941_));
  INV_X1     g14918(.I(new_n15941_), .ZN(new_n15942_));
  NOR2_X1    g14919(.A1(new_n15933_), .A2(new_n15942_), .ZN(new_n15943_));
  INV_X1     g14920(.I(new_n15933_), .ZN(new_n15944_));
  NOR2_X1    g14921(.A1(new_n15944_), .A2(new_n15941_), .ZN(new_n15945_));
  NOR2_X1    g14922(.A1(new_n15945_), .A2(new_n15943_), .ZN(new_n15946_));
  NOR2_X1    g14923(.A1(new_n15946_), .A2(new_n15931_), .ZN(new_n15947_));
  INV_X1     g14924(.I(new_n15931_), .ZN(new_n15948_));
  NOR3_X1    g14925(.A1(new_n15945_), .A2(new_n15948_), .A3(new_n15943_), .ZN(new_n15949_));
  NOR2_X1    g14926(.A1(new_n15947_), .A2(new_n15949_), .ZN(new_n15950_));
  OAI21_X1   g14927(.A1(new_n15765_), .A2(new_n15762_), .B(new_n15670_), .ZN(new_n15951_));
  INV_X1     g14928(.I(new_n15951_), .ZN(new_n15952_));
  AOI21_X1   g14929(.A1(new_n15591_), .A2(new_n15666_), .B(new_n15653_), .ZN(new_n15953_));
  NOR2_X1    g14930(.A1(new_n8092_), .A2(new_n8103_), .ZN(new_n15954_));
  NOR2_X1    g14931(.A1(new_n15954_), .A2(new_n15618_), .ZN(new_n15955_));
  NAND2_X1   g14932(.A1(new_n8033_), .A2(new_n8013_), .ZN(new_n15956_));
  NAND2_X1   g14933(.A1(new_n8026_), .A2(new_n8018_), .ZN(new_n15957_));
  NAND3_X1   g14934(.A1(new_n15956_), .A2(new_n15957_), .A3(new_n15599_), .ZN(new_n15958_));
  INV_X1     g14935(.I(new_n15958_), .ZN(new_n15959_));
  XOR2_X1    g14936(.A1(new_n15623_), .A2(new_n15626_), .Z(new_n15960_));
  NAND3_X1   g14937(.A1(new_n15959_), .A2(new_n15960_), .A3(new_n15627_), .ZN(new_n15961_));
  NAND2_X1   g14938(.A1(new_n15623_), .A2(new_n15626_), .ZN(new_n15962_));
  AOI21_X1   g14939(.A1(new_n15961_), .A2(new_n15962_), .B(new_n15955_), .ZN(new_n15963_));
  NAND3_X1   g14940(.A1(new_n15961_), .A2(new_n15955_), .A3(new_n15962_), .ZN(new_n15964_));
  INV_X1     g14941(.I(new_n15964_), .ZN(new_n15965_));
  NOR2_X1    g14942(.A1(new_n15965_), .A2(new_n15963_), .ZN(new_n15966_));
  INV_X1     g14943(.I(new_n15966_), .ZN(new_n15967_));
  NOR2_X1    g14944(.A1(new_n15643_), .A2(new_n15642_), .ZN(new_n15968_));
  OAI21_X1   g14945(.A1(new_n15966_), .A2(new_n15968_), .B(new_n15641_), .ZN(new_n15969_));
  AOI21_X1   g14946(.A1(new_n15966_), .A2(new_n15968_), .B(new_n15651_), .ZN(new_n15970_));
  AOI22_X1   g14947(.A1(new_n15970_), .A2(new_n15969_), .B1(new_n15953_), .B2(new_n15967_), .ZN(new_n15971_));
  NAND2_X1   g14948(.A1(new_n15563_), .A2(new_n15564_), .ZN(new_n15972_));
  NOR2_X1    g14949(.A1(new_n15972_), .A2(new_n15568_), .ZN(new_n15973_));
  XOR2_X1    g14950(.A1(new_n15557_), .A2(new_n15560_), .Z(new_n15974_));
  NAND2_X1   g14951(.A1(new_n7987_), .A2(new_n7939_), .ZN(new_n15975_));
  XNOR2_X1   g14952(.A1(new_n15533_), .A2(new_n15532_), .ZN(new_n15976_));
  NOR4_X1    g14953(.A1(new_n15976_), .A2(new_n15975_), .A3(new_n15551_), .A4(new_n15522_), .ZN(new_n15977_));
  NAND2_X1   g14954(.A1(new_n15975_), .A2(new_n15522_), .ZN(new_n15978_));
  NAND4_X1   g14955(.A1(new_n15977_), .A2(new_n15972_), .A3(new_n15974_), .A4(new_n15978_), .ZN(new_n15979_));
  NOR2_X1    g14956(.A1(new_n15979_), .A2(new_n15973_), .ZN(new_n15980_));
  INV_X1     g14957(.I(new_n15980_), .ZN(new_n15981_));
  INV_X1     g14958(.I(new_n15584_), .ZN(new_n15982_));
  NOR2_X1    g14959(.A1(new_n15982_), .A2(new_n15582_), .ZN(new_n15983_));
  NAND2_X1   g14960(.A1(new_n15523_), .A2(new_n15532_), .ZN(new_n15984_));
  NAND3_X1   g14961(.A1(new_n7987_), .A2(new_n7939_), .A3(new_n15533_), .ZN(new_n15985_));
  NAND2_X1   g14962(.A1(new_n15984_), .A2(new_n15985_), .ZN(new_n15986_));
  NOR2_X1    g14963(.A1(new_n15533_), .A2(new_n15532_), .ZN(new_n15987_));
  NAND2_X1   g14964(.A1(new_n15568_), .A2(new_n15557_), .ZN(new_n15988_));
  NAND2_X1   g14965(.A1(new_n15972_), .A2(new_n15560_), .ZN(new_n15989_));
  NAND2_X1   g14966(.A1(new_n15989_), .A2(new_n15988_), .ZN(new_n15990_));
  NOR2_X1    g14967(.A1(new_n15557_), .A2(new_n15560_), .ZN(new_n15991_));
  NOR4_X1    g14968(.A1(new_n15990_), .A2(new_n15986_), .A3(new_n15987_), .A4(new_n15991_), .ZN(new_n15992_));
  INV_X1     g14969(.I(new_n15992_), .ZN(new_n15993_));
  NOR2_X1    g14970(.A1(new_n15983_), .A2(new_n15993_), .ZN(new_n15994_));
  NAND2_X1   g14971(.A1(new_n15660_), .A2(new_n15584_), .ZN(new_n15995_));
  NOR2_X1    g14972(.A1(new_n15995_), .A2(new_n15992_), .ZN(new_n15996_));
  OAI21_X1   g14973(.A1(new_n15996_), .A2(new_n15994_), .B(new_n15981_), .ZN(new_n15997_));
  NAND2_X1   g14974(.A1(new_n15995_), .A2(new_n15992_), .ZN(new_n15998_));
  NAND2_X1   g14975(.A1(new_n15983_), .A2(new_n15993_), .ZN(new_n15999_));
  NAND3_X1   g14976(.A1(new_n15998_), .A2(new_n15999_), .A3(new_n15980_), .ZN(new_n16000_));
  AOI21_X1   g14977(.A1(new_n15997_), .A2(new_n16000_), .B(new_n15971_), .ZN(new_n16001_));
  INV_X1     g14978(.I(new_n15971_), .ZN(new_n16002_));
  AOI21_X1   g14979(.A1(new_n15998_), .A2(new_n15999_), .B(new_n15980_), .ZN(new_n16003_));
  NOR3_X1    g14980(.A1(new_n15996_), .A2(new_n15994_), .A3(new_n15981_), .ZN(new_n16004_));
  NOR3_X1    g14981(.A1(new_n16002_), .A2(new_n16004_), .A3(new_n16003_), .ZN(new_n16005_));
  OAI21_X1   g14982(.A1(new_n16001_), .A2(new_n16005_), .B(new_n15952_), .ZN(new_n16006_));
  AOI21_X1   g14983(.A1(new_n16000_), .A2(new_n15997_), .B(new_n16002_), .ZN(new_n16007_));
  NOR3_X1    g14984(.A1(new_n16003_), .A2(new_n16004_), .A3(new_n15971_), .ZN(new_n16008_));
  OAI21_X1   g14985(.A1(new_n16007_), .A2(new_n16008_), .B(new_n15951_), .ZN(new_n16009_));
  NAND2_X1   g14986(.A1(new_n16006_), .A2(new_n16009_), .ZN(new_n16010_));
  NAND2_X1   g14987(.A1(new_n16010_), .A2(new_n15950_), .ZN(new_n16011_));
  INV_X1     g14988(.I(new_n15950_), .ZN(new_n16012_));
  NAND3_X1   g14989(.A1(new_n16012_), .A2(new_n16006_), .A3(new_n16009_), .ZN(new_n16013_));
  NAND2_X1   g14990(.A1(new_n16011_), .A2(new_n16013_), .ZN(new_n16014_));
  OAI22_X1   g14991(.A1(new_n15788_), .A2(new_n15784_), .B1(new_n15503_), .B2(new_n15507_), .ZN(new_n16015_));
  NAND3_X1   g14992(.A1(new_n15778_), .A2(new_n15508_), .A3(new_n15771_), .ZN(new_n16016_));
  NAND2_X1   g14993(.A1(new_n15769_), .A2(new_n15792_), .ZN(new_n16017_));
  NAND3_X1   g14994(.A1(new_n15782_), .A2(new_n15761_), .A3(new_n15768_), .ZN(new_n16018_));
  NAND2_X1   g14995(.A1(new_n16017_), .A2(new_n16018_), .ZN(new_n16019_));
  NAND2_X1   g14996(.A1(new_n16016_), .A2(new_n16019_), .ZN(new_n16020_));
  NOR2_X1    g14997(.A1(new_n15792_), .A2(new_n15750_), .ZN(new_n16021_));
  AOI21_X1   g14998(.A1(new_n15656_), .A2(new_n15670_), .B(new_n15672_), .ZN(new_n16022_));
  NOR3_X1    g14999(.A1(new_n15765_), .A2(new_n15762_), .A3(new_n15763_), .ZN(new_n16023_));
  NOR2_X1    g15000(.A1(new_n16022_), .A2(new_n16023_), .ZN(new_n16024_));
  AOI21_X1   g15001(.A1(new_n15792_), .A2(new_n15750_), .B(new_n16024_), .ZN(new_n16025_));
  NOR2_X1    g15002(.A1(new_n16025_), .A2(new_n16021_), .ZN(new_n16026_));
  INV_X1     g15003(.I(new_n16026_), .ZN(new_n16027_));
  NAND3_X1   g15004(.A1(new_n16020_), .A2(new_n16015_), .A3(new_n16027_), .ZN(new_n16028_));
  INV_X1     g15005(.I(new_n16015_), .ZN(new_n16029_));
  NOR2_X1    g15006(.A1(new_n15788_), .A2(new_n15784_), .ZN(new_n16030_));
  AOI22_X1   g15007(.A1(new_n16030_), .A2(new_n15508_), .B1(new_n16017_), .B2(new_n16018_), .ZN(new_n16031_));
  OAI21_X1   g15008(.A1(new_n16031_), .A2(new_n16029_), .B(new_n16026_), .ZN(new_n16032_));
  AOI21_X1   g15009(.A1(new_n16032_), .A2(new_n16028_), .B(new_n16014_), .ZN(new_n16033_));
  INV_X1     g15010(.I(new_n16014_), .ZN(new_n16034_));
  NOR3_X1    g15011(.A1(new_n16031_), .A2(new_n16029_), .A3(new_n16026_), .ZN(new_n16035_));
  AOI21_X1   g15012(.A1(new_n16020_), .A2(new_n16015_), .B(new_n16027_), .ZN(new_n16036_));
  NOR3_X1    g15013(.A1(new_n16035_), .A2(new_n16036_), .A3(new_n16034_), .ZN(new_n16037_));
  OAI21_X1   g15014(.A1(new_n16037_), .A2(new_n16033_), .B(new_n15919_), .ZN(new_n16038_));
  OAI21_X1   g15015(.A1(new_n16035_), .A2(new_n16036_), .B(new_n16034_), .ZN(new_n16039_));
  NAND3_X1   g15016(.A1(new_n16032_), .A2(new_n16028_), .A3(new_n16014_), .ZN(new_n16040_));
  NAND3_X1   g15017(.A1(new_n16039_), .A2(new_n16040_), .A3(new_n15918_), .ZN(new_n16041_));
  AOI21_X1   g15018(.A1(new_n15335_), .A2(new_n15343_), .B(new_n15810_), .ZN(new_n16042_));
  AOI21_X1   g15019(.A1(new_n14968_), .A2(new_n15329_), .B(new_n15321_), .ZN(new_n16043_));
  AOI21_X1   g15020(.A1(new_n15298_), .A2(new_n15299_), .B(new_n15314_), .ZN(new_n16044_));
  NOR2_X1    g15021(.A1(new_n12682_), .A2(new_n12699_), .ZN(new_n16045_));
  NAND2_X1   g15022(.A1(new_n12692_), .A2(new_n12613_), .ZN(new_n16046_));
  INV_X1     g15023(.I(new_n16046_), .ZN(new_n16047_));
  NOR2_X1    g15024(.A1(new_n15262_), .A2(new_n15215_), .ZN(new_n16048_));
  XOR2_X1    g15025(.A1(new_n15246_), .A2(new_n15250_), .Z(new_n16049_));
  XOR2_X1    g15026(.A1(new_n15227_), .A2(new_n15229_), .Z(new_n16050_));
  AND2_X2    g15027(.A1(new_n16049_), .A2(new_n16050_), .Z(new_n16051_));
  NAND4_X1   g15028(.A1(new_n16051_), .A2(new_n16045_), .A3(new_n16048_), .A4(new_n16047_), .ZN(new_n16052_));
  NAND2_X1   g15029(.A1(new_n12684_), .A2(new_n12637_), .ZN(new_n16053_));
  NAND2_X1   g15030(.A1(new_n15215_), .A2(new_n16053_), .ZN(new_n16054_));
  AOI22_X1   g15031(.A1(new_n15261_), .A2(new_n15238_), .B1(new_n12692_), .B2(new_n12613_), .ZN(new_n16055_));
  INV_X1     g15032(.I(new_n16055_), .ZN(new_n16056_));
  NAND2_X1   g15033(.A1(new_n16056_), .A2(new_n16054_), .ZN(new_n16057_));
  NOR2_X1    g15034(.A1(new_n16052_), .A2(new_n16057_), .ZN(new_n16058_));
  NOR2_X1    g15035(.A1(new_n16045_), .A2(new_n15233_), .ZN(new_n16059_));
  NAND2_X1   g15036(.A1(new_n15227_), .A2(new_n15229_), .ZN(new_n16060_));
  AOI21_X1   g15037(.A1(new_n16059_), .A2(new_n16060_), .B(new_n15230_), .ZN(new_n16061_));
  NAND2_X1   g15038(.A1(new_n15246_), .A2(new_n15250_), .ZN(new_n16062_));
  AOI21_X1   g15039(.A1(new_n16055_), .A2(new_n16062_), .B(new_n15251_), .ZN(new_n16063_));
  NOR2_X1    g15040(.A1(new_n16061_), .A2(new_n16063_), .ZN(new_n16064_));
  OAI21_X1   g15041(.A1(new_n15210_), .A2(new_n15278_), .B(new_n16064_), .ZN(new_n16065_));
  INV_X1     g15042(.I(new_n16060_), .ZN(new_n16066_));
  OAI21_X1   g15043(.A1(new_n16054_), .A2(new_n16066_), .B(new_n15224_), .ZN(new_n16067_));
  INV_X1     g15044(.I(new_n16063_), .ZN(new_n16068_));
  NAND2_X1   g15045(.A1(new_n16068_), .A2(new_n16067_), .ZN(new_n16069_));
  NAND3_X1   g15046(.A1(new_n16069_), .A2(new_n15276_), .A3(new_n15293_), .ZN(new_n16070_));
  AOI21_X1   g15047(.A1(new_n16070_), .A2(new_n16065_), .B(new_n16058_), .ZN(new_n16071_));
  NAND4_X1   g15048(.A1(new_n16048_), .A2(new_n16045_), .A3(new_n16049_), .A4(new_n16050_), .ZN(new_n16072_));
  OR3_X2     g15049(.A1(new_n16072_), .A2(new_n16046_), .A3(new_n16057_), .Z(new_n16073_));
  AOI21_X1   g15050(.A1(new_n15276_), .A2(new_n15293_), .B(new_n16069_), .ZN(new_n16074_));
  NOR3_X1    g15051(.A1(new_n15210_), .A2(new_n15278_), .A3(new_n16064_), .ZN(new_n16075_));
  NOR3_X1    g15052(.A1(new_n16074_), .A2(new_n16075_), .A3(new_n16073_), .ZN(new_n16076_));
  NOR2_X1    g15053(.A1(new_n16076_), .A2(new_n16071_), .ZN(new_n16077_));
  NAND2_X1   g15054(.A1(new_n12847_), .A2(new_n12830_), .ZN(new_n16078_));
  INV_X1     g15055(.I(new_n16078_), .ZN(new_n16079_));
  NOR2_X1    g15056(.A1(new_n12757_), .A2(new_n12840_), .ZN(new_n16080_));
  NOR2_X1    g15057(.A1(new_n15172_), .A2(new_n15166_), .ZN(new_n16081_));
  NOR2_X1    g15058(.A1(new_n15178_), .A2(new_n15174_), .ZN(new_n16082_));
  XNOR2_X1   g15059(.A1(new_n16082_), .A2(new_n16081_), .ZN(new_n16083_));
  XNOR2_X1   g15060(.A1(new_n15140_), .A2(new_n15144_), .ZN(new_n16084_));
  NOR4_X1    g15061(.A1(new_n16083_), .A2(new_n15156_), .A3(new_n15164_), .A4(new_n16084_), .ZN(new_n16085_));
  AOI22_X1   g15062(.A1(new_n15155_), .A2(new_n15132_), .B1(new_n12847_), .B2(new_n12830_), .ZN(new_n16086_));
  AOI22_X1   g15063(.A1(new_n12718_), .A2(new_n12759_), .B1(new_n15163_), .B2(new_n15161_), .ZN(new_n16087_));
  NOR2_X1    g15064(.A1(new_n16086_), .A2(new_n16087_), .ZN(new_n16088_));
  NAND4_X1   g15065(.A1(new_n16085_), .A2(new_n16079_), .A3(new_n16080_), .A4(new_n16088_), .ZN(new_n16089_));
  NAND2_X1   g15066(.A1(new_n15156_), .A2(new_n16078_), .ZN(new_n16090_));
  NAND2_X1   g15067(.A1(new_n15140_), .A2(new_n15144_), .ZN(new_n16091_));
  INV_X1     g15068(.I(new_n16091_), .ZN(new_n16092_));
  OAI21_X1   g15069(.A1(new_n16090_), .A2(new_n16092_), .B(new_n15151_), .ZN(new_n16093_));
  OAI22_X1   g15070(.A1(new_n15190_), .A2(new_n15188_), .B1(new_n12757_), .B2(new_n12840_), .ZN(new_n16094_));
  NAND2_X1   g15071(.A1(new_n16082_), .A2(new_n16081_), .ZN(new_n16095_));
  INV_X1     g15072(.I(new_n16095_), .ZN(new_n16096_));
  OAI21_X1   g15073(.A1(new_n16094_), .A2(new_n16096_), .B(new_n15179_), .ZN(new_n16097_));
  NAND2_X1   g15074(.A1(new_n16093_), .A2(new_n16097_), .ZN(new_n16098_));
  AOI21_X1   g15075(.A1(new_n15131_), .A2(new_n15207_), .B(new_n16098_), .ZN(new_n16099_));
  AOI21_X1   g15076(.A1(new_n16086_), .A2(new_n16091_), .B(new_n15145_), .ZN(new_n16100_));
  AOI21_X1   g15077(.A1(new_n16087_), .A2(new_n16095_), .B(new_n15185_), .ZN(new_n16101_));
  NOR2_X1    g15078(.A1(new_n16100_), .A2(new_n16101_), .ZN(new_n16102_));
  NOR3_X1    g15079(.A1(new_n15205_), .A2(new_n15286_), .A3(new_n16102_), .ZN(new_n16103_));
  OAI21_X1   g15080(.A1(new_n16099_), .A2(new_n16103_), .B(new_n16089_), .ZN(new_n16104_));
  INV_X1     g15081(.I(new_n16089_), .ZN(new_n16105_));
  OAI21_X1   g15082(.A1(new_n15205_), .A2(new_n15286_), .B(new_n16102_), .ZN(new_n16106_));
  NAND3_X1   g15083(.A1(new_n15131_), .A2(new_n16098_), .A3(new_n15207_), .ZN(new_n16107_));
  NAND3_X1   g15084(.A1(new_n16107_), .A2(new_n16106_), .A3(new_n16105_), .ZN(new_n16108_));
  NAND2_X1   g15085(.A1(new_n16104_), .A2(new_n16108_), .ZN(new_n16109_));
  NAND2_X1   g15086(.A1(new_n16077_), .A2(new_n16109_), .ZN(new_n16110_));
  OAI21_X1   g15087(.A1(new_n16074_), .A2(new_n16075_), .B(new_n16073_), .ZN(new_n16111_));
  NAND3_X1   g15088(.A1(new_n16070_), .A2(new_n16065_), .A3(new_n16058_), .ZN(new_n16112_));
  NAND2_X1   g15089(.A1(new_n16111_), .A2(new_n16112_), .ZN(new_n16113_));
  AOI21_X1   g15090(.A1(new_n16107_), .A2(new_n16106_), .B(new_n16105_), .ZN(new_n16114_));
  NOR3_X1    g15091(.A1(new_n16099_), .A2(new_n16103_), .A3(new_n16089_), .ZN(new_n16115_));
  NOR2_X1    g15092(.A1(new_n16114_), .A2(new_n16115_), .ZN(new_n16116_));
  NAND2_X1   g15093(.A1(new_n16116_), .A2(new_n16113_), .ZN(new_n16117_));
  AOI21_X1   g15094(.A1(new_n16110_), .A2(new_n16117_), .B(new_n16044_), .ZN(new_n16118_));
  OAI21_X1   g15095(.A1(new_n15130_), .A2(new_n15313_), .B(new_n15300_), .ZN(new_n16119_));
  NAND2_X1   g15096(.A1(new_n16109_), .A2(new_n16113_), .ZN(new_n16120_));
  NAND4_X1   g15097(.A1(new_n16111_), .A2(new_n16104_), .A3(new_n16108_), .A4(new_n16112_), .ZN(new_n16121_));
  AOI21_X1   g15098(.A1(new_n16120_), .A2(new_n16121_), .B(new_n16119_), .ZN(new_n16122_));
  NOR2_X1    g15099(.A1(new_n16118_), .A2(new_n16122_), .ZN(new_n16123_));
  NAND2_X1   g15100(.A1(new_n15127_), .A2(new_n15126_), .ZN(new_n16124_));
  NOR2_X1    g15101(.A1(new_n13005_), .A2(new_n12957_), .ZN(new_n16125_));
  NAND2_X1   g15102(.A1(new_n13012_), .A2(new_n12936_), .ZN(new_n16126_));
  NAND2_X1   g15103(.A1(new_n16126_), .A2(new_n15093_), .ZN(new_n16127_));
  XOR2_X1    g15104(.A1(new_n15082_), .A2(new_n15078_), .Z(new_n16128_));
  XOR2_X1    g15105(.A1(new_n15052_), .A2(new_n15055_), .Z(new_n16129_));
  AND4_X2    g15106(.A1(new_n15049_), .A2(new_n16129_), .A3(new_n15074_), .A4(new_n16128_), .Z(new_n16130_));
  NAND2_X1   g15107(.A1(new_n13019_), .A2(new_n13003_), .ZN(new_n16131_));
  AOI21_X1   g15108(.A1(new_n16131_), .A2(new_n15048_), .B(new_n16126_), .ZN(new_n16132_));
  NAND4_X1   g15109(.A1(new_n16130_), .A2(new_n16125_), .A3(new_n16127_), .A4(new_n16132_), .ZN(new_n16133_));
  NOR2_X1    g15110(.A1(new_n15060_), .A2(new_n15063_), .ZN(new_n16134_));
  AOI21_X1   g15111(.A1(new_n15049_), .A2(new_n15060_), .B(new_n16134_), .ZN(new_n16135_));
  OAI21_X1   g15112(.A1(new_n16131_), .A2(new_n15055_), .B(new_n16135_), .ZN(new_n16136_));
  INV_X1     g15113(.I(new_n16136_), .ZN(new_n16137_));
  NOR4_X1    g15114(.A1(new_n15087_), .A2(new_n15089_), .A3(new_n15075_), .A4(new_n15079_), .ZN(new_n16138_));
  OAI21_X1   g15115(.A1(new_n16127_), .A2(new_n16138_), .B(new_n15090_), .ZN(new_n16139_));
  NAND2_X1   g15116(.A1(new_n16137_), .A2(new_n16139_), .ZN(new_n16140_));
  AOI21_X1   g15117(.A1(new_n15106_), .A2(new_n15108_), .B(new_n16140_), .ZN(new_n16141_));
  INV_X1     g15118(.I(new_n15108_), .ZN(new_n16142_));
  INV_X1     g15119(.I(new_n16139_), .ZN(new_n16143_));
  NOR2_X1    g15120(.A1(new_n16143_), .A2(new_n16136_), .ZN(new_n16144_));
  NOR3_X1    g15121(.A1(new_n16142_), .A2(new_n15121_), .A3(new_n16144_), .ZN(new_n16145_));
  OAI21_X1   g15122(.A1(new_n16145_), .A2(new_n16141_), .B(new_n16133_), .ZN(new_n16146_));
  INV_X1     g15123(.I(new_n16133_), .ZN(new_n16147_));
  OAI21_X1   g15124(.A1(new_n16142_), .A2(new_n15121_), .B(new_n16144_), .ZN(new_n16148_));
  NAND3_X1   g15125(.A1(new_n15106_), .A2(new_n16140_), .A3(new_n15108_), .ZN(new_n16149_));
  NAND3_X1   g15126(.A1(new_n16148_), .A2(new_n16149_), .A3(new_n16147_), .ZN(new_n16150_));
  NAND2_X1   g15127(.A1(new_n15036_), .A2(new_n15038_), .ZN(new_n16151_));
  NAND2_X1   g15128(.A1(new_n13148_), .A2(new_n14973_), .ZN(new_n16152_));
  AOI21_X1   g15129(.A1(new_n16152_), .A2(new_n13052_), .B(new_n13058_), .ZN(new_n16153_));
  NAND2_X1   g15130(.A1(new_n13158_), .A2(new_n13139_), .ZN(new_n16154_));
  XOR2_X1    g15131(.A1(new_n14986_), .A2(new_n14977_), .Z(new_n16155_));
  XOR2_X1    g15132(.A1(new_n15012_), .A2(new_n15009_), .Z(new_n16156_));
  NAND3_X1   g15133(.A1(new_n16156_), .A2(new_n14973_), .A3(new_n15006_), .ZN(new_n16157_));
  OR3_X2     g15134(.A1(new_n16157_), .A2(new_n16154_), .A3(new_n16155_), .Z(new_n16158_));
  NAND2_X1   g15135(.A1(new_n16154_), .A2(new_n15022_), .ZN(new_n16159_));
  NAND3_X1   g15136(.A1(new_n16159_), .A2(new_n13071_), .A3(new_n13073_), .ZN(new_n16160_));
  NOR3_X1    g15137(.A1(new_n16158_), .A2(new_n16153_), .A3(new_n16160_), .ZN(new_n16161_));
  INV_X1     g15138(.I(new_n16161_), .ZN(new_n16162_));
  NOR2_X1    g15139(.A1(new_n16153_), .A2(new_n14987_), .ZN(new_n16163_));
  NOR3_X1    g15140(.A1(new_n14977_), .A2(new_n14978_), .A3(new_n14980_), .ZN(new_n16164_));
  INV_X1     g15141(.I(new_n16159_), .ZN(new_n16165_));
  NAND2_X1   g15142(.A1(new_n15012_), .A2(new_n15009_), .ZN(new_n16166_));
  AOI21_X1   g15143(.A1(new_n16165_), .A2(new_n16166_), .B(new_n15013_), .ZN(new_n16167_));
  NOR2_X1    g15144(.A1(new_n16151_), .A2(new_n16162_), .ZN(new_n16168_));
  NAND3_X1   g15145(.A1(new_n16146_), .A2(new_n16168_), .A3(new_n16150_), .ZN(new_n16169_));
  AOI21_X1   g15146(.A1(new_n16148_), .A2(new_n16149_), .B(new_n16147_), .ZN(new_n16170_));
  NOR3_X1    g15147(.A1(new_n16145_), .A2(new_n16141_), .A3(new_n16133_), .ZN(new_n16171_));
  INV_X1     g15148(.I(new_n15038_), .ZN(new_n16172_));
  NOR2_X1    g15149(.A1(new_n14970_), .A2(new_n16172_), .ZN(new_n16173_));
  NAND2_X1   g15150(.A1(new_n16173_), .A2(new_n16161_), .ZN(new_n16174_));
  OAI21_X1   g15151(.A1(new_n16171_), .A2(new_n16170_), .B(new_n16174_), .ZN(new_n16175_));
  AOI22_X1   g15152(.A1(new_n16124_), .A2(new_n15128_), .B1(new_n16169_), .B2(new_n16175_), .ZN(new_n16176_));
  OAI21_X1   g15153(.A1(new_n14969_), .A2(new_n15307_), .B(new_n15128_), .ZN(new_n16177_));
  OAI21_X1   g15154(.A1(new_n16171_), .A2(new_n16170_), .B(new_n16168_), .ZN(new_n16178_));
  NAND3_X1   g15155(.A1(new_n16146_), .A2(new_n16174_), .A3(new_n16150_), .ZN(new_n16179_));
  AOI21_X1   g15156(.A1(new_n16178_), .A2(new_n16179_), .B(new_n16177_), .ZN(new_n16180_));
  OAI21_X1   g15157(.A1(new_n16176_), .A2(new_n16180_), .B(new_n16123_), .ZN(new_n16181_));
  NOR2_X1    g15158(.A1(new_n16116_), .A2(new_n16113_), .ZN(new_n16182_));
  NOR2_X1    g15159(.A1(new_n16077_), .A2(new_n16109_), .ZN(new_n16183_));
  OAI21_X1   g15160(.A1(new_n16183_), .A2(new_n16182_), .B(new_n16119_), .ZN(new_n16184_));
  NOR2_X1    g15161(.A1(new_n16116_), .A2(new_n16077_), .ZN(new_n16185_));
  NOR4_X1    g15162(.A1(new_n16076_), .A2(new_n16114_), .A3(new_n16115_), .A4(new_n16071_), .ZN(new_n16186_));
  OAI21_X1   g15163(.A1(new_n16185_), .A2(new_n16186_), .B(new_n16044_), .ZN(new_n16187_));
  NAND2_X1   g15164(.A1(new_n16184_), .A2(new_n16187_), .ZN(new_n16188_));
  NAND2_X1   g15165(.A1(new_n16175_), .A2(new_n16169_), .ZN(new_n16189_));
  NAND2_X1   g15166(.A1(new_n16189_), .A2(new_n16177_), .ZN(new_n16190_));
  AOI21_X1   g15167(.A1(new_n15126_), .A2(new_n15127_), .B(new_n15308_), .ZN(new_n16191_));
  NAND2_X1   g15168(.A1(new_n16178_), .A2(new_n16179_), .ZN(new_n16192_));
  NAND2_X1   g15169(.A1(new_n16192_), .A2(new_n16191_), .ZN(new_n16193_));
  NAND3_X1   g15170(.A1(new_n16188_), .A2(new_n16190_), .A3(new_n16193_), .ZN(new_n16194_));
  AOI21_X1   g15171(.A1(new_n16181_), .A2(new_n16194_), .B(new_n16043_), .ZN(new_n16195_));
  OAI21_X1   g15172(.A1(new_n15319_), .A2(new_n15320_), .B(new_n15330_), .ZN(new_n16196_));
  OAI22_X1   g15173(.A1(new_n16180_), .A2(new_n16176_), .B1(new_n16118_), .B2(new_n16122_), .ZN(new_n16197_));
  NAND3_X1   g15174(.A1(new_n16123_), .A2(new_n16190_), .A3(new_n16193_), .ZN(new_n16198_));
  AOI21_X1   g15175(.A1(new_n16197_), .A2(new_n16198_), .B(new_n16196_), .ZN(new_n16199_));
  NOR2_X1    g15176(.A1(new_n16195_), .A2(new_n16199_), .ZN(new_n16200_));
  OAI21_X1   g15177(.A1(new_n14964_), .A2(new_n14965_), .B(new_n15341_), .ZN(new_n16201_));
  OAI21_X1   g15178(.A1(new_n14958_), .A2(new_n14957_), .B(new_n14942_), .ZN(new_n16202_));
  NAND2_X1   g15179(.A1(new_n13270_), .A2(new_n13225_), .ZN(new_n16203_));
  NOR2_X1    g15180(.A1(new_n13300_), .A2(new_n13344_), .ZN(new_n16204_));
  NOR2_X1    g15181(.A1(new_n14857_), .A2(new_n14907_), .ZN(new_n16205_));
  XOR2_X1    g15182(.A1(new_n14894_), .A2(new_n14898_), .Z(new_n16206_));
  NOR2_X1    g15183(.A1(new_n14861_), .A2(new_n14859_), .ZN(new_n16207_));
  NOR2_X1    g15184(.A1(new_n14867_), .A2(new_n14863_), .ZN(new_n16208_));
  XOR2_X1    g15185(.A1(new_n16207_), .A2(new_n16208_), .Z(new_n16209_));
  NAND4_X1   g15186(.A1(new_n16209_), .A2(new_n16205_), .A3(new_n16206_), .A4(new_n16204_), .ZN(new_n16210_));
  OAI21_X1   g15187(.A1(new_n13300_), .A2(new_n13344_), .B(new_n14857_), .ZN(new_n16211_));
  NAND2_X1   g15188(.A1(new_n16203_), .A2(new_n14907_), .ZN(new_n16212_));
  NAND2_X1   g15189(.A1(new_n16211_), .A2(new_n16212_), .ZN(new_n16213_));
  NOR3_X1    g15190(.A1(new_n16210_), .A2(new_n16213_), .A3(new_n16203_), .ZN(new_n16214_));
  INV_X1     g15191(.I(new_n16214_), .ZN(new_n16215_));
  AOI21_X1   g15192(.A1(new_n16207_), .A2(new_n16208_), .B(new_n16211_), .ZN(new_n16216_));
  AOI21_X1   g15193(.A1(new_n14894_), .A2(new_n14898_), .B(new_n16212_), .ZN(new_n16217_));
  OAI22_X1   g15194(.A1(new_n14874_), .A2(new_n16216_), .B1(new_n16217_), .B2(new_n14899_), .ZN(new_n16218_));
  AOI21_X1   g15195(.A1(new_n14921_), .A2(new_n14935_), .B(new_n16218_), .ZN(new_n16219_));
  NAND2_X1   g15196(.A1(new_n14921_), .A2(new_n14935_), .ZN(new_n16220_));
  NOR2_X1    g15197(.A1(new_n14877_), .A2(new_n16204_), .ZN(new_n16221_));
  NAND2_X1   g15198(.A1(new_n16207_), .A2(new_n16208_), .ZN(new_n16222_));
  AOI21_X1   g15199(.A1(new_n16221_), .A2(new_n16222_), .B(new_n14874_), .ZN(new_n16223_));
  NOR2_X1    g15200(.A1(new_n13268_), .A2(new_n13352_), .ZN(new_n16224_));
  NOR2_X1    g15201(.A1(new_n14886_), .A2(new_n16224_), .ZN(new_n16225_));
  NAND2_X1   g15202(.A1(new_n14894_), .A2(new_n14898_), .ZN(new_n16226_));
  AOI21_X1   g15203(.A1(new_n16225_), .A2(new_n16226_), .B(new_n14899_), .ZN(new_n16227_));
  NOR2_X1    g15204(.A1(new_n16223_), .A2(new_n16227_), .ZN(new_n16228_));
  NOR2_X1    g15205(.A1(new_n16220_), .A2(new_n16228_), .ZN(new_n16229_));
  OAI21_X1   g15206(.A1(new_n16229_), .A2(new_n16219_), .B(new_n16215_), .ZN(new_n16230_));
  NAND2_X1   g15207(.A1(new_n16220_), .A2(new_n16228_), .ZN(new_n16231_));
  NAND3_X1   g15208(.A1(new_n16218_), .A2(new_n14921_), .A3(new_n14935_), .ZN(new_n16232_));
  NAND3_X1   g15209(.A1(new_n16231_), .A2(new_n16232_), .A3(new_n16214_), .ZN(new_n16233_));
  NAND2_X1   g15210(.A1(new_n14847_), .A2(new_n14849_), .ZN(new_n16234_));
  AOI21_X1   g15211(.A1(new_n13409_), .A2(new_n14789_), .B(new_n13395_), .ZN(new_n16235_));
  NOR2_X1    g15212(.A1(new_n16235_), .A2(new_n13386_), .ZN(new_n16236_));
  NOR2_X1    g15213(.A1(new_n13501_), .A2(new_n13481_), .ZN(new_n16237_));
  XOR2_X1    g15214(.A1(new_n14801_), .A2(new_n14800_), .Z(new_n16238_));
  XOR2_X1    g15215(.A1(new_n14823_), .A2(new_n14820_), .Z(new_n16239_));
  AND3_X2    g15216(.A1(new_n16239_), .A2(new_n14789_), .A3(new_n14817_), .Z(new_n16240_));
  NAND3_X1   g15217(.A1(new_n16240_), .A2(new_n16237_), .A3(new_n16238_), .ZN(new_n16241_));
  AOI21_X1   g15218(.A1(new_n13483_), .A2(new_n13421_), .B(new_n14817_), .ZN(new_n16242_));
  OR3_X2     g15219(.A1(new_n16242_), .A2(new_n13409_), .A3(new_n13411_), .Z(new_n16243_));
  NOR3_X1    g15220(.A1(new_n16241_), .A2(new_n16243_), .A3(new_n16236_), .ZN(new_n16244_));
  INV_X1     g15221(.I(new_n16244_), .ZN(new_n16245_));
  OAI21_X1   g15222(.A1(new_n16235_), .A2(new_n13386_), .B(new_n14798_), .ZN(new_n16246_));
  INV_X1     g15223(.I(new_n16246_), .ZN(new_n16247_));
  NOR3_X1    g15224(.A1(new_n14794_), .A2(new_n14797_), .A3(new_n14795_), .ZN(new_n16248_));
  OAI21_X1   g15225(.A1(new_n14826_), .A2(new_n14829_), .B(new_n16242_), .ZN(new_n16249_));
  NAND2_X1   g15226(.A1(new_n16249_), .A2(new_n14830_), .ZN(new_n16250_));
  INV_X1     g15227(.I(new_n16250_), .ZN(new_n16251_));
  NOR2_X1    g15228(.A1(new_n16234_), .A2(new_n16245_), .ZN(new_n16252_));
  NAND3_X1   g15229(.A1(new_n16252_), .A2(new_n16230_), .A3(new_n16233_), .ZN(new_n16253_));
  AOI21_X1   g15230(.A1(new_n16231_), .A2(new_n16232_), .B(new_n16214_), .ZN(new_n16254_));
  NOR3_X1    g15231(.A1(new_n16229_), .A2(new_n16219_), .A3(new_n16215_), .ZN(new_n16255_));
  NOR2_X1    g15232(.A1(new_n14844_), .A2(new_n14808_), .ZN(new_n16256_));
  NOR2_X1    g15233(.A1(new_n14786_), .A2(new_n16256_), .ZN(new_n16257_));
  NAND2_X1   g15234(.A1(new_n16257_), .A2(new_n16244_), .ZN(new_n16258_));
  OAI21_X1   g15235(.A1(new_n16255_), .A2(new_n16254_), .B(new_n16258_), .ZN(new_n16259_));
  NAND2_X1   g15236(.A1(new_n16259_), .A2(new_n16253_), .ZN(new_n16260_));
  NAND2_X1   g15237(.A1(new_n16260_), .A2(new_n16202_), .ZN(new_n16261_));
  AOI21_X1   g15238(.A1(new_n14940_), .A2(new_n14941_), .B(new_n14959_), .ZN(new_n16262_));
  OAI21_X1   g15239(.A1(new_n16254_), .A2(new_n16255_), .B(new_n16252_), .ZN(new_n16263_));
  NAND3_X1   g15240(.A1(new_n16230_), .A2(new_n16258_), .A3(new_n16233_), .ZN(new_n16264_));
  NAND2_X1   g15241(.A1(new_n16263_), .A2(new_n16264_), .ZN(new_n16265_));
  NAND2_X1   g15242(.A1(new_n16265_), .A2(new_n16262_), .ZN(new_n16266_));
  NAND2_X1   g15243(.A1(new_n16266_), .A2(new_n16261_), .ZN(new_n16267_));
  NAND2_X1   g15244(.A1(new_n14950_), .A2(new_n14616_), .ZN(new_n16268_));
  NAND2_X1   g15245(.A1(new_n13709_), .A2(new_n13694_), .ZN(new_n16269_));
  NAND2_X1   g15246(.A1(new_n13622_), .A2(new_n13702_), .ZN(new_n16270_));
  NAND2_X1   g15247(.A1(new_n16270_), .A2(new_n14720_), .ZN(new_n16271_));
  INV_X1     g15248(.I(new_n16271_), .ZN(new_n16272_));
  NOR2_X1    g15249(.A1(new_n14728_), .A2(new_n14721_), .ZN(new_n16273_));
  NOR2_X1    g15250(.A1(new_n14734_), .A2(new_n14730_), .ZN(new_n16274_));
  XOR2_X1    g15251(.A1(new_n16274_), .A2(new_n16273_), .Z(new_n16275_));
  XOR2_X1    g15252(.A1(new_n14696_), .A2(new_n14700_), .Z(new_n16276_));
  NAND4_X1   g15253(.A1(new_n16276_), .A2(new_n16275_), .A3(new_n14712_), .A4(new_n14743_), .ZN(new_n16277_));
  NOR2_X1    g15254(.A1(new_n13696_), .A2(new_n13648_), .ZN(new_n16278_));
  INV_X1     g15255(.I(new_n16270_), .ZN(new_n16279_));
  OAI21_X1   g15256(.A1(new_n16278_), .A2(new_n14712_), .B(new_n16279_), .ZN(new_n16280_));
  NOR4_X1    g15257(.A1(new_n16280_), .A2(new_n16277_), .A3(new_n16269_), .A4(new_n16272_), .ZN(new_n16281_));
  INV_X1     g15258(.I(new_n16281_), .ZN(new_n16282_));
  NAND2_X1   g15259(.A1(new_n16278_), .A2(new_n14700_), .ZN(new_n16283_));
  NOR2_X1    g15260(.A1(new_n14693_), .A2(new_n14705_), .ZN(new_n16284_));
  NOR2_X1    g15261(.A1(new_n14696_), .A2(new_n14700_), .ZN(new_n16285_));
  NOR2_X1    g15262(.A1(new_n16284_), .A2(new_n16285_), .ZN(new_n16286_));
  NOR4_X1    g15263(.A1(new_n14734_), .A2(new_n14728_), .A3(new_n14721_), .A4(new_n14730_), .ZN(new_n16287_));
  OAI21_X1   g15264(.A1(new_n16271_), .A2(new_n16287_), .B(new_n14735_), .ZN(new_n16288_));
  NAND3_X1   g15265(.A1(new_n16288_), .A2(new_n16283_), .A3(new_n16286_), .ZN(new_n16289_));
  AOI21_X1   g15266(.A1(new_n14767_), .A2(new_n14758_), .B(new_n16289_), .ZN(new_n16290_));
  NOR3_X1    g15267(.A1(new_n14747_), .A2(new_n14750_), .A3(new_n14749_), .ZN(new_n16291_));
  INV_X1     g15268(.I(new_n16289_), .ZN(new_n16292_));
  NOR3_X1    g15269(.A1(new_n14756_), .A2(new_n16292_), .A3(new_n16291_), .ZN(new_n16293_));
  OAI21_X1   g15270(.A1(new_n16290_), .A2(new_n16293_), .B(new_n16282_), .ZN(new_n16294_));
  OAI21_X1   g15271(.A1(new_n14756_), .A2(new_n16291_), .B(new_n16292_), .ZN(new_n16295_));
  NAND4_X1   g15272(.A1(new_n14685_), .A2(new_n14758_), .A3(new_n13864_), .A4(new_n16289_), .ZN(new_n16296_));
  NAND3_X1   g15273(.A1(new_n16295_), .A2(new_n16296_), .A3(new_n16281_), .ZN(new_n16297_));
  NAND2_X1   g15274(.A1(new_n14777_), .A2(new_n14683_), .ZN(new_n16298_));
  AOI21_X1   g15275(.A1(new_n13757_), .A2(new_n14620_), .B(new_n13741_), .ZN(new_n16299_));
  NAND2_X1   g15276(.A1(new_n13836_), .A2(new_n13838_), .ZN(new_n16300_));
  NOR2_X1    g15277(.A1(new_n14635_), .A2(new_n14627_), .ZN(new_n16301_));
  XNOR2_X1   g15278(.A1(new_n16301_), .A2(new_n14625_), .ZN(new_n16302_));
  NOR2_X1    g15279(.A1(new_n13846_), .A2(new_n13825_), .ZN(new_n16303_));
  XNOR2_X1   g15280(.A1(new_n14662_), .A2(new_n14657_), .ZN(new_n16304_));
  NAND4_X1   g15281(.A1(new_n16303_), .A2(new_n16304_), .A3(new_n14620_), .A4(new_n14653_), .ZN(new_n16305_));
  NOR2_X1    g15282(.A1(new_n16303_), .A2(new_n14653_), .ZN(new_n16306_));
  NOR4_X1    g15283(.A1(new_n16305_), .A2(new_n16300_), .A3(new_n16306_), .A4(new_n16302_), .ZN(new_n16307_));
  OAI21_X1   g15284(.A1(new_n13730_), .A2(new_n16299_), .B(new_n16307_), .ZN(new_n16308_));
  NOR2_X1    g15285(.A1(new_n16299_), .A2(new_n13730_), .ZN(new_n16309_));
  NOR2_X1    g15286(.A1(new_n16309_), .A2(new_n14632_), .ZN(new_n16310_));
  NOR4_X1    g15287(.A1(new_n14634_), .A2(new_n14635_), .A3(new_n14621_), .A4(new_n14627_), .ZN(new_n16311_));
  NOR2_X1    g15288(.A1(new_n14658_), .A2(new_n14662_), .ZN(new_n16312_));
  OR3_X2     g15289(.A1(new_n16303_), .A2(new_n14653_), .A3(new_n16312_), .Z(new_n16313_));
  NAND2_X1   g15290(.A1(new_n16313_), .A2(new_n14663_), .ZN(new_n16314_));
  INV_X1     g15291(.I(new_n16314_), .ZN(new_n16315_));
  NOR2_X1    g15292(.A1(new_n16298_), .A2(new_n16308_), .ZN(new_n16316_));
  NAND3_X1   g15293(.A1(new_n16294_), .A2(new_n16316_), .A3(new_n16297_), .ZN(new_n16317_));
  AOI21_X1   g15294(.A1(new_n16295_), .A2(new_n16296_), .B(new_n16281_), .ZN(new_n16318_));
  NOR3_X1    g15295(.A1(new_n16290_), .A2(new_n16293_), .A3(new_n16282_), .ZN(new_n16319_));
  INV_X1     g15296(.I(new_n14683_), .ZN(new_n16320_));
  NOR2_X1    g15297(.A1(new_n16320_), .A2(new_n14679_), .ZN(new_n16321_));
  OR2_X2     g15298(.A1(new_n16306_), .A2(new_n16300_), .Z(new_n16322_));
  NOR4_X1    g15299(.A1(new_n16322_), .A2(new_n16309_), .A3(new_n16302_), .A4(new_n16305_), .ZN(new_n16323_));
  NAND2_X1   g15300(.A1(new_n16321_), .A2(new_n16323_), .ZN(new_n16324_));
  OAI21_X1   g15301(.A1(new_n16319_), .A2(new_n16318_), .B(new_n16324_), .ZN(new_n16325_));
  AOI22_X1   g15302(.A1(new_n16268_), .A2(new_n14951_), .B1(new_n16317_), .B2(new_n16325_), .ZN(new_n16326_));
  OAI21_X1   g15303(.A1(new_n14773_), .A2(new_n14780_), .B(new_n14951_), .ZN(new_n16327_));
  OAI21_X1   g15304(.A1(new_n16319_), .A2(new_n16318_), .B(new_n16316_), .ZN(new_n16328_));
  NAND3_X1   g15305(.A1(new_n16294_), .A2(new_n16324_), .A3(new_n16297_), .ZN(new_n16329_));
  AOI21_X1   g15306(.A1(new_n16328_), .A2(new_n16329_), .B(new_n16327_), .ZN(new_n16330_));
  NOR2_X1    g15307(.A1(new_n16330_), .A2(new_n16326_), .ZN(new_n16331_));
  NOR2_X1    g15308(.A1(new_n16331_), .A2(new_n16267_), .ZN(new_n16332_));
  NAND2_X1   g15309(.A1(new_n14941_), .A2(new_n14940_), .ZN(new_n16333_));
  AOI22_X1   g15310(.A1(new_n16333_), .A2(new_n14942_), .B1(new_n16253_), .B2(new_n16259_), .ZN(new_n16334_));
  AOI21_X1   g15311(.A1(new_n16230_), .A2(new_n16233_), .B(new_n16258_), .ZN(new_n16335_));
  NOR3_X1    g15312(.A1(new_n16252_), .A2(new_n16255_), .A3(new_n16254_), .ZN(new_n16336_));
  NOR2_X1    g15313(.A1(new_n16335_), .A2(new_n16336_), .ZN(new_n16337_));
  NOR2_X1    g15314(.A1(new_n16337_), .A2(new_n16202_), .ZN(new_n16338_));
  NOR2_X1    g15315(.A1(new_n16338_), .A2(new_n16334_), .ZN(new_n16339_));
  NAND2_X1   g15316(.A1(new_n16325_), .A2(new_n16317_), .ZN(new_n16340_));
  NAND2_X1   g15317(.A1(new_n16340_), .A2(new_n16327_), .ZN(new_n16341_));
  AOI21_X1   g15318(.A1(new_n14616_), .A2(new_n14950_), .B(new_n14781_), .ZN(new_n16342_));
  NAND2_X1   g15319(.A1(new_n16328_), .A2(new_n16329_), .ZN(new_n16343_));
  NAND2_X1   g15320(.A1(new_n16343_), .A2(new_n16342_), .ZN(new_n16344_));
  NAND2_X1   g15321(.A1(new_n16344_), .A2(new_n16341_), .ZN(new_n16345_));
  NOR2_X1    g15322(.A1(new_n16345_), .A2(new_n16339_), .ZN(new_n16346_));
  OAI21_X1   g15323(.A1(new_n16332_), .A2(new_n16346_), .B(new_n16201_), .ZN(new_n16347_));
  AOI21_X1   g15324(.A1(new_n14615_), .A2(new_n15340_), .B(new_n14966_), .ZN(new_n16348_));
  AOI22_X1   g15325(.A1(new_n16341_), .A2(new_n16344_), .B1(new_n16266_), .B2(new_n16261_), .ZN(new_n16349_));
  NOR4_X1    g15326(.A1(new_n16330_), .A2(new_n16338_), .A3(new_n16326_), .A4(new_n16334_), .ZN(new_n16350_));
  OAI21_X1   g15327(.A1(new_n16349_), .A2(new_n16350_), .B(new_n16348_), .ZN(new_n16351_));
  NAND2_X1   g15328(.A1(new_n16347_), .A2(new_n16351_), .ZN(new_n16352_));
  NAND2_X1   g15329(.A1(new_n16352_), .A2(new_n16200_), .ZN(new_n16353_));
  AOI21_X1   g15330(.A1(new_n16190_), .A2(new_n16193_), .B(new_n16188_), .ZN(new_n16354_));
  NOR3_X1    g15331(.A1(new_n16123_), .A2(new_n16180_), .A3(new_n16176_), .ZN(new_n16355_));
  OAI21_X1   g15332(.A1(new_n16354_), .A2(new_n16355_), .B(new_n16196_), .ZN(new_n16356_));
  AOI22_X1   g15333(.A1(new_n16193_), .A2(new_n16190_), .B1(new_n16184_), .B2(new_n16187_), .ZN(new_n16357_));
  NOR4_X1    g15334(.A1(new_n16180_), .A2(new_n16118_), .A3(new_n16176_), .A4(new_n16122_), .ZN(new_n16358_));
  OAI21_X1   g15335(.A1(new_n16357_), .A2(new_n16358_), .B(new_n16043_), .ZN(new_n16359_));
  NAND2_X1   g15336(.A1(new_n16359_), .A2(new_n16356_), .ZN(new_n16360_));
  NAND2_X1   g15337(.A1(new_n16345_), .A2(new_n16339_), .ZN(new_n16361_));
  NAND2_X1   g15338(.A1(new_n16331_), .A2(new_n16267_), .ZN(new_n16362_));
  AOI21_X1   g15339(.A1(new_n16362_), .A2(new_n16361_), .B(new_n16348_), .ZN(new_n16363_));
  OAI22_X1   g15340(.A1(new_n16330_), .A2(new_n16326_), .B1(new_n16338_), .B2(new_n16334_), .ZN(new_n16364_));
  NAND4_X1   g15341(.A1(new_n16341_), .A2(new_n16344_), .A3(new_n16266_), .A4(new_n16261_), .ZN(new_n16365_));
  AOI21_X1   g15342(.A1(new_n16364_), .A2(new_n16365_), .B(new_n16201_), .ZN(new_n16366_));
  NOR2_X1    g15343(.A1(new_n16363_), .A2(new_n16366_), .ZN(new_n16367_));
  NAND2_X1   g15344(.A1(new_n16367_), .A2(new_n16360_), .ZN(new_n16368_));
  AOI21_X1   g15345(.A1(new_n16368_), .A2(new_n16353_), .B(new_n16042_), .ZN(new_n16369_));
  OAI21_X1   g15346(.A1(new_n14614_), .A2(new_n15811_), .B(new_n15336_), .ZN(new_n16370_));
  NAND4_X1   g15347(.A1(new_n16347_), .A2(new_n16351_), .A3(new_n16359_), .A4(new_n16356_), .ZN(new_n16371_));
  OAI22_X1   g15348(.A1(new_n16363_), .A2(new_n16366_), .B1(new_n16195_), .B2(new_n16199_), .ZN(new_n16372_));
  AOI21_X1   g15349(.A1(new_n16371_), .A2(new_n16372_), .B(new_n16370_), .ZN(new_n16373_));
  NOR2_X1    g15350(.A1(new_n16369_), .A2(new_n16373_), .ZN(new_n16374_));
  NAND3_X1   g15351(.A1(new_n16038_), .A2(new_n16041_), .A3(new_n16374_), .ZN(new_n16375_));
  AOI21_X1   g15352(.A1(new_n16039_), .A2(new_n16040_), .B(new_n15918_), .ZN(new_n16376_));
  NOR3_X1    g15353(.A1(new_n16037_), .A2(new_n16033_), .A3(new_n15919_), .ZN(new_n16377_));
  NOR2_X1    g15354(.A1(new_n16367_), .A2(new_n16360_), .ZN(new_n16378_));
  NOR2_X1    g15355(.A1(new_n16352_), .A2(new_n16200_), .ZN(new_n16379_));
  OAI21_X1   g15356(.A1(new_n16378_), .A2(new_n16379_), .B(new_n16370_), .ZN(new_n16380_));
  NOR4_X1    g15357(.A1(new_n16363_), .A2(new_n16366_), .A3(new_n16195_), .A4(new_n16199_), .ZN(new_n16381_));
  AOI22_X1   g15358(.A1(new_n16347_), .A2(new_n16351_), .B1(new_n16359_), .B2(new_n16356_), .ZN(new_n16382_));
  OAI21_X1   g15359(.A1(new_n16381_), .A2(new_n16382_), .B(new_n16042_), .ZN(new_n16383_));
  NAND2_X1   g15360(.A1(new_n16380_), .A2(new_n16383_), .ZN(new_n16384_));
  OAI21_X1   g15361(.A1(new_n16377_), .A2(new_n16376_), .B(new_n16384_), .ZN(new_n16385_));
  NAND2_X1   g15362(.A1(new_n16385_), .A2(new_n16375_), .ZN(new_n16386_));
  OAI21_X1   g15363(.A1(new_n15832_), .A2(new_n14612_), .B(new_n15816_), .ZN(new_n16387_));
  AOI21_X1   g15364(.A1(new_n14595_), .A2(new_n14270_), .B(new_n14593_), .ZN(new_n16388_));
  INV_X1     g15365(.I(new_n16388_), .ZN(new_n16389_));
  NAND2_X1   g15366(.A1(new_n14562_), .A2(new_n14545_), .ZN(new_n16390_));
  INV_X1     g15367(.I(new_n16390_), .ZN(new_n16391_));
  NOR2_X1    g15368(.A1(new_n4284_), .A2(new_n4325_), .ZN(new_n16392_));
  NAND2_X1   g15369(.A1(new_n14523_), .A2(new_n14520_), .ZN(new_n16393_));
  NAND2_X1   g15370(.A1(new_n14527_), .A2(new_n14524_), .ZN(new_n16394_));
  XNOR2_X1   g15371(.A1(new_n16394_), .A2(new_n16393_), .ZN(new_n16395_));
  XNOR2_X1   g15372(.A1(new_n14505_), .A2(new_n14500_), .ZN(new_n16396_));
  NOR4_X1    g15373(.A1(new_n16396_), .A2(new_n16395_), .A3(new_n14494_), .A4(new_n14518_), .ZN(new_n16397_));
  NOR2_X1    g15374(.A1(new_n14519_), .A2(new_n16392_), .ZN(new_n16398_));
  NOR2_X1    g15375(.A1(new_n14495_), .A2(new_n14493_), .ZN(new_n16399_));
  NOR2_X1    g15376(.A1(new_n16398_), .A2(new_n16399_), .ZN(new_n16400_));
  NAND4_X1   g15377(.A1(new_n16397_), .A2(new_n16400_), .A3(new_n14495_), .A4(new_n16392_), .ZN(new_n16401_));
  NOR2_X1    g15378(.A1(new_n16399_), .A2(new_n14508_), .ZN(new_n16402_));
  NOR2_X1    g15379(.A1(new_n14505_), .A2(new_n14500_), .ZN(new_n16403_));
  INV_X1     g15380(.I(new_n14528_), .ZN(new_n16404_));
  OAI21_X1   g15381(.A1(new_n14519_), .A2(new_n16392_), .B(new_n16404_), .ZN(new_n16405_));
  NAND4_X1   g15382(.A1(new_n14527_), .A2(new_n14523_), .A3(new_n14520_), .A4(new_n14524_), .ZN(new_n16406_));
  NAND2_X1   g15383(.A1(new_n16405_), .A2(new_n16406_), .ZN(new_n16407_));
  NOR3_X1    g15384(.A1(new_n16407_), .A2(new_n16402_), .A3(new_n16403_), .ZN(new_n16408_));
  NAND2_X1   g15385(.A1(new_n16401_), .A2(new_n16408_), .ZN(new_n16409_));
  INV_X1     g15386(.I(new_n16409_), .ZN(new_n16410_));
  NOR2_X1    g15387(.A1(new_n16401_), .A2(new_n16408_), .ZN(new_n16411_));
  NOR2_X1    g15388(.A1(new_n16410_), .A2(new_n16411_), .ZN(new_n16412_));
  NOR2_X1    g15389(.A1(new_n16412_), .A2(new_n16391_), .ZN(new_n16413_));
  INV_X1     g15390(.I(new_n16411_), .ZN(new_n16414_));
  NAND2_X1   g15391(.A1(new_n16414_), .A2(new_n16409_), .ZN(new_n16415_));
  NOR2_X1    g15392(.A1(new_n16415_), .A2(new_n16390_), .ZN(new_n16416_));
  NOR2_X1    g15393(.A1(new_n16413_), .A2(new_n16416_), .ZN(new_n16417_));
  INV_X1     g15394(.I(new_n16417_), .ZN(new_n16418_));
  NAND2_X1   g15395(.A1(new_n14486_), .A2(new_n14422_), .ZN(new_n16419_));
  NOR2_X1    g15396(.A1(new_n14455_), .A2(new_n14426_), .ZN(new_n16420_));
  INV_X1     g15397(.I(new_n14460_), .ZN(new_n16421_));
  NAND2_X1   g15398(.A1(new_n16421_), .A2(new_n14456_), .ZN(new_n16422_));
  NOR2_X1    g15399(.A1(new_n4093_), .A2(new_n14463_), .ZN(new_n16423_));
  NAND2_X1   g15400(.A1(new_n4416_), .A2(new_n16423_), .ZN(new_n16424_));
  NAND2_X1   g15401(.A1(new_n16424_), .A2(new_n14461_), .ZN(new_n16425_));
  XOR2_X1    g15402(.A1(new_n16422_), .A2(new_n16425_), .Z(new_n16426_));
  XNOR2_X1   g15403(.A1(new_n14438_), .A2(new_n14434_), .ZN(new_n16427_));
  NAND4_X1   g15404(.A1(new_n16426_), .A2(new_n16420_), .A3(new_n16427_), .A4(new_n14437_), .ZN(new_n16428_));
  NAND2_X1   g15405(.A1(new_n14455_), .A2(new_n14470_), .ZN(new_n16429_));
  NAND2_X1   g15406(.A1(new_n14428_), .A2(new_n14426_), .ZN(new_n16430_));
  NAND2_X1   g15407(.A1(new_n16429_), .A2(new_n16430_), .ZN(new_n16431_));
  NOR3_X1    g15408(.A1(new_n16428_), .A2(new_n14470_), .A3(new_n16431_), .ZN(new_n16432_));
  NAND2_X1   g15409(.A1(new_n16430_), .A2(new_n14440_), .ZN(new_n16433_));
  NOR2_X1    g15410(.A1(new_n14439_), .A2(new_n14438_), .ZN(new_n16434_));
  INV_X1     g15411(.I(new_n16434_), .ZN(new_n16435_));
  NAND2_X1   g15412(.A1(new_n16433_), .A2(new_n16435_), .ZN(new_n16436_));
  NAND2_X1   g15413(.A1(new_n16429_), .A2(new_n14465_), .ZN(new_n16437_));
  NOR2_X1    g15414(.A1(new_n16422_), .A2(new_n16425_), .ZN(new_n16438_));
  INV_X1     g15415(.I(new_n16438_), .ZN(new_n16439_));
  NAND2_X1   g15416(.A1(new_n16437_), .A2(new_n16439_), .ZN(new_n16440_));
  NOR3_X1    g15417(.A1(new_n16432_), .A2(new_n16436_), .A3(new_n16440_), .ZN(new_n16441_));
  INV_X1     g15418(.I(new_n16432_), .ZN(new_n16442_));
  NOR2_X1    g15419(.A1(new_n16440_), .A2(new_n16436_), .ZN(new_n16443_));
  NOR2_X1    g15420(.A1(new_n16442_), .A2(new_n16443_), .ZN(new_n16444_));
  OAI21_X1   g15421(.A1(new_n16444_), .A2(new_n16441_), .B(new_n16419_), .ZN(new_n16445_));
  NOR2_X1    g15422(.A1(new_n14555_), .A2(new_n14484_), .ZN(new_n16446_));
  NAND2_X1   g15423(.A1(new_n16442_), .A2(new_n16443_), .ZN(new_n16447_));
  OAI21_X1   g15424(.A1(new_n16440_), .A2(new_n16436_), .B(new_n16432_), .ZN(new_n16448_));
  NAND3_X1   g15425(.A1(new_n16447_), .A2(new_n16446_), .A3(new_n16448_), .ZN(new_n16449_));
  NAND2_X1   g15426(.A1(new_n16445_), .A2(new_n16449_), .ZN(new_n16450_));
  AOI21_X1   g15427(.A1(new_n14567_), .A2(new_n14568_), .B(new_n14582_), .ZN(new_n16451_));
  NOR2_X1    g15428(.A1(new_n16451_), .A2(new_n16450_), .ZN(new_n16452_));
  NAND2_X1   g15429(.A1(new_n16451_), .A2(new_n16450_), .ZN(new_n16453_));
  INV_X1     g15430(.I(new_n16453_), .ZN(new_n16454_));
  OAI21_X1   g15431(.A1(new_n16454_), .A2(new_n16452_), .B(new_n16418_), .ZN(new_n16455_));
  AOI21_X1   g15432(.A1(new_n16447_), .A2(new_n16448_), .B(new_n16446_), .ZN(new_n16456_));
  NOR3_X1    g15433(.A1(new_n16444_), .A2(new_n16419_), .A3(new_n16441_), .ZN(new_n16457_));
  NOR2_X1    g15434(.A1(new_n16456_), .A2(new_n16457_), .ZN(new_n16458_));
  NOR2_X1    g15435(.A1(new_n16451_), .A2(new_n16458_), .ZN(new_n16459_));
  NAND2_X1   g15436(.A1(new_n16451_), .A2(new_n16458_), .ZN(new_n16460_));
  INV_X1     g15437(.I(new_n16460_), .ZN(new_n16461_));
  OAI21_X1   g15438(.A1(new_n16461_), .A2(new_n16459_), .B(new_n16417_), .ZN(new_n16462_));
  NAND2_X1   g15439(.A1(new_n16455_), .A2(new_n16462_), .ZN(new_n16463_));
  NOR2_X1    g15440(.A1(new_n14410_), .A2(new_n14393_), .ZN(new_n16464_));
  INV_X1     g15441(.I(new_n16464_), .ZN(new_n16465_));
  NOR2_X1    g15442(.A1(new_n14365_), .A2(new_n14342_), .ZN(new_n16466_));
  NAND2_X1   g15443(.A1(new_n14370_), .A2(new_n14367_), .ZN(new_n16467_));
  NAND2_X1   g15444(.A1(new_n14374_), .A2(new_n14371_), .ZN(new_n16468_));
  XOR2_X1    g15445(.A1(new_n16468_), .A2(new_n16467_), .Z(new_n16469_));
  NAND2_X1   g15446(.A1(new_n14347_), .A2(new_n14345_), .ZN(new_n16470_));
  NAND2_X1   g15447(.A1(new_n14351_), .A2(new_n14348_), .ZN(new_n16471_));
  XOR2_X1    g15448(.A1(new_n16470_), .A2(new_n16471_), .Z(new_n16472_));
  AND4_X2    g15449(.A1(new_n14343_), .A2(new_n16466_), .A3(new_n16469_), .A4(new_n16472_), .Z(new_n16473_));
  NAND2_X1   g15450(.A1(new_n14365_), .A2(new_n14378_), .ZN(new_n16474_));
  OAI21_X1   g15451(.A1(new_n4566_), .A2(new_n4598_), .B(new_n14342_), .ZN(new_n16475_));
  AND2_X2    g15452(.A1(new_n16475_), .A2(new_n16474_), .Z(new_n16476_));
  NAND3_X1   g15453(.A1(new_n16473_), .A2(new_n16476_), .A3(new_n14366_), .ZN(new_n16477_));
  NAND2_X1   g15454(.A1(new_n16475_), .A2(new_n14353_), .ZN(new_n16478_));
  NOR2_X1    g15455(.A1(new_n16470_), .A2(new_n16471_), .ZN(new_n16479_));
  INV_X1     g15456(.I(new_n16479_), .ZN(new_n16480_));
  NAND2_X1   g15457(.A1(new_n16478_), .A2(new_n16480_), .ZN(new_n16481_));
  NAND2_X1   g15458(.A1(new_n16474_), .A2(new_n14376_), .ZN(new_n16482_));
  NAND4_X1   g15459(.A1(new_n14374_), .A2(new_n14370_), .A3(new_n14367_), .A4(new_n14371_), .ZN(new_n16483_));
  NAND2_X1   g15460(.A1(new_n16482_), .A2(new_n16483_), .ZN(new_n16484_));
  NOR2_X1    g15461(.A1(new_n16481_), .A2(new_n16484_), .ZN(new_n16485_));
  NAND2_X1   g15462(.A1(new_n16477_), .A2(new_n16485_), .ZN(new_n16486_));
  INV_X1     g15463(.I(new_n16486_), .ZN(new_n16487_));
  NOR2_X1    g15464(.A1(new_n16477_), .A2(new_n16485_), .ZN(new_n16488_));
  OAI21_X1   g15465(.A1(new_n16487_), .A2(new_n16488_), .B(new_n16465_), .ZN(new_n16489_));
  INV_X1     g15466(.I(new_n16488_), .ZN(new_n16490_));
  NAND3_X1   g15467(.A1(new_n16490_), .A2(new_n16486_), .A3(new_n16464_), .ZN(new_n16491_));
  NAND2_X1   g15468(.A1(new_n16489_), .A2(new_n16491_), .ZN(new_n16492_));
  NOR2_X1    g15469(.A1(new_n14335_), .A2(new_n14274_), .ZN(new_n16493_));
  INV_X1     g15470(.I(new_n16493_), .ZN(new_n16494_));
  NAND2_X1   g15471(.A1(new_n14294_), .A2(new_n14302_), .ZN(new_n16495_));
  XNOR2_X1   g15472(.A1(new_n14314_), .A2(new_n14315_), .ZN(new_n16496_));
  NAND2_X1   g15473(.A1(new_n14283_), .A2(new_n14281_), .ZN(new_n16497_));
  NAND2_X1   g15474(.A1(new_n14287_), .A2(new_n14284_), .ZN(new_n16498_));
  XNOR2_X1   g15475(.A1(new_n16497_), .A2(new_n16498_), .ZN(new_n16499_));
  NOR4_X1    g15476(.A1(new_n16495_), .A2(new_n14291_), .A3(new_n16496_), .A4(new_n16499_), .ZN(new_n16500_));
  NOR2_X1    g15477(.A1(new_n14313_), .A2(new_n14302_), .ZN(new_n16501_));
  AOI21_X1   g15478(.A1(new_n14278_), .A2(new_n14291_), .B(new_n16501_), .ZN(new_n16502_));
  NAND3_X1   g15479(.A1(new_n16500_), .A2(new_n14313_), .A3(new_n16502_), .ZN(new_n16503_));
  OAI21_X1   g15480(.A1(new_n14294_), .A2(new_n14279_), .B(new_n14289_), .ZN(new_n16504_));
  NAND4_X1   g15481(.A1(new_n14283_), .A2(new_n14287_), .A3(new_n14281_), .A4(new_n14284_), .ZN(new_n16505_));
  AND2_X2    g15482(.A1(new_n16504_), .A2(new_n16505_), .Z(new_n16506_));
  OAI21_X1   g15483(.A1(new_n14313_), .A2(new_n14302_), .B(new_n14316_), .ZN(new_n16507_));
  NAND4_X1   g15484(.A1(new_n14306_), .A2(new_n14310_), .A3(new_n14303_), .A4(new_n14307_), .ZN(new_n16508_));
  NAND2_X1   g15485(.A1(new_n16507_), .A2(new_n16508_), .ZN(new_n16509_));
  INV_X1     g15486(.I(new_n16509_), .ZN(new_n16510_));
  NAND3_X1   g15487(.A1(new_n16503_), .A2(new_n16506_), .A3(new_n16510_), .ZN(new_n16511_));
  INV_X1     g15488(.I(new_n16511_), .ZN(new_n16512_));
  AOI21_X1   g15489(.A1(new_n16510_), .A2(new_n16506_), .B(new_n16503_), .ZN(new_n16513_));
  OAI21_X1   g15490(.A1(new_n16512_), .A2(new_n16513_), .B(new_n16494_), .ZN(new_n16514_));
  INV_X1     g15491(.I(new_n16503_), .ZN(new_n16515_));
  NAND2_X1   g15492(.A1(new_n16506_), .A2(new_n16510_), .ZN(new_n16516_));
  NAND2_X1   g15493(.A1(new_n16515_), .A2(new_n16516_), .ZN(new_n16517_));
  NAND3_X1   g15494(.A1(new_n16517_), .A2(new_n16493_), .A3(new_n16511_), .ZN(new_n16518_));
  NAND2_X1   g15495(.A1(new_n16514_), .A2(new_n16518_), .ZN(new_n16519_));
  INV_X1     g15496(.I(new_n14417_), .ZN(new_n16520_));
  AOI22_X1   g15497(.A1(new_n14412_), .A2(new_n14337_), .B1(new_n14272_), .B2(new_n4776_), .ZN(new_n16521_));
  NOR2_X1    g15498(.A1(new_n16521_), .A2(new_n16520_), .ZN(new_n16522_));
  NOR2_X1    g15499(.A1(new_n16522_), .A2(new_n16519_), .ZN(new_n16523_));
  AOI21_X1   g15500(.A1(new_n16517_), .A2(new_n16511_), .B(new_n16493_), .ZN(new_n16524_));
  NOR3_X1    g15501(.A1(new_n16512_), .A2(new_n16494_), .A3(new_n16513_), .ZN(new_n16525_));
  NOR2_X1    g15502(.A1(new_n16525_), .A2(new_n16524_), .ZN(new_n16526_));
  NOR3_X1    g15503(.A1(new_n16521_), .A2(new_n16526_), .A3(new_n16520_), .ZN(new_n16527_));
  OAI21_X1   g15504(.A1(new_n16523_), .A2(new_n16527_), .B(new_n16492_), .ZN(new_n16528_));
  INV_X1     g15505(.I(new_n16492_), .ZN(new_n16529_));
  NAND2_X1   g15506(.A1(new_n14273_), .A2(new_n14416_), .ZN(new_n16530_));
  AOI21_X1   g15507(.A1(new_n16530_), .A2(new_n14417_), .B(new_n16526_), .ZN(new_n16531_));
  NOR3_X1    g15508(.A1(new_n16521_), .A2(new_n16519_), .A3(new_n16520_), .ZN(new_n16532_));
  OAI21_X1   g15509(.A1(new_n16531_), .A2(new_n16532_), .B(new_n16529_), .ZN(new_n16533_));
  NAND2_X1   g15510(.A1(new_n16528_), .A2(new_n16533_), .ZN(new_n16534_));
  AOI21_X1   g15511(.A1(new_n14271_), .A2(new_n14604_), .B(new_n14589_), .ZN(new_n16535_));
  NOR2_X1    g15512(.A1(new_n16534_), .A2(new_n16535_), .ZN(new_n16536_));
  NAND2_X1   g15513(.A1(new_n16530_), .A2(new_n14417_), .ZN(new_n16537_));
  NAND2_X1   g15514(.A1(new_n16537_), .A2(new_n16526_), .ZN(new_n16538_));
  NAND3_X1   g15515(.A1(new_n16530_), .A2(new_n16519_), .A3(new_n14417_), .ZN(new_n16539_));
  NAND2_X1   g15516(.A1(new_n16538_), .A2(new_n16539_), .ZN(new_n16540_));
  OAI21_X1   g15517(.A1(new_n16521_), .A2(new_n16520_), .B(new_n16519_), .ZN(new_n16541_));
  NAND3_X1   g15518(.A1(new_n16530_), .A2(new_n16526_), .A3(new_n14417_), .ZN(new_n16542_));
  AOI21_X1   g15519(.A1(new_n16541_), .A2(new_n16542_), .B(new_n16492_), .ZN(new_n16543_));
  AOI21_X1   g15520(.A1(new_n16540_), .A2(new_n16492_), .B(new_n16543_), .ZN(new_n16544_));
  OAI21_X1   g15521(.A1(new_n14588_), .A2(new_n14587_), .B(new_n14605_), .ZN(new_n16545_));
  NOR2_X1    g15522(.A1(new_n16545_), .A2(new_n16544_), .ZN(new_n16546_));
  OAI21_X1   g15523(.A1(new_n16546_), .A2(new_n16536_), .B(new_n16463_), .ZN(new_n16547_));
  OAI21_X1   g15524(.A1(new_n14421_), .A2(new_n14581_), .B(new_n14569_), .ZN(new_n16548_));
  NAND2_X1   g15525(.A1(new_n16548_), .A2(new_n16458_), .ZN(new_n16549_));
  AOI21_X1   g15526(.A1(new_n16549_), .A2(new_n16453_), .B(new_n16417_), .ZN(new_n16550_));
  NOR2_X1    g15527(.A1(new_n14581_), .A2(new_n14421_), .ZN(new_n16551_));
  OAI21_X1   g15528(.A1(new_n16551_), .A2(new_n14582_), .B(new_n16450_), .ZN(new_n16552_));
  AOI21_X1   g15529(.A1(new_n16552_), .A2(new_n16460_), .B(new_n16418_), .ZN(new_n16553_));
  NOR2_X1    g15530(.A1(new_n16550_), .A2(new_n16553_), .ZN(new_n16554_));
  NOR2_X1    g15531(.A1(new_n16544_), .A2(new_n16535_), .ZN(new_n16555_));
  NOR2_X1    g15532(.A1(new_n16545_), .A2(new_n16534_), .ZN(new_n16556_));
  OAI21_X1   g15533(.A1(new_n16556_), .A2(new_n16555_), .B(new_n16554_), .ZN(new_n16557_));
  NAND2_X1   g15534(.A1(new_n16547_), .A2(new_n16557_), .ZN(new_n16558_));
  NAND2_X1   g15535(.A1(new_n14115_), .A2(new_n14254_), .ZN(new_n16559_));
  OAI21_X1   g15536(.A1(new_n14113_), .A2(new_n14255_), .B(new_n16559_), .ZN(new_n16560_));
  NOR2_X1    g15537(.A1(new_n14246_), .A2(new_n14228_), .ZN(new_n16561_));
  NOR2_X1    g15538(.A1(new_n14203_), .A2(new_n14179_), .ZN(new_n16562_));
  XOR2_X1    g15539(.A1(new_n14210_), .A2(new_n14207_), .Z(new_n16563_));
  NAND2_X1   g15540(.A1(new_n14185_), .A2(new_n14182_), .ZN(new_n16564_));
  NAND2_X1   g15541(.A1(new_n14189_), .A2(new_n14186_), .ZN(new_n16565_));
  XOR2_X1    g15542(.A1(new_n16564_), .A2(new_n16565_), .Z(new_n16566_));
  NAND4_X1   g15543(.A1(new_n16566_), .A2(new_n16562_), .A3(new_n14192_), .A4(new_n16563_), .ZN(new_n16567_));
  NAND2_X1   g15544(.A1(new_n14213_), .A2(new_n14203_), .ZN(new_n16568_));
  NAND2_X1   g15545(.A1(new_n14181_), .A2(new_n14179_), .ZN(new_n16569_));
  NAND2_X1   g15546(.A1(new_n16569_), .A2(new_n16568_), .ZN(new_n16570_));
  NOR3_X1    g15547(.A1(new_n16567_), .A2(new_n16570_), .A3(new_n14213_), .ZN(new_n16571_));
  INV_X1     g15548(.I(new_n16571_), .ZN(new_n16572_));
  AOI21_X1   g15549(.A1(new_n14181_), .A2(new_n14179_), .B(new_n14190_), .ZN(new_n16573_));
  NAND4_X1   g15550(.A1(new_n14185_), .A2(new_n14182_), .A3(new_n14186_), .A4(new_n14189_), .ZN(new_n16574_));
  INV_X1     g15551(.I(new_n16574_), .ZN(new_n16575_));
  NOR2_X1    g15552(.A1(new_n16573_), .A2(new_n16575_), .ZN(new_n16576_));
  INV_X1     g15553(.I(new_n16576_), .ZN(new_n16577_));
  AOI21_X1   g15554(.A1(new_n14213_), .A2(new_n14203_), .B(new_n14214_), .ZN(new_n16578_));
  NOR2_X1    g15555(.A1(new_n14210_), .A2(new_n14207_), .ZN(new_n16579_));
  NOR2_X1    g15556(.A1(new_n16578_), .A2(new_n16579_), .ZN(new_n16580_));
  INV_X1     g15557(.I(new_n16580_), .ZN(new_n16581_));
  NOR2_X1    g15558(.A1(new_n16577_), .A2(new_n16581_), .ZN(new_n16582_));
  NAND2_X1   g15559(.A1(new_n16572_), .A2(new_n16582_), .ZN(new_n16583_));
  NOR2_X1    g15560(.A1(new_n16572_), .A2(new_n16582_), .ZN(new_n16584_));
  INV_X1     g15561(.I(new_n16584_), .ZN(new_n16585_));
  AOI21_X1   g15562(.A1(new_n16585_), .A2(new_n16583_), .B(new_n16561_), .ZN(new_n16586_));
  NAND3_X1   g15563(.A1(new_n16585_), .A2(new_n16561_), .A3(new_n16583_), .ZN(new_n16587_));
  INV_X1     g15564(.I(new_n16587_), .ZN(new_n16588_));
  NOR2_X1    g15565(.A1(new_n16588_), .A2(new_n16586_), .ZN(new_n16589_));
  INV_X1     g15566(.I(new_n16589_), .ZN(new_n16590_));
  NAND2_X1   g15567(.A1(new_n14128_), .A2(new_n14126_), .ZN(new_n16591_));
  NAND2_X1   g15568(.A1(new_n14123_), .A2(new_n16591_), .ZN(new_n16592_));
  NAND2_X1   g15569(.A1(new_n14131_), .A2(new_n14129_), .ZN(new_n16593_));
  NAND2_X1   g15570(.A1(new_n14134_), .A2(new_n16593_), .ZN(new_n16594_));
  NAND2_X1   g15571(.A1(new_n16592_), .A2(new_n16594_), .ZN(new_n16595_));
  NOR2_X1    g15572(.A1(new_n16591_), .A2(new_n16593_), .ZN(new_n16596_));
  NOR2_X1    g15573(.A1(new_n16595_), .A2(new_n16596_), .ZN(new_n16597_));
  NAND2_X1   g15574(.A1(new_n14145_), .A2(new_n14151_), .ZN(new_n16598_));
  NAND2_X1   g15575(.A1(new_n14147_), .A2(new_n14154_), .ZN(new_n16599_));
  NAND2_X1   g15576(.A1(new_n16599_), .A2(new_n16598_), .ZN(new_n16600_));
  NOR2_X1    g15577(.A1(new_n14151_), .A2(new_n14154_), .ZN(new_n16601_));
  NOR2_X1    g15578(.A1(new_n16600_), .A2(new_n16601_), .ZN(new_n16602_));
  XOR2_X1    g15579(.A1(new_n16597_), .A2(new_n16602_), .Z(new_n16603_));
  NOR2_X1    g15580(.A1(new_n14239_), .A2(new_n14117_), .ZN(new_n16604_));
  NOR2_X1    g15581(.A1(new_n14147_), .A2(new_n14145_), .ZN(new_n16605_));
  XOR2_X1    g15582(.A1(new_n14151_), .A2(new_n14154_), .Z(new_n16606_));
  XOR2_X1    g15583(.A1(new_n16591_), .A2(new_n16593_), .Z(new_n16607_));
  NAND4_X1   g15584(.A1(new_n16607_), .A2(new_n16606_), .A3(new_n14123_), .A4(new_n14145_), .ZN(new_n16608_));
  OAI21_X1   g15585(.A1(new_n14123_), .A2(new_n14134_), .B(new_n14147_), .ZN(new_n16609_));
  NOR4_X1    g15586(.A1(new_n16608_), .A2(new_n14124_), .A3(new_n16605_), .A4(new_n16609_), .ZN(new_n16610_));
  OAI21_X1   g15587(.A1(new_n16604_), .A2(new_n16610_), .B(new_n16603_), .ZN(new_n16611_));
  AOI21_X1   g15588(.A1(new_n14250_), .A2(new_n14251_), .B(new_n14260_), .ZN(new_n16612_));
  NOR2_X1    g15589(.A1(new_n16612_), .A2(new_n16611_), .ZN(new_n16613_));
  INV_X1     g15590(.I(new_n16611_), .ZN(new_n16614_));
  OAI21_X1   g15591(.A1(new_n14259_), .A2(new_n14116_), .B(new_n14252_), .ZN(new_n16615_));
  NOR2_X1    g15592(.A1(new_n16615_), .A2(new_n16614_), .ZN(new_n16616_));
  OAI21_X1   g15593(.A1(new_n16616_), .A2(new_n16613_), .B(new_n16590_), .ZN(new_n16617_));
  NOR2_X1    g15594(.A1(new_n16612_), .A2(new_n16614_), .ZN(new_n16618_));
  NOR2_X1    g15595(.A1(new_n16615_), .A2(new_n16611_), .ZN(new_n16619_));
  OAI21_X1   g15596(.A1(new_n16619_), .A2(new_n16618_), .B(new_n16589_), .ZN(new_n16620_));
  NAND2_X1   g15597(.A1(new_n16617_), .A2(new_n16620_), .ZN(new_n16621_));
  AOI21_X1   g15598(.A1(new_n14108_), .A2(new_n14099_), .B(new_n14101_), .ZN(new_n16622_));
  OAI21_X1   g15599(.A1(new_n13992_), .A2(new_n14000_), .B(new_n13991_), .ZN(new_n16623_));
  XNOR2_X1   g15600(.A1(new_n13990_), .A2(new_n13988_), .ZN(new_n16624_));
  INV_X1     g15601(.I(new_n14000_), .ZN(new_n16625_));
  NOR2_X1    g15602(.A1(new_n16624_), .A2(new_n16625_), .ZN(new_n16626_));
  XNOR2_X1   g15603(.A1(new_n14011_), .A2(new_n14015_), .ZN(new_n16627_));
  NOR2_X1    g15604(.A1(new_n16627_), .A2(new_n14006_), .ZN(new_n16628_));
  NAND4_X1   g15605(.A1(new_n16626_), .A2(new_n13992_), .A3(new_n16628_), .A4(new_n14007_), .ZN(new_n16629_));
  OAI21_X1   g15606(.A1(new_n5055_), .A2(new_n5087_), .B(new_n14006_), .ZN(new_n16630_));
  INV_X1     g15607(.I(new_n16630_), .ZN(new_n16631_));
  NOR3_X1    g15608(.A1(new_n16629_), .A2(new_n16623_), .A3(new_n16631_), .ZN(new_n16632_));
  NOR2_X1    g15609(.A1(new_n14024_), .A2(new_n14001_), .ZN(new_n16633_));
  NOR2_X1    g15610(.A1(new_n14011_), .A2(new_n14015_), .ZN(new_n16634_));
  AOI21_X1   g15611(.A1(new_n16630_), .A2(new_n14016_), .B(new_n16634_), .ZN(new_n16635_));
  NAND2_X1   g15612(.A1(new_n14000_), .A2(new_n13988_), .ZN(new_n16636_));
  NAND2_X1   g15613(.A1(new_n13992_), .A2(new_n13990_), .ZN(new_n16637_));
  NOR2_X1    g15614(.A1(new_n13990_), .A2(new_n13988_), .ZN(new_n16638_));
  INV_X1     g15615(.I(new_n16638_), .ZN(new_n16639_));
  NAND4_X1   g15616(.A1(new_n16635_), .A2(new_n16637_), .A3(new_n16636_), .A4(new_n16639_), .ZN(new_n16640_));
  INV_X1     g15617(.I(new_n16640_), .ZN(new_n16641_));
  OAI21_X1   g15618(.A1(new_n16633_), .A2(new_n14002_), .B(new_n16641_), .ZN(new_n16642_));
  NAND3_X1   g15619(.A1(new_n14030_), .A2(new_n14020_), .A3(new_n14023_), .ZN(new_n16643_));
  NAND3_X1   g15620(.A1(new_n14027_), .A2(new_n16643_), .A3(new_n16640_), .ZN(new_n16644_));
  AOI21_X1   g15621(.A1(new_n16642_), .A2(new_n16644_), .B(new_n16632_), .ZN(new_n16645_));
  INV_X1     g15622(.I(new_n16632_), .ZN(new_n16646_));
  AOI21_X1   g15623(.A1(new_n14027_), .A2(new_n16643_), .B(new_n16640_), .ZN(new_n16647_));
  NOR3_X1    g15624(.A1(new_n16633_), .A2(new_n16641_), .A3(new_n14002_), .ZN(new_n16648_));
  NOR3_X1    g15625(.A1(new_n16648_), .A2(new_n16647_), .A3(new_n16646_), .ZN(new_n16649_));
  NAND2_X1   g15626(.A1(new_n14042_), .A2(new_n14054_), .ZN(new_n16650_));
  NAND2_X1   g15627(.A1(new_n14053_), .A2(new_n14055_), .ZN(new_n16651_));
  NAND2_X1   g15628(.A1(new_n16651_), .A2(new_n16650_), .ZN(new_n16652_));
  NOR2_X1    g15629(.A1(new_n14054_), .A2(new_n14055_), .ZN(new_n16653_));
  NOR2_X1    g15630(.A1(new_n16652_), .A2(new_n16653_), .ZN(new_n16654_));
  NAND2_X1   g15631(.A1(new_n14067_), .A2(new_n14072_), .ZN(new_n16655_));
  NAND2_X1   g15632(.A1(new_n14078_), .A2(new_n14076_), .ZN(new_n16656_));
  NAND2_X1   g15633(.A1(new_n14080_), .A2(new_n14079_), .ZN(new_n16657_));
  NAND3_X1   g15634(.A1(new_n16657_), .A2(new_n16655_), .A3(new_n16656_), .ZN(new_n16658_));
  XOR2_X1    g15635(.A1(new_n16654_), .A2(new_n16658_), .Z(new_n16659_));
  OAI21_X1   g15636(.A1(new_n14063_), .A2(new_n14092_), .B(new_n14037_), .ZN(new_n16660_));
  NOR2_X1    g15637(.A1(new_n14067_), .A2(new_n14078_), .ZN(new_n16661_));
  XOR2_X1    g15638(.A1(new_n14076_), .A2(new_n14072_), .Z(new_n16662_));
  XOR2_X1    g15639(.A1(new_n14054_), .A2(new_n14055_), .Z(new_n16663_));
  NAND4_X1   g15640(.A1(new_n16662_), .A2(new_n14042_), .A3(new_n14067_), .A4(new_n16663_), .ZN(new_n16664_));
  AOI21_X1   g15641(.A1(new_n14059_), .A2(new_n14043_), .B(new_n14068_), .ZN(new_n16665_));
  INV_X1     g15642(.I(new_n16665_), .ZN(new_n16666_));
  NOR4_X1    g15643(.A1(new_n16664_), .A2(new_n14043_), .A3(new_n16661_), .A4(new_n16666_), .ZN(new_n16667_));
  INV_X1     g15644(.I(new_n16667_), .ZN(new_n16668_));
  AOI21_X1   g15645(.A1(new_n16668_), .A2(new_n16660_), .B(new_n16659_), .ZN(new_n16669_));
  NOR3_X1    g15646(.A1(new_n16645_), .A2(new_n16649_), .A3(new_n16669_), .ZN(new_n16670_));
  OAI21_X1   g15647(.A1(new_n16648_), .A2(new_n16647_), .B(new_n16646_), .ZN(new_n16671_));
  NAND3_X1   g15648(.A1(new_n16642_), .A2(new_n16644_), .A3(new_n16632_), .ZN(new_n16672_));
  INV_X1     g15649(.I(new_n16669_), .ZN(new_n16673_));
  AOI21_X1   g15650(.A1(new_n16671_), .A2(new_n16672_), .B(new_n16673_), .ZN(new_n16674_));
  NOR2_X1    g15651(.A1(new_n16674_), .A2(new_n16670_), .ZN(new_n16675_));
  NOR2_X1    g15652(.A1(new_n16675_), .A2(new_n16622_), .ZN(new_n16676_));
  INV_X1     g15653(.I(new_n14101_), .ZN(new_n16677_));
  NAND2_X1   g15654(.A1(new_n14108_), .A2(new_n14099_), .ZN(new_n16678_));
  NAND2_X1   g15655(.A1(new_n16678_), .A2(new_n16677_), .ZN(new_n16679_));
  AOI21_X1   g15656(.A1(new_n16671_), .A2(new_n16672_), .B(new_n16669_), .ZN(new_n16680_));
  NOR3_X1    g15657(.A1(new_n16645_), .A2(new_n16649_), .A3(new_n16673_), .ZN(new_n16681_));
  NOR2_X1    g15658(.A1(new_n16680_), .A2(new_n16681_), .ZN(new_n16682_));
  NOR2_X1    g15659(.A1(new_n16679_), .A2(new_n16682_), .ZN(new_n16683_));
  NOR2_X1    g15660(.A1(new_n16683_), .A2(new_n16676_), .ZN(new_n16684_));
  NOR2_X1    g15661(.A1(new_n16621_), .A2(new_n16684_), .ZN(new_n16685_));
  NAND2_X1   g15662(.A1(new_n16615_), .A2(new_n16614_), .ZN(new_n16686_));
  NAND2_X1   g15663(.A1(new_n16612_), .A2(new_n16611_), .ZN(new_n16687_));
  AOI21_X1   g15664(.A1(new_n16686_), .A2(new_n16687_), .B(new_n16589_), .ZN(new_n16688_));
  NAND2_X1   g15665(.A1(new_n16615_), .A2(new_n16611_), .ZN(new_n16689_));
  NAND2_X1   g15666(.A1(new_n16612_), .A2(new_n16614_), .ZN(new_n16690_));
  AOI21_X1   g15667(.A1(new_n16689_), .A2(new_n16690_), .B(new_n16590_), .ZN(new_n16691_));
  NOR2_X1    g15668(.A1(new_n16691_), .A2(new_n16688_), .ZN(new_n16692_));
  NOR2_X1    g15669(.A1(new_n14100_), .A2(new_n14035_), .ZN(new_n16693_));
  OAI22_X1   g15670(.A1(new_n16693_), .A2(new_n14101_), .B1(new_n16670_), .B2(new_n16674_), .ZN(new_n16694_));
  OAI21_X1   g15671(.A1(new_n16680_), .A2(new_n16681_), .B(new_n16622_), .ZN(new_n16695_));
  NAND2_X1   g15672(.A1(new_n16694_), .A2(new_n16695_), .ZN(new_n16696_));
  NOR2_X1    g15673(.A1(new_n16696_), .A2(new_n16692_), .ZN(new_n16697_));
  OAI21_X1   g15674(.A1(new_n16697_), .A2(new_n16685_), .B(new_n16560_), .ZN(new_n16698_));
  INV_X1     g15675(.I(new_n14113_), .ZN(new_n16699_));
  NAND3_X1   g15676(.A1(new_n14262_), .A2(new_n5341_), .A3(new_n14114_), .ZN(new_n16700_));
  AOI21_X1   g15677(.A1(new_n16699_), .A2(new_n16700_), .B(new_n14263_), .ZN(new_n16701_));
  AOI22_X1   g15678(.A1(new_n16694_), .A2(new_n16695_), .B1(new_n16617_), .B2(new_n16620_), .ZN(new_n16702_));
  NOR4_X1    g15679(.A1(new_n16683_), .A2(new_n16691_), .A3(new_n16688_), .A4(new_n16676_), .ZN(new_n16703_));
  OAI21_X1   g15680(.A1(new_n16702_), .A2(new_n16703_), .B(new_n16701_), .ZN(new_n16704_));
  AOI21_X1   g15681(.A1(new_n16698_), .A2(new_n16704_), .B(new_n16558_), .ZN(new_n16705_));
  NAND2_X1   g15682(.A1(new_n16698_), .A2(new_n16704_), .ZN(new_n16706_));
  AOI21_X1   g15683(.A1(new_n16547_), .A2(new_n16557_), .B(new_n16706_), .ZN(new_n16707_));
  OAI21_X1   g15684(.A1(new_n16705_), .A2(new_n16707_), .B(new_n16389_), .ZN(new_n16708_));
  NAND2_X1   g15685(.A1(new_n16545_), .A2(new_n16544_), .ZN(new_n16709_));
  NAND2_X1   g15686(.A1(new_n16534_), .A2(new_n16535_), .ZN(new_n16710_));
  AOI21_X1   g15687(.A1(new_n16709_), .A2(new_n16710_), .B(new_n16554_), .ZN(new_n16711_));
  NAND2_X1   g15688(.A1(new_n16545_), .A2(new_n16534_), .ZN(new_n16712_));
  NAND2_X1   g15689(.A1(new_n16544_), .A2(new_n16535_), .ZN(new_n16713_));
  AOI21_X1   g15690(.A1(new_n16712_), .A2(new_n16713_), .B(new_n16463_), .ZN(new_n16714_));
  NAND2_X1   g15691(.A1(new_n16696_), .A2(new_n16692_), .ZN(new_n16715_));
  NAND2_X1   g15692(.A1(new_n16621_), .A2(new_n16684_), .ZN(new_n16716_));
  AOI21_X1   g15693(.A1(new_n16715_), .A2(new_n16716_), .B(new_n16701_), .ZN(new_n16717_));
  OAI22_X1   g15694(.A1(new_n16676_), .A2(new_n16683_), .B1(new_n16691_), .B2(new_n16688_), .ZN(new_n16718_));
  NAND4_X1   g15695(.A1(new_n16617_), .A2(new_n16694_), .A3(new_n16695_), .A4(new_n16620_), .ZN(new_n16719_));
  AOI21_X1   g15696(.A1(new_n16718_), .A2(new_n16719_), .B(new_n16560_), .ZN(new_n16720_));
  NOR4_X1    g15697(.A1(new_n16711_), .A2(new_n16714_), .A3(new_n16717_), .A4(new_n16720_), .ZN(new_n16721_));
  AOI22_X1   g15698(.A1(new_n16547_), .A2(new_n16557_), .B1(new_n16698_), .B2(new_n16704_), .ZN(new_n16722_));
  OAI21_X1   g15699(.A1(new_n16722_), .A2(new_n16721_), .B(new_n16388_), .ZN(new_n16723_));
  NAND2_X1   g15700(.A1(new_n16708_), .A2(new_n16723_), .ZN(new_n16724_));
  XOR2_X1    g15701(.A1(new_n16724_), .A2(new_n16387_), .Z(new_n16725_));
  NAND2_X1   g15702(.A1(new_n16725_), .A2(new_n16386_), .ZN(new_n16726_));
  INV_X1     g15703(.I(new_n16386_), .ZN(new_n16727_));
  AOI21_X1   g15704(.A1(new_n15817_), .A2(new_n14613_), .B(new_n15831_), .ZN(new_n16728_));
  XOR2_X1    g15705(.A1(new_n16724_), .A2(new_n16728_), .Z(new_n16729_));
  NAND2_X1   g15706(.A1(new_n16729_), .A2(new_n16727_), .ZN(new_n16730_));
  NAND3_X1   g15707(.A1(new_n16730_), .A2(new_n16726_), .A3(new_n15854_), .ZN(new_n16731_));
  NOR2_X1    g15708(.A1(new_n15830_), .A2(new_n15845_), .ZN(new_n16732_));
  NAND2_X1   g15709(.A1(new_n15830_), .A2(new_n15845_), .ZN(new_n16733_));
  NOR2_X1    g15710(.A1(new_n14610_), .A2(new_n15833_), .ZN(new_n16734_));
  AOI21_X1   g15711(.A1(new_n16733_), .A2(new_n16734_), .B(new_n16732_), .ZN(new_n16735_));
  XOR2_X1    g15712(.A1(new_n16724_), .A2(new_n16728_), .Z(new_n16736_));
  NOR2_X1    g15713(.A1(new_n16736_), .A2(new_n16727_), .ZN(new_n16737_));
  XOR2_X1    g15714(.A1(new_n16724_), .A2(new_n16387_), .Z(new_n16738_));
  NOR2_X1    g15715(.A1(new_n16738_), .A2(new_n16386_), .ZN(new_n16739_));
  OAI21_X1   g15716(.A1(new_n16737_), .A2(new_n16739_), .B(new_n16735_), .ZN(new_n16740_));
  AOI21_X1   g15717(.A1(new_n16740_), .A2(new_n16731_), .B(new_n15849_), .ZN(new_n16741_));
  NOR3_X1    g15718(.A1(new_n16377_), .A2(new_n16376_), .A3(new_n16384_), .ZN(new_n16742_));
  AOI21_X1   g15719(.A1(new_n16038_), .A2(new_n16041_), .B(new_n16374_), .ZN(new_n16743_));
  NOR2_X1    g15720(.A1(new_n16743_), .A2(new_n16728_), .ZN(new_n16744_));
  NOR2_X1    g15721(.A1(new_n16744_), .A2(new_n16742_), .ZN(new_n16745_));
  AOI21_X1   g15722(.A1(new_n16370_), .A2(new_n16372_), .B(new_n16381_), .ZN(new_n16746_));
  OAI21_X1   g15723(.A1(new_n16348_), .A2(new_n16349_), .B(new_n16365_), .ZN(new_n16747_));
  INV_X1     g15724(.I(new_n16310_), .ZN(new_n16748_));
  INV_X1     g15725(.I(new_n16311_), .ZN(new_n16749_));
  NAND3_X1   g15726(.A1(new_n16315_), .A2(new_n16748_), .A3(new_n16749_), .ZN(new_n16750_));
  NAND2_X1   g15727(.A1(new_n16748_), .A2(new_n16749_), .ZN(new_n16751_));
  NAND2_X1   g15728(.A1(new_n16751_), .A2(new_n16314_), .ZN(new_n16752_));
  OAI22_X1   g15729(.A1(new_n16750_), .A2(new_n16308_), .B1(new_n16298_), .B2(new_n16752_), .ZN(new_n16753_));
  INV_X1     g15730(.I(new_n16751_), .ZN(new_n16754_));
  NAND2_X1   g15731(.A1(new_n16754_), .A2(new_n16315_), .ZN(new_n16755_));
  NAND2_X1   g15732(.A1(new_n16755_), .A2(new_n16752_), .ZN(new_n16756_));
  NAND2_X1   g15733(.A1(new_n14767_), .A2(new_n14758_), .ZN(new_n16757_));
  NAND2_X1   g15734(.A1(new_n16283_), .A2(new_n16286_), .ZN(new_n16758_));
  XOR2_X1    g15735(.A1(new_n16758_), .A2(new_n16288_), .Z(new_n16759_));
  NOR4_X1    g15736(.A1(new_n16757_), .A2(new_n16759_), .A3(new_n16308_), .A4(new_n16282_), .ZN(new_n16760_));
  AOI21_X1   g15737(.A1(new_n14767_), .A2(new_n14758_), .B(new_n16281_), .ZN(new_n16761_));
  NOR2_X1    g15738(.A1(new_n16298_), .A2(new_n16761_), .ZN(new_n16762_));
  NAND4_X1   g15739(.A1(new_n16753_), .A2(new_n16756_), .A3(new_n16760_), .A4(new_n16762_), .ZN(new_n16763_));
  NOR2_X1    g15740(.A1(new_n16312_), .A2(new_n16311_), .ZN(new_n16764_));
  OAI21_X1   g15741(.A1(new_n16306_), .A2(new_n14666_), .B(new_n16764_), .ZN(new_n16765_));
  OAI22_X1   g15742(.A1(new_n16321_), .A2(new_n16323_), .B1(new_n16310_), .B2(new_n16765_), .ZN(new_n16766_));
  NAND2_X1   g15743(.A1(new_n16315_), .A2(new_n16751_), .ZN(new_n16767_));
  INV_X1     g15744(.I(new_n16758_), .ZN(new_n16768_));
  NOR2_X1    g15745(.A1(new_n16274_), .A2(new_n16273_), .ZN(new_n16769_));
  NOR2_X1    g15746(.A1(new_n16768_), .A2(new_n16288_), .ZN(new_n16770_));
  AOI21_X1   g15747(.A1(new_n16770_), .A2(new_n16769_), .B(new_n16281_), .ZN(new_n16771_));
  NOR2_X1    g15748(.A1(new_n16771_), .A2(new_n16757_), .ZN(new_n16772_));
  NAND3_X1   g15749(.A1(new_n16766_), .A2(new_n16767_), .A3(new_n16772_), .ZN(new_n16773_));
  AOI21_X1   g15750(.A1(new_n16342_), .A2(new_n16329_), .B(new_n16773_), .ZN(new_n16774_));
  NOR3_X1    g15751(.A1(new_n16319_), .A2(new_n16318_), .A3(new_n16316_), .ZN(new_n16775_));
  NOR2_X1    g15752(.A1(new_n16765_), .A2(new_n16310_), .ZN(new_n16776_));
  AOI21_X1   g15753(.A1(new_n16298_), .A2(new_n16308_), .B(new_n16776_), .ZN(new_n16777_));
  INV_X1     g15754(.I(new_n16767_), .ZN(new_n16778_));
  NOR4_X1    g15755(.A1(new_n16777_), .A2(new_n16778_), .A3(new_n16757_), .A4(new_n16771_), .ZN(new_n16779_));
  NOR3_X1    g15756(.A1(new_n16327_), .A2(new_n16775_), .A3(new_n16779_), .ZN(new_n16780_));
  OAI21_X1   g15757(.A1(new_n16774_), .A2(new_n16780_), .B(new_n16763_), .ZN(new_n16781_));
  INV_X1     g15758(.I(new_n16763_), .ZN(new_n16782_));
  OAI21_X1   g15759(.A1(new_n16327_), .A2(new_n16775_), .B(new_n16779_), .ZN(new_n16783_));
  NAND4_X1   g15760(.A1(new_n16268_), .A2(new_n14951_), .A3(new_n16773_), .A4(new_n16329_), .ZN(new_n16784_));
  NAND3_X1   g15761(.A1(new_n16783_), .A2(new_n16784_), .A3(new_n16782_), .ZN(new_n16785_));
  NAND2_X1   g15762(.A1(new_n16781_), .A2(new_n16785_), .ZN(new_n16786_));
  INV_X1     g15763(.I(new_n16248_), .ZN(new_n16787_));
  NAND2_X1   g15764(.A1(new_n16246_), .A2(new_n16787_), .ZN(new_n16788_));
  INV_X1     g15765(.I(new_n16788_), .ZN(new_n16789_));
  NOR2_X1    g15766(.A1(new_n16251_), .A2(new_n16789_), .ZN(new_n16790_));
  INV_X1     g15767(.I(new_n16790_), .ZN(new_n16791_));
  NOR3_X1    g15768(.A1(new_n16250_), .A2(new_n16247_), .A3(new_n16248_), .ZN(new_n16792_));
  NAND2_X1   g15769(.A1(new_n16244_), .A2(new_n16792_), .ZN(new_n16793_));
  OAI21_X1   g15770(.A1(new_n16791_), .A2(new_n16234_), .B(new_n16793_), .ZN(new_n16794_));
  NAND2_X1   g15771(.A1(new_n16220_), .A2(new_n16215_), .ZN(new_n16795_));
  NOR2_X1    g15772(.A1(new_n16250_), .A2(new_n16788_), .ZN(new_n16796_));
  NOR2_X1    g15773(.A1(new_n16790_), .A2(new_n16796_), .ZN(new_n16797_));
  XOR2_X1    g15774(.A1(new_n16223_), .A2(new_n16227_), .Z(new_n16798_));
  NAND3_X1   g15775(.A1(new_n16798_), .A2(new_n16244_), .A3(new_n16214_), .ZN(new_n16799_));
  NOR3_X1    g15776(.A1(new_n16797_), .A2(new_n16799_), .A3(new_n16220_), .ZN(new_n16800_));
  NAND4_X1   g15777(.A1(new_n16800_), .A2(new_n16794_), .A3(new_n16257_), .A4(new_n16795_), .ZN(new_n16801_));
  INV_X1     g15778(.I(new_n16801_), .ZN(new_n16802_));
  AOI21_X1   g15779(.A1(new_n14820_), .A2(new_n14823_), .B(new_n16248_), .ZN(new_n16803_));
  OAI21_X1   g15780(.A1(new_n16242_), .A2(new_n14824_), .B(new_n16803_), .ZN(new_n16804_));
  NOR2_X1    g15781(.A1(new_n16247_), .A2(new_n16804_), .ZN(new_n16805_));
  AOI21_X1   g15782(.A1(new_n16234_), .A2(new_n16245_), .B(new_n16805_), .ZN(new_n16806_));
  NOR2_X1    g15783(.A1(new_n16789_), .A2(new_n16250_), .ZN(new_n16807_));
  OAI22_X1   g15784(.A1(new_n16207_), .A2(new_n14898_), .B1(new_n16208_), .B2(new_n14894_), .ZN(new_n16808_));
  OAI21_X1   g15785(.A1(new_n16221_), .A2(new_n14874_), .B(new_n16808_), .ZN(new_n16809_));
  AOI21_X1   g15786(.A1(new_n14904_), .A2(new_n16212_), .B(new_n16809_), .ZN(new_n16810_));
  NOR4_X1    g15787(.A1(new_n16216_), .A2(new_n16217_), .A3(new_n14874_), .A4(new_n14899_), .ZN(new_n16811_));
  AOI21_X1   g15788(.A1(new_n16811_), .A2(new_n16810_), .B(new_n16214_), .ZN(new_n16812_));
  NOR2_X1    g15789(.A1(new_n16812_), .A2(new_n16220_), .ZN(new_n16813_));
  INV_X1     g15790(.I(new_n16813_), .ZN(new_n16814_));
  NOR3_X1    g15791(.A1(new_n16806_), .A2(new_n16814_), .A3(new_n16807_), .ZN(new_n16815_));
  OAI21_X1   g15792(.A1(new_n16202_), .A2(new_n16336_), .B(new_n16815_), .ZN(new_n16816_));
  OAI22_X1   g15793(.A1(new_n16257_), .A2(new_n16244_), .B1(new_n16247_), .B2(new_n16804_), .ZN(new_n16817_));
  INV_X1     g15794(.I(new_n16807_), .ZN(new_n16818_));
  NAND3_X1   g15795(.A1(new_n16817_), .A2(new_n16818_), .A3(new_n16813_), .ZN(new_n16819_));
  NAND4_X1   g15796(.A1(new_n16333_), .A2(new_n14942_), .A3(new_n16264_), .A4(new_n16819_), .ZN(new_n16820_));
  AOI21_X1   g15797(.A1(new_n16816_), .A2(new_n16820_), .B(new_n16802_), .ZN(new_n16821_));
  AOI21_X1   g15798(.A1(new_n16262_), .A2(new_n16264_), .B(new_n16819_), .ZN(new_n16822_));
  NOR3_X1    g15799(.A1(new_n16202_), .A2(new_n16336_), .A3(new_n16815_), .ZN(new_n16823_));
  NOR3_X1    g15800(.A1(new_n16822_), .A2(new_n16823_), .A3(new_n16801_), .ZN(new_n16824_));
  NOR2_X1    g15801(.A1(new_n16824_), .A2(new_n16821_), .ZN(new_n16825_));
  NOR2_X1    g15802(.A1(new_n16825_), .A2(new_n16786_), .ZN(new_n16826_));
  AOI21_X1   g15803(.A1(new_n16783_), .A2(new_n16784_), .B(new_n16782_), .ZN(new_n16827_));
  NOR3_X1    g15804(.A1(new_n16774_), .A2(new_n16780_), .A3(new_n16763_), .ZN(new_n16828_));
  NOR2_X1    g15805(.A1(new_n16828_), .A2(new_n16827_), .ZN(new_n16829_));
  OAI21_X1   g15806(.A1(new_n16822_), .A2(new_n16823_), .B(new_n16801_), .ZN(new_n16830_));
  NAND3_X1   g15807(.A1(new_n16816_), .A2(new_n16820_), .A3(new_n16802_), .ZN(new_n16831_));
  NAND2_X1   g15808(.A1(new_n16830_), .A2(new_n16831_), .ZN(new_n16832_));
  NOR2_X1    g15809(.A1(new_n16829_), .A2(new_n16832_), .ZN(new_n16833_));
  OAI21_X1   g15810(.A1(new_n16826_), .A2(new_n16833_), .B(new_n16747_), .ZN(new_n16834_));
  AOI21_X1   g15811(.A1(new_n16201_), .A2(new_n16364_), .B(new_n16350_), .ZN(new_n16835_));
  NOR2_X1    g15812(.A1(new_n16829_), .A2(new_n16825_), .ZN(new_n16836_));
  NOR4_X1    g15813(.A1(new_n16827_), .A2(new_n16828_), .A3(new_n16824_), .A4(new_n16821_), .ZN(new_n16837_));
  OAI21_X1   g15814(.A1(new_n16836_), .A2(new_n16837_), .B(new_n16835_), .ZN(new_n16838_));
  OAI21_X1   g15815(.A1(new_n16043_), .A2(new_n16357_), .B(new_n16198_), .ZN(new_n16839_));
  INV_X1     g15816(.I(new_n16163_), .ZN(new_n16840_));
  INV_X1     g15817(.I(new_n16164_), .ZN(new_n16841_));
  NAND4_X1   g15818(.A1(new_n16161_), .A2(new_n16840_), .A3(new_n16841_), .A4(new_n16167_), .ZN(new_n16842_));
  NOR2_X1    g15819(.A1(new_n16163_), .A2(new_n16164_), .ZN(new_n16843_));
  NOR2_X1    g15820(.A1(new_n16843_), .A2(new_n16167_), .ZN(new_n16844_));
  NAND2_X1   g15821(.A1(new_n16173_), .A2(new_n16844_), .ZN(new_n16845_));
  NAND2_X1   g15822(.A1(new_n16845_), .A2(new_n16842_), .ZN(new_n16846_));
  NAND2_X1   g15823(.A1(new_n15106_), .A2(new_n15108_), .ZN(new_n16847_));
  INV_X1     g15824(.I(new_n16167_), .ZN(new_n16848_));
  INV_X1     g15825(.I(new_n16843_), .ZN(new_n16849_));
  NOR2_X1    g15826(.A1(new_n16849_), .A2(new_n16848_), .ZN(new_n16850_));
  NOR2_X1    g15827(.A1(new_n16850_), .A2(new_n16844_), .ZN(new_n16851_));
  XNOR2_X1   g15828(.A1(new_n16139_), .A2(new_n16136_), .ZN(new_n16852_));
  NAND3_X1   g15829(.A1(new_n16852_), .A2(new_n16147_), .A3(new_n16161_), .ZN(new_n16853_));
  NOR3_X1    g15830(.A1(new_n16851_), .A2(new_n16847_), .A3(new_n16853_), .ZN(new_n16854_));
  NAND2_X1   g15831(.A1(new_n16847_), .A2(new_n16133_), .ZN(new_n16855_));
  NAND4_X1   g15832(.A1(new_n16854_), .A2(new_n16846_), .A3(new_n16173_), .A4(new_n16855_), .ZN(new_n16856_));
  NAND2_X1   g15833(.A1(new_n16159_), .A2(new_n15019_), .ZN(new_n16857_));
  AOI21_X1   g15834(.A1(new_n15009_), .A2(new_n15012_), .B(new_n16164_), .ZN(new_n16858_));
  NAND2_X1   g15835(.A1(new_n16857_), .A2(new_n16858_), .ZN(new_n16859_));
  OAI22_X1   g15836(.A1(new_n16173_), .A2(new_n16161_), .B1(new_n16163_), .B2(new_n16859_), .ZN(new_n16860_));
  NOR2_X1    g15837(.A1(new_n16848_), .A2(new_n16843_), .ZN(new_n16861_));
  INV_X1     g15838(.I(new_n16861_), .ZN(new_n16862_));
  OR2_X2     g15839(.A1(new_n15082_), .A2(new_n15078_), .Z(new_n16864_));
  NAND2_X1   g15840(.A1(new_n16143_), .A2(new_n16136_), .ZN(new_n16865_));
  NOR2_X1    g15841(.A1(new_n16865_), .A2(new_n16864_), .ZN(new_n16866_));
  NOR2_X1    g15842(.A1(new_n16866_), .A2(new_n16147_), .ZN(new_n16867_));
  NOR2_X1    g15843(.A1(new_n16867_), .A2(new_n16847_), .ZN(new_n16868_));
  NAND3_X1   g15844(.A1(new_n16860_), .A2(new_n16868_), .A3(new_n16862_), .ZN(new_n16869_));
  AOI21_X1   g15845(.A1(new_n16191_), .A2(new_n16179_), .B(new_n16869_), .ZN(new_n16870_));
  INV_X1     g15846(.I(new_n16179_), .ZN(new_n16871_));
  INV_X1     g15847(.I(new_n16859_), .ZN(new_n16872_));
  AOI22_X1   g15848(.A1(new_n16151_), .A2(new_n16162_), .B1(new_n16840_), .B2(new_n16872_), .ZN(new_n16873_));
  NOR4_X1    g15849(.A1(new_n16873_), .A2(new_n16847_), .A3(new_n16861_), .A4(new_n16867_), .ZN(new_n16874_));
  NOR3_X1    g15850(.A1(new_n16871_), .A2(new_n16177_), .A3(new_n16874_), .ZN(new_n16875_));
  OAI21_X1   g15851(.A1(new_n16870_), .A2(new_n16875_), .B(new_n16856_), .ZN(new_n16876_));
  INV_X1     g15852(.I(new_n16856_), .ZN(new_n16877_));
  OAI21_X1   g15853(.A1(new_n16871_), .A2(new_n16177_), .B(new_n16874_), .ZN(new_n16878_));
  NAND4_X1   g15854(.A1(new_n16124_), .A2(new_n15128_), .A3(new_n16869_), .A4(new_n16179_), .ZN(new_n16879_));
  NAND3_X1   g15855(.A1(new_n16878_), .A2(new_n16877_), .A3(new_n16879_), .ZN(new_n16880_));
  NOR2_X1    g15856(.A1(new_n15210_), .A2(new_n15278_), .ZN(new_n16881_));
  NOR2_X1    g15857(.A1(new_n15205_), .A2(new_n15286_), .ZN(new_n16882_));
  XOR2_X1    g15858(.A1(new_n16061_), .A2(new_n16063_), .Z(new_n16883_));
  XOR2_X1    g15859(.A1(new_n16097_), .A2(new_n16100_), .Z(new_n16884_));
  NOR3_X1    g15860(.A1(new_n16884_), .A2(new_n16073_), .A3(new_n16089_), .ZN(new_n16885_));
  NAND4_X1   g15861(.A1(new_n16885_), .A2(new_n16881_), .A3(new_n16882_), .A4(new_n16883_), .ZN(new_n16886_));
  OAI22_X1   g15862(.A1(new_n16105_), .A2(new_n16882_), .B1(new_n16881_), .B2(new_n16058_), .ZN(new_n16887_));
  NOR2_X1    g15863(.A1(new_n16886_), .A2(new_n16887_), .ZN(new_n16888_));
  INV_X1     g15864(.I(new_n16888_), .ZN(new_n16889_));
  NOR2_X1    g15865(.A1(new_n16087_), .A2(new_n15185_), .ZN(new_n16890_));
  NAND2_X1   g15866(.A1(new_n16095_), .A2(new_n15144_), .ZN(new_n16891_));
  OAI21_X1   g15867(.A1(new_n16095_), .A2(new_n15144_), .B(new_n15140_), .ZN(new_n16892_));
  AND3_X2    g15868(.A1(new_n16086_), .A2(new_n16891_), .A3(new_n16892_), .Z(new_n16893_));
  AOI22_X1   g15869(.A1(new_n16882_), .A2(new_n16893_), .B1(new_n16105_), .B2(new_n16890_), .ZN(new_n16894_));
  NAND2_X1   g15870(.A1(new_n16100_), .A2(new_n16101_), .ZN(new_n16895_));
  NOR4_X1    g15871(.A1(new_n16052_), .A2(new_n15251_), .A3(new_n16059_), .A4(new_n16055_), .ZN(new_n16896_));
  NAND2_X1   g15872(.A1(new_n16062_), .A2(new_n15229_), .ZN(new_n16897_));
  OAI21_X1   g15873(.A1(new_n16062_), .A2(new_n15229_), .B(new_n15227_), .ZN(new_n16898_));
  NAND2_X1   g15874(.A1(new_n16898_), .A2(new_n16897_), .ZN(new_n16899_));
  NOR4_X1    g15875(.A1(new_n15210_), .A2(new_n15278_), .A3(new_n16054_), .A4(new_n16899_), .ZN(new_n16900_));
  NOR2_X1    g15876(.A1(new_n16068_), .A2(new_n16067_), .ZN(new_n16901_));
  NOR3_X1    g15877(.A1(new_n16900_), .A2(new_n16896_), .A3(new_n16901_), .ZN(new_n16902_));
  NAND3_X1   g15878(.A1(new_n16894_), .A2(new_n16902_), .A3(new_n16895_), .ZN(new_n16903_));
  AOI21_X1   g15879(.A1(new_n16044_), .A2(new_n16121_), .B(new_n16903_), .ZN(new_n16904_));
  AND3_X2    g15880(.A1(new_n16894_), .A2(new_n16902_), .A3(new_n16895_), .Z(new_n16905_));
  NOR3_X1    g15881(.A1(new_n16119_), .A2(new_n16905_), .A3(new_n16186_), .ZN(new_n16906_));
  OAI21_X1   g15882(.A1(new_n16906_), .A2(new_n16904_), .B(new_n16889_), .ZN(new_n16907_));
  OAI21_X1   g15883(.A1(new_n16119_), .A2(new_n16186_), .B(new_n16905_), .ZN(new_n16908_));
  NAND3_X1   g15884(.A1(new_n16044_), .A2(new_n16121_), .A3(new_n16903_), .ZN(new_n16909_));
  NAND3_X1   g15885(.A1(new_n16908_), .A2(new_n16909_), .A3(new_n16888_), .ZN(new_n16910_));
  NAND2_X1   g15886(.A1(new_n16907_), .A2(new_n16910_), .ZN(new_n16911_));
  NAND3_X1   g15887(.A1(new_n16911_), .A2(new_n16876_), .A3(new_n16880_), .ZN(new_n16912_));
  INV_X1     g15888(.I(new_n16912_), .ZN(new_n16913_));
  AOI21_X1   g15889(.A1(new_n16876_), .A2(new_n16880_), .B(new_n16911_), .ZN(new_n16914_));
  OAI21_X1   g15890(.A1(new_n16913_), .A2(new_n16914_), .B(new_n16839_), .ZN(new_n16915_));
  AOI21_X1   g15891(.A1(new_n16196_), .A2(new_n16197_), .B(new_n16358_), .ZN(new_n16916_));
  AOI21_X1   g15892(.A1(new_n16908_), .A2(new_n16909_), .B(new_n16888_), .ZN(new_n16917_));
  NOR3_X1    g15893(.A1(new_n16906_), .A2(new_n16904_), .A3(new_n16889_), .ZN(new_n16918_));
  NOR2_X1    g15894(.A1(new_n16918_), .A2(new_n16917_), .ZN(new_n16919_));
  AOI21_X1   g15895(.A1(new_n16876_), .A2(new_n16880_), .B(new_n16919_), .ZN(new_n16920_));
  AOI21_X1   g15896(.A1(new_n16878_), .A2(new_n16879_), .B(new_n16877_), .ZN(new_n16921_));
  NOR3_X1    g15897(.A1(new_n16870_), .A2(new_n16875_), .A3(new_n16856_), .ZN(new_n16922_));
  NOR3_X1    g15898(.A1(new_n16922_), .A2(new_n16911_), .A3(new_n16921_), .ZN(new_n16923_));
  OAI21_X1   g15899(.A1(new_n16920_), .A2(new_n16923_), .B(new_n16916_), .ZN(new_n16924_));
  NAND2_X1   g15900(.A1(new_n16915_), .A2(new_n16924_), .ZN(new_n16925_));
  NAND3_X1   g15901(.A1(new_n16925_), .A2(new_n16834_), .A3(new_n16838_), .ZN(new_n16926_));
  NAND2_X1   g15902(.A1(new_n16834_), .A2(new_n16838_), .ZN(new_n16927_));
  NAND3_X1   g15903(.A1(new_n16927_), .A2(new_n16915_), .A3(new_n16924_), .ZN(new_n16928_));
  AOI21_X1   g15904(.A1(new_n16928_), .A2(new_n16926_), .B(new_n16746_), .ZN(new_n16929_));
  OAI21_X1   g15905(.A1(new_n16042_), .A2(new_n16382_), .B(new_n16371_), .ZN(new_n16930_));
  NAND4_X1   g15906(.A1(new_n16834_), .A2(new_n16838_), .A3(new_n16915_), .A4(new_n16924_), .ZN(new_n16931_));
  NAND2_X1   g15907(.A1(new_n16829_), .A2(new_n16832_), .ZN(new_n16932_));
  NAND2_X1   g15908(.A1(new_n16825_), .A2(new_n16786_), .ZN(new_n16933_));
  AOI21_X1   g15909(.A1(new_n16933_), .A2(new_n16932_), .B(new_n16835_), .ZN(new_n16934_));
  NAND2_X1   g15910(.A1(new_n16786_), .A2(new_n16832_), .ZN(new_n16935_));
  NAND4_X1   g15911(.A1(new_n16781_), .A2(new_n16830_), .A3(new_n16785_), .A4(new_n16831_), .ZN(new_n16936_));
  AOI21_X1   g15912(.A1(new_n16935_), .A2(new_n16936_), .B(new_n16747_), .ZN(new_n16937_));
  NAND2_X1   g15913(.A1(new_n16196_), .A2(new_n16197_), .ZN(new_n16938_));
  OAI21_X1   g15914(.A1(new_n16921_), .A2(new_n16922_), .B(new_n16919_), .ZN(new_n16939_));
  AOI22_X1   g15915(.A1(new_n16939_), .A2(new_n16912_), .B1(new_n16938_), .B2(new_n16198_), .ZN(new_n16940_));
  OAI21_X1   g15916(.A1(new_n16921_), .A2(new_n16922_), .B(new_n16911_), .ZN(new_n16941_));
  NAND3_X1   g15917(.A1(new_n16919_), .A2(new_n16876_), .A3(new_n16880_), .ZN(new_n16942_));
  AOI21_X1   g15918(.A1(new_n16941_), .A2(new_n16942_), .B(new_n16839_), .ZN(new_n16943_));
  OAI22_X1   g15919(.A1(new_n16934_), .A2(new_n16937_), .B1(new_n16943_), .B2(new_n16940_), .ZN(new_n16944_));
  AOI21_X1   g15920(.A1(new_n16931_), .A2(new_n16944_), .B(new_n16930_), .ZN(new_n16945_));
  NOR2_X1    g15921(.A1(new_n16929_), .A2(new_n16945_), .ZN(new_n16946_));
  NOR2_X1    g15922(.A1(new_n16031_), .A2(new_n16029_), .ZN(new_n16947_));
  NOR2_X1    g15923(.A1(new_n15919_), .A2(new_n16947_), .ZN(new_n16948_));
  NAND2_X1   g15924(.A1(new_n16014_), .A2(new_n16026_), .ZN(new_n16949_));
  NAND3_X1   g15925(.A1(new_n16027_), .A2(new_n16011_), .A3(new_n16013_), .ZN(new_n16950_));
  AOI22_X1   g15926(.A1(new_n15919_), .A2(new_n16947_), .B1(new_n16949_), .B2(new_n16950_), .ZN(new_n16951_));
  NOR2_X1    g15927(.A1(new_n16951_), .A2(new_n16948_), .ZN(new_n16952_));
  INV_X1     g15928(.I(new_n16952_), .ZN(new_n16953_));
  NOR2_X1    g15929(.A1(new_n15986_), .A2(new_n15987_), .ZN(new_n16954_));
  NOR2_X1    g15930(.A1(new_n15990_), .A2(new_n15991_), .ZN(new_n16955_));
  XNOR2_X1   g15931(.A1(new_n16955_), .A2(new_n16954_), .ZN(new_n16956_));
  NOR2_X1    g15932(.A1(new_n15983_), .A2(new_n15980_), .ZN(new_n16957_));
  NOR2_X1    g15933(.A1(new_n16956_), .A2(new_n16957_), .ZN(new_n16958_));
  NOR2_X1    g15934(.A1(new_n16955_), .A2(new_n16954_), .ZN(new_n16959_));
  NOR2_X1    g15935(.A1(new_n16959_), .A2(new_n15992_), .ZN(new_n16960_));
  NOR2_X1    g15936(.A1(new_n16960_), .A2(new_n15980_), .ZN(new_n16961_));
  NAND3_X1   g15937(.A1(new_n16002_), .A2(new_n15983_), .A3(new_n16961_), .ZN(new_n16962_));
  NOR2_X1    g15938(.A1(new_n16962_), .A2(new_n16958_), .ZN(new_n16963_));
  NOR4_X1    g15939(.A1(new_n15557_), .A2(new_n15560_), .A3(new_n15533_), .A4(new_n15532_), .ZN(new_n16964_));
  NAND4_X1   g15940(.A1(new_n15980_), .A2(new_n15986_), .A3(new_n15990_), .A4(new_n16964_), .ZN(new_n16965_));
  AOI21_X1   g15941(.A1(new_n16965_), .A2(new_n15660_), .B(new_n15584_), .ZN(new_n16966_));
  NOR2_X1    g15942(.A1(new_n16966_), .A2(new_n16959_), .ZN(new_n16967_));
  INV_X1     g15943(.I(new_n15953_), .ZN(new_n16968_));
  OAI21_X1   g15944(.A1(new_n15954_), .A2(new_n15618_), .B(new_n15627_), .ZN(new_n16969_));
  OAI21_X1   g15945(.A1(new_n15623_), .A2(new_n15626_), .B(new_n16969_), .ZN(new_n16970_));
  NAND2_X1   g15946(.A1(new_n16970_), .A2(new_n15959_), .ZN(new_n16971_));
  NOR2_X1    g15947(.A1(new_n16970_), .A2(new_n15959_), .ZN(new_n16972_));
  OAI21_X1   g15948(.A1(new_n16968_), .A2(new_n16972_), .B(new_n16971_), .ZN(new_n16973_));
  INV_X1     g15949(.I(new_n16973_), .ZN(new_n16974_));
  NAND2_X1   g15950(.A1(new_n16967_), .A2(new_n16974_), .ZN(new_n16975_));
  INV_X1     g15951(.I(new_n16975_), .ZN(new_n16976_));
  OAI21_X1   g15952(.A1(new_n15951_), .A2(new_n16008_), .B(new_n16976_), .ZN(new_n16977_));
  NOR2_X1    g15953(.A1(new_n16008_), .A2(new_n15951_), .ZN(new_n16978_));
  NAND2_X1   g15954(.A1(new_n16978_), .A2(new_n16975_), .ZN(new_n16979_));
  AOI21_X1   g15955(.A1(new_n16977_), .A2(new_n16979_), .B(new_n16963_), .ZN(new_n16980_));
  NAND3_X1   g15956(.A1(new_n16977_), .A2(new_n16979_), .A3(new_n16963_), .ZN(new_n16981_));
  INV_X1     g15957(.I(new_n16981_), .ZN(new_n16982_));
  NOR3_X1    g15958(.A1(new_n15936_), .A2(new_n15924_), .A3(new_n15925_), .ZN(new_n16984_));
  NOR2_X1    g15959(.A1(new_n15931_), .A2(new_n15940_), .ZN(new_n16985_));
  AOI21_X1   g15960(.A1(new_n15944_), .A2(new_n16985_), .B(new_n16984_), .ZN(new_n16986_));
  INV_X1     g15961(.I(new_n16986_), .ZN(new_n16987_));
  NOR3_X1    g15962(.A1(new_n16982_), .A2(new_n16980_), .A3(new_n16987_), .ZN(new_n16988_));
  INV_X1     g15963(.I(new_n16988_), .ZN(new_n16989_));
  INV_X1     g15964(.I(new_n16001_), .ZN(new_n16990_));
  NAND3_X1   g15965(.A1(new_n15997_), .A2(new_n16000_), .A3(new_n15971_), .ZN(new_n16991_));
  AOI21_X1   g15966(.A1(new_n16990_), .A2(new_n16991_), .B(new_n15951_), .ZN(new_n16992_));
  OAI21_X1   g15967(.A1(new_n16026_), .A2(new_n15950_), .B(new_n16009_), .ZN(new_n16993_));
  NOR2_X1    g15968(.A1(new_n16010_), .A2(new_n15950_), .ZN(new_n16994_));
  AOI21_X1   g15969(.A1(new_n16993_), .A2(new_n16992_), .B(new_n16994_), .ZN(new_n16995_));
  XOR2_X1    g15970(.A1(new_n16967_), .A2(new_n16973_), .Z(new_n16996_));
  NOR2_X1    g15971(.A1(new_n16963_), .A2(new_n16978_), .ZN(new_n16997_));
  NOR2_X1    g15972(.A1(new_n16997_), .A2(new_n16996_), .ZN(new_n16998_));
  INV_X1     g15973(.I(new_n16978_), .ZN(new_n16999_));
  INV_X1     g15974(.I(new_n16996_), .ZN(new_n17000_));
  OAI21_X1   g15975(.A1(new_n16956_), .A2(new_n16957_), .B(new_n16962_), .ZN(new_n17001_));
  NAND3_X1   g15976(.A1(new_n17000_), .A2(new_n16999_), .A3(new_n17001_), .ZN(new_n17002_));
  NAND3_X1   g15977(.A1(new_n17002_), .A2(new_n16998_), .A3(new_n16987_), .ZN(new_n17003_));
  NOR2_X1    g15978(.A1(new_n16995_), .A2(new_n17003_), .ZN(new_n17004_));
  INV_X1     g15979(.I(new_n17002_), .ZN(new_n17005_));
  NAND2_X1   g15980(.A1(new_n15782_), .A2(new_n15759_), .ZN(new_n17006_));
  OAI21_X1   g15981(.A1(new_n15762_), .A2(new_n15763_), .B(new_n15765_), .ZN(new_n17007_));
  NAND3_X1   g15982(.A1(new_n15672_), .A2(new_n15656_), .A3(new_n15670_), .ZN(new_n17008_));
  NAND2_X1   g15983(.A1(new_n17007_), .A2(new_n17008_), .ZN(new_n17009_));
  OAI21_X1   g15984(.A1(new_n15782_), .A2(new_n15759_), .B(new_n17009_), .ZN(new_n17010_));
  AOI21_X1   g15985(.A1(new_n17010_), .A2(new_n17006_), .B(new_n16006_), .ZN(new_n17011_));
  NAND3_X1   g15986(.A1(new_n17010_), .A2(new_n17006_), .A3(new_n16006_), .ZN(new_n17012_));
  NOR2_X1    g15987(.A1(new_n16009_), .A2(new_n15950_), .ZN(new_n17013_));
  AOI21_X1   g15988(.A1(new_n17012_), .A2(new_n17013_), .B(new_n17011_), .ZN(new_n17014_));
  NOR3_X1    g15989(.A1(new_n17014_), .A2(new_n16986_), .A3(new_n17005_), .ZN(new_n17015_));
  OAI21_X1   g15990(.A1(new_n16025_), .A2(new_n16021_), .B(new_n16992_), .ZN(new_n17016_));
  NOR3_X1    g15991(.A1(new_n16025_), .A2(new_n16021_), .A3(new_n16992_), .ZN(new_n17017_));
  INV_X1     g15992(.I(new_n17013_), .ZN(new_n17018_));
  OAI21_X1   g15993(.A1(new_n17017_), .A2(new_n17018_), .B(new_n17016_), .ZN(new_n17019_));
  AOI21_X1   g15994(.A1(new_n17019_), .A2(new_n16987_), .B(new_n17002_), .ZN(new_n17020_));
  OAI21_X1   g15995(.A1(new_n17020_), .A2(new_n17015_), .B(new_n16998_), .ZN(new_n17021_));
  NAND4_X1   g15996(.A1(new_n15909_), .A2(new_n15879_), .A3(new_n15882_), .A4(new_n15912_), .ZN(new_n17022_));
  NAND3_X1   g15997(.A1(new_n17022_), .A2(new_n15855_), .A3(new_n15506_), .ZN(new_n17023_));
  INV_X1     g15998(.I(new_n17023_), .ZN(new_n17024_));
  NAND2_X1   g15999(.A1(new_n15871_), .A2(new_n15434_), .ZN(new_n17025_));
  NAND2_X1   g16000(.A1(new_n15873_), .A2(new_n15465_), .ZN(new_n17026_));
  XOR2_X1    g16001(.A1(new_n17025_), .A2(new_n17026_), .Z(new_n17027_));
  XNOR2_X1   g16002(.A1(new_n15904_), .A2(new_n15899_), .ZN(new_n17028_));
  NOR3_X1    g16003(.A1(new_n17028_), .A2(new_n15867_), .A3(new_n15896_), .ZN(new_n17029_));
  NAND4_X1   g16004(.A1(new_n17029_), .A2(new_n15868_), .A3(new_n15897_), .A4(new_n17027_), .ZN(new_n17030_));
  OAI22_X1   g16005(.A1(new_n15868_), .A2(new_n15866_), .B1(new_n15897_), .B2(new_n15895_), .ZN(new_n17031_));
  NOR2_X1    g16006(.A1(new_n17030_), .A2(new_n17031_), .ZN(new_n17032_));
  AOI22_X1   g16007(.A1(new_n15902_), .A2(new_n15363_), .B1(new_n15364_), .B2(new_n15887_), .ZN(new_n17033_));
  OAI21_X1   g16008(.A1(new_n15900_), .A2(new_n15393_), .B(new_n17033_), .ZN(new_n17034_));
  AOI21_X1   g16009(.A1(new_n15896_), .A2(new_n15907_), .B(new_n17034_), .ZN(new_n17035_));
  NAND2_X1   g16010(.A1(new_n15893_), .A2(new_n15365_), .ZN(new_n17036_));
  NOR2_X1    g16011(.A1(new_n17035_), .A2(new_n17036_), .ZN(new_n17037_));
  NOR2_X1    g16012(.A1(new_n15904_), .A2(new_n15899_), .ZN(new_n17038_));
  NOR2_X1    g16013(.A1(new_n17037_), .A2(new_n17038_), .ZN(new_n17039_));
  NAND2_X1   g16014(.A1(new_n15867_), .A2(new_n15877_), .ZN(new_n17040_));
  OAI22_X1   g16015(.A1(new_n15859_), .A2(new_n15459_), .B1(new_n15437_), .B2(new_n15454_), .ZN(new_n17041_));
  AOI21_X1   g16016(.A1(new_n15864_), .A2(new_n15465_), .B(new_n17041_), .ZN(new_n17042_));
  NOR2_X1    g16017(.A1(new_n15869_), .A2(new_n15438_), .ZN(new_n17043_));
  INV_X1     g16018(.I(new_n17043_), .ZN(new_n17044_));
  AOI21_X1   g16019(.A1(new_n17040_), .A2(new_n17042_), .B(new_n17044_), .ZN(new_n17045_));
  NOR2_X1    g16020(.A1(new_n17025_), .A2(new_n17026_), .ZN(new_n17046_));
  NOR2_X1    g16021(.A1(new_n17045_), .A2(new_n17046_), .ZN(new_n17047_));
  NAND2_X1   g16022(.A1(new_n17047_), .A2(new_n17039_), .ZN(new_n17048_));
  XOR2_X1    g16023(.A1(new_n17048_), .A2(new_n17032_), .Z(new_n17049_));
  XOR2_X1    g16024(.A1(new_n17049_), .A2(new_n17024_), .Z(new_n17050_));
  NAND2_X1   g16025(.A1(new_n17021_), .A2(new_n17050_), .ZN(new_n17051_));
  NAND3_X1   g16026(.A1(new_n17051_), .A2(new_n16989_), .A3(new_n17004_), .ZN(new_n17052_));
  INV_X1     g16027(.I(new_n16998_), .ZN(new_n17053_));
  NAND3_X1   g16028(.A1(new_n17019_), .A2(new_n16987_), .A3(new_n17002_), .ZN(new_n17054_));
  OAI21_X1   g16029(.A1(new_n17014_), .A2(new_n16986_), .B(new_n17005_), .ZN(new_n17055_));
  AOI21_X1   g16030(.A1(new_n17055_), .A2(new_n17054_), .B(new_n17053_), .ZN(new_n17056_));
  XOR2_X1    g16031(.A1(new_n17049_), .A2(new_n17023_), .Z(new_n17057_));
  OAI21_X1   g16032(.A1(new_n17056_), .A2(new_n17057_), .B(new_n17004_), .ZN(new_n17058_));
  NAND2_X1   g16033(.A1(new_n17058_), .A2(new_n16988_), .ZN(new_n17059_));
  NAND3_X1   g16034(.A1(new_n17059_), .A2(new_n17052_), .A3(new_n16953_), .ZN(new_n17060_));
  NOR2_X1    g16035(.A1(new_n17058_), .A2(new_n16988_), .ZN(new_n17061_));
  AOI21_X1   g16036(.A1(new_n17051_), .A2(new_n17004_), .B(new_n16989_), .ZN(new_n17062_));
  OAI21_X1   g16037(.A1(new_n17061_), .A2(new_n17062_), .B(new_n16952_), .ZN(new_n17063_));
  AOI21_X1   g16038(.A1(new_n17063_), .A2(new_n17060_), .B(new_n16946_), .ZN(new_n17064_));
  INV_X1     g16039(.I(new_n16946_), .ZN(new_n17065_));
  OAI21_X1   g16040(.A1(new_n17061_), .A2(new_n17062_), .B(new_n16953_), .ZN(new_n17066_));
  NAND3_X1   g16041(.A1(new_n17059_), .A2(new_n17052_), .A3(new_n16952_), .ZN(new_n17067_));
  AOI21_X1   g16042(.A1(new_n17066_), .A2(new_n17067_), .B(new_n17065_), .ZN(new_n17068_));
  NOR2_X1    g16043(.A1(new_n17064_), .A2(new_n17068_), .ZN(new_n17069_));
  INV_X1     g16044(.I(new_n17069_), .ZN(new_n17070_));
  NAND2_X1   g16045(.A1(new_n15854_), .A2(new_n16724_), .ZN(new_n17071_));
  NOR3_X1    g16046(.A1(new_n16742_), .A2(new_n16743_), .A3(new_n16728_), .ZN(new_n17072_));
  AOI21_X1   g16047(.A1(new_n16385_), .A2(new_n16375_), .B(new_n16387_), .ZN(new_n17073_));
  OAI22_X1   g16048(.A1(new_n15854_), .A2(new_n16724_), .B1(new_n17072_), .B2(new_n17073_), .ZN(new_n17074_));
  OAI22_X1   g16049(.A1(new_n16711_), .A2(new_n16714_), .B1(new_n16717_), .B2(new_n16720_), .ZN(new_n17075_));
  AOI21_X1   g16050(.A1(new_n16389_), .A2(new_n17075_), .B(new_n16721_), .ZN(new_n17076_));
  OAI21_X1   g16051(.A1(new_n16701_), .A2(new_n16702_), .B(new_n16719_), .ZN(new_n17077_));
  INV_X1     g16052(.I(new_n16659_), .ZN(new_n17078_));
  INV_X1     g16053(.I(new_n16660_), .ZN(new_n17079_));
  NOR2_X1    g16054(.A1(new_n16633_), .A2(new_n14002_), .ZN(new_n17080_));
  NAND3_X1   g16055(.A1(new_n16637_), .A2(new_n16636_), .A3(new_n16639_), .ZN(new_n17081_));
  XNOR2_X1   g16056(.A1(new_n17081_), .A2(new_n16635_), .ZN(new_n17082_));
  AND3_X2    g16057(.A1(new_n17080_), .A2(new_n16632_), .A3(new_n17082_), .Z(new_n17083_));
  NAND4_X1   g16058(.A1(new_n17083_), .A2(new_n17078_), .A3(new_n17079_), .A4(new_n16667_), .ZN(new_n17084_));
  INV_X1     g16059(.I(new_n16681_), .ZN(new_n17085_));
  NAND2_X1   g16060(.A1(new_n16668_), .A2(new_n16660_), .ZN(new_n17086_));
  NAND2_X1   g16061(.A1(new_n16655_), .A2(new_n16656_), .ZN(new_n17087_));
  NOR2_X1    g16062(.A1(new_n14076_), .A2(new_n14072_), .ZN(new_n17088_));
  NAND4_X1   g16063(.A1(new_n17087_), .A2(new_n16652_), .A3(new_n16653_), .A4(new_n17088_), .ZN(new_n17089_));
  OAI21_X1   g16064(.A1(new_n16652_), .A2(new_n16653_), .B(new_n16658_), .ZN(new_n17090_));
  INV_X1     g16065(.I(new_n17090_), .ZN(new_n17091_));
  AOI21_X1   g16066(.A1(new_n17086_), .A2(new_n17089_), .B(new_n17091_), .ZN(new_n17092_));
  NAND2_X1   g16067(.A1(new_n16637_), .A2(new_n16636_), .ZN(new_n17093_));
  NOR3_X1    g16068(.A1(new_n16639_), .A2(new_n14011_), .A3(new_n14015_), .ZN(new_n17094_));
  NAND4_X1   g16069(.A1(new_n17093_), .A2(new_n14016_), .A3(new_n16630_), .A4(new_n17094_), .ZN(new_n17095_));
  INV_X1     g16070(.I(new_n16635_), .ZN(new_n17096_));
  NAND2_X1   g16071(.A1(new_n17096_), .A2(new_n17081_), .ZN(new_n17097_));
  NOR2_X1    g16072(.A1(new_n17097_), .A2(new_n17095_), .ZN(new_n17098_));
  NOR2_X1    g16073(.A1(new_n17080_), .A2(new_n17098_), .ZN(new_n17099_));
  NOR2_X1    g16074(.A1(new_n17099_), .A2(new_n16646_), .ZN(new_n17100_));
  NAND2_X1   g16075(.A1(new_n17100_), .A2(new_n17092_), .ZN(new_n17101_));
  AOI21_X1   g16076(.A1(new_n16622_), .A2(new_n17085_), .B(new_n17101_), .ZN(new_n17102_));
  NAND3_X1   g16077(.A1(new_n16622_), .A2(new_n17085_), .A3(new_n17101_), .ZN(new_n17103_));
  INV_X1     g16078(.I(new_n17103_), .ZN(new_n17104_));
  OAI21_X1   g16079(.A1(new_n17104_), .A2(new_n17102_), .B(new_n17084_), .ZN(new_n17105_));
  INV_X1     g16080(.I(new_n17084_), .ZN(new_n17106_));
  INV_X1     g16081(.I(new_n17101_), .ZN(new_n17107_));
  OAI21_X1   g16082(.A1(new_n16679_), .A2(new_n16681_), .B(new_n17107_), .ZN(new_n17108_));
  NAND3_X1   g16083(.A1(new_n17108_), .A2(new_n17103_), .A3(new_n17106_), .ZN(new_n17109_));
  NAND2_X1   g16084(.A1(new_n14171_), .A2(new_n14118_), .ZN(new_n17110_));
  INV_X1     g16085(.I(new_n16610_), .ZN(new_n17111_));
  NAND2_X1   g16086(.A1(new_n17110_), .A2(new_n17111_), .ZN(new_n17112_));
  NAND2_X1   g16087(.A1(new_n17112_), .A2(new_n16603_), .ZN(new_n17113_));
  NAND3_X1   g16088(.A1(new_n16603_), .A2(new_n16604_), .A3(new_n16610_), .ZN(new_n17114_));
  NOR2_X1    g16089(.A1(new_n16561_), .A2(new_n16571_), .ZN(new_n17115_));
  XOR2_X1    g16090(.A1(new_n16576_), .A2(new_n16580_), .Z(new_n17116_));
  NAND3_X1   g16091(.A1(new_n16561_), .A2(new_n16571_), .A3(new_n17116_), .ZN(new_n17117_));
  NOR4_X1    g16092(.A1(new_n17113_), .A2(new_n17114_), .A3(new_n17115_), .A4(new_n17117_), .ZN(new_n17118_));
  INV_X1     g16093(.I(new_n17118_), .ZN(new_n17119_));
  NAND2_X1   g16094(.A1(new_n14230_), .A2(new_n14174_), .ZN(new_n17120_));
  INV_X1     g16095(.I(new_n16583_), .ZN(new_n17121_));
  OAI21_X1   g16096(.A1(new_n17121_), .A2(new_n16584_), .B(new_n17120_), .ZN(new_n17122_));
  NAND3_X1   g16097(.A1(new_n16614_), .A2(new_n17122_), .A3(new_n16587_), .ZN(new_n17123_));
  NOR4_X1    g16098(.A1(new_n14151_), .A2(new_n16591_), .A3(new_n16593_), .A4(new_n14154_), .ZN(new_n17124_));
  NAND3_X1   g16099(.A1(new_n16595_), .A2(new_n16600_), .A3(new_n17124_), .ZN(new_n17125_));
  INV_X1     g16100(.I(new_n17125_), .ZN(new_n17126_));
  AOI21_X1   g16101(.A1(new_n17111_), .A2(new_n17110_), .B(new_n17126_), .ZN(new_n17127_));
  NOR2_X1    g16102(.A1(new_n16597_), .A2(new_n16602_), .ZN(new_n17128_));
  NOR2_X1    g16103(.A1(new_n17127_), .A2(new_n17128_), .ZN(new_n17129_));
  NAND4_X1   g16104(.A1(new_n16573_), .A2(new_n16578_), .A3(new_n16575_), .A4(new_n16579_), .ZN(new_n17130_));
  INV_X1     g16105(.I(new_n17130_), .ZN(new_n17131_));
  OAI21_X1   g16106(.A1(new_n16561_), .A2(new_n17131_), .B(new_n16571_), .ZN(new_n17132_));
  INV_X1     g16107(.I(new_n17132_), .ZN(new_n17133_));
  NAND2_X1   g16108(.A1(new_n17129_), .A2(new_n17133_), .ZN(new_n17134_));
  AOI21_X1   g16109(.A1(new_n16612_), .A2(new_n17123_), .B(new_n17134_), .ZN(new_n17135_));
  NOR3_X1    g16110(.A1(new_n16588_), .A2(new_n16586_), .A3(new_n16611_), .ZN(new_n17136_));
  INV_X1     g16111(.I(new_n17129_), .ZN(new_n17137_));
  NOR2_X1    g16112(.A1(new_n17137_), .A2(new_n17132_), .ZN(new_n17138_));
  NOR3_X1    g16113(.A1(new_n17136_), .A2(new_n17138_), .A3(new_n16615_), .ZN(new_n17139_));
  OAI21_X1   g16114(.A1(new_n17139_), .A2(new_n17135_), .B(new_n17119_), .ZN(new_n17140_));
  OAI21_X1   g16115(.A1(new_n17136_), .A2(new_n16615_), .B(new_n17138_), .ZN(new_n17141_));
  NAND3_X1   g16116(.A1(new_n16612_), .A2(new_n17123_), .A3(new_n17134_), .ZN(new_n17142_));
  NAND3_X1   g16117(.A1(new_n17141_), .A2(new_n17142_), .A3(new_n17118_), .ZN(new_n17143_));
  NAND2_X1   g16118(.A1(new_n17143_), .A2(new_n17140_), .ZN(new_n17144_));
  NAND3_X1   g16119(.A1(new_n17105_), .A2(new_n17144_), .A3(new_n17109_), .ZN(new_n17145_));
  AOI21_X1   g16120(.A1(new_n17108_), .A2(new_n17103_), .B(new_n17106_), .ZN(new_n17146_));
  NOR3_X1    g16121(.A1(new_n17104_), .A2(new_n17102_), .A3(new_n17084_), .ZN(new_n17147_));
  AOI21_X1   g16122(.A1(new_n17141_), .A2(new_n17142_), .B(new_n17118_), .ZN(new_n17148_));
  NOR3_X1    g16123(.A1(new_n17139_), .A2(new_n17135_), .A3(new_n17119_), .ZN(new_n17149_));
  NOR2_X1    g16124(.A1(new_n17148_), .A2(new_n17149_), .ZN(new_n17150_));
  OAI21_X1   g16125(.A1(new_n17147_), .A2(new_n17146_), .B(new_n17150_), .ZN(new_n17151_));
  NAND2_X1   g16126(.A1(new_n17151_), .A2(new_n17145_), .ZN(new_n17152_));
  NAND2_X1   g16127(.A1(new_n17152_), .A2(new_n17077_), .ZN(new_n17153_));
  AOI21_X1   g16128(.A1(new_n16718_), .A2(new_n16560_), .B(new_n16703_), .ZN(new_n17154_));
  OAI21_X1   g16129(.A1(new_n17147_), .A2(new_n17146_), .B(new_n17144_), .ZN(new_n17155_));
  NAND3_X1   g16130(.A1(new_n17105_), .A2(new_n17150_), .A3(new_n17109_), .ZN(new_n17156_));
  NAND2_X1   g16131(.A1(new_n17155_), .A2(new_n17156_), .ZN(new_n17157_));
  NAND2_X1   g16132(.A1(new_n17157_), .A2(new_n17154_), .ZN(new_n17158_));
  NAND2_X1   g16133(.A1(new_n17158_), .A2(new_n17153_), .ZN(new_n17159_));
  OAI21_X1   g16134(.A1(new_n16545_), .A2(new_n16544_), .B(new_n16554_), .ZN(new_n17160_));
  XOR2_X1    g16135(.A1(new_n16481_), .A2(new_n16484_), .Z(new_n17161_));
  XOR2_X1    g16136(.A1(new_n16506_), .A2(new_n16509_), .Z(new_n17162_));
  NOR3_X1    g16137(.A1(new_n17162_), .A2(new_n16477_), .A3(new_n16503_), .ZN(new_n17163_));
  NAND4_X1   g16138(.A1(new_n17163_), .A2(new_n16464_), .A3(new_n16493_), .A4(new_n17161_), .ZN(new_n17164_));
  NAND2_X1   g16139(.A1(new_n16465_), .A2(new_n16477_), .ZN(new_n17165_));
  NAND2_X1   g16140(.A1(new_n16494_), .A2(new_n16503_), .ZN(new_n17166_));
  NAND2_X1   g16141(.A1(new_n17165_), .A2(new_n17166_), .ZN(new_n17167_));
  NOR2_X1    g16142(.A1(new_n17164_), .A2(new_n17167_), .ZN(new_n17168_));
  NOR2_X1    g16143(.A1(new_n16492_), .A2(new_n16519_), .ZN(new_n17169_));
  INV_X1     g16144(.I(new_n16477_), .ZN(new_n17170_));
  NOR4_X1    g16145(.A1(new_n16504_), .A2(new_n16505_), .A3(new_n16507_), .A4(new_n16508_), .ZN(new_n17171_));
  OR2_X2     g16146(.A1(new_n16493_), .A2(new_n17171_), .Z(new_n17172_));
  NOR4_X1    g16147(.A1(new_n16478_), .A2(new_n16482_), .A3(new_n16480_), .A4(new_n16483_), .ZN(new_n17173_));
  OR2_X2     g16148(.A1(new_n16464_), .A2(new_n17173_), .Z(new_n17174_));
  NAND4_X1   g16149(.A1(new_n17174_), .A2(new_n17172_), .A3(new_n17170_), .A4(new_n16515_), .ZN(new_n17175_));
  INV_X1     g16150(.I(new_n17175_), .ZN(new_n17176_));
  OAI21_X1   g16151(.A1(new_n17169_), .A2(new_n16537_), .B(new_n17176_), .ZN(new_n17177_));
  NAND3_X1   g16152(.A1(new_n16526_), .A2(new_n16489_), .A3(new_n16491_), .ZN(new_n17178_));
  NAND3_X1   g16153(.A1(new_n16522_), .A2(new_n17178_), .A3(new_n17175_), .ZN(new_n17179_));
  AOI21_X1   g16154(.A1(new_n17177_), .A2(new_n17179_), .B(new_n17168_), .ZN(new_n17180_));
  INV_X1     g16155(.I(new_n17168_), .ZN(new_n17181_));
  AOI21_X1   g16156(.A1(new_n16522_), .A2(new_n17178_), .B(new_n17175_), .ZN(new_n17182_));
  NOR3_X1    g16157(.A1(new_n17169_), .A2(new_n16537_), .A3(new_n17176_), .ZN(new_n17183_));
  NOR3_X1    g16158(.A1(new_n17182_), .A2(new_n17183_), .A3(new_n17181_), .ZN(new_n17184_));
  NOR2_X1    g16159(.A1(new_n17184_), .A2(new_n17180_), .ZN(new_n17185_));
  NOR2_X1    g16160(.A1(new_n16402_), .A2(new_n16403_), .ZN(new_n17186_));
  XNOR2_X1   g16161(.A1(new_n17186_), .A2(new_n16407_), .ZN(new_n17187_));
  XNOR2_X1   g16162(.A1(new_n16440_), .A2(new_n16436_), .ZN(new_n17188_));
  NOR3_X1    g16163(.A1(new_n17188_), .A2(new_n16401_), .A3(new_n16442_), .ZN(new_n17189_));
  NAND4_X1   g16164(.A1(new_n17189_), .A2(new_n16391_), .A3(new_n16446_), .A4(new_n17187_), .ZN(new_n17190_));
  NAND2_X1   g16165(.A1(new_n16390_), .A2(new_n16401_), .ZN(new_n17191_));
  NAND2_X1   g16166(.A1(new_n16419_), .A2(new_n16442_), .ZN(new_n17192_));
  NAND2_X1   g16167(.A1(new_n17192_), .A2(new_n17191_), .ZN(new_n17193_));
  NOR2_X1    g16168(.A1(new_n17190_), .A2(new_n17193_), .ZN(new_n17194_));
  INV_X1     g16169(.I(new_n17194_), .ZN(new_n17195_));
  NAND2_X1   g16170(.A1(new_n16415_), .A2(new_n16390_), .ZN(new_n17196_));
  NAND2_X1   g16171(.A1(new_n16412_), .A2(new_n16391_), .ZN(new_n17197_));
  NAND3_X1   g16172(.A1(new_n16458_), .A2(new_n17197_), .A3(new_n17196_), .ZN(new_n17198_));
  NOR4_X1    g16173(.A1(new_n16437_), .A2(new_n16433_), .A3(new_n16435_), .A4(new_n16439_), .ZN(new_n17199_));
  OAI21_X1   g16174(.A1(new_n16446_), .A2(new_n17199_), .B(new_n16432_), .ZN(new_n17200_));
  INV_X1     g16175(.I(new_n16401_), .ZN(new_n17201_));
  INV_X1     g16176(.I(new_n16402_), .ZN(new_n17202_));
  INV_X1     g16177(.I(new_n16403_), .ZN(new_n17203_));
  NOR4_X1    g16178(.A1(new_n17202_), .A2(new_n17203_), .A3(new_n16405_), .A4(new_n16406_), .ZN(new_n17204_));
  OAI21_X1   g16179(.A1(new_n16391_), .A2(new_n17204_), .B(new_n17201_), .ZN(new_n17205_));
  NOR2_X1    g16180(.A1(new_n17205_), .A2(new_n17200_), .ZN(new_n17206_));
  INV_X1     g16181(.I(new_n17206_), .ZN(new_n17207_));
  AOI21_X1   g16182(.A1(new_n17198_), .A2(new_n16451_), .B(new_n17207_), .ZN(new_n17208_));
  NOR3_X1    g16183(.A1(new_n16450_), .A2(new_n16413_), .A3(new_n16416_), .ZN(new_n17209_));
  NOR3_X1    g16184(.A1(new_n16548_), .A2(new_n17209_), .A3(new_n17206_), .ZN(new_n17210_));
  OAI21_X1   g16185(.A1(new_n17210_), .A2(new_n17208_), .B(new_n17195_), .ZN(new_n17211_));
  OAI21_X1   g16186(.A1(new_n16548_), .A2(new_n17209_), .B(new_n17206_), .ZN(new_n17212_));
  NAND3_X1   g16187(.A1(new_n17198_), .A2(new_n17207_), .A3(new_n16451_), .ZN(new_n17213_));
  NAND3_X1   g16188(.A1(new_n17212_), .A2(new_n17213_), .A3(new_n17194_), .ZN(new_n17214_));
  NAND2_X1   g16189(.A1(new_n17211_), .A2(new_n17214_), .ZN(new_n17215_));
  NAND2_X1   g16190(.A1(new_n17185_), .A2(new_n17215_), .ZN(new_n17216_));
  OAI21_X1   g16191(.A1(new_n17182_), .A2(new_n17183_), .B(new_n17181_), .ZN(new_n17217_));
  NAND3_X1   g16192(.A1(new_n17177_), .A2(new_n17179_), .A3(new_n17168_), .ZN(new_n17218_));
  NAND2_X1   g16193(.A1(new_n17217_), .A2(new_n17218_), .ZN(new_n17219_));
  AOI21_X1   g16194(.A1(new_n17212_), .A2(new_n17213_), .B(new_n17194_), .ZN(new_n17220_));
  NOR3_X1    g16195(.A1(new_n17210_), .A2(new_n17208_), .A3(new_n17195_), .ZN(new_n17221_));
  NOR2_X1    g16196(.A1(new_n17221_), .A2(new_n17220_), .ZN(new_n17222_));
  NAND2_X1   g16197(.A1(new_n17219_), .A2(new_n17222_), .ZN(new_n17223_));
  AOI22_X1   g16198(.A1(new_n17223_), .A2(new_n17216_), .B1(new_n17160_), .B2(new_n16709_), .ZN(new_n17224_));
  NAND2_X1   g16199(.A1(new_n17160_), .A2(new_n16709_), .ZN(new_n17225_));
  AOI22_X1   g16200(.A1(new_n17217_), .A2(new_n17218_), .B1(new_n17211_), .B2(new_n17214_), .ZN(new_n17226_));
  NOR4_X1    g16201(.A1(new_n17180_), .A2(new_n17184_), .A3(new_n17221_), .A4(new_n17220_), .ZN(new_n17227_));
  NOR2_X1    g16202(.A1(new_n17227_), .A2(new_n17226_), .ZN(new_n17228_));
  NOR2_X1    g16203(.A1(new_n17225_), .A2(new_n17228_), .ZN(new_n17229_));
  NOR2_X1    g16204(.A1(new_n17229_), .A2(new_n17224_), .ZN(new_n17230_));
  XOR2_X1    g16205(.A1(new_n17159_), .A2(new_n17230_), .Z(new_n17231_));
  AOI21_X1   g16206(.A1(new_n17145_), .A2(new_n17151_), .B(new_n17154_), .ZN(new_n17232_));
  AOI21_X1   g16207(.A1(new_n17155_), .A2(new_n17156_), .B(new_n17077_), .ZN(new_n17233_));
  NOR4_X1    g16208(.A1(new_n17229_), .A2(new_n17233_), .A3(new_n17232_), .A4(new_n17224_), .ZN(new_n17234_));
  AOI21_X1   g16209(.A1(new_n16534_), .A2(new_n16535_), .B(new_n16463_), .ZN(new_n17235_));
  NOR2_X1    g16210(.A1(new_n17219_), .A2(new_n17222_), .ZN(new_n17236_));
  NOR2_X1    g16211(.A1(new_n17185_), .A2(new_n17215_), .ZN(new_n17237_));
  OAI22_X1   g16212(.A1(new_n17235_), .A2(new_n16536_), .B1(new_n17236_), .B2(new_n17237_), .ZN(new_n17238_));
  NAND2_X1   g16213(.A1(new_n17215_), .A2(new_n17219_), .ZN(new_n17239_));
  NAND4_X1   g16214(.A1(new_n17217_), .A2(new_n17218_), .A3(new_n17211_), .A4(new_n17214_), .ZN(new_n17240_));
  NAND2_X1   g16215(.A1(new_n17239_), .A2(new_n17240_), .ZN(new_n17241_));
  NAND3_X1   g16216(.A1(new_n17241_), .A2(new_n16709_), .A3(new_n17160_), .ZN(new_n17242_));
  AOI22_X1   g16217(.A1(new_n17153_), .A2(new_n17158_), .B1(new_n17242_), .B2(new_n17238_), .ZN(new_n17243_));
  OAI21_X1   g16218(.A1(new_n17234_), .A2(new_n17243_), .B(new_n17076_), .ZN(new_n17244_));
  OAI21_X1   g16219(.A1(new_n17231_), .A2(new_n17076_), .B(new_n17244_), .ZN(new_n17245_));
  NAND3_X1   g16220(.A1(new_n17074_), .A2(new_n17071_), .A3(new_n17245_), .ZN(new_n17246_));
  AOI21_X1   g16221(.A1(new_n17074_), .A2(new_n17071_), .B(new_n17245_), .ZN(new_n17247_));
  INV_X1     g16222(.I(new_n17247_), .ZN(new_n17248_));
  AOI21_X1   g16223(.A1(new_n17248_), .A2(new_n17246_), .B(new_n17070_), .ZN(new_n17249_));
  INV_X1     g16224(.I(new_n17246_), .ZN(new_n17250_));
  NOR3_X1    g16225(.A1(new_n17250_), .A2(new_n17069_), .A3(new_n17247_), .ZN(new_n17251_));
  OAI21_X1   g16226(.A1(new_n17249_), .A2(new_n17251_), .B(new_n16745_), .ZN(new_n17252_));
  NAND2_X1   g16227(.A1(new_n16385_), .A2(new_n16387_), .ZN(new_n17253_));
  NAND2_X1   g16228(.A1(new_n17253_), .A2(new_n16375_), .ZN(new_n17254_));
  OAI21_X1   g16229(.A1(new_n17250_), .A2(new_n17247_), .B(new_n17069_), .ZN(new_n17255_));
  NAND3_X1   g16230(.A1(new_n17248_), .A2(new_n17070_), .A3(new_n17246_), .ZN(new_n17256_));
  NAND3_X1   g16231(.A1(new_n17256_), .A2(new_n17255_), .A3(new_n17254_), .ZN(new_n17257_));
  AOI21_X1   g16232(.A1(new_n17252_), .A2(new_n17257_), .B(new_n16741_), .ZN(new_n17258_));
  INV_X1     g16233(.I(new_n15849_), .ZN(new_n17259_));
  NOR3_X1    g16234(.A1(new_n16737_), .A2(new_n16739_), .A3(new_n16735_), .ZN(new_n17260_));
  AOI21_X1   g16235(.A1(new_n16730_), .A2(new_n16726_), .B(new_n15854_), .ZN(new_n17261_));
  OAI21_X1   g16236(.A1(new_n17261_), .A2(new_n17260_), .B(new_n17259_), .ZN(new_n17262_));
  AOI21_X1   g16237(.A1(new_n17256_), .A2(new_n17255_), .B(new_n17254_), .ZN(new_n17263_));
  NOR3_X1    g16238(.A1(new_n17249_), .A2(new_n17251_), .A3(new_n16745_), .ZN(new_n17264_));
  NOR3_X1    g16239(.A1(new_n17263_), .A2(new_n17264_), .A3(new_n17262_), .ZN(new_n17265_));
  AOI21_X1   g16240(.A1(new_n16730_), .A2(new_n16726_), .B(new_n16735_), .ZN(new_n17266_));
  NOR3_X1    g16241(.A1(new_n16737_), .A2(new_n16739_), .A3(new_n15854_), .ZN(new_n17267_));
  OAI21_X1   g16242(.A1(new_n17266_), .A2(new_n17267_), .B(new_n17259_), .ZN(new_n17268_));
  OAI21_X1   g16243(.A1(new_n17261_), .A2(new_n17260_), .B(new_n15849_), .ZN(new_n17269_));
  INV_X1     g16244(.I(new_n13955_), .ZN(new_n17270_));
  NAND2_X1   g16245(.A1(new_n15846_), .A2(new_n13986_), .ZN(new_n17271_));
  NAND3_X1   g16246(.A1(new_n15819_), .A2(new_n15834_), .A3(new_n15845_), .ZN(new_n17272_));
  AOI21_X1   g16247(.A1(new_n17271_), .A2(new_n17272_), .B(new_n17270_), .ZN(new_n17273_));
  AOI21_X1   g16248(.A1(new_n15847_), .A2(new_n15835_), .B(new_n13955_), .ZN(new_n17274_));
  INV_X1     g16249(.I(new_n13952_), .ZN(new_n17275_));
  INV_X1     g16250(.I(new_n13953_), .ZN(new_n17276_));
  NOR2_X1    g16251(.A1(new_n17275_), .A2(new_n17276_), .ZN(new_n17277_));
  XNOR2_X1   g16252(.A1(new_n17277_), .A2(new_n13939_), .ZN(new_n17278_));
  NAND2_X1   g16253(.A1(new_n13983_), .A2(new_n13952_), .ZN(new_n17279_));
  NAND3_X1   g16254(.A1(new_n13942_), .A2(new_n17279_), .A3(new_n17277_), .ZN(new_n17280_));
  INV_X1     g16255(.I(new_n17280_), .ZN(new_n17281_));
  AOI21_X1   g16256(.A1(new_n13942_), .A2(new_n17279_), .B(new_n17277_), .ZN(new_n17282_));
  OAI21_X1   g16257(.A1(new_n17281_), .A2(new_n17282_), .B(new_n13939_), .ZN(new_n17283_));
  INV_X1     g16258(.I(new_n17282_), .ZN(new_n17284_));
  NAND3_X1   g16259(.A1(new_n17284_), .A2(new_n13940_), .A3(new_n17280_), .ZN(new_n17285_));
  NAND2_X1   g16260(.A1(new_n17285_), .A2(new_n17283_), .ZN(new_n17286_));
  OAI22_X1   g16261(.A1(new_n17273_), .A2(new_n17274_), .B1(new_n17286_), .B2(new_n17278_), .ZN(new_n17287_));
  NAND3_X1   g16262(.A1(new_n17268_), .A2(new_n17269_), .A3(new_n17287_), .ZN(new_n17288_));
  OAI21_X1   g16263(.A1(new_n17265_), .A2(new_n17258_), .B(new_n17288_), .ZN(new_n17289_));
  NOR3_X1    g16264(.A1(new_n16995_), .A2(new_n16988_), .A3(new_n17003_), .ZN(new_n17290_));
  OAI21_X1   g16265(.A1(new_n16951_), .A2(new_n16948_), .B(new_n17290_), .ZN(new_n17291_));
  NOR3_X1    g16266(.A1(new_n16951_), .A2(new_n17290_), .A3(new_n16948_), .ZN(new_n17292_));
  NAND2_X1   g16267(.A1(new_n17056_), .A2(new_n17057_), .ZN(new_n17293_));
  OAI21_X1   g16268(.A1(new_n17292_), .A2(new_n17293_), .B(new_n17291_), .ZN(new_n17294_));
  NOR3_X1    g16269(.A1(new_n17005_), .A2(new_n16998_), .A3(new_n16987_), .ZN(new_n17295_));
  NOR3_X1    g16270(.A1(new_n16982_), .A2(new_n16980_), .A3(new_n16986_), .ZN(new_n17296_));
  NAND2_X1   g16271(.A1(new_n17046_), .A2(new_n17038_), .ZN(new_n17297_));
  INV_X1     g16272(.I(new_n17297_), .ZN(new_n17298_));
  AND3_X2    g16273(.A1(new_n17045_), .A2(new_n17037_), .A3(new_n17298_), .Z(new_n17299_));
  OAI21_X1   g16274(.A1(new_n17030_), .A2(new_n17031_), .B(new_n17039_), .ZN(new_n17300_));
  INV_X1     g16275(.I(new_n17300_), .ZN(new_n17301_));
  AOI22_X1   g16276(.A1(new_n17301_), .A2(new_n17023_), .B1(new_n17047_), .B2(new_n17299_), .ZN(new_n17302_));
  NOR2_X1    g16277(.A1(new_n16968_), .A2(new_n16972_), .ZN(new_n17303_));
  OAI21_X1   g16278(.A1(new_n16954_), .A2(new_n16955_), .B(new_n16971_), .ZN(new_n17304_));
  NOR3_X1    g16279(.A1(new_n16966_), .A2(new_n17303_), .A3(new_n17304_), .ZN(new_n17305_));
  NOR2_X1    g16280(.A1(new_n16997_), .A2(new_n17305_), .ZN(new_n17306_));
  NOR2_X1    g16281(.A1(new_n16967_), .A2(new_n16974_), .ZN(new_n17307_));
  NOR3_X1    g16282(.A1(new_n17302_), .A2(new_n17306_), .A3(new_n17307_), .ZN(new_n17308_));
  OAI21_X1   g16283(.A1(new_n17296_), .A2(new_n17019_), .B(new_n17308_), .ZN(new_n17309_));
  INV_X1     g16284(.I(new_n16980_), .ZN(new_n17310_));
  NAND3_X1   g16285(.A1(new_n17310_), .A2(new_n16981_), .A3(new_n16987_), .ZN(new_n17311_));
  NAND4_X1   g16286(.A1(new_n17047_), .A2(new_n17037_), .A3(new_n17045_), .A4(new_n17298_), .ZN(new_n17312_));
  OAI21_X1   g16287(.A1(new_n17024_), .A2(new_n17300_), .B(new_n17312_), .ZN(new_n17313_));
  INV_X1     g16288(.I(new_n17306_), .ZN(new_n17314_));
  INV_X1     g16289(.I(new_n17307_), .ZN(new_n17315_));
  NAND3_X1   g16290(.A1(new_n17313_), .A2(new_n17314_), .A3(new_n17315_), .ZN(new_n17316_));
  NAND3_X1   g16291(.A1(new_n17316_), .A2(new_n17014_), .A3(new_n17311_), .ZN(new_n17317_));
  AOI21_X1   g16292(.A1(new_n17309_), .A2(new_n17317_), .B(new_n17295_), .ZN(new_n17318_));
  INV_X1     g16293(.I(new_n17295_), .ZN(new_n17319_));
  AOI21_X1   g16294(.A1(new_n17014_), .A2(new_n17311_), .B(new_n17316_), .ZN(new_n17320_));
  NOR3_X1    g16295(.A1(new_n17308_), .A2(new_n17296_), .A3(new_n17019_), .ZN(new_n17321_));
  NOR3_X1    g16296(.A1(new_n17320_), .A2(new_n17319_), .A3(new_n17321_), .ZN(new_n17322_));
  NOR2_X1    g16297(.A1(new_n17322_), .A2(new_n17318_), .ZN(new_n17323_));
  AOI22_X1   g16298(.A1(new_n16834_), .A2(new_n16838_), .B1(new_n16915_), .B2(new_n16924_), .ZN(new_n17324_));
  OAI21_X1   g16299(.A1(new_n16746_), .A2(new_n17324_), .B(new_n16931_), .ZN(new_n17325_));
  NOR2_X1    g16300(.A1(new_n16119_), .A2(new_n16186_), .ZN(new_n17326_));
  INV_X1     g16301(.I(new_n17326_), .ZN(new_n17327_));
  NOR2_X1    g16302(.A1(new_n16871_), .A2(new_n16177_), .ZN(new_n17328_));
  NOR2_X1    g16303(.A1(new_n16873_), .A2(new_n16861_), .ZN(new_n17329_));
  XOR2_X1    g16304(.A1(new_n17329_), .A2(new_n16868_), .Z(new_n17330_));
  AND2_X2    g16305(.A1(new_n16894_), .A2(new_n16895_), .Z(new_n17331_));
  XOR2_X1    g16306(.A1(new_n17331_), .A2(new_n16902_), .Z(new_n17332_));
  NOR2_X1    g16307(.A1(new_n16856_), .A2(new_n16889_), .ZN(new_n17333_));
  NAND4_X1   g16308(.A1(new_n17330_), .A2(new_n17332_), .A3(new_n17333_), .A4(new_n17328_), .ZN(new_n17334_));
  NOR2_X1    g16309(.A1(new_n17328_), .A2(new_n16877_), .ZN(new_n17335_));
  NOR2_X1    g16310(.A1(new_n17326_), .A2(new_n16888_), .ZN(new_n17336_));
  NOR4_X1    g16311(.A1(new_n17334_), .A2(new_n17327_), .A3(new_n17335_), .A4(new_n17336_), .ZN(new_n17337_));
  INV_X1     g16312(.I(new_n17337_), .ZN(new_n17338_));
  NAND2_X1   g16313(.A1(new_n16855_), .A2(new_n16864_), .ZN(new_n17339_));
  NOR2_X1    g16314(.A1(new_n16856_), .A2(new_n17339_), .ZN(new_n17340_));
  NAND2_X1   g16315(.A1(new_n17329_), .A2(new_n16865_), .ZN(new_n17341_));
  NOR3_X1    g16316(.A1(new_n17341_), .A2(new_n16871_), .A3(new_n16177_), .ZN(new_n17342_));
  NOR2_X1    g16317(.A1(new_n17342_), .A2(new_n17340_), .ZN(new_n17343_));
  NOR2_X1    g16318(.A1(new_n17329_), .A2(new_n16868_), .ZN(new_n17344_));
  INV_X1     g16319(.I(new_n17344_), .ZN(new_n17345_));
  NOR2_X1    g16320(.A1(new_n16900_), .A2(new_n16896_), .ZN(new_n17346_));
  INV_X1     g16321(.I(new_n16901_), .ZN(new_n17347_));
  NOR4_X1    g16322(.A1(new_n16894_), .A2(new_n17346_), .A3(new_n16895_), .A4(new_n17347_), .ZN(new_n17348_));
  INV_X1     g16323(.I(new_n17348_), .ZN(new_n17349_));
  OAI21_X1   g16324(.A1(new_n17326_), .A2(new_n16888_), .B(new_n17349_), .ZN(new_n17350_));
  OR2_X2     g16325(.A1(new_n17331_), .A2(new_n16902_), .Z(new_n17351_));
  NAND4_X1   g16326(.A1(new_n17343_), .A2(new_n17345_), .A3(new_n17350_), .A4(new_n17351_), .ZN(new_n17352_));
  AOI21_X1   g16327(.A1(new_n16916_), .A2(new_n16942_), .B(new_n17352_), .ZN(new_n17353_));
  NAND2_X1   g16328(.A1(new_n17350_), .A2(new_n17351_), .ZN(new_n17354_));
  NOR4_X1    g16329(.A1(new_n17354_), .A2(new_n17340_), .A3(new_n17342_), .A4(new_n17344_), .ZN(new_n17355_));
  NOR3_X1    g16330(.A1(new_n16839_), .A2(new_n16923_), .A3(new_n17355_), .ZN(new_n17356_));
  OAI21_X1   g16331(.A1(new_n17356_), .A2(new_n17353_), .B(new_n17338_), .ZN(new_n17357_));
  OAI21_X1   g16332(.A1(new_n16839_), .A2(new_n16923_), .B(new_n17355_), .ZN(new_n17358_));
  NAND3_X1   g16333(.A1(new_n16916_), .A2(new_n16942_), .A3(new_n17352_), .ZN(new_n17359_));
  NAND3_X1   g16334(.A1(new_n17358_), .A2(new_n17359_), .A3(new_n17337_), .ZN(new_n17360_));
  NAND2_X1   g16335(.A1(new_n17357_), .A2(new_n17360_), .ZN(new_n17361_));
  NOR2_X1    g16336(.A1(new_n16202_), .A2(new_n16336_), .ZN(new_n17362_));
  NAND2_X1   g16337(.A1(new_n16342_), .A2(new_n16329_), .ZN(new_n17363_));
  NOR2_X1    g16338(.A1(new_n16777_), .A2(new_n16778_), .ZN(new_n17364_));
  XNOR2_X1   g16339(.A1(new_n17364_), .A2(new_n16772_), .ZN(new_n17365_));
  NOR2_X1    g16340(.A1(new_n16806_), .A2(new_n16807_), .ZN(new_n17366_));
  XOR2_X1    g16341(.A1(new_n17366_), .A2(new_n16814_), .Z(new_n17367_));
  NAND2_X1   g16342(.A1(new_n16782_), .A2(new_n16802_), .ZN(new_n17368_));
  NOR4_X1    g16343(.A1(new_n17368_), .A2(new_n17365_), .A3(new_n17367_), .A4(new_n17363_), .ZN(new_n17369_));
  NOR2_X1    g16344(.A1(new_n17362_), .A2(new_n16802_), .ZN(new_n17370_));
  AOI21_X1   g16345(.A1(new_n16763_), .A2(new_n17363_), .B(new_n17370_), .ZN(new_n17371_));
  NAND3_X1   g16346(.A1(new_n17371_), .A2(new_n17369_), .A3(new_n17362_), .ZN(new_n17372_));
  INV_X1     g16347(.I(new_n17372_), .ZN(new_n17373_));
  NOR2_X1    g16348(.A1(new_n16761_), .A2(new_n16769_), .ZN(new_n17374_));
  NAND2_X1   g16349(.A1(new_n16782_), .A2(new_n17374_), .ZN(new_n17375_));
  NOR2_X1    g16350(.A1(new_n16327_), .A2(new_n16775_), .ZN(new_n17376_));
  NOR3_X1    g16351(.A1(new_n16777_), .A2(new_n16778_), .A3(new_n16770_), .ZN(new_n17377_));
  NAND2_X1   g16352(.A1(new_n17376_), .A2(new_n17377_), .ZN(new_n17378_));
  OAI22_X1   g16353(.A1(new_n16777_), .A2(new_n16778_), .B1(new_n16757_), .B2(new_n16771_), .ZN(new_n17379_));
  NAND3_X1   g16354(.A1(new_n17378_), .A2(new_n17375_), .A3(new_n17379_), .ZN(new_n17380_));
  INV_X1     g16355(.I(new_n16795_), .ZN(new_n17381_));
  NOR3_X1    g16356(.A1(new_n16801_), .A2(new_n17381_), .A3(new_n16810_), .ZN(new_n17382_));
  INV_X1     g16357(.I(new_n17382_), .ZN(new_n17383_));
  NAND2_X1   g16358(.A1(new_n16817_), .A2(new_n16818_), .ZN(new_n17384_));
  NOR2_X1    g16359(.A1(new_n17384_), .A2(new_n16811_), .ZN(new_n17385_));
  NAND3_X1   g16360(.A1(new_n17385_), .A2(new_n16262_), .A3(new_n16264_), .ZN(new_n17386_));
  NOR2_X1    g16361(.A1(new_n17366_), .A2(new_n16813_), .ZN(new_n17387_));
  INV_X1     g16362(.I(new_n17387_), .ZN(new_n17388_));
  NAND3_X1   g16363(.A1(new_n17383_), .A2(new_n17386_), .A3(new_n17388_), .ZN(new_n17389_));
  NOR2_X1    g16364(.A1(new_n17380_), .A2(new_n17389_), .ZN(new_n17390_));
  OAI21_X1   g16365(.A1(new_n16747_), .A2(new_n16837_), .B(new_n17390_), .ZN(new_n17391_));
  NAND2_X1   g16366(.A1(new_n16201_), .A2(new_n16364_), .ZN(new_n17392_));
  AOI22_X1   g16367(.A1(new_n17376_), .A2(new_n17377_), .B1(new_n16782_), .B2(new_n17374_), .ZN(new_n17393_));
  NOR4_X1    g16368(.A1(new_n16202_), .A2(new_n16336_), .A3(new_n17384_), .A4(new_n16811_), .ZN(new_n17394_));
  NOR3_X1    g16369(.A1(new_n17394_), .A2(new_n17382_), .A3(new_n17387_), .ZN(new_n17395_));
  NAND3_X1   g16370(.A1(new_n17395_), .A2(new_n17393_), .A3(new_n17379_), .ZN(new_n17396_));
  NAND4_X1   g16371(.A1(new_n17392_), .A2(new_n16936_), .A3(new_n16365_), .A4(new_n17396_), .ZN(new_n17397_));
  AOI21_X1   g16372(.A1(new_n17391_), .A2(new_n17397_), .B(new_n17373_), .ZN(new_n17398_));
  AOI21_X1   g16373(.A1(new_n16835_), .A2(new_n16936_), .B(new_n17396_), .ZN(new_n17399_));
  NOR3_X1    g16374(.A1(new_n16747_), .A2(new_n16837_), .A3(new_n17390_), .ZN(new_n17400_));
  NOR3_X1    g16375(.A1(new_n17400_), .A2(new_n17399_), .A3(new_n17372_), .ZN(new_n17401_));
  NOR2_X1    g16376(.A1(new_n17401_), .A2(new_n17398_), .ZN(new_n17402_));
  NOR2_X1    g16377(.A1(new_n17402_), .A2(new_n17361_), .ZN(new_n17403_));
  AOI21_X1   g16378(.A1(new_n17358_), .A2(new_n17359_), .B(new_n17337_), .ZN(new_n17404_));
  NOR3_X1    g16379(.A1(new_n17356_), .A2(new_n17353_), .A3(new_n17338_), .ZN(new_n17405_));
  NOR2_X1    g16380(.A1(new_n17405_), .A2(new_n17404_), .ZN(new_n17406_));
  OAI21_X1   g16381(.A1(new_n17400_), .A2(new_n17399_), .B(new_n17372_), .ZN(new_n17407_));
  NAND3_X1   g16382(.A1(new_n17391_), .A2(new_n17397_), .A3(new_n17373_), .ZN(new_n17408_));
  NAND2_X1   g16383(.A1(new_n17407_), .A2(new_n17408_), .ZN(new_n17409_));
  NOR2_X1    g16384(.A1(new_n17409_), .A2(new_n17406_), .ZN(new_n17410_));
  OAI21_X1   g16385(.A1(new_n17410_), .A2(new_n17403_), .B(new_n17325_), .ZN(new_n17411_));
  NOR4_X1    g16386(.A1(new_n16934_), .A2(new_n16937_), .A3(new_n16943_), .A4(new_n16940_), .ZN(new_n17412_));
  AOI21_X1   g16387(.A1(new_n16930_), .A2(new_n16944_), .B(new_n17412_), .ZN(new_n17413_));
  NOR2_X1    g16388(.A1(new_n17402_), .A2(new_n17406_), .ZN(new_n17414_));
  NOR2_X1    g16389(.A1(new_n17409_), .A2(new_n17361_), .ZN(new_n17415_));
  OAI21_X1   g16390(.A1(new_n17414_), .A2(new_n17415_), .B(new_n17413_), .ZN(new_n17416_));
  AOI21_X1   g16391(.A1(new_n17411_), .A2(new_n17416_), .B(new_n17323_), .ZN(new_n17417_));
  OAI21_X1   g16392(.A1(new_n17320_), .A2(new_n17321_), .B(new_n17319_), .ZN(new_n17418_));
  NAND3_X1   g16393(.A1(new_n17309_), .A2(new_n17317_), .A3(new_n17295_), .ZN(new_n17419_));
  NAND2_X1   g16394(.A1(new_n17418_), .A2(new_n17419_), .ZN(new_n17420_));
  NAND2_X1   g16395(.A1(new_n17409_), .A2(new_n17406_), .ZN(new_n17421_));
  NAND2_X1   g16396(.A1(new_n17402_), .A2(new_n17361_), .ZN(new_n17422_));
  AOI21_X1   g16397(.A1(new_n17421_), .A2(new_n17422_), .B(new_n17413_), .ZN(new_n17423_));
  NAND2_X1   g16398(.A1(new_n17409_), .A2(new_n17361_), .ZN(new_n17424_));
  NAND2_X1   g16399(.A1(new_n17402_), .A2(new_n17406_), .ZN(new_n17425_));
  AOI21_X1   g16400(.A1(new_n17425_), .A2(new_n17424_), .B(new_n17325_), .ZN(new_n17426_));
  NOR3_X1    g16401(.A1(new_n17423_), .A2(new_n17426_), .A3(new_n17420_), .ZN(new_n17427_));
  OAI21_X1   g16402(.A1(new_n17427_), .A2(new_n17417_), .B(new_n17294_), .ZN(new_n17428_));
  INV_X1     g16403(.I(new_n17291_), .ZN(new_n17429_));
  NOR2_X1    g16404(.A1(new_n17292_), .A2(new_n17293_), .ZN(new_n17430_));
  NOR2_X1    g16405(.A1(new_n17430_), .A2(new_n17429_), .ZN(new_n17431_));
  AOI21_X1   g16406(.A1(new_n17411_), .A2(new_n17416_), .B(new_n17420_), .ZN(new_n17432_));
  NOR3_X1    g16407(.A1(new_n17423_), .A2(new_n17426_), .A3(new_n17323_), .ZN(new_n17433_));
  OAI21_X1   g16408(.A1(new_n17433_), .A2(new_n17432_), .B(new_n17431_), .ZN(new_n17434_));
  NAND2_X1   g16409(.A1(new_n17428_), .A2(new_n17434_), .ZN(new_n17435_));
  NAND4_X1   g16410(.A1(new_n17158_), .A2(new_n17242_), .A3(new_n17153_), .A4(new_n17238_), .ZN(new_n17436_));
  OAI21_X1   g16411(.A1(new_n17076_), .A2(new_n17243_), .B(new_n17436_), .ZN(new_n17437_));
  NOR2_X1    g16412(.A1(new_n16548_), .A2(new_n17209_), .ZN(new_n17438_));
  NAND2_X1   g16413(.A1(new_n17172_), .A2(new_n16515_), .ZN(new_n17439_));
  NAND2_X1   g16414(.A1(new_n17174_), .A2(new_n17170_), .ZN(new_n17440_));
  XNOR2_X1   g16415(.A1(new_n17440_), .A2(new_n17439_), .ZN(new_n17441_));
  XOR2_X1    g16416(.A1(new_n17205_), .A2(new_n17200_), .Z(new_n17442_));
  NAND3_X1   g16417(.A1(new_n17442_), .A2(new_n17168_), .A3(new_n17194_), .ZN(new_n17443_));
  NOR4_X1    g16418(.A1(new_n17443_), .A2(new_n16537_), .A3(new_n17441_), .A4(new_n17169_), .ZN(new_n17444_));
  NOR2_X1    g16419(.A1(new_n17169_), .A2(new_n16537_), .ZN(new_n17445_));
  NOR2_X1    g16420(.A1(new_n17445_), .A2(new_n17168_), .ZN(new_n17446_));
  NOR2_X1    g16421(.A1(new_n17438_), .A2(new_n17194_), .ZN(new_n17447_));
  NOR2_X1    g16422(.A1(new_n17446_), .A2(new_n17447_), .ZN(new_n17448_));
  NAND3_X1   g16423(.A1(new_n17448_), .A2(new_n17444_), .A3(new_n17438_), .ZN(new_n17449_));
  INV_X1     g16424(.I(new_n17449_), .ZN(new_n17450_));
  NAND3_X1   g16425(.A1(new_n17160_), .A2(new_n16709_), .A3(new_n17240_), .ZN(new_n17451_));
  OR4_X2     g16426(.A1(new_n16504_), .A2(new_n16507_), .A3(new_n16505_), .A4(new_n16508_), .Z(new_n17452_));
  OAI22_X1   g16427(.A1(new_n16504_), .A2(new_n16508_), .B1(new_n16505_), .B2(new_n16507_), .ZN(new_n17453_));
  OR4_X2     g16428(.A1(new_n16478_), .A2(new_n16482_), .A3(new_n16480_), .A4(new_n16483_), .Z(new_n17454_));
  OAI22_X1   g16429(.A1(new_n16478_), .A2(new_n16483_), .B1(new_n16482_), .B2(new_n16480_), .ZN(new_n17455_));
  AND4_X2    g16430(.A1(new_n17452_), .A2(new_n17454_), .A3(new_n17453_), .A4(new_n17455_), .Z(new_n17456_));
  NAND3_X1   g16431(.A1(new_n17165_), .A2(new_n17166_), .A3(new_n17456_), .ZN(new_n17457_));
  NAND2_X1   g16432(.A1(new_n17440_), .A2(new_n17439_), .ZN(new_n17458_));
  NOR2_X1    g16433(.A1(new_n17458_), .A2(new_n17457_), .ZN(new_n17459_));
  OAI21_X1   g16434(.A1(new_n17445_), .A2(new_n17459_), .B(new_n17168_), .ZN(new_n17460_));
  OR4_X2     g16435(.A1(new_n16433_), .A2(new_n16437_), .A3(new_n16435_), .A4(new_n16439_), .Z(new_n17461_));
  OAI22_X1   g16436(.A1(new_n16437_), .A2(new_n16435_), .B1(new_n16433_), .B2(new_n16439_), .ZN(new_n17462_));
  OR4_X2     g16437(.A1(new_n17202_), .A2(new_n16405_), .A3(new_n17203_), .A4(new_n16406_), .Z(new_n17463_));
  OAI22_X1   g16438(.A1(new_n17202_), .A2(new_n16406_), .B1(new_n17203_), .B2(new_n16405_), .ZN(new_n17464_));
  AND4_X2    g16439(.A1(new_n17461_), .A2(new_n17463_), .A3(new_n17462_), .A4(new_n17464_), .Z(new_n17465_));
  NAND3_X1   g16440(.A1(new_n17465_), .A2(new_n17191_), .A3(new_n17192_), .ZN(new_n17466_));
  NAND2_X1   g16441(.A1(new_n17205_), .A2(new_n17200_), .ZN(new_n17467_));
  OAI22_X1   g16442(.A1(new_n16548_), .A2(new_n17209_), .B1(new_n17466_), .B2(new_n17467_), .ZN(new_n17468_));
  NAND2_X1   g16443(.A1(new_n17468_), .A2(new_n17194_), .ZN(new_n17469_));
  NOR2_X1    g16444(.A1(new_n17469_), .A2(new_n17460_), .ZN(new_n17470_));
  NAND2_X1   g16445(.A1(new_n17451_), .A2(new_n17470_), .ZN(new_n17471_));
  NOR2_X1    g16446(.A1(new_n17235_), .A2(new_n16536_), .ZN(new_n17472_));
  INV_X1     g16447(.I(new_n17470_), .ZN(new_n17473_));
  NAND3_X1   g16448(.A1(new_n17472_), .A2(new_n17240_), .A3(new_n17473_), .ZN(new_n17474_));
  AOI21_X1   g16449(.A1(new_n17474_), .A2(new_n17471_), .B(new_n17450_), .ZN(new_n17475_));
  AOI21_X1   g16450(.A1(new_n17472_), .A2(new_n17240_), .B(new_n17473_), .ZN(new_n17476_));
  NOR2_X1    g16451(.A1(new_n17451_), .A2(new_n17470_), .ZN(new_n17477_));
  NOR3_X1    g16452(.A1(new_n17476_), .A2(new_n17477_), .A3(new_n17449_), .ZN(new_n17478_));
  NAND2_X1   g16453(.A1(new_n16622_), .A2(new_n17085_), .ZN(new_n17479_));
  INV_X1     g16454(.I(new_n17479_), .ZN(new_n17480_));
  NAND2_X1   g16455(.A1(new_n17479_), .A2(new_n17084_), .ZN(new_n17481_));
  NOR2_X1    g16456(.A1(new_n17136_), .A2(new_n16615_), .ZN(new_n17482_));
  INV_X1     g16457(.I(new_n17482_), .ZN(new_n17483_));
  NAND2_X1   g16458(.A1(new_n17483_), .A2(new_n17119_), .ZN(new_n17484_));
  XNOR2_X1   g16459(.A1(new_n17100_), .A2(new_n17092_), .ZN(new_n17485_));
  XOR2_X1    g16460(.A1(new_n17129_), .A2(new_n17132_), .Z(new_n17486_));
  NAND2_X1   g16461(.A1(new_n17106_), .A2(new_n17118_), .ZN(new_n17487_));
  NOR4_X1    g16462(.A1(new_n17487_), .A2(new_n17483_), .A3(new_n17485_), .A4(new_n17486_), .ZN(new_n17488_));
  NAND4_X1   g16463(.A1(new_n17488_), .A2(new_n17480_), .A3(new_n17481_), .A4(new_n17484_), .ZN(new_n17489_));
  INV_X1     g16464(.I(new_n17489_), .ZN(new_n17490_));
  NOR3_X1    g16465(.A1(new_n17147_), .A2(new_n17144_), .A3(new_n17146_), .ZN(new_n17491_));
  AOI21_X1   g16466(.A1(new_n17096_), .A2(new_n17081_), .B(new_n17095_), .ZN(new_n17492_));
  AOI21_X1   g16467(.A1(new_n17092_), .A2(new_n17492_), .B(new_n16632_), .ZN(new_n17493_));
  NOR3_X1    g16468(.A1(new_n17493_), .A2(new_n14002_), .A3(new_n16633_), .ZN(new_n17494_));
  NOR2_X1    g16469(.A1(new_n17100_), .A2(new_n17092_), .ZN(new_n17495_));
  AOI22_X1   g16470(.A1(new_n16622_), .A2(new_n17085_), .B1(new_n17494_), .B2(new_n17495_), .ZN(new_n17496_));
  INV_X1     g16471(.I(new_n16578_), .ZN(new_n17497_));
  NAND3_X1   g16472(.A1(new_n16573_), .A2(new_n16575_), .A3(new_n16579_), .ZN(new_n17498_));
  AND2_X2    g16473(.A1(new_n16573_), .A2(new_n16579_), .Z(new_n17499_));
  NOR4_X1    g16474(.A1(new_n17499_), .A2(new_n16575_), .A3(new_n17497_), .A4(new_n17498_), .ZN(new_n17500_));
  NAND2_X1   g16475(.A1(new_n17129_), .A2(new_n17500_), .ZN(new_n17501_));
  AOI21_X1   g16476(.A1(new_n17501_), .A2(new_n17120_), .B(new_n16572_), .ZN(new_n17502_));
  NOR2_X1    g16477(.A1(new_n17129_), .A2(new_n17133_), .ZN(new_n17503_));
  AOI21_X1   g16478(.A1(new_n17502_), .A2(new_n17503_), .B(new_n17482_), .ZN(new_n17504_));
  NOR4_X1    g16479(.A1(new_n17504_), .A2(new_n17084_), .A3(new_n17119_), .A4(new_n17496_), .ZN(new_n17505_));
  OAI21_X1   g16480(.A1(new_n17077_), .A2(new_n17491_), .B(new_n17505_), .ZN(new_n17506_));
  INV_X1     g16481(.I(new_n17505_), .ZN(new_n17507_));
  NAND3_X1   g16482(.A1(new_n17154_), .A2(new_n17156_), .A3(new_n17507_), .ZN(new_n17508_));
  AOI21_X1   g16483(.A1(new_n17506_), .A2(new_n17508_), .B(new_n17490_), .ZN(new_n17509_));
  AOI21_X1   g16484(.A1(new_n17154_), .A2(new_n17156_), .B(new_n17507_), .ZN(new_n17510_));
  NOR3_X1    g16485(.A1(new_n17077_), .A2(new_n17491_), .A3(new_n17505_), .ZN(new_n17511_));
  NOR3_X1    g16486(.A1(new_n17511_), .A2(new_n17510_), .A3(new_n17489_), .ZN(new_n17512_));
  NOR2_X1    g16487(.A1(new_n17512_), .A2(new_n17509_), .ZN(new_n17513_));
  NOR3_X1    g16488(.A1(new_n17513_), .A2(new_n17478_), .A3(new_n17475_), .ZN(new_n17514_));
  OAI21_X1   g16489(.A1(new_n17476_), .A2(new_n17477_), .B(new_n17449_), .ZN(new_n17515_));
  NAND3_X1   g16490(.A1(new_n17474_), .A2(new_n17471_), .A3(new_n17450_), .ZN(new_n17516_));
  OAI21_X1   g16491(.A1(new_n17511_), .A2(new_n17510_), .B(new_n17489_), .ZN(new_n17517_));
  NAND3_X1   g16492(.A1(new_n17506_), .A2(new_n17508_), .A3(new_n17490_), .ZN(new_n17518_));
  NAND2_X1   g16493(.A1(new_n17517_), .A2(new_n17518_), .ZN(new_n17519_));
  AOI21_X1   g16494(.A1(new_n17515_), .A2(new_n17516_), .B(new_n17519_), .ZN(new_n17520_));
  OAI21_X1   g16495(.A1(new_n17520_), .A2(new_n17514_), .B(new_n17437_), .ZN(new_n17521_));
  NAND4_X1   g16496(.A1(new_n16547_), .A2(new_n16557_), .A3(new_n16698_), .A4(new_n16704_), .ZN(new_n17522_));
  OAI21_X1   g16497(.A1(new_n16388_), .A2(new_n16722_), .B(new_n17522_), .ZN(new_n17523_));
  OAI22_X1   g16498(.A1(new_n17229_), .A2(new_n17224_), .B1(new_n17233_), .B2(new_n17232_), .ZN(new_n17524_));
  AOI21_X1   g16499(.A1(new_n17523_), .A2(new_n17524_), .B(new_n17234_), .ZN(new_n17525_));
  AOI21_X1   g16500(.A1(new_n17515_), .A2(new_n17516_), .B(new_n17513_), .ZN(new_n17526_));
  NOR3_X1    g16501(.A1(new_n17478_), .A2(new_n17519_), .A3(new_n17475_), .ZN(new_n17527_));
  OAI21_X1   g16502(.A1(new_n17526_), .A2(new_n17527_), .B(new_n17525_), .ZN(new_n17528_));
  NAND2_X1   g16503(.A1(new_n17521_), .A2(new_n17528_), .ZN(new_n17529_));
  NAND2_X1   g16504(.A1(new_n17063_), .A2(new_n17060_), .ZN(new_n17530_));
  AOI21_X1   g16505(.A1(new_n17253_), .A2(new_n16375_), .B(new_n16946_), .ZN(new_n17531_));
  NAND3_X1   g16506(.A1(new_n17253_), .A2(new_n16375_), .A3(new_n16946_), .ZN(new_n17532_));
  AOI21_X1   g16507(.A1(new_n17530_), .A2(new_n17532_), .B(new_n17531_), .ZN(new_n17533_));
  NOR2_X1    g16508(.A1(new_n17533_), .A2(new_n17529_), .ZN(new_n17534_));
  NAND3_X1   g16509(.A1(new_n17519_), .A2(new_n17515_), .A3(new_n17516_), .ZN(new_n17535_));
  OAI21_X1   g16510(.A1(new_n17475_), .A2(new_n17478_), .B(new_n17513_), .ZN(new_n17536_));
  AOI21_X1   g16511(.A1(new_n17536_), .A2(new_n17535_), .B(new_n17525_), .ZN(new_n17537_));
  OAI21_X1   g16512(.A1(new_n17475_), .A2(new_n17478_), .B(new_n17519_), .ZN(new_n17538_));
  NAND3_X1   g16513(.A1(new_n17513_), .A2(new_n17515_), .A3(new_n17516_), .ZN(new_n17539_));
  AOI21_X1   g16514(.A1(new_n17538_), .A2(new_n17539_), .B(new_n17437_), .ZN(new_n17540_));
  NOR2_X1    g16515(.A1(new_n17540_), .A2(new_n17537_), .ZN(new_n17541_));
  NOR3_X1    g16516(.A1(new_n17061_), .A2(new_n17062_), .A3(new_n16952_), .ZN(new_n17542_));
  AOI21_X1   g16517(.A1(new_n17059_), .A2(new_n17052_), .B(new_n16953_), .ZN(new_n17543_));
  NOR2_X1    g16518(.A1(new_n17542_), .A2(new_n17543_), .ZN(new_n17544_));
  OAI21_X1   g16519(.A1(new_n16744_), .A2(new_n16742_), .B(new_n17065_), .ZN(new_n17545_));
  NOR3_X1    g16520(.A1(new_n16744_), .A2(new_n16742_), .A3(new_n17065_), .ZN(new_n17546_));
  OAI21_X1   g16521(.A1(new_n17544_), .A2(new_n17546_), .B(new_n17545_), .ZN(new_n17547_));
  NOR2_X1    g16522(.A1(new_n17547_), .A2(new_n17541_), .ZN(new_n17548_));
  OAI21_X1   g16523(.A1(new_n17534_), .A2(new_n17548_), .B(new_n17435_), .ZN(new_n17549_));
  OAI21_X1   g16524(.A1(new_n17423_), .A2(new_n17426_), .B(new_n17420_), .ZN(new_n17550_));
  NAND3_X1   g16525(.A1(new_n17411_), .A2(new_n17416_), .A3(new_n17323_), .ZN(new_n17551_));
  AOI21_X1   g16526(.A1(new_n17550_), .A2(new_n17551_), .B(new_n17431_), .ZN(new_n17552_));
  OAI21_X1   g16527(.A1(new_n17423_), .A2(new_n17426_), .B(new_n17323_), .ZN(new_n17553_));
  NAND3_X1   g16528(.A1(new_n17411_), .A2(new_n17416_), .A3(new_n17420_), .ZN(new_n17554_));
  AOI21_X1   g16529(.A1(new_n17553_), .A2(new_n17554_), .B(new_n17294_), .ZN(new_n17555_));
  NOR2_X1    g16530(.A1(new_n17552_), .A2(new_n17555_), .ZN(new_n17556_));
  NOR2_X1    g16531(.A1(new_n17533_), .A2(new_n17541_), .ZN(new_n17557_));
  NOR2_X1    g16532(.A1(new_n17529_), .A2(new_n17547_), .ZN(new_n17558_));
  OAI21_X1   g16533(.A1(new_n17558_), .A2(new_n17557_), .B(new_n17556_), .ZN(new_n17559_));
  NAND2_X1   g16534(.A1(new_n17549_), .A2(new_n17559_), .ZN(new_n17560_));
  XNOR2_X1   g16535(.A1(new_n17159_), .A2(new_n17230_), .ZN(new_n17561_));
  AOI21_X1   g16536(.A1(new_n17436_), .A2(new_n17524_), .B(new_n17523_), .ZN(new_n17562_));
  AOI21_X1   g16537(.A1(new_n17561_), .A2(new_n17523_), .B(new_n17562_), .ZN(new_n17563_));
  AOI21_X1   g16538(.A1(new_n17074_), .A2(new_n17071_), .B(new_n17563_), .ZN(new_n17564_));
  NAND3_X1   g16539(.A1(new_n17074_), .A2(new_n17071_), .A3(new_n17563_), .ZN(new_n17565_));
  OAI21_X1   g16540(.A1(new_n17542_), .A2(new_n17543_), .B(new_n17065_), .ZN(new_n17566_));
  AOI21_X1   g16541(.A1(new_n17059_), .A2(new_n17052_), .B(new_n16952_), .ZN(new_n17567_));
  NOR3_X1    g16542(.A1(new_n17061_), .A2(new_n17062_), .A3(new_n16953_), .ZN(new_n17568_));
  OAI21_X1   g16543(.A1(new_n17568_), .A2(new_n17567_), .B(new_n16946_), .ZN(new_n17569_));
  NAND3_X1   g16544(.A1(new_n17566_), .A2(new_n17569_), .A3(new_n17254_), .ZN(new_n17570_));
  OAI21_X1   g16545(.A1(new_n17064_), .A2(new_n17068_), .B(new_n16745_), .ZN(new_n17571_));
  NAND2_X1   g16546(.A1(new_n17570_), .A2(new_n17571_), .ZN(new_n17572_));
  AOI21_X1   g16547(.A1(new_n17572_), .A2(new_n17565_), .B(new_n17564_), .ZN(new_n17573_));
  NOR2_X1    g16548(.A1(new_n17560_), .A2(new_n17573_), .ZN(new_n17574_));
  NAND2_X1   g16549(.A1(new_n17547_), .A2(new_n17541_), .ZN(new_n17575_));
  NAND2_X1   g16550(.A1(new_n17533_), .A2(new_n17529_), .ZN(new_n17576_));
  AOI21_X1   g16551(.A1(new_n17576_), .A2(new_n17575_), .B(new_n17556_), .ZN(new_n17577_));
  NAND2_X1   g16552(.A1(new_n17529_), .A2(new_n17547_), .ZN(new_n17578_));
  NAND2_X1   g16553(.A1(new_n17533_), .A2(new_n17541_), .ZN(new_n17579_));
  AOI21_X1   g16554(.A1(new_n17578_), .A2(new_n17579_), .B(new_n17435_), .ZN(new_n17580_));
  NOR2_X1    g16555(.A1(new_n17577_), .A2(new_n17580_), .ZN(new_n17581_));
  XOR2_X1    g16556(.A1(new_n16558_), .A2(new_n16706_), .Z(new_n17582_));
  INV_X1     g16557(.I(new_n16723_), .ZN(new_n17583_));
  AOI21_X1   g16558(.A1(new_n17582_), .A2(new_n16389_), .B(new_n17583_), .ZN(new_n17584_));
  NOR2_X1    g16559(.A1(new_n16735_), .A2(new_n17584_), .ZN(new_n17585_));
  NAND3_X1   g16560(.A1(new_n16385_), .A2(new_n16375_), .A3(new_n16387_), .ZN(new_n17586_));
  OAI21_X1   g16561(.A1(new_n16742_), .A2(new_n16743_), .B(new_n16728_), .ZN(new_n17587_));
  AOI22_X1   g16562(.A1(new_n16735_), .A2(new_n17584_), .B1(new_n17586_), .B2(new_n17587_), .ZN(new_n17588_));
  OAI21_X1   g16563(.A1(new_n17588_), .A2(new_n17585_), .B(new_n17245_), .ZN(new_n17589_));
  NOR3_X1    g16564(.A1(new_n17588_), .A2(new_n17585_), .A3(new_n17245_), .ZN(new_n17590_));
  NOR3_X1    g16565(.A1(new_n17064_), .A2(new_n17068_), .A3(new_n16745_), .ZN(new_n17591_));
  AOI21_X1   g16566(.A1(new_n17566_), .A2(new_n17569_), .B(new_n17254_), .ZN(new_n17592_));
  NOR2_X1    g16567(.A1(new_n17592_), .A2(new_n17591_), .ZN(new_n17593_));
  OAI21_X1   g16568(.A1(new_n17590_), .A2(new_n17593_), .B(new_n17589_), .ZN(new_n17594_));
  NOR2_X1    g16569(.A1(new_n17581_), .A2(new_n17594_), .ZN(new_n17595_));
  NOR2_X1    g16570(.A1(new_n17595_), .A2(new_n17574_), .ZN(new_n17596_));
  AOI21_X1   g16571(.A1(new_n17252_), .A2(new_n17257_), .B(new_n17262_), .ZN(new_n17597_));
  NAND2_X1   g16572(.A1(new_n17596_), .A2(new_n17597_), .ZN(new_n17598_));
  XOR2_X1    g16573(.A1(new_n17560_), .A2(new_n17594_), .Z(new_n17599_));
  OAI21_X1   g16574(.A1(new_n17263_), .A2(new_n17264_), .B(new_n16741_), .ZN(new_n17600_));
  NAND2_X1   g16575(.A1(new_n17599_), .A2(new_n17600_), .ZN(new_n17601_));
  AOI21_X1   g16576(.A1(new_n17601_), .A2(new_n17598_), .B(new_n17289_), .ZN(new_n17602_));
  NAND2_X1   g16577(.A1(new_n17599_), .A2(new_n17597_), .ZN(new_n17603_));
  NAND2_X1   g16578(.A1(new_n17411_), .A2(new_n17416_), .ZN(new_n17604_));
  NAND2_X1   g16579(.A1(new_n17547_), .A2(new_n17604_), .ZN(new_n17605_));
  XOR2_X1    g16580(.A1(new_n17294_), .A2(new_n17420_), .Z(new_n17606_));
  OAI21_X1   g16581(.A1(new_n17547_), .A2(new_n17604_), .B(new_n17606_), .ZN(new_n17607_));
  NAND2_X1   g16582(.A1(new_n17607_), .A2(new_n17605_), .ZN(new_n17608_));
  XOR2_X1    g16583(.A1(new_n17308_), .A2(new_n17295_), .Z(new_n17609_));
  NAND4_X1   g16584(.A1(new_n17294_), .A2(new_n17014_), .A3(new_n17311_), .A4(new_n17609_), .ZN(new_n17612_));
  NOR2_X1    g16585(.A1(new_n16747_), .A2(new_n16837_), .ZN(new_n17613_));
  INV_X1     g16586(.I(new_n17613_), .ZN(new_n17614_));
  NOR2_X1    g16587(.A1(new_n17394_), .A2(new_n17382_), .ZN(new_n17615_));
  NOR4_X1    g16588(.A1(new_n17393_), .A2(new_n17615_), .A3(new_n17379_), .A4(new_n17388_), .ZN(new_n17616_));
  AOI21_X1   g16589(.A1(new_n17614_), .A2(new_n17372_), .B(new_n17616_), .ZN(new_n17617_));
  INV_X1     g16590(.I(new_n17380_), .ZN(new_n17618_));
  NOR2_X1    g16591(.A1(new_n17618_), .A2(new_n17395_), .ZN(new_n17619_));
  NOR2_X1    g16592(.A1(new_n17617_), .A2(new_n17619_), .ZN(new_n17620_));
  OR4_X2     g16593(.A1(new_n17343_), .A2(new_n17345_), .A3(new_n17350_), .A4(new_n17351_), .Z(new_n17621_));
  NAND2_X1   g16594(.A1(new_n16916_), .A2(new_n16942_), .ZN(new_n17622_));
  NAND2_X1   g16595(.A1(new_n17622_), .A2(new_n17338_), .ZN(new_n17623_));
  NAND2_X1   g16596(.A1(new_n17623_), .A2(new_n17621_), .ZN(new_n17624_));
  NAND2_X1   g16597(.A1(new_n17343_), .A2(new_n17345_), .ZN(new_n17625_));
  NAND2_X1   g16598(.A1(new_n17625_), .A2(new_n17354_), .ZN(new_n17626_));
  NAND2_X1   g16599(.A1(new_n17624_), .A2(new_n17626_), .ZN(new_n17627_));
  XOR2_X1    g16600(.A1(new_n17620_), .A2(new_n17627_), .Z(new_n17628_));
  INV_X1     g16601(.I(new_n17628_), .ZN(new_n17629_));
  NAND2_X1   g16602(.A1(new_n17425_), .A2(new_n17413_), .ZN(new_n17630_));
  NAND2_X1   g16603(.A1(new_n17614_), .A2(new_n17372_), .ZN(new_n17631_));
  XOR2_X1    g16604(.A1(new_n17625_), .A2(new_n17354_), .Z(new_n17632_));
  XOR2_X1    g16605(.A1(new_n17380_), .A2(new_n17389_), .Z(new_n17633_));
  NAND4_X1   g16606(.A1(new_n17632_), .A2(new_n17633_), .A3(new_n17337_), .A4(new_n17373_), .ZN(new_n17634_));
  NOR2_X1    g16607(.A1(new_n17634_), .A2(new_n17622_), .ZN(new_n17635_));
  NAND4_X1   g16608(.A1(new_n17635_), .A2(new_n17613_), .A3(new_n17631_), .A4(new_n17623_), .ZN(new_n17636_));
  NAND2_X1   g16609(.A1(new_n17630_), .A2(new_n17636_), .ZN(new_n17637_));
  NAND2_X1   g16610(.A1(new_n17629_), .A2(new_n17637_), .ZN(new_n17638_));
  NOR3_X1    g16611(.A1(new_n17628_), .A2(new_n17630_), .A3(new_n17636_), .ZN(new_n17639_));
  INV_X1     g16612(.I(new_n17639_), .ZN(new_n17640_));
  NOR2_X1    g16613(.A1(new_n17640_), .A2(new_n17638_), .ZN(new_n17641_));
  XOR2_X1    g16614(.A1(new_n17641_), .A2(new_n17612_), .Z(new_n17642_));
  NOR2_X1    g16615(.A1(new_n17573_), .A2(new_n17541_), .ZN(new_n17643_));
  NOR2_X1    g16616(.A1(new_n17533_), .A2(new_n17435_), .ZN(new_n17644_));
  NOR2_X1    g16617(.A1(new_n17547_), .A2(new_n17556_), .ZN(new_n17645_));
  NOR2_X1    g16618(.A1(new_n17644_), .A2(new_n17645_), .ZN(new_n17646_));
  AOI21_X1   g16619(.A1(new_n17573_), .A2(new_n17541_), .B(new_n17646_), .ZN(new_n17647_));
  INV_X1     g16620(.I(new_n17451_), .ZN(new_n17648_));
  NAND2_X1   g16621(.A1(new_n17154_), .A2(new_n17156_), .ZN(new_n17649_));
  INV_X1     g16622(.I(new_n17649_), .ZN(new_n17650_));
  NOR2_X1    g16623(.A1(new_n17496_), .A2(new_n17084_), .ZN(new_n17651_));
  NOR2_X1    g16624(.A1(new_n17504_), .A2(new_n17119_), .ZN(new_n17652_));
  XOR2_X1    g16625(.A1(new_n17652_), .A2(new_n17651_), .Z(new_n17653_));
  XNOR2_X1   g16626(.A1(new_n17469_), .A2(new_n17460_), .ZN(new_n17654_));
  NOR3_X1    g16627(.A1(new_n17654_), .A2(new_n17449_), .A3(new_n17489_), .ZN(new_n17655_));
  NAND4_X1   g16628(.A1(new_n17650_), .A2(new_n17648_), .A3(new_n17653_), .A4(new_n17655_), .ZN(new_n17656_));
  NOR2_X1    g16629(.A1(new_n17648_), .A2(new_n17450_), .ZN(new_n17657_));
  NOR2_X1    g16630(.A1(new_n17650_), .A2(new_n17490_), .ZN(new_n17658_));
  NOR3_X1    g16631(.A1(new_n17656_), .A2(new_n17657_), .A3(new_n17658_), .ZN(new_n17659_));
  NAND2_X1   g16632(.A1(new_n17539_), .A2(new_n17525_), .ZN(new_n17660_));
  NAND2_X1   g16633(.A1(new_n17495_), .A2(new_n17503_), .ZN(new_n17661_));
  NOR3_X1    g16634(.A1(new_n17661_), .A2(new_n17494_), .A3(new_n17502_), .ZN(new_n17662_));
  AND3_X2    g16635(.A1(new_n17484_), .A2(new_n17481_), .A3(new_n17662_), .Z(new_n17663_));
  INV_X1     g16636(.I(new_n17663_), .ZN(new_n17664_));
  NOR3_X1    g16637(.A1(new_n17664_), .A2(new_n17651_), .A3(new_n17652_), .ZN(new_n17665_));
  OAI21_X1   g16638(.A1(new_n17650_), .A2(new_n17665_), .B(new_n17490_), .ZN(new_n17666_));
  INV_X1     g16639(.I(new_n17458_), .ZN(new_n17667_));
  INV_X1     g16640(.I(new_n17467_), .ZN(new_n17668_));
  NAND4_X1   g16641(.A1(new_n17667_), .A2(new_n17457_), .A3(new_n17466_), .A4(new_n17668_), .ZN(new_n17669_));
  OR3_X2     g16642(.A1(new_n17446_), .A2(new_n17447_), .A3(new_n17669_), .Z(new_n17670_));
  NAND2_X1   g16643(.A1(new_n17469_), .A2(new_n17460_), .ZN(new_n17671_));
  NOR2_X1    g16644(.A1(new_n17670_), .A2(new_n17671_), .ZN(new_n17672_));
  OAI21_X1   g16645(.A1(new_n17648_), .A2(new_n17672_), .B(new_n17450_), .ZN(new_n17673_));
  NOR2_X1    g16646(.A1(new_n17666_), .A2(new_n17673_), .ZN(new_n17674_));
  XOR2_X1    g16647(.A1(new_n17660_), .A2(new_n17674_), .Z(new_n17675_));
  XOR2_X1    g16648(.A1(new_n17675_), .A2(new_n17659_), .Z(new_n17676_));
  NOR3_X1    g16649(.A1(new_n17647_), .A2(new_n17643_), .A3(new_n17676_), .ZN(new_n17677_));
  NAND2_X1   g16650(.A1(new_n17594_), .A2(new_n17529_), .ZN(new_n17678_));
  NAND2_X1   g16651(.A1(new_n17547_), .A2(new_n17556_), .ZN(new_n17679_));
  NAND2_X1   g16652(.A1(new_n17533_), .A2(new_n17435_), .ZN(new_n17680_));
  NAND2_X1   g16653(.A1(new_n17680_), .A2(new_n17679_), .ZN(new_n17681_));
  OAI21_X1   g16654(.A1(new_n17594_), .A2(new_n17529_), .B(new_n17681_), .ZN(new_n17682_));
  INV_X1     g16655(.I(new_n17659_), .ZN(new_n17683_));
  XOR2_X1    g16656(.A1(new_n17675_), .A2(new_n17683_), .Z(new_n17684_));
  AOI21_X1   g16657(.A1(new_n17682_), .A2(new_n17678_), .B(new_n17684_), .ZN(new_n17685_));
  OAI21_X1   g16658(.A1(new_n17685_), .A2(new_n17677_), .B(new_n17642_), .ZN(new_n17686_));
  INV_X1     g16659(.I(new_n17642_), .ZN(new_n17687_));
  NAND3_X1   g16660(.A1(new_n17682_), .A2(new_n17678_), .A3(new_n17684_), .ZN(new_n17688_));
  OAI21_X1   g16661(.A1(new_n17647_), .A2(new_n17643_), .B(new_n17676_), .ZN(new_n17689_));
  NAND3_X1   g16662(.A1(new_n17688_), .A2(new_n17689_), .A3(new_n17687_), .ZN(new_n17690_));
  AOI21_X1   g16663(.A1(new_n17686_), .A2(new_n17690_), .B(new_n17608_), .ZN(new_n17691_));
  INV_X1     g16664(.I(new_n17608_), .ZN(new_n17692_));
  AOI21_X1   g16665(.A1(new_n17688_), .A2(new_n17689_), .B(new_n17687_), .ZN(new_n17693_));
  NOR3_X1    g16666(.A1(new_n17685_), .A2(new_n17677_), .A3(new_n17642_), .ZN(new_n17694_));
  NOR3_X1    g16667(.A1(new_n17693_), .A2(new_n17694_), .A3(new_n17692_), .ZN(new_n17695_));
  OAI21_X1   g16668(.A1(new_n17695_), .A2(new_n17691_), .B(new_n17603_), .ZN(new_n17696_));
  NOR2_X1    g16669(.A1(new_n17596_), .A2(new_n17600_), .ZN(new_n17697_));
  OAI21_X1   g16670(.A1(new_n17693_), .A2(new_n17694_), .B(new_n17692_), .ZN(new_n17698_));
  NAND3_X1   g16671(.A1(new_n17686_), .A2(new_n17690_), .A3(new_n17608_), .ZN(new_n17699_));
  NAND3_X1   g16672(.A1(new_n17698_), .A2(new_n17699_), .A3(new_n17697_), .ZN(new_n17700_));
  AOI21_X1   g16673(.A1(new_n17696_), .A2(new_n17700_), .B(new_n17602_), .ZN(new_n17701_));
  OAI21_X1   g16674(.A1(new_n17263_), .A2(new_n17264_), .B(new_n17262_), .ZN(new_n17702_));
  NAND3_X1   g16675(.A1(new_n17252_), .A2(new_n17257_), .A3(new_n16741_), .ZN(new_n17703_));
  OAI21_X1   g16676(.A1(new_n16737_), .A2(new_n16739_), .B(new_n15854_), .ZN(new_n17704_));
  NAND3_X1   g16677(.A1(new_n16730_), .A2(new_n16726_), .A3(new_n16735_), .ZN(new_n17705_));
  AOI21_X1   g16678(.A1(new_n17704_), .A2(new_n17705_), .B(new_n15849_), .ZN(new_n17706_));
  AOI21_X1   g16679(.A1(new_n16740_), .A2(new_n16731_), .B(new_n17259_), .ZN(new_n17707_));
  NOR2_X1    g16680(.A1(new_n17706_), .A2(new_n17707_), .ZN(new_n17708_));
  AOI22_X1   g16681(.A1(new_n17702_), .A2(new_n17703_), .B1(new_n17708_), .B2(new_n17287_), .ZN(new_n17709_));
  NOR2_X1    g16682(.A1(new_n17599_), .A2(new_n17600_), .ZN(new_n17710_));
  NOR2_X1    g16683(.A1(new_n17596_), .A2(new_n17597_), .ZN(new_n17711_));
  OAI21_X1   g16684(.A1(new_n17710_), .A2(new_n17711_), .B(new_n17709_), .ZN(new_n17712_));
  AOI21_X1   g16685(.A1(new_n17698_), .A2(new_n17699_), .B(new_n17697_), .ZN(new_n17713_));
  NOR3_X1    g16686(.A1(new_n17695_), .A2(new_n17691_), .A3(new_n17603_), .ZN(new_n17714_));
  NOR3_X1    g16687(.A1(new_n17714_), .A2(new_n17713_), .A3(new_n17712_), .ZN(new_n17715_));
  NOR2_X1    g16688(.A1(new_n17710_), .A2(new_n17711_), .ZN(new_n17716_));
  NAND3_X1   g16689(.A1(new_n17702_), .A2(new_n17703_), .A3(new_n17708_), .ZN(new_n17717_));
  OR2_X2     g16690(.A1(new_n17273_), .A2(new_n17274_), .Z(new_n17718_));
  AND3_X2    g16691(.A1(new_n13949_), .A2(new_n13948_), .A3(new_n13950_), .Z(new_n17719_));
  NOR2_X1    g16692(.A1(new_n17719_), .A2(new_n13951_), .ZN(new_n17720_));
  XNOR2_X1   g16693(.A1(new_n17720_), .A2(\A[1000] ), .ZN(new_n17721_));
  NOR2_X1    g16694(.A1(new_n17278_), .A2(new_n17721_), .ZN(new_n17722_));
  NAND2_X1   g16695(.A1(new_n17718_), .A2(new_n17722_), .ZN(new_n17723_));
  INV_X1     g16696(.I(new_n17278_), .ZN(new_n17724_));
  NOR2_X1    g16697(.A1(new_n17724_), .A2(new_n17721_), .ZN(new_n17725_));
  NAND3_X1   g16698(.A1(new_n17723_), .A2(new_n17286_), .A3(new_n17725_), .ZN(new_n17726_));
  NAND2_X1   g16699(.A1(new_n17286_), .A2(new_n17725_), .ZN(new_n17727_));
  NAND3_X1   g16700(.A1(new_n17718_), .A2(new_n17722_), .A3(new_n17727_), .ZN(new_n17728_));
  AOI21_X1   g16701(.A1(new_n17726_), .A2(new_n17728_), .B(new_n17287_), .ZN(new_n17729_));
  NAND2_X1   g16702(.A1(new_n17729_), .A2(new_n17717_), .ZN(new_n17730_));
  OAI21_X1   g16703(.A1(new_n17709_), .A2(new_n17716_), .B(new_n17730_), .ZN(new_n17731_));
  OAI21_X1   g16704(.A1(new_n17715_), .A2(new_n17701_), .B(new_n17731_), .ZN(new_n17732_));
  NOR2_X1    g16705(.A1(new_n17716_), .A2(new_n17709_), .ZN(new_n17733_));
  NAND4_X1   g16706(.A1(new_n17696_), .A2(new_n17700_), .A3(new_n17712_), .A4(new_n17730_), .ZN(new_n17734_));
  NAND2_X1   g16707(.A1(new_n17734_), .A2(new_n17733_), .ZN(new_n17735_));
  AOI21_X1   g16708(.A1(new_n17696_), .A2(new_n17700_), .B(new_n17712_), .ZN(new_n17736_));
  NAND2_X1   g16709(.A1(new_n17698_), .A2(new_n17699_), .ZN(new_n17737_));
  NAND3_X1   g16710(.A1(new_n17682_), .A2(new_n17678_), .A3(new_n17608_), .ZN(new_n17738_));
  OAI21_X1   g16711(.A1(new_n17647_), .A2(new_n17643_), .B(new_n17692_), .ZN(new_n17739_));
  NAND3_X1   g16712(.A1(new_n17738_), .A2(new_n17739_), .A3(new_n17642_), .ZN(new_n17740_));
  NAND2_X1   g16713(.A1(new_n17740_), .A2(new_n17684_), .ZN(new_n17741_));
  XOR2_X1    g16714(.A1(new_n17608_), .A2(new_n17642_), .Z(new_n17742_));
  NAND2_X1   g16715(.A1(new_n17742_), .A2(new_n17684_), .ZN(new_n17743_));
  NOR3_X1    g16716(.A1(new_n17640_), .A2(new_n17638_), .A3(new_n17612_), .ZN(new_n17744_));
  NAND3_X1   g16717(.A1(new_n17609_), .A2(new_n17014_), .A3(new_n17311_), .ZN(new_n17745_));
  INV_X1     g16718(.I(new_n17627_), .ZN(new_n17746_));
  NOR2_X1    g16719(.A1(new_n17431_), .A2(new_n17745_), .ZN(new_n17751_));
  INV_X1     g16720(.I(new_n17751_), .ZN(new_n17752_));
  NOR2_X1    g16721(.A1(new_n17431_), .A2(new_n17745_), .ZN(new_n17753_));
  INV_X1     g16722(.I(new_n17753_), .ZN(new_n17754_));
  NOR3_X1    g16723(.A1(new_n17626_), .A2(new_n17618_), .A3(new_n17395_), .ZN(new_n17755_));
  NAND2_X1   g16724(.A1(new_n17617_), .A2(new_n17755_), .ZN(new_n17756_));
  OAI21_X1   g16725(.A1(new_n17624_), .A2(new_n17756_), .B(new_n17637_), .ZN(new_n17757_));
  NOR2_X1    g16726(.A1(new_n17746_), .A2(new_n17620_), .ZN(new_n17758_));
  INV_X1     g16727(.I(new_n17758_), .ZN(new_n17759_));
  NAND2_X1   g16728(.A1(new_n17757_), .A2(new_n17759_), .ZN(new_n17760_));
  NOR2_X1    g16729(.A1(new_n17754_), .A2(new_n17758_), .ZN(new_n17761_));
  AOI22_X1   g16730(.A1(new_n17761_), .A2(new_n17757_), .B1(new_n17760_), .B2(new_n17754_), .ZN(new_n17762_));
  INV_X1     g16731(.I(new_n17658_), .ZN(new_n17763_));
  NAND4_X1   g16732(.A1(new_n17664_), .A2(new_n17460_), .A3(new_n17469_), .A4(new_n17670_), .ZN(new_n17764_));
  NOR4_X1    g16733(.A1(new_n17657_), .A2(new_n17651_), .A3(new_n17652_), .A4(new_n17764_), .ZN(new_n17765_));
  NAND4_X1   g16734(.A1(new_n17765_), .A2(new_n17763_), .A3(new_n17666_), .A4(new_n17673_), .ZN(new_n17766_));
  AOI21_X1   g16735(.A1(new_n17660_), .A2(new_n17766_), .B(new_n17683_), .ZN(new_n17767_));
  INV_X1     g16736(.I(new_n17767_), .ZN(new_n17768_));
  NOR2_X1    g16737(.A1(new_n17762_), .A2(new_n17768_), .ZN(new_n17769_));
  NAND2_X1   g16738(.A1(new_n17769_), .A2(new_n17752_), .ZN(new_n17770_));
  OAI21_X1   g16739(.A1(new_n17762_), .A2(new_n17768_), .B(new_n17751_), .ZN(new_n17771_));
  NAND2_X1   g16740(.A1(new_n17770_), .A2(new_n17771_), .ZN(new_n17772_));
  NAND2_X1   g16741(.A1(new_n17772_), .A2(new_n17744_), .ZN(new_n17773_));
  INV_X1     g16742(.I(new_n17773_), .ZN(new_n17774_));
  OAI21_X1   g16743(.A1(new_n17741_), .A2(new_n17743_), .B(new_n17774_), .ZN(new_n17775_));
  NAND4_X1   g16744(.A1(new_n17740_), .A2(new_n17684_), .A3(new_n17742_), .A4(new_n17773_), .ZN(new_n17776_));
  AOI22_X1   g16745(.A1(new_n17737_), .A2(new_n17697_), .B1(new_n17775_), .B2(new_n17776_), .ZN(new_n17777_));
  OAI21_X1   g16746(.A1(new_n17695_), .A2(new_n17691_), .B(new_n17697_), .ZN(new_n17778_));
  NAND2_X1   g16747(.A1(new_n17682_), .A2(new_n17678_), .ZN(new_n17779_));
  AOI21_X1   g16748(.A1(new_n17779_), .A2(new_n17692_), .B(new_n17687_), .ZN(new_n17780_));
  AOI21_X1   g16749(.A1(new_n17780_), .A2(new_n17738_), .B(new_n17676_), .ZN(new_n17781_));
  INV_X1     g16750(.I(new_n17743_), .ZN(new_n17782_));
  AOI21_X1   g16751(.A1(new_n17781_), .A2(new_n17782_), .B(new_n17773_), .ZN(new_n17783_));
  INV_X1     g16752(.I(new_n17776_), .ZN(new_n17784_));
  NOR3_X1    g16753(.A1(new_n17778_), .A2(new_n17783_), .A3(new_n17784_), .ZN(new_n17785_));
  NOR3_X1    g16754(.A1(new_n17736_), .A2(new_n17785_), .A3(new_n17777_), .ZN(new_n17786_));
  NOR3_X1    g16755(.A1(new_n17786_), .A2(new_n17732_), .A3(new_n17735_), .ZN(new_n17787_));
  OAI21_X1   g16756(.A1(new_n17777_), .A2(new_n17785_), .B(new_n17736_), .ZN(new_n17788_));
  AOI21_X1   g16757(.A1(new_n17698_), .A2(new_n17699_), .B(new_n17603_), .ZN(new_n17789_));
  NAND2_X1   g16758(.A1(new_n17775_), .A2(new_n17776_), .ZN(new_n17790_));
  NOR2_X1    g16759(.A1(new_n17744_), .A2(new_n17751_), .ZN(new_n17791_));
  NAND2_X1   g16760(.A1(new_n17791_), .A2(new_n17753_), .ZN(new_n17792_));
  NOR2_X1    g16761(.A1(new_n17757_), .A2(new_n17759_), .ZN(new_n17793_));
  OAI21_X1   g16762(.A1(new_n17791_), .A2(new_n17753_), .B(new_n17793_), .ZN(new_n17794_));
  NAND2_X1   g16763(.A1(new_n17794_), .A2(new_n17792_), .ZN(new_n17795_));
  INV_X1     g16764(.I(new_n17795_), .ZN(new_n17796_));
  OAI21_X1   g16765(.A1(new_n17781_), .A2(new_n17782_), .B(new_n17774_), .ZN(new_n17797_));
  NAND3_X1   g16766(.A1(new_n17741_), .A2(new_n17743_), .A3(new_n17773_), .ZN(new_n17798_));
  NAND2_X1   g16767(.A1(new_n17797_), .A2(new_n17798_), .ZN(new_n17799_));
  INV_X1     g16768(.I(new_n17799_), .ZN(new_n17800_));
  NAND3_X1   g16769(.A1(new_n17800_), .A2(new_n17789_), .A3(new_n17790_), .ZN(new_n17801_));
  NAND2_X1   g16770(.A1(new_n17790_), .A2(new_n17789_), .ZN(new_n17802_));
  NAND2_X1   g16771(.A1(new_n17802_), .A2(new_n17799_), .ZN(new_n17803_));
  AOI21_X1   g16772(.A1(new_n17801_), .A2(new_n17803_), .B(new_n17788_), .ZN(new_n17804_));
  AOI21_X1   g16773(.A1(new_n17735_), .A2(new_n17786_), .B(new_n17732_), .ZN(new_n17805_));
  OAI21_X1   g16774(.A1(new_n17787_), .A2(new_n17804_), .B(new_n17805_), .ZN(new_n17806_));
  NOR2_X1    g16775(.A1(new_n17714_), .A2(new_n17713_), .ZN(new_n17807_));
  OAI22_X1   g16776(.A1(new_n17777_), .A2(new_n17785_), .B1(new_n17807_), .B2(new_n17712_), .ZN(new_n17808_));
  NAND2_X1   g16777(.A1(new_n17790_), .A2(new_n17778_), .ZN(new_n17809_));
  NOR2_X1    g16778(.A1(new_n17783_), .A2(new_n17784_), .ZN(new_n17810_));
  NAND2_X1   g16779(.A1(new_n17810_), .A2(new_n17789_), .ZN(new_n17811_));
  NAND3_X1   g16780(.A1(new_n17811_), .A2(new_n17809_), .A3(new_n17736_), .ZN(new_n17812_));
  NAND2_X1   g16781(.A1(new_n17808_), .A2(new_n17812_), .ZN(new_n17813_));
  NAND2_X1   g16782(.A1(new_n17802_), .A2(new_n17800_), .ZN(new_n17814_));
  NOR2_X1    g16783(.A1(new_n17781_), .A2(new_n17782_), .ZN(new_n17815_));
  NAND2_X1   g16784(.A1(new_n17815_), .A2(new_n17773_), .ZN(new_n17816_));
  NOR2_X1    g16785(.A1(new_n17816_), .A2(new_n17796_), .ZN(new_n17817_));
  AOI21_X1   g16786(.A1(new_n17815_), .A2(new_n17773_), .B(new_n17795_), .ZN(new_n17818_));
  NAND4_X1   g16787(.A1(new_n17697_), .A2(new_n17782_), .A3(new_n17774_), .A4(new_n17795_), .ZN(new_n17819_));
  NOR3_X1    g16788(.A1(new_n17819_), .A2(new_n17815_), .A3(new_n17741_), .ZN(new_n17820_));
  NAND4_X1   g16789(.A1(new_n17820_), .A2(new_n17737_), .A3(new_n17773_), .A4(new_n17815_), .ZN(new_n17821_));
  NOR4_X1    g16790(.A1(new_n17821_), .A2(new_n17802_), .A3(new_n17800_), .A4(new_n17818_), .ZN(new_n17822_));
  NAND4_X1   g16791(.A1(new_n17813_), .A2(new_n17814_), .A3(new_n17817_), .A4(new_n17822_), .ZN(new_n17823_));
  NOR4_X1    g16792(.A1(new_n17802_), .A2(new_n17800_), .A3(new_n17796_), .A4(new_n17816_), .ZN(new_n17824_));
  NAND2_X1   g16793(.A1(new_n17804_), .A2(new_n17824_), .ZN(new_n17825_));
  AOI21_X1   g16794(.A1(new_n17806_), .A2(new_n17823_), .B(new_n17825_), .ZN(maj));
endmodule


