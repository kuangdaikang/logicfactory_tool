// Benchmark "apex6" written by ABC on Fri Feb 25 15:13:02 2022

module apex6 ( 
    PSRW, VFIN, PFIN, INFIN, VYBB0, VYBB1, VZZZE, PYBB0, PYBB1, PYBB2,
    PYBB3, PYBB4, PYBB5, PYBB6, PYBB7, PYBB8, PZZZE, INYBB0, INYBB1,
    INYBB2, INYBB3, INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, INZZZE, MMERR,
    ESRSUM, CBT0, CBT1, CBT2, SLAD0, SLAD1, SLAD2, SLAD3, PSYNC, RPTEN,
    ICLR, STW_N, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3, P1ZZZ4, P1ZZZ5, P1ZZZ6,
    P1ZZZ7, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3, P2ZZZ4, P2ZZZ5, P2ZZZ6, P2ZZZ7,
    I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3, I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, I2ZZZ0,
    I2ZZZ1, I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, I2ZZZ7, TXMESS_N, RYZ,
    COMPPAR, RPTWIN, XZFR0, XZFR1, XZFS, RXZ0, RXZ1, OFS2, OFS1, A, B, C,
    QPR0, QPR1, QPR2, QPR3, QPR4, AXZ0, AXZ1, V1ZZZ0, V1ZZZ1, V1ZZZ2,
    V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3,
    V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, TXWRD0, TXWRD1, TXWRD2, TXWRD3, TXWRD4,
    TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, TXWRD10, TXWRD11, TXWRD12,
    TXWRD13, TXWRD14, TXWRD15, XZ320, XZ321, XZ322, XZ323, XZ324, XZ160_N,
    XZ161, XZ162, XZ163, ENWIN,
    SBUFF, STW_F, TD_P, FSESR_P, P1ZZZ0_P, P1ZZZ1_P, P1ZZZ2_P, P1ZZZ3_P,
    P1ZZZ4_P, P1ZZZ5_P, P1ZZZ6_P, P1ZZZ7_P, P2ZZZ0_P, P2ZZZ1_P, P2ZZZ2_P,
    P2ZZZ3_P, P2ZZZ4_P, P2ZZZ5_P, P2ZZZ6_P, P2ZZZ7_P, I1ZZZ0_P, I1ZZZ1_P,
    I1ZZZ2_P, I1ZZZ3_P, I1ZZZ4_P, I1ZZZ5_P, I1ZZZ6_P, I1ZZZ7_P, I2ZZZ0_P,
    I2ZZZ1_P, I2ZZZ2_P, I2ZZZ3_P, I2ZZZ4_P, I2ZZZ5_P, I2ZZZ6_P, I2ZZZ7_P,
    TXMESS_F, RYZ_P, COMPPAR_P, RPTWIN_P, XZFR0_P, XZFR1_P, XZFS_P, RXZ0_P,
    RXZ1_P, OFS2_P, OFS1_P, A_P, B_P, C_P, QPR0_P, QPR1_P, QPR2_P, QPR3_P,
    QPR4_P, AXZ0_P, AXZ1_P, V1ZZZ0_P, V1ZZZ1_P, V1ZZZ2_P, V1ZZZ3_P,
    V1ZZZ4_P, V1ZZZ5_P, V1ZZZ6_P, V1ZZZ7_P, V2ZZZ0_P, V2ZZZ1_P, V2ZZZ2_P,
    V2ZZZ3_P, V2ZZZ4_P, V2ZZZ5_P, V2ZZZ6_P, V2ZZZ7_P, TXWRD0_P, TXWRD1_P,
    TXWRD2_P, TXWRD3_P, TXWRD4_P, TXWRD5_P, TXWRD6_P, TXWRD7_P, TXWRD8_P,
    TXWRD9_P, TXWRD10_P, TXWRD11_P, TXWRD12_P, TXWRD13_P, TXWRD14_P,
    TXWRD15_P, XZ320_P, XZ321_P, XZ322_P, XZ323_P, XZ324_P, XZ160_F,
    XZ161_P, XZ162_P, XZ163_P, ENWIN_P  );
  input  PSRW, VFIN, PFIN, INFIN, VYBB0, VYBB1, VZZZE, PYBB0, PYBB1,
    PYBB2, PYBB3, PYBB4, PYBB5, PYBB6, PYBB7, PYBB8, PZZZE, INYBB0, INYBB1,
    INYBB2, INYBB3, INYBB4, INYBB5, INYBB6, INYBB7, INYBB8, INZZZE, MMERR,
    ESRSUM, CBT0, CBT1, CBT2, SLAD0, SLAD1, SLAD2, SLAD3, PSYNC, RPTEN,
    ICLR, STW_N, P1ZZZ0, P1ZZZ1, P1ZZZ2, P1ZZZ3, P1ZZZ4, P1ZZZ5, P1ZZZ6,
    P1ZZZ7, P2ZZZ0, P2ZZZ1, P2ZZZ2, P2ZZZ3, P2ZZZ4, P2ZZZ5, P2ZZZ6, P2ZZZ7,
    I1ZZZ0, I1ZZZ1, I1ZZZ2, I1ZZZ3, I1ZZZ4, I1ZZZ5, I1ZZZ6, I1ZZZ7, I2ZZZ0,
    I2ZZZ1, I2ZZZ2, I2ZZZ3, I2ZZZ4, I2ZZZ5, I2ZZZ6, I2ZZZ7, TXMESS_N, RYZ,
    COMPPAR, RPTWIN, XZFR0, XZFR1, XZFS, RXZ0, RXZ1, OFS2, OFS1, A, B, C,
    QPR0, QPR1, QPR2, QPR3, QPR4, AXZ0, AXZ1, V1ZZZ0, V1ZZZ1, V1ZZZ2,
    V1ZZZ3, V1ZZZ4, V1ZZZ5, V1ZZZ6, V1ZZZ7, V2ZZZ0, V2ZZZ1, V2ZZZ2, V2ZZZ3,
    V2ZZZ4, V2ZZZ5, V2ZZZ6, V2ZZZ7, TXWRD0, TXWRD1, TXWRD2, TXWRD3, TXWRD4,
    TXWRD5, TXWRD6, TXWRD7, TXWRD8, TXWRD9, TXWRD10, TXWRD11, TXWRD12,
    TXWRD13, TXWRD14, TXWRD15, XZ320, XZ321, XZ322, XZ323, XZ324, XZ160_N,
    XZ161, XZ162, XZ163, ENWIN;
  output SBUFF, STW_F, TD_P, FSESR_P, P1ZZZ0_P, P1ZZZ1_P, P1ZZZ2_P, P1ZZZ3_P,
    P1ZZZ4_P, P1ZZZ5_P, P1ZZZ6_P, P1ZZZ7_P, P2ZZZ0_P, P2ZZZ1_P, P2ZZZ2_P,
    P2ZZZ3_P, P2ZZZ4_P, P2ZZZ5_P, P2ZZZ6_P, P2ZZZ7_P, I1ZZZ0_P, I1ZZZ1_P,
    I1ZZZ2_P, I1ZZZ3_P, I1ZZZ4_P, I1ZZZ5_P, I1ZZZ6_P, I1ZZZ7_P, I2ZZZ0_P,
    I2ZZZ1_P, I2ZZZ2_P, I2ZZZ3_P, I2ZZZ4_P, I2ZZZ5_P, I2ZZZ6_P, I2ZZZ7_P,
    TXMESS_F, RYZ_P, COMPPAR_P, RPTWIN_P, XZFR0_P, XZFR1_P, XZFS_P, RXZ0_P,
    RXZ1_P, OFS2_P, OFS1_P, A_P, B_P, C_P, QPR0_P, QPR1_P, QPR2_P, QPR3_P,
    QPR4_P, AXZ0_P, AXZ1_P, V1ZZZ0_P, V1ZZZ1_P, V1ZZZ2_P, V1ZZZ3_P,
    V1ZZZ4_P, V1ZZZ5_P, V1ZZZ6_P, V1ZZZ7_P, V2ZZZ0_P, V2ZZZ1_P, V2ZZZ2_P,
    V2ZZZ3_P, V2ZZZ4_P, V2ZZZ5_P, V2ZZZ6_P, V2ZZZ7_P, TXWRD0_P, TXWRD1_P,
    TXWRD2_P, TXWRD3_P, TXWRD4_P, TXWRD5_P, TXWRD6_P, TXWRD7_P, TXWRD8_P,
    TXWRD9_P, TXWRD10_P, TXWRD11_P, TXWRD12_P, TXWRD13_P, TXWRD14_P,
    TXWRD15_P, XZ320_P, XZ321_P, XZ322_P, XZ323_P, XZ324_P, XZ160_F,
    XZ161_P, XZ162_P, XZ163_P, ENWIN_P;
  wire new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_,
    new_n242_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n288_, new_n289_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n297_, new_n298_, new_n300_, new_n301_,
    new_n303_, new_n304_, new_n306_, new_n307_, new_n309_, new_n310_,
    new_n312_, new_n313_, new_n315_, new_n316_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n324_, new_n325_, new_n327_,
    new_n328_, new_n330_, new_n331_, new_n333_, new_n334_, new_n336_,
    new_n337_, new_n339_, new_n340_, new_n342_, new_n343_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n351_, new_n352_,
    new_n354_, new_n355_, new_n357_, new_n358_, new_n360_, new_n361_,
    new_n363_, new_n364_, new_n366_, new_n367_, new_n369_, new_n370_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n378_,
    new_n379_, new_n381_, new_n382_, new_n384_, new_n385_, new_n387_,
    new_n388_, new_n390_, new_n391_, new_n393_, new_n394_, new_n396_,
    new_n397_, new_n399_, new_n400_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_;
  assign SBUFF = ~TXMESS_N | RPTWIN;
  assign new_n236_ = ~PFIN & ~INFIN;
  assign new_n237_ = ~TXMESS_N & AXZ0;
  assign new_n238_ = AXZ1 & new_n237_;
  assign new_n239_ = A & new_n238_;
  assign new_n240_ = ~STW_N & ~new_n239_;
  assign new_n241_ = new_n236_ & ~new_n240_;
  assign new_n242_ = ~VFIN & new_n241_;
  assign STW_F = RYZ | new_n242_;
  assign new_n244_ = SLAD2 & QPR0;
  assign new_n245_ = SLAD3 & ~QPR0;
  assign new_n246_ = ~new_n244_ & ~new_n245_;
  assign new_n247_ = SLAD1 & ~QPR0;
  assign new_n248_ = SLAD0 & QPR0;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = QPR2 & ~new_n249_;
  assign new_n251_ = ~QPR1 & new_n250_;
  assign new_n252_ = ~QPR2 & ~new_n246_;
  assign new_n253_ = QPR1 & new_n252_;
  assign new_n254_ = ~new_n251_ & ~new_n253_;
  assign new_n255_ = ESRSUM & ~AXZ0;
  assign new_n256_ = ~COMPPAR & AXZ0;
  assign new_n257_ = ~new_n255_ & ~new_n256_;
  assign new_n258_ = AXZ1 & ~new_n257_;
  assign new_n259_ = AXZ0 & ~AXZ1;
  assign new_n260_ = ~MMERR & new_n259_;
  assign new_n261_ = ~new_n258_ & ~new_n260_;
  assign new_n262_ = ~B & ~C;
  assign new_n263_ = ~AXZ0 & ~AXZ1;
  assign new_n264_ = A & ~new_n263_;
  assign new_n265_ = A & ~new_n261_;
  assign new_n266_ = TXWRD0 & ~new_n264_;
  assign new_n267_ = ~new_n262_ & new_n266_;
  assign new_n268_ = ~new_n265_ & ~new_n267_;
  assign new_n269_ = new_n262_ & ~new_n264_;
  assign new_n270_ = ~RPTWIN & new_n269_;
  assign new_n271_ = SBUFF & ~new_n270_;
  assign new_n272_ = RXZ0 & ~RXZ1;
  assign new_n273_ = ~ESRSUM & new_n272_;
  assign new_n274_ = ~RXZ0 & RXZ1;
  assign new_n275_ = ESRSUM & new_n274_;
  assign new_n276_ = ~new_n273_ & ~new_n275_;
  assign new_n277_ = RPTEN & ~new_n276_;
  assign new_n278_ = RPTWIN & new_n277_;
  assign new_n279_ = ~TXMESS_N & ~new_n268_;
  assign new_n280_ = ~RPTWIN & new_n279_;
  assign new_n281_ = ~QPR3 & ~new_n254_;
  assign new_n282_ = ~QPR4 & ~new_n271_;
  assign new_n283_ = new_n281_ & new_n282_;
  assign new_n284_ = ~new_n280_ & ~new_n283_;
  assign new_n285_ = ~new_n278_ & new_n284_;
  assign TD_P = ~RYZ & ~new_n285_;
  assign OFS2_P = ~ICLR & OFS1;
  assign new_n288_ = OFS2 & OFS2_P;
  assign new_n289_ = ~ICLR & XZFR1;
  assign FSESR_P = new_n288_ | new_n289_;
  assign new_n291_ = PYBB0 & ~PZZZE;
  assign new_n292_ = ~RYZ & ~new_n291_;
  assign new_n293_ = ~RYZ & new_n291_;
  assign new_n294_ = P1ZZZ0 & new_n292_;
  assign new_n295_ = PYBB1 & new_n293_;
  assign P1ZZZ0_P = new_n294_ | new_n295_;
  assign new_n297_ = P1ZZZ1 & new_n292_;
  assign new_n298_ = PYBB2 & new_n293_;
  assign P1ZZZ1_P = new_n297_ | new_n298_;
  assign new_n300_ = P1ZZZ2 & new_n292_;
  assign new_n301_ = PYBB3 & new_n293_;
  assign P1ZZZ2_P = new_n300_ | new_n301_;
  assign new_n303_ = P1ZZZ3 & new_n292_;
  assign new_n304_ = PYBB4 & new_n293_;
  assign P1ZZZ3_P = new_n303_ | new_n304_;
  assign new_n306_ = P1ZZZ4 & new_n292_;
  assign new_n307_ = PYBB5 & new_n293_;
  assign P1ZZZ4_P = new_n306_ | new_n307_;
  assign new_n309_ = P1ZZZ5 & new_n292_;
  assign new_n310_ = PYBB6 & new_n293_;
  assign P1ZZZ5_P = new_n309_ | new_n310_;
  assign new_n312_ = P1ZZZ6 & new_n292_;
  assign new_n313_ = PYBB7 & new_n293_;
  assign P1ZZZ6_P = new_n312_ | new_n313_;
  assign new_n315_ = P1ZZZ7 & new_n292_;
  assign new_n316_ = PYBB8 & new_n293_;
  assign P1ZZZ7_P = new_n315_ | new_n316_;
  assign new_n318_ = PYBB0 & PZZZE;
  assign new_n319_ = ~RYZ & ~new_n318_;
  assign new_n320_ = ~RYZ & new_n318_;
  assign new_n321_ = P2ZZZ0 & new_n319_;
  assign new_n322_ = PYBB1 & new_n320_;
  assign P2ZZZ0_P = new_n321_ | new_n322_;
  assign new_n324_ = P2ZZZ1 & new_n319_;
  assign new_n325_ = PYBB2 & new_n320_;
  assign P2ZZZ1_P = new_n324_ | new_n325_;
  assign new_n327_ = P2ZZZ2 & new_n319_;
  assign new_n328_ = PYBB3 & new_n320_;
  assign P2ZZZ2_P = new_n327_ | new_n328_;
  assign new_n330_ = P2ZZZ3 & new_n319_;
  assign new_n331_ = PYBB4 & new_n320_;
  assign P2ZZZ3_P = new_n330_ | new_n331_;
  assign new_n333_ = P2ZZZ4 & new_n319_;
  assign new_n334_ = PYBB5 & new_n320_;
  assign P2ZZZ4_P = new_n333_ | new_n334_;
  assign new_n336_ = P2ZZZ5 & new_n319_;
  assign new_n337_ = PYBB6 & new_n320_;
  assign P2ZZZ5_P = new_n336_ | new_n337_;
  assign new_n339_ = P2ZZZ6 & new_n319_;
  assign new_n340_ = PYBB7 & new_n320_;
  assign P2ZZZ6_P = new_n339_ | new_n340_;
  assign new_n342_ = P2ZZZ7 & new_n319_;
  assign new_n343_ = PYBB8 & new_n320_;
  assign P2ZZZ7_P = new_n342_ | new_n343_;
  assign new_n345_ = INYBB0 & ~INZZZE;
  assign new_n346_ = ~RYZ & ~new_n345_;
  assign new_n347_ = ~RYZ & new_n345_;
  assign new_n348_ = I1ZZZ0 & new_n346_;
  assign new_n349_ = INYBB1 & new_n347_;
  assign I1ZZZ0_P = new_n348_ | new_n349_;
  assign new_n351_ = I1ZZZ1 & new_n346_;
  assign new_n352_ = INYBB2 & new_n347_;
  assign I1ZZZ1_P = new_n351_ | new_n352_;
  assign new_n354_ = I1ZZZ2 & new_n346_;
  assign new_n355_ = INYBB3 & new_n347_;
  assign I1ZZZ2_P = new_n354_ | new_n355_;
  assign new_n357_ = I1ZZZ3 & new_n346_;
  assign new_n358_ = INYBB4 & new_n347_;
  assign I1ZZZ3_P = new_n357_ | new_n358_;
  assign new_n360_ = I1ZZZ4 & new_n346_;
  assign new_n361_ = INYBB5 & new_n347_;
  assign I1ZZZ4_P = new_n360_ | new_n361_;
  assign new_n363_ = I1ZZZ5 & new_n346_;
  assign new_n364_ = INYBB6 & new_n347_;
  assign I1ZZZ5_P = new_n363_ | new_n364_;
  assign new_n366_ = I1ZZZ6 & new_n346_;
  assign new_n367_ = INYBB7 & new_n347_;
  assign I1ZZZ6_P = new_n366_ | new_n367_;
  assign new_n369_ = I1ZZZ7 & new_n346_;
  assign new_n370_ = INYBB8 & new_n347_;
  assign I1ZZZ7_P = new_n369_ | new_n370_;
  assign new_n372_ = INYBB0 & INZZZE;
  assign new_n373_ = ~RYZ & ~new_n372_;
  assign new_n374_ = ~RYZ & new_n372_;
  assign new_n375_ = I2ZZZ0 & new_n373_;
  assign new_n376_ = INYBB1 & new_n374_;
  assign I2ZZZ0_P = new_n375_ | new_n376_;
  assign new_n378_ = I2ZZZ1 & new_n373_;
  assign new_n379_ = INYBB2 & new_n374_;
  assign I2ZZZ1_P = new_n378_ | new_n379_;
  assign new_n381_ = I2ZZZ2 & new_n373_;
  assign new_n382_ = INYBB3 & new_n374_;
  assign I2ZZZ2_P = new_n381_ | new_n382_;
  assign new_n384_ = I2ZZZ3 & new_n373_;
  assign new_n385_ = INYBB4 & new_n374_;
  assign I2ZZZ3_P = new_n384_ | new_n385_;
  assign new_n387_ = I2ZZZ4 & new_n373_;
  assign new_n388_ = INYBB5 & new_n374_;
  assign I2ZZZ4_P = new_n387_ | new_n388_;
  assign new_n390_ = I2ZZZ5 & new_n373_;
  assign new_n391_ = INYBB6 & new_n374_;
  assign I2ZZZ5_P = new_n390_ | new_n391_;
  assign new_n393_ = I2ZZZ6 & new_n373_;
  assign new_n394_ = INYBB7 & new_n374_;
  assign I2ZZZ6_P = new_n393_ | new_n394_;
  assign new_n396_ = I2ZZZ7 & new_n373_;
  assign new_n397_ = INYBB8 & new_n374_;
  assign I2ZZZ7_P = new_n396_ | new_n397_;
  assign new_n399_ = ~VFIN & TXMESS_N;
  assign new_n400_ = new_n236_ & new_n399_;
  assign TXMESS_F = RYZ | new_n400_;
  assign RYZ_P = ICLR | new_n239_;
  assign new_n403_ = TXWRD0 & ~new_n262_;
  assign new_n404_ = ~QPR4 & ~new_n254_;
  assign new_n405_ = ~QPR3 & new_n262_;
  assign new_n406_ = new_n404_ & new_n405_;
  assign new_n407_ = ~new_n403_ & ~new_n406_;
  assign new_n408_ = ESRSUM & AXZ1;
  assign new_n409_ = ~MMERR & AXZ0;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = ~ESRSUM & AXZ1;
  assign new_n412_ = MMERR & AXZ0;
  assign new_n413_ = ~new_n411_ & ~new_n412_;
  assign new_n414_ = COMPPAR & ~new_n413_;
  assign new_n415_ = ~TXMESS_N & ~COMPPAR;
  assign new_n416_ = ~new_n410_ & new_n415_;
  assign new_n417_ = ~new_n414_ & ~new_n416_;
  assign new_n418_ = ~new_n238_ & new_n417_;
  assign new_n419_ = ~new_n264_ & new_n407_;
  assign new_n420_ = ~TXMESS_N & ~new_n419_;
  assign new_n421_ = COMPPAR & ~new_n420_;
  assign new_n422_ = A & ~new_n418_;
  assign new_n423_ = ~new_n264_ & ~new_n407_;
  assign new_n424_ = new_n415_ & new_n423_;
  assign new_n425_ = ~new_n422_ & ~new_n424_;
  assign new_n426_ = ~new_n421_ & new_n425_;
  assign COMPPAR_P = ~RYZ & ~new_n426_;
  assign new_n428_ = RXZ0 & RXZ1;
  assign new_n429_ = PSYNC & XZFS;
  assign new_n430_ = ~SLAD2 & ~SLAD3;
  assign new_n431_ = new_n429_ & new_n430_;
  assign new_n432_ = XZ321 & XZ322;
  assign new_n433_ = XZ320 & XZ323;
  assign new_n434_ = new_n432_ & new_n433_;
  assign new_n435_ = ~SLAD3 & ~XZ163;
  assign new_n436_ = SLAD3 & XZ163;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = ~SLAD2 & ~XZ162;
  assign new_n439_ = SLAD2 & XZ162;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~new_n437_ & ~new_n440_;
  assign new_n442_ = ~SLAD1 & ~XZ161;
  assign new_n443_ = SLAD1 & XZ161;
  assign new_n444_ = ~new_n442_ & ~new_n443_;
  assign new_n445_ = ~SLAD0 & XZ160_N;
  assign new_n446_ = SLAD0 & ~XZ160_N;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = XZ324 & ENWIN;
  assign new_n449_ = new_n434_ & new_n448_;
  assign new_n450_ = new_n441_ & new_n449_;
  assign new_n451_ = ~new_n444_ & new_n450_;
  assign new_n452_ = ~new_n447_ & new_n451_;
  assign new_n453_ = RPTWIN & ~new_n428_;
  assign new_n454_ = ~SLAD1 & new_n431_;
  assign new_n455_ = ~SLAD0 & new_n454_;
  assign new_n456_ = ~new_n453_ & ~new_n455_;
  assign new_n457_ = ~new_n452_ & new_n456_;
  assign RPTWIN_P = ~RYZ & ~new_n457_;
  assign new_n459_ = XZ323 & XZ324;
  assign new_n460_ = new_n432_ & new_n459_;
  assign new_n461_ = ~XZ163 & new_n460_;
  assign new_n462_ = XZ160_N & ~XZ161;
  assign new_n463_ = ~XZ162 & new_n462_;
  assign new_n464_ = new_n461_ & new_n463_;
  assign new_n465_ = ~PSYNC & ~ICLR;
  assign XZ320_P = ~XZ320 & new_n465_;
  assign new_n467_ = ~new_n464_ & new_n465_;
  assign new_n468_ = ~XZ320_P & ~new_n467_;
  assign new_n469_ = XZ320 & new_n465_;
  assign new_n470_ = XZFR0 & ~new_n468_;
  assign new_n471_ = new_n464_ & new_n469_;
  assign new_n472_ = ~XZFR0 & new_n471_;
  assign XZFR0_P = new_n470_ | new_n472_;
  assign new_n474_ = ~XZFR0 & new_n465_;
  assign new_n475_ = new_n468_ & ~new_n474_;
  assign new_n476_ = XZFR1 & ~new_n475_;
  assign new_n477_ = XZFR0 & ~XZFR1;
  assign new_n478_ = new_n471_ & new_n477_;
  assign XZFR1_P = new_n476_ | new_n478_;
  assign OFS1_P = PSYNC & ~ICLR;
  assign new_n481_ = ~ICLR & XZFS;
  assign new_n482_ = ~OFS1_P & ~new_n481_;
  assign new_n483_ = OFS2 & OFS1;
  assign new_n484_ = PSRW & ~new_n482_;
  assign XZFS_P = ~new_n483_ & new_n484_;
  assign new_n486_ = ~RPTWIN & ~new_n452_;
  assign new_n487_ = ~ICLR & ~new_n486_;
  assign new_n488_ = ~SLAD0 & XZFS;
  assign new_n489_ = OFS1_P & new_n488_;
  assign new_n490_ = ~SLAD1 & new_n430_;
  assign new_n491_ = new_n489_ & new_n490_;
  assign new_n492_ = ~new_n487_ & ~new_n491_;
  assign new_n493_ = ~SLAD2 & XZ162;
  assign new_n494_ = XZ163 & ~new_n493_;
  assign new_n495_ = XZ320 & new_n494_;
  assign new_n496_ = ~SLAD3 & XZ163;
  assign new_n497_ = XZ162 & ~new_n496_;
  assign new_n498_ = XZ320 & new_n497_;
  assign new_n499_ = ~SLAD0 & ~XZ160_N;
  assign new_n500_ = new_n460_ & ~new_n499_;
  assign new_n501_ = ~new_n493_ & ~new_n496_;
  assign new_n502_ = XZ320 & new_n501_;
  assign new_n503_ = XZ161 & ENWIN;
  assign new_n504_ = new_n500_ & new_n502_;
  assign new_n505_ = new_n503_ & new_n504_;
  assign new_n506_ = ~SLAD1 & XZ161;
  assign new_n507_ = ENWIN & ~new_n506_;
  assign new_n508_ = new_n500_ & new_n507_;
  assign new_n509_ = ~XZ160_N & new_n460_;
  assign new_n510_ = new_n507_ & new_n509_;
  assign new_n511_ = new_n502_ & new_n510_;
  assign new_n512_ = ~XZFS & ~new_n502_;
  assign new_n513_ = SLAD0 & ~new_n511_;
  assign new_n514_ = ~new_n431_ & ~new_n508_;
  assign new_n515_ = ~new_n513_ & ~new_n514_;
  assign new_n516_ = ~new_n512_ & new_n515_;
  assign new_n517_ = ~PSYNC & ~new_n501_;
  assign new_n518_ = SLAD3 & ~new_n495_;
  assign new_n519_ = ~new_n517_ & ~new_n518_;
  assign new_n520_ = SLAD2 & ~new_n498_;
  assign new_n521_ = SLAD1 & ~new_n505_;
  assign new_n522_ = ~new_n520_ & ~new_n521_;
  assign new_n523_ = new_n519_ & new_n522_;
  assign new_n524_ = new_n516_ & new_n523_;
  assign new_n525_ = ~ICLR & ~new_n524_;
  assign new_n526_ = ~XZ320_P & ~new_n525_;
  assign new_n527_ = ~RXZ0 & ~new_n492_;
  assign new_n528_ = RXZ0 & ~new_n526_;
  assign new_n529_ = ~RPTWIN & new_n528_;
  assign RXZ0_P = new_n527_ | new_n529_;
  assign new_n531_ = ~ICLR & ~RXZ0;
  assign new_n532_ = ~RPTWIN & ~new_n526_;
  assign new_n533_ = ~new_n531_ & ~new_n532_;
  assign new_n534_ = RXZ1 & ~new_n533_;
  assign new_n535_ = ~RXZ1 & ~new_n492_;
  assign new_n536_ = RXZ0 & new_n535_;
  assign RXZ1_P = new_n534_ | new_n536_;
  assign new_n538_ = QPR0 & ~QPR1;
  assign new_n539_ = QPR2 & new_n538_;
  assign new_n540_ = CBT2 & ~QPR4;
  assign new_n541_ = B & ~QPR4;
  assign new_n542_ = ~QPR3 & ~new_n540_;
  assign new_n543_ = QPR3 & new_n541_;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = new_n539_ & ~new_n544_;
  assign new_n546_ = ~TXMESS_N & new_n545_;
  assign new_n547_ = ~A & ~new_n546_;
  assign A_P = ~RYZ & ~new_n547_;
  assign new_n549_ = ~CBT0 & ~CBT1;
  assign new_n550_ = CBT2 & ~new_n549_;
  assign new_n551_ = ~QPR4 & new_n539_;
  assign new_n552_ = ~QPR3 & ~new_n550_;
  assign new_n553_ = ~TXMESS_N & ~new_n552_;
  assign new_n554_ = new_n551_ & new_n553_;
  assign new_n555_ = B & ~new_n554_;
  assign new_n556_ = ~B & new_n539_;
  assign new_n557_ = new_n550_ & new_n556_;
  assign new_n558_ = ~TXMESS_N & ~QPR4;
  assign new_n559_ = ~QPR3 & new_n558_;
  assign new_n560_ = new_n557_ & new_n559_;
  assign new_n561_ = ~new_n555_ & ~new_n560_;
  assign B_P = ~RYZ & ~new_n561_;
  assign new_n563_ = CBT2 & new_n549_;
  assign new_n564_ = ~TXMESS_N & ~QPR3;
  assign new_n565_ = ~QPR4 & ~new_n563_;
  assign new_n566_ = new_n539_ & ~new_n565_;
  assign new_n567_ = new_n564_ & new_n566_;
  assign new_n568_ = ~C & new_n567_;
  assign new_n569_ = C & ~new_n567_;
  assign new_n570_ = ~new_n568_ & ~new_n569_;
  assign C_P = ~RYZ & ~new_n570_;
  assign new_n572_ = QPR0 & new_n400_;
  assign new_n573_ = ~RYZ & new_n572_;
  assign new_n574_ = ~QPR0 & ~TXMESS_F;
  assign QPR0_P = new_n573_ | new_n574_;
  assign new_n576_ = QPR0 & ~new_n400_;
  assign new_n577_ = ~RYZ & ~new_n576_;
  assign new_n578_ = QPR1 & new_n577_;
  assign new_n579_ = ~QPR1 & ~TXMESS_F;
  assign new_n580_ = QPR0 & new_n579_;
  assign QPR1_P = new_n578_ | new_n580_;
  assign new_n582_ = QPR1 & new_n576_;
  assign new_n583_ = QPR0 & QPR1;
  assign new_n584_ = ~TXMESS_F & new_n583_;
  assign new_n585_ = ~QPR2 & new_n584_;
  assign new_n586_ = ~RYZ & ~new_n582_;
  assign new_n587_ = QPR2 & new_n586_;
  assign QPR2_P = new_n585_ | new_n587_;
  assign new_n589_ = QPR2 & new_n582_;
  assign new_n590_ = ~QPR3 & new_n584_;
  assign new_n591_ = QPR2 & new_n590_;
  assign new_n592_ = ~RYZ & ~new_n589_;
  assign new_n593_ = QPR3 & new_n592_;
  assign QPR3_P = new_n591_ | new_n593_;
  assign new_n595_ = QPR3 & new_n589_;
  assign new_n596_ = ~RYZ & QPR4;
  assign new_n597_ = ~new_n595_ & new_n596_;
  assign new_n598_ = QPR2 & QPR3;
  assign new_n599_ = ~QPR4 & new_n584_;
  assign new_n600_ = new_n598_ & new_n599_;
  assign QPR4_P = new_n597_ | new_n600_;
  assign new_n602_ = ~A & ~new_n545_;
  assign new_n603_ = ~TXMESS_N & ~new_n602_;
  assign new_n604_ = ~AXZ0 & new_n603_;
  assign new_n605_ = AXZ0 & ~new_n603_;
  assign new_n606_ = ~new_n604_ & ~new_n605_;
  assign AXZ0_P = ~RYZ & ~new_n606_;
  assign new_n608_ = AXZ0 & new_n603_;
  assign new_n609_ = AXZ1 & ~new_n608_;
  assign new_n610_ = new_n259_ & new_n603_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign AXZ1_P = ~RYZ & ~new_n611_;
  assign new_n613_ = VYBB0 & ~VZZZE;
  assign new_n614_ = ~RYZ & ~new_n613_;
  assign new_n615_ = ~RYZ & new_n613_;
  assign new_n616_ = V1ZZZ1 & new_n615_;
  assign new_n617_ = V1ZZZ0 & new_n614_;
  assign V1ZZZ0_P = new_n616_ | new_n617_;
  assign new_n619_ = V1ZZZ2 & new_n615_;
  assign new_n620_ = V1ZZZ1 & new_n614_;
  assign V1ZZZ1_P = new_n619_ | new_n620_;
  assign new_n622_ = V1ZZZ3 & new_n615_;
  assign new_n623_ = V1ZZZ2 & new_n614_;
  assign V1ZZZ2_P = new_n622_ | new_n623_;
  assign new_n625_ = V1ZZZ4 & new_n615_;
  assign new_n626_ = V1ZZZ3 & new_n614_;
  assign V1ZZZ3_P = new_n625_ | new_n626_;
  assign new_n628_ = V1ZZZ5 & new_n615_;
  assign new_n629_ = V1ZZZ4 & new_n614_;
  assign V1ZZZ4_P = new_n628_ | new_n629_;
  assign new_n631_ = V1ZZZ6 & new_n615_;
  assign new_n632_ = V1ZZZ5 & new_n614_;
  assign V1ZZZ5_P = new_n631_ | new_n632_;
  assign new_n634_ = V1ZZZ7 & new_n615_;
  assign new_n635_ = V1ZZZ6 & new_n614_;
  assign V1ZZZ6_P = new_n634_ | new_n635_;
  assign new_n637_ = V1ZZZ7 & new_n614_;
  assign new_n638_ = VYBB1 & new_n615_;
  assign V1ZZZ7_P = new_n637_ | new_n638_;
  assign new_n640_ = VYBB0 & VZZZE;
  assign new_n641_ = ~RYZ & ~new_n640_;
  assign new_n642_ = ~RYZ & new_n640_;
  assign new_n643_ = V2ZZZ1 & new_n642_;
  assign new_n644_ = V2ZZZ0 & new_n641_;
  assign V2ZZZ0_P = new_n643_ | new_n644_;
  assign new_n646_ = V2ZZZ2 & new_n642_;
  assign new_n647_ = V2ZZZ1 & new_n641_;
  assign V2ZZZ1_P = new_n646_ | new_n647_;
  assign new_n649_ = V2ZZZ3 & new_n642_;
  assign new_n650_ = V2ZZZ2 & new_n641_;
  assign V2ZZZ2_P = new_n649_ | new_n650_;
  assign new_n652_ = V2ZZZ4 & new_n642_;
  assign new_n653_ = V2ZZZ3 & new_n641_;
  assign V2ZZZ3_P = new_n652_ | new_n653_;
  assign new_n655_ = V2ZZZ5 & new_n642_;
  assign new_n656_ = V2ZZZ4 & new_n641_;
  assign V2ZZZ4_P = new_n655_ | new_n656_;
  assign new_n658_ = V2ZZZ6 & new_n642_;
  assign new_n659_ = V2ZZZ5 & new_n641_;
  assign V2ZZZ5_P = new_n658_ | new_n659_;
  assign new_n661_ = V2ZZZ7 & new_n642_;
  assign new_n662_ = V2ZZZ6 & new_n641_;
  assign V2ZZZ6_P = new_n661_ | new_n662_;
  assign new_n664_ = V2ZZZ7 & new_n641_;
  assign new_n665_ = VYBB1 & new_n642_;
  assign V2ZZZ7_P = new_n664_ | new_n665_;
  assign new_n667_ = PFIN & ~INFIN;
  assign new_n668_ = ~TXMESS_N & ~new_n262_;
  assign new_n669_ = ~VFIN & ~new_n668_;
  assign new_n670_ = ~VFIN & new_n668_;
  assign new_n671_ = TXWRD1 & new_n670_;
  assign new_n672_ = VFIN & V1ZZZ0;
  assign new_n673_ = TXWRD0 & new_n669_;
  assign new_n674_ = ~new_n672_ & ~new_n673_;
  assign new_n675_ = ~new_n671_ & new_n674_;
  assign new_n676_ = P1ZZZ0 & new_n667_;
  assign new_n677_ = INFIN & I1ZZZ0;
  assign new_n678_ = new_n236_ & ~new_n675_;
  assign new_n679_ = ~new_n677_ & ~new_n678_;
  assign new_n680_ = ~new_n676_ & new_n679_;
  assign TXWRD0_P = ~RYZ & ~new_n680_;
  assign new_n682_ = ~INFIN & ~RYZ;
  assign new_n683_ = INFIN & ~RYZ;
  assign new_n684_ = ~PFIN & new_n669_;
  assign new_n685_ = ~PFIN & new_n670_;
  assign new_n686_ = VFIN & ~PFIN;
  assign new_n687_ = V1ZZZ1 & new_n686_;
  assign new_n688_ = TXWRD2 & new_n685_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = PFIN & P1ZZZ1;
  assign new_n691_ = TXWRD1 & new_n684_;
  assign new_n692_ = ~new_n690_ & ~new_n691_;
  assign new_n693_ = new_n689_ & new_n692_;
  assign new_n694_ = I1ZZZ1 & new_n683_;
  assign new_n695_ = new_n682_ & ~new_n693_;
  assign TXWRD1_P = new_n694_ | new_n695_;
  assign new_n697_ = V1ZZZ2 & new_n686_;
  assign new_n698_ = TXWRD3 & new_n685_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign new_n700_ = PFIN & P1ZZZ2;
  assign new_n701_ = TXWRD2 & new_n684_;
  assign new_n702_ = ~new_n700_ & ~new_n701_;
  assign new_n703_ = new_n699_ & new_n702_;
  assign new_n704_ = I1ZZZ2 & new_n683_;
  assign new_n705_ = new_n682_ & ~new_n703_;
  assign TXWRD2_P = new_n704_ | new_n705_;
  assign new_n707_ = PFIN & new_n682_;
  assign new_n708_ = TXWRD4 & new_n670_;
  assign new_n709_ = VFIN & V1ZZZ3;
  assign new_n710_ = TXWRD3 & new_n669_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = ~new_n708_ & new_n711_;
  assign new_n713_ = ~PFIN & new_n682_;
  assign new_n714_ = ~new_n712_ & new_n713_;
  assign new_n715_ = I1ZZZ3 & new_n683_;
  assign new_n716_ = P1ZZZ3 & new_n707_;
  assign new_n717_ = ~new_n715_ & ~new_n716_;
  assign TXWRD3_P = new_n714_ | ~new_n717_;
  assign new_n719_ = TXWRD5 & new_n670_;
  assign new_n720_ = VFIN & V1ZZZ4;
  assign new_n721_ = TXWRD4 & new_n669_;
  assign new_n722_ = ~new_n720_ & ~new_n721_;
  assign new_n723_ = ~new_n719_ & new_n722_;
  assign new_n724_ = new_n713_ & ~new_n723_;
  assign new_n725_ = I1ZZZ4 & new_n683_;
  assign new_n726_ = P1ZZZ4 & new_n707_;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign TXWRD4_P = new_n724_ | ~new_n727_;
  assign new_n729_ = TXWRD6 & new_n670_;
  assign new_n730_ = VFIN & V1ZZZ5;
  assign new_n731_ = TXWRD5 & new_n669_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = ~new_n729_ & new_n732_;
  assign new_n734_ = new_n713_ & ~new_n733_;
  assign new_n735_ = I1ZZZ5 & new_n683_;
  assign new_n736_ = P1ZZZ5 & new_n707_;
  assign new_n737_ = ~new_n735_ & ~new_n736_;
  assign TXWRD5_P = new_n734_ | ~new_n737_;
  assign new_n739_ = TXWRD7 & new_n670_;
  assign new_n740_ = VFIN & V1ZZZ6;
  assign new_n741_ = TXWRD6 & new_n669_;
  assign new_n742_ = ~new_n740_ & ~new_n741_;
  assign new_n743_ = ~new_n739_ & new_n742_;
  assign new_n744_ = new_n713_ & ~new_n743_;
  assign new_n745_ = I1ZZZ6 & new_n683_;
  assign new_n746_ = P1ZZZ6 & new_n707_;
  assign new_n747_ = ~new_n745_ & ~new_n746_;
  assign TXWRD6_P = new_n744_ | ~new_n747_;
  assign new_n749_ = TXWRD8 & new_n670_;
  assign new_n750_ = VFIN & V1ZZZ7;
  assign new_n751_ = TXWRD7 & new_n669_;
  assign new_n752_ = ~new_n750_ & ~new_n751_;
  assign new_n753_ = ~new_n749_ & new_n752_;
  assign new_n754_ = P1ZZZ7 & new_n667_;
  assign new_n755_ = new_n236_ & ~new_n753_;
  assign new_n756_ = INFIN & I1ZZZ7;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign new_n758_ = ~new_n754_ & new_n757_;
  assign TXWRD7_P = ~RYZ & ~new_n758_;
  assign new_n760_ = TXWRD9 & new_n670_;
  assign new_n761_ = VFIN & V2ZZZ0;
  assign new_n762_ = TXWRD8 & new_n669_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = ~new_n760_ & new_n763_;
  assign new_n765_ = new_n713_ & ~new_n764_;
  assign new_n766_ = I2ZZZ0 & new_n683_;
  assign new_n767_ = P2ZZZ0 & new_n707_;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign TXWRD8_P = new_n765_ | ~new_n768_;
  assign new_n770_ = V2ZZZ1 & new_n686_;
  assign new_n771_ = TXWRD10 & new_n685_;
  assign new_n772_ = ~new_n770_ & ~new_n771_;
  assign new_n773_ = PFIN & P2ZZZ1;
  assign new_n774_ = TXWRD9 & new_n684_;
  assign new_n775_ = ~new_n773_ & ~new_n774_;
  assign new_n776_ = new_n772_ & new_n775_;
  assign new_n777_ = I2ZZZ1 & new_n683_;
  assign new_n778_ = new_n682_ & ~new_n776_;
  assign TXWRD9_P = new_n777_ | new_n778_;
  assign new_n780_ = TXWRD11 & new_n670_;
  assign new_n781_ = VFIN & V2ZZZ2;
  assign new_n782_ = TXWRD10 & new_n669_;
  assign new_n783_ = ~new_n781_ & ~new_n782_;
  assign new_n784_ = ~new_n780_ & new_n783_;
  assign new_n785_ = INFIN & I2ZZZ2;
  assign new_n786_ = P2ZZZ2 & new_n667_;
  assign new_n787_ = new_n236_ & ~new_n784_;
  assign new_n788_ = ~new_n786_ & ~new_n787_;
  assign new_n789_ = ~new_n785_ & new_n788_;
  assign TXWRD10_P = ~RYZ & ~new_n789_;
  assign new_n791_ = TXWRD12 & new_n670_;
  assign new_n792_ = VFIN & V2ZZZ3;
  assign new_n793_ = TXWRD11 & new_n669_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = ~new_n791_ & new_n794_;
  assign new_n796_ = INFIN & I2ZZZ3;
  assign new_n797_ = P2ZZZ3 & new_n667_;
  assign new_n798_ = new_n236_ & ~new_n795_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = ~new_n796_ & new_n799_;
  assign TXWRD11_P = ~RYZ & ~new_n800_;
  assign new_n802_ = TXWRD13 & new_n670_;
  assign new_n803_ = VFIN & V2ZZZ4;
  assign new_n804_ = TXWRD12 & new_n669_;
  assign new_n805_ = ~new_n803_ & ~new_n804_;
  assign new_n806_ = ~new_n802_ & new_n805_;
  assign new_n807_ = INFIN & I2ZZZ4;
  assign new_n808_ = P2ZZZ4 & new_n667_;
  assign new_n809_ = new_n236_ & ~new_n806_;
  assign new_n810_ = ~new_n808_ & ~new_n809_;
  assign new_n811_ = ~new_n807_ & new_n810_;
  assign TXWRD12_P = ~RYZ & ~new_n811_;
  assign new_n813_ = TXWRD14 & new_n670_;
  assign new_n814_ = VFIN & V2ZZZ5;
  assign new_n815_ = TXWRD13 & new_n669_;
  assign new_n816_ = ~new_n814_ & ~new_n815_;
  assign new_n817_ = ~new_n813_ & new_n816_;
  assign new_n818_ = new_n713_ & ~new_n817_;
  assign new_n819_ = P2ZZZ5 & new_n707_;
  assign new_n820_ = I2ZZZ5 & new_n683_;
  assign new_n821_ = ~new_n819_ & ~new_n820_;
  assign TXWRD13_P = new_n818_ | ~new_n821_;
  assign new_n823_ = TXWRD15 & new_n670_;
  assign new_n824_ = VFIN & V2ZZZ6;
  assign new_n825_ = TXWRD14 & new_n669_;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = ~new_n823_ & new_n826_;
  assign new_n828_ = I2ZZZ6 & new_n683_;
  assign new_n829_ = P2ZZZ6 & new_n707_;
  assign new_n830_ = ~new_n828_ & ~new_n829_;
  assign new_n831_ = new_n713_ & ~new_n827_;
  assign TXWRD14_P = ~new_n830_ | new_n831_;
  assign new_n833_ = V2ZZZ7 & new_n686_;
  assign new_n834_ = PFIN & P2ZZZ7;
  assign new_n835_ = TXWRD15 & new_n684_;
  assign new_n836_ = ~new_n834_ & ~new_n835_;
  assign new_n837_ = ~new_n833_ & new_n836_;
  assign new_n838_ = I2ZZZ7 & new_n683_;
  assign new_n839_ = new_n682_ & ~new_n837_;
  assign TXWRD15_P = new_n838_ | new_n839_;
  assign new_n841_ = ~XZ321 & new_n469_;
  assign new_n842_ = XZ321 & XZ320_P;
  assign XZ321_P = new_n841_ | new_n842_;
  assign new_n844_ = ~XZ321 & new_n465_;
  assign new_n845_ = ~XZ320_P & ~new_n844_;
  assign new_n846_ = XZ322 & ~new_n845_;
  assign new_n847_ = ~XZ322 & new_n469_;
  assign new_n848_ = XZ321 & new_n847_;
  assign XZ322_P = new_n846_ | new_n848_;
  assign new_n850_ = ~XZ322 & new_n465_;
  assign new_n851_ = new_n845_ & ~new_n850_;
  assign new_n852_ = new_n432_ & new_n469_;
  assign new_n853_ = ~XZ323 & new_n852_;
  assign new_n854_ = XZ323 & ~new_n851_;
  assign XZ323_P = new_n853_ | new_n854_;
  assign new_n856_ = XZ322 & XZ323;
  assign new_n857_ = new_n465_ & ~new_n856_;
  assign new_n858_ = new_n845_ & ~new_n857_;
  assign new_n859_ = new_n434_ & new_n465_;
  assign new_n860_ = ~XZ324 & new_n859_;
  assign new_n861_ = XZ324 & ~new_n858_;
  assign XZ324_P = new_n860_ | new_n861_;
  assign new_n863_ = ~new_n460_ & new_n465_;
  assign new_n864_ = ~XZ320_P & ~new_n863_;
  assign new_n865_ = XZ160_N & ~new_n864_;
  assign new_n866_ = new_n469_ & new_n509_;
  assign XZ160_F = new_n865_ | new_n866_;
  assign new_n868_ = new_n465_ & ~new_n509_;
  assign new_n869_ = ~XZ320_P & ~new_n868_;
  assign new_n870_ = XZ161 & ~new_n869_;
  assign new_n871_ = ~XZ161 & new_n866_;
  assign XZ161_P = new_n870_ | new_n871_;
  assign new_n873_ = XZ320 & XZ161;
  assign new_n874_ = new_n509_ & new_n873_;
  assign new_n875_ = ~XZ161 & new_n465_;
  assign new_n876_ = new_n869_ & ~new_n875_;
  assign new_n877_ = XZ162 & ~new_n876_;
  assign new_n878_ = ~XZ162 & new_n465_;
  assign new_n879_ = new_n874_ & new_n878_;
  assign XZ162_P = new_n877_ | new_n879_;
  assign new_n881_ = XZ161 & XZ162;
  assign new_n882_ = new_n465_ & ~new_n881_;
  assign new_n883_ = new_n869_ & ~new_n882_;
  assign new_n884_ = XZ163 & ~new_n883_;
  assign new_n885_ = XZ162 & new_n874_;
  assign new_n886_ = ~XZ163 & new_n465_;
  assign new_n887_ = new_n885_ & new_n886_;
  assign XZ163_P = new_n884_ | new_n887_;
  assign new_n889_ = XZFS & OFS1_P;
  assign new_n890_ = ~ICLR & ENWIN;
  assign new_n891_ = ~new_n889_ & ~new_n890_;
  assign new_n892_ = PSRW & ~new_n891_;
  assign ENWIN_P = ~new_n483_ & new_n892_;
endmodule


