// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:33 2022

module t1  ( 
    v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15,
    v16, v17, v18, v19, v20,
    \v21.0 , \v21.1 , \v21.2 , \v21.3 , \v21.4 , \v21.5 , \v21.6 , \v21.7 ,
    \v21.8 , \v21.9 , \v21.10 , \v21.11 , \v21.12 , \v21.13 , \v21.14 ,
    \v21.15 , \v21.16 , \v21.17 , \v21.18 , \v21.19 , \v21.20 , \v21.21 ,
    \v21.22   );
  input  v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14,
    v15, v16, v17, v18, v19, v20;
  output \v21.0 , \v21.1 , \v21.2 , \v21.3 , \v21.4 , \v21.5 , \v21.6 ,
    \v21.7 , \v21.8 , \v21.9 , \v21.10 , \v21.11 , \v21.12 , \v21.13 ,
    \v21.14 , \v21.15 , \v21.16 , \v21.17 , \v21.18 , \v21.19 , \v21.20 ,
    \v21.21 , \v21.22 ;
  wire new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n133_,
    new_n134_, new_n135_, new_n136_, new_n137_, new_n138_, new_n139_,
    new_n140_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n240_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n357_, new_n358_, new_n359_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n366_, new_n367_,
    new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_;
  assign new_n45_ = v6 & ~v15;
  assign new_n46_ = v3 & new_n45_;
  assign new_n47_ = ~v15 & ~new_n46_;
  assign new_n48_ = v20 & ~new_n47_;
  assign new_n49_ = v15 & ~v20;
  assign new_n50_ = ~new_n48_ & ~new_n49_;
  assign new_n51_ = v19 & ~new_n50_;
  assign new_n52_ = v15 & ~v19;
  assign new_n53_ = ~new_n51_ & ~new_n52_;
  assign new_n54_ = ~v17 & ~new_n53_;
  assign new_n55_ = v15 & v17;
  assign new_n56_ = ~new_n54_ & ~new_n55_;
  assign new_n57_ = ~v4 & ~new_n56_;
  assign new_n58_ = v4 & v15;
  assign new_n59_ = ~new_n57_ & ~new_n58_;
  assign new_n60_ = v18 & ~new_n59_;
  assign new_n61_ = ~v17 & v19;
  assign new_n62_ = ~v17 & ~new_n61_;
  assign new_n63_ = ~v17 & ~v19;
  assign new_n64_ = new_n62_ & ~new_n63_;
  assign new_n65_ = ~v18 & ~new_n64_;
  assign new_n66_ = v15 & new_n65_;
  assign new_n67_ = ~new_n60_ & ~new_n66_;
  assign new_n68_ = ~v16 & ~new_n67_;
  assign new_n69_ = ~v4 & ~v18;
  assign new_n70_ = ~v4 & ~new_n69_;
  assign new_n71_ = v18 & ~v19;
  assign new_n72_ = ~v4 & new_n71_;
  assign new_n73_ = new_n70_ & ~new_n72_;
  assign new_n74_ = ~v4 & v18;
  assign new_n75_ = v19 & ~v20;
  assign new_n76_ = new_n74_ & new_n75_;
  assign new_n77_ = new_n73_ & ~new_n76_;
  assign new_n78_ = v16 & ~new_n77_;
  assign new_n79_ = v15 & new_n78_;
  assign new_n80_ = ~new_n68_ & ~new_n79_;
  assign \v21.0  = ~v0 & ~new_n80_;
  assign new_n82_ = v6 & ~v7;
  assign new_n83_ = v6 & ~new_n82_;
  assign new_n84_ = v20 & ~new_n83_;
  assign new_n85_ = ~v16 & new_n84_;
  assign new_n86_ = v3 & new_n85_;
  assign new_n87_ = v16 & ~v20;
  assign new_n88_ = ~new_n86_ & ~new_n87_;
  assign new_n89_ = v19 & ~new_n88_;
  assign new_n90_ = v16 & ~v19;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = v18 & ~new_n91_;
  assign new_n93_ = v16 & ~v18;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ~v15 & ~new_n94_;
  assign new_n96_ = ~v16 & v20;
  assign new_n97_ = ~new_n87_ & ~new_n96_;
  assign new_n98_ = v19 & ~new_n97_;
  assign new_n99_ = ~new_n90_ & ~new_n98_;
  assign new_n100_ = v18 & ~new_n99_;
  assign new_n101_ = ~new_n93_ & ~new_n100_;
  assign new_n102_ = v15 & ~new_n101_;
  assign new_n103_ = ~new_n95_ & ~new_n102_;
  assign new_n104_ = ~v4 & ~new_n103_;
  assign new_n105_ = v4 & v16;
  assign new_n106_ = ~new_n104_ & ~new_n105_;
  assign new_n107_ = ~v17 & ~new_n106_;
  assign new_n108_ = v17 & ~new_n77_;
  assign new_n109_ = v16 & new_n108_;
  assign new_n110_ = ~new_n107_ & ~new_n109_;
  assign \v21.1  = ~v0 & ~new_n110_;
  assign new_n112_ = v3 & v6;
  assign new_n113_ = v3 & ~new_n112_;
  assign new_n114_ = v20 & ~new_n113_;
  assign new_n115_ = ~v17 & new_n114_;
  assign new_n116_ = v17 & ~v20;
  assign new_n117_ = ~new_n115_ & ~new_n116_;
  assign new_n118_ = v19 & ~new_n117_;
  assign new_n119_ = v17 & ~v19;
  assign new_n120_ = ~new_n118_ & ~new_n119_;
  assign new_n121_ = v18 & ~new_n120_;
  assign new_n122_ = v17 & ~v18;
  assign new_n123_ = ~new_n121_ & ~new_n122_;
  assign new_n124_ = ~v4 & ~new_n123_;
  assign new_n125_ = v4 & v17;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign new_n127_ = ~v16 & ~new_n126_;
  assign new_n128_ = ~new_n109_ & ~new_n127_;
  assign new_n129_ = ~v15 & ~new_n128_;
  assign new_n130_ = v15 & new_n108_;
  assign new_n131_ = ~new_n129_ & ~new_n130_;
  assign \v21.2  = ~v0 & ~new_n131_;
  assign new_n133_ = ~v4 & ~v19;
  assign new_n134_ = ~v4 & ~new_n133_;
  assign new_n135_ = ~v4 & new_n75_;
  assign new_n136_ = new_n134_ & ~new_n135_;
  assign new_n137_ = v18 & ~new_n136_;
  assign new_n138_ = v19 & v20;
  assign new_n139_ = new_n69_ & new_n138_;
  assign new_n140_ = ~new_n137_ & ~new_n139_;
  assign \v21.3  = ~v0 & ~new_n140_;
  assign new_n142_ = ~v4 & ~v20;
  assign new_n143_ = ~v4 & ~new_n142_;
  assign new_n144_ = v19 & ~new_n143_;
  assign new_n145_ = ~v19 & v20;
  assign new_n146_ = ~v4 & new_n145_;
  assign new_n147_ = ~new_n144_ & ~new_n146_;
  assign \v21.4  = ~v0 & ~new_n147_;
  assign new_n149_ = v4 & v20;
  assign new_n150_ = ~v4 & new_n87_;
  assign new_n151_ = ~new_n149_ & ~new_n150_;
  assign new_n152_ = ~v4 & ~v16;
  assign new_n153_ = new_n116_ & new_n152_;
  assign new_n154_ = new_n151_ & ~new_n153_;
  assign new_n155_ = v18 & ~v20;
  assign new_n156_ = ~v17 & new_n155_;
  assign new_n157_ = new_n152_ & new_n156_;
  assign new_n158_ = new_n154_ & ~new_n157_;
  assign new_n159_ = ~v4 & v19;
  assign new_n160_ = v19 & ~new_n159_;
  assign new_n161_ = ~v20 & ~new_n160_;
  assign new_n162_ = ~v18 & new_n161_;
  assign new_n163_ = ~v17 & new_n162_;
  assign new_n164_ = ~v16 & new_n163_;
  assign new_n165_ = new_n158_ & ~new_n164_;
  assign \v21.5  = ~v0 & ~new_n165_;
  assign new_n167_ = v2 & ~v15;
  assign new_n168_ = ~v1 & new_n167_;
  assign new_n169_ = ~v3 & ~new_n168_;
  assign new_n170_ = ~v16 & ~new_n169_;
  assign new_n171_ = ~v1 & v2;
  assign new_n172_ = ~v3 & ~new_n171_;
  assign new_n173_ = v17 & ~new_n172_;
  assign new_n174_ = v16 & new_n173_;
  assign new_n175_ = ~v15 & new_n174_;
  assign new_n176_ = ~new_n170_ & ~new_n175_;
  assign new_n177_ = ~v15 & ~v17;
  assign new_n178_ = ~v15 & ~new_n177_;
  assign new_n179_ = ~v18 & ~new_n178_;
  assign new_n180_ = v16 & new_n179_;
  assign new_n181_ = v3 & new_n180_;
  assign new_n182_ = new_n176_ & ~new_n181_;
  assign new_n183_ = ~v19 & ~new_n178_;
  assign new_n184_ = v18 & new_n183_;
  assign new_n185_ = v16 & new_n184_;
  assign new_n186_ = v3 & new_n185_;
  assign new_n187_ = new_n182_ & ~new_n186_;
  assign new_n188_ = v16 & ~new_n178_;
  assign new_n189_ = v3 & new_n188_;
  assign new_n190_ = v1 & v2;
  assign new_n191_ = ~v16 & ~v17;
  assign new_n192_ = ~v15 & new_n191_;
  assign new_n193_ = new_n190_ & new_n192_;
  assign new_n194_ = ~new_n189_ & ~new_n193_;
  assign new_n195_ = ~v20 & ~new_n194_;
  assign new_n196_ = v19 & new_n195_;
  assign new_n197_ = v18 & new_n196_;
  assign new_n198_ = new_n187_ & ~new_n197_;
  assign \v21.6  = ~v0 & ~new_n198_;
  assign new_n200_ = ~v9 & v16;
  assign new_n201_ = ~v8 & new_n200_;
  assign new_n202_ = v16 & ~new_n201_;
  assign new_n203_ = ~v9 & v13;
  assign new_n204_ = v15 & v16;
  assign new_n205_ = new_n203_ & new_n204_;
  assign new_n206_ = new_n202_ & ~new_n205_;
  assign new_n207_ = ~v18 & ~new_n206_;
  assign new_n208_ = ~v20 & ~new_n206_;
  assign new_n209_ = ~v19 & new_n208_;
  assign new_n210_ = v18 & new_n209_;
  assign new_n211_ = ~new_n207_ & ~new_n210_;
  assign new_n212_ = ~v17 & ~new_n211_;
  assign new_n213_ = v13 & v16;
  assign new_n214_ = v8 & ~new_n213_;
  assign new_n215_ = ~v19 & ~v20;
  assign new_n216_ = v18 & new_n215_;
  assign new_n217_ = v18 & ~new_n216_;
  assign new_n218_ = ~new_n214_ & ~new_n217_;
  assign new_n219_ = v17 & new_n218_;
  assign new_n220_ = v15 & new_n219_;
  assign new_n221_ = ~v9 & new_n220_;
  assign \v21.7  = new_n212_ | new_n221_;
  assign new_n223_ = v9 & v16;
  assign new_n224_ = ~v8 & new_n223_;
  assign new_n225_ = v16 & ~new_n224_;
  assign new_n226_ = ~new_n205_ & new_n225_;
  assign new_n227_ = ~v18 & ~new_n226_;
  assign new_n228_ = ~v20 & ~new_n226_;
  assign new_n229_ = ~v19 & new_n228_;
  assign new_n230_ = v18 & new_n229_;
  assign new_n231_ = ~new_n227_ & ~new_n230_;
  assign new_n232_ = ~v17 & ~new_n231_;
  assign new_n233_ = ~v8 & v9;
  assign new_n234_ = ~v9 & new_n213_;
  assign new_n235_ = ~new_n233_ & ~new_n234_;
  assign new_n236_ = ~new_n217_ & ~new_n235_;
  assign new_n237_ = v17 & new_n236_;
  assign new_n238_ = v15 & new_n237_;
  assign \v21.8  = new_n232_ | new_n238_;
  assign new_n240_ = v8 & new_n200_;
  assign new_n241_ = v16 & ~new_n240_;
  assign new_n242_ = ~new_n205_ & new_n241_;
  assign new_n243_ = ~v18 & ~new_n242_;
  assign new_n244_ = ~v20 & ~new_n242_;
  assign new_n245_ = ~v19 & new_n244_;
  assign new_n246_ = v18 & new_n245_;
  assign new_n247_ = ~new_n243_ & ~new_n246_;
  assign new_n248_ = ~v17 & ~new_n247_;
  assign new_n249_ = ~v8 & ~new_n213_;
  assign new_n250_ = ~new_n217_ & ~new_n249_;
  assign new_n251_ = v17 & new_n250_;
  assign new_n252_ = v15 & new_n251_;
  assign new_n253_ = ~v9 & new_n252_;
  assign \v21.9  = new_n248_ | new_n253_;
  assign new_n255_ = v8 & new_n223_;
  assign new_n256_ = v16 & ~new_n255_;
  assign new_n257_ = ~new_n205_ & new_n256_;
  assign new_n258_ = ~v18 & ~new_n257_;
  assign new_n259_ = ~v20 & ~new_n257_;
  assign new_n260_ = ~v19 & new_n259_;
  assign new_n261_ = v18 & new_n260_;
  assign new_n262_ = ~new_n258_ & ~new_n261_;
  assign new_n263_ = ~v17 & ~new_n262_;
  assign new_n264_ = v8 & v9;
  assign new_n265_ = ~new_n234_ & ~new_n264_;
  assign new_n266_ = ~new_n217_ & ~new_n265_;
  assign new_n267_ = v17 & new_n266_;
  assign new_n268_ = v15 & new_n267_;
  assign \v21.10  = new_n263_ | new_n268_;
  assign new_n270_ = ~v16 & v17;
  assign new_n271_ = ~v16 & ~new_n270_;
  assign new_n272_ = ~v17 & ~v18;
  assign new_n273_ = ~v16 & new_n272_;
  assign new_n274_ = new_n271_ & ~new_n273_;
  assign new_n275_ = v18 & v19;
  assign new_n276_ = new_n191_ & new_n275_;
  assign new_n277_ = new_n274_ & ~new_n276_;
  assign new_n278_ = new_n191_ & new_n216_;
  assign \v21.11  = ~new_n277_ | new_n278_;
  assign new_n280_ = ~v18 & v19;
  assign new_n281_ = ~v18 & ~new_n280_;
  assign new_n282_ = ~v11 & v16;
  assign new_n283_ = ~v10 & new_n282_;
  assign new_n284_ = v16 & ~new_n283_;
  assign new_n285_ = ~new_n205_ & new_n284_;
  assign new_n286_ = ~new_n281_ & ~new_n285_;
  assign new_n287_ = ~v17 & new_n286_;
  assign new_n288_ = ~v10 & ~v11;
  assign new_n289_ = ~new_n234_ & ~new_n288_;
  assign new_n290_ = ~new_n281_ & ~new_n289_;
  assign new_n291_ = v17 & new_n290_;
  assign new_n292_ = v15 & new_n291_;
  assign \v21.12  = new_n287_ | new_n292_;
  assign new_n294_ = v11 & v16;
  assign new_n295_ = ~v10 & new_n294_;
  assign new_n296_ = v16 & ~new_n295_;
  assign new_n297_ = ~new_n205_ & new_n296_;
  assign new_n298_ = ~new_n281_ & ~new_n297_;
  assign new_n299_ = ~v17 & new_n298_;
  assign new_n300_ = ~v10 & v11;
  assign new_n301_ = ~new_n234_ & ~new_n300_;
  assign new_n302_ = ~new_n281_ & ~new_n301_;
  assign new_n303_ = v17 & new_n302_;
  assign new_n304_ = v15 & new_n303_;
  assign \v21.13  = new_n299_ | new_n304_;
  assign new_n306_ = v10 & new_n282_;
  assign new_n307_ = v16 & ~new_n306_;
  assign new_n308_ = ~new_n205_ & new_n307_;
  assign new_n309_ = ~new_n281_ & ~new_n308_;
  assign new_n310_ = ~v17 & new_n309_;
  assign new_n311_ = v10 & ~v11;
  assign new_n312_ = ~new_n234_ & ~new_n311_;
  assign new_n313_ = ~new_n281_ & ~new_n312_;
  assign new_n314_ = v17 & new_n313_;
  assign new_n315_ = v15 & new_n314_;
  assign \v21.14  = new_n310_ | new_n315_;
  assign new_n317_ = v10 & new_n294_;
  assign new_n318_ = v16 & ~new_n317_;
  assign new_n319_ = ~new_n205_ & new_n318_;
  assign new_n320_ = ~new_n281_ & ~new_n319_;
  assign new_n321_ = ~v17 & new_n320_;
  assign new_n322_ = v10 & v11;
  assign new_n323_ = ~new_n234_ & ~new_n322_;
  assign new_n324_ = ~new_n281_ & ~new_n323_;
  assign new_n325_ = v17 & new_n324_;
  assign new_n326_ = v15 & new_n325_;
  assign \v21.15  = new_n321_ | new_n326_;
  assign new_n328_ = ~v5 & ~v17;
  assign new_n329_ = ~v12 & new_n55_;
  assign new_n330_ = ~new_n328_ & ~new_n329_;
  assign new_n331_ = ~v16 & ~new_n330_;
  assign new_n332_ = v16 & ~v17;
  assign new_n333_ = ~v12 & ~v15;
  assign new_n334_ = new_n332_ & new_n333_;
  assign new_n335_ = ~new_n331_ & ~new_n334_;
  assign \v21.16  = ~new_n281_ & ~new_n335_;
  assign new_n337_ = v5 & ~v17;
  assign new_n338_ = v12 & new_n55_;
  assign new_n339_ = ~new_n337_ & ~new_n338_;
  assign new_n340_ = ~v16 & ~new_n339_;
  assign new_n341_ = v12 & ~v15;
  assign new_n342_ = new_n332_ & new_n341_;
  assign new_n343_ = ~new_n340_ & ~new_n342_;
  assign \v21.17  = ~new_n281_ & ~new_n343_;
  assign new_n345_ = ~new_n61_ & ~new_n119_;
  assign new_n346_ = ~v16 & v18;
  assign new_n347_ = ~new_n93_ & ~new_n346_;
  assign new_n348_ = ~new_n345_ & ~new_n347_;
  assign new_n349_ = ~new_n71_ & ~new_n280_;
  assign new_n350_ = v16 & ~new_n349_;
  assign new_n351_ = ~v16 & ~v18;
  assign new_n352_ = ~new_n350_ & ~new_n351_;
  assign new_n353_ = v17 & ~new_n352_;
  assign new_n354_ = v16 & new_n63_;
  assign new_n355_ = ~new_n353_ & ~new_n354_;
  assign \v21.18  = new_n348_ | ~new_n355_;
  assign new_n357_ = v15 & new_n270_;
  assign new_n358_ = ~v15 & new_n332_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign \v21.19  = ~new_n349_ & ~new_n359_;
  assign new_n361_ = v18 & ~new_n71_;
  assign new_n362_ = v18 & new_n75_;
  assign new_n363_ = new_n361_ & ~new_n362_;
  assign new_n364_ = v16 & ~new_n363_;
  assign \v21.20  = v15 & new_n364_;
  assign new_n366_ = ~v12 & ~v14;
  assign new_n367_ = ~v14 & ~new_n366_;
  assign new_n368_ = ~new_n349_ & ~new_n367_;
  assign new_n369_ = ~v18 & new_n145_;
  assign new_n370_ = ~new_n362_ & ~new_n369_;
  assign new_n371_ = ~new_n367_ & ~new_n370_;
  assign new_n372_ = ~new_n368_ & ~new_n371_;
  assign new_n373_ = v16 & ~new_n372_;
  assign \v21.21  = v15 & new_n373_;
  assign new_n375_ = v12 & ~v14;
  assign new_n376_ = ~v14 & ~new_n375_;
  assign new_n377_ = ~new_n349_ & ~new_n376_;
  assign new_n378_ = ~new_n370_ & ~new_n376_;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_ = v16 & ~new_n379_;
  assign \v21.22  = v15 & new_n380_;
endmodule


