// Benchmark "source.pla" written by ABC on Fri Feb 25 15:12:45 2022

module ex5  ( 
    v0, v1, v2, v3, v4, v5, v6, v7,
    \v8.0 , \v8.1 , \v8.2 , \v8.3 , \v8.4 , \v8.5 , \v8.6 , \v8.7 , \v8.8 ,
    \v8.9 , \v8.10 , \v8.11 , \v8.12 , \v8.13 , \v8.14 , \v8.15 , \v8.16 ,
    \v8.17 , \v8.18 , \v8.19 , \v8.20 , \v8.21 , \v8.22 , \v8.23 , \v8.24 ,
    \v8.25 , \v8.26 , \v8.27 , \v8.28 , \v8.29 , \v8.30 , \v8.31 , \v8.32 ,
    \v8.33 , \v8.34 , \v8.35 , \v8.36 , \v8.37 , \v8.38 , \v8.39 , \v8.40 ,
    \v8.41 , \v8.42 , \v8.43 , \v8.44 , \v8.45 , \v8.46 , \v8.47 , \v8.48 ,
    \v8.49 , \v8.50 , \v8.51 , \v8.52 , \v8.53 , \v8.54 , \v8.55 , \v8.56 ,
    \v8.57 , \v8.58 , \v8.59 , \v8.60 , \v8.61 , \v8.62   );
  input  v0, v1, v2, v3, v4, v5, v6, v7;
  output \v8.0 , \v8.1 , \v8.2 , \v8.3 , \v8.4 , \v8.5 , \v8.6 , \v8.7 ,
    \v8.8 , \v8.9 , \v8.10 , \v8.11 , \v8.12 , \v8.13 , \v8.14 , \v8.15 ,
    \v8.16 , \v8.17 , \v8.18 , \v8.19 , \v8.20 , \v8.21 , \v8.22 , \v8.23 ,
    \v8.24 , \v8.25 , \v8.26 , \v8.27 , \v8.28 , \v8.29 , \v8.30 , \v8.31 ,
    \v8.32 , \v8.33 , \v8.34 , \v8.35 , \v8.36 , \v8.37 , \v8.38 , \v8.39 ,
    \v8.40 , \v8.41 , \v8.42 , \v8.43 , \v8.44 , \v8.45 , \v8.46 , \v8.47 ,
    \v8.48 , \v8.49 , \v8.50 , \v8.51 , \v8.52 , \v8.53 , \v8.54 , \v8.55 ,
    \v8.56 , \v8.57 , \v8.58 , \v8.59 , \v8.60 , \v8.61 , \v8.62 ;
  wire new_n72_, new_n74_, new_n76_, new_n77_, new_n80_, new_n81_, new_n82_,
    new_n84_, new_n86_, new_n87_, new_n88_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n117_, new_n118_, new_n119_, new_n120_, new_n121_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n152_, new_n153_, new_n154_, new_n156_, new_n157_, new_n158_,
    new_n160_, new_n161_, new_n162_, new_n164_, new_n165_, new_n166_,
    new_n168_, new_n169_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n176_, new_n177_, new_n178_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n186_, new_n187_, new_n189_, new_n190_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n202_, new_n204_, new_n205_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_;
  assign new_n72_ = ~v5 & ~v6;
  assign \v8.0  = ~v4 & new_n72_;
  assign new_n74_ = ~v6 & ~v7;
  assign \v8.1  = ~v5 & new_n74_;
  assign new_n76_ = v5 & new_n74_;
  assign new_n77_ = ~v4 & new_n76_;
  assign \v8.2  = ~v3 & new_n77_;
  assign \v8.3  = v3 & new_n77_;
  assign new_n80_ = v6 & ~v7;
  assign new_n81_ = ~v5 & new_n80_;
  assign new_n82_ = ~v4 & new_n81_;
  assign \v8.4  = v3 & new_n82_;
  assign new_n84_ = v5 & new_n80_;
  assign \v8.5  = ~v4 & new_n84_;
  assign new_n86_ = v3 & \v8.0 ;
  assign new_n87_ = v2 & new_n86_;
  assign new_n88_ = ~v1 & new_n87_;
  assign \v8.6  = ~v0 & new_n88_;
  assign new_n90_ = ~v0 & v1;
  assign new_n91_ = ~v2 & new_n90_;
  assign new_n92_ = ~v3 & new_n91_;
  assign new_n93_ = ~v4 & new_n92_;
  assign new_n94_ = v5 & new_n93_;
  assign new_n95_ = v6 & new_n94_;
  assign \v8.7  = v7 & new_n95_;
  assign new_n97_ = v0 & v1;
  assign new_n98_ = v2 & new_n97_;
  assign new_n99_ = ~v3 & new_n98_;
  assign new_n100_ = ~v4 & new_n99_;
  assign new_n101_ = v5 & new_n100_;
  assign new_n102_ = v6 & new_n101_;
  assign \v8.8  = v7 & new_n102_;
  assign new_n104_ = ~v0 & ~v1;
  assign new_n105_ = v2 & new_n104_;
  assign new_n106_ = ~v3 & new_n105_;
  assign new_n107_ = ~v4 & new_n106_;
  assign new_n108_ = ~v5 & new_n107_;
  assign new_n109_ = v6 & new_n108_;
  assign \v8.9  = v7 & new_n109_;
  assign new_n111_ = v6 & v7;
  assign new_n112_ = v5 & new_n111_;
  assign new_n113_ = ~v4 & new_n112_;
  assign new_n114_ = v2 & new_n113_;
  assign new_n115_ = v1 & new_n114_;
  assign \v8.10  = ~v0 & new_n115_;
  assign new_n117_ = ~v2 & new_n97_;
  assign new_n118_ = ~v3 & new_n117_;
  assign new_n119_ = ~v4 & new_n118_;
  assign new_n120_ = v5 & new_n119_;
  assign new_n121_ = v6 & new_n120_;
  assign \v8.11  = v7 & new_n121_;
  assign new_n123_ = v0 & ~v1;
  assign new_n124_ = v2 & new_n123_;
  assign new_n125_ = ~v3 & new_n124_;
  assign new_n126_ = ~v4 & new_n125_;
  assign new_n127_ = v5 & new_n126_;
  assign new_n128_ = v6 & new_n127_;
  assign \v8.12  = v7 & new_n128_;
  assign new_n130_ = v3 & new_n91_;
  assign new_n131_ = ~v4 & new_n130_;
  assign new_n132_ = v5 & new_n131_;
  assign new_n133_ = v6 & new_n132_;
  assign \v8.13  = v7 & new_n133_;
  assign new_n135_ = ~v2 & new_n123_;
  assign new_n136_ = v3 & new_n135_;
  assign new_n137_ = ~v4 & new_n136_;
  assign new_n138_ = v5 & new_n137_;
  assign new_n139_ = v6 & new_n138_;
  assign \v8.14  = v7 & new_n139_;
  assign new_n141_ = v2 & new_n90_;
  assign new_n142_ = v3 & new_n141_;
  assign new_n143_ = ~v4 & new_n142_;
  assign new_n144_ = v5 & new_n143_;
  assign new_n145_ = v6 & new_n144_;
  assign \v8.15  = v7 & new_n145_;
  assign new_n147_ = v3 & new_n117_;
  assign new_n148_ = ~v4 & new_n147_;
  assign new_n149_ = v5 & new_n148_;
  assign new_n150_ = v6 & new_n149_;
  assign \v8.16  = v7 & new_n150_;
  assign new_n152_ = v4 & ~v5;
  assign new_n153_ = ~v2 & new_n152_;
  assign new_n154_ = ~v1 & new_n153_;
  assign \v8.17  = v0 & new_n154_;
  assign new_n156_ = v3 & new_n152_;
  assign new_n157_ = v2 & new_n156_;
  assign new_n158_ = ~v1 & new_n157_;
  assign \v8.18  = ~v0 & new_n158_;
  assign new_n160_ = ~v3 & v4;
  assign new_n161_ = ~v2 & new_n160_;
  assign new_n162_ = ~v1 & new_n161_;
  assign \v8.19  = ~v0 & new_n162_;
  assign new_n164_ = ~v3 & \v8.0 ;
  assign new_n165_ = ~v2 & new_n164_;
  assign new_n166_ = ~v1 & new_n165_;
  assign \v8.20  = v0 & new_n166_;
  assign new_n168_ = ~v2 & new_n86_;
  assign new_n169_ = ~v1 & new_n168_;
  assign \v8.21  = v0 & new_n169_;
  assign new_n171_ = ~v5 & new_n111_;
  assign new_n172_ = ~v4 & new_n171_;
  assign new_n173_ = ~v2 & new_n172_;
  assign new_n174_ = ~v1 & new_n173_;
  assign \v8.22  = v0 & new_n174_;
  assign new_n176_ = v3 & v5;
  assign new_n177_ = ~v2 & new_n176_;
  assign new_n178_ = ~v1 & new_n177_;
  assign \v8.23  = ~v0 & new_n178_;
  assign new_n180_ = ~v2 & new_n104_;
  assign new_n181_ = ~v3 & new_n180_;
  assign new_n182_ = ~v4 & new_n181_;
  assign new_n183_ = ~v5 & new_n182_;
  assign new_n184_ = v6 & new_n183_;
  assign \v8.24  = ~v7 & new_n184_;
  assign new_n186_ = ~v5 & new_n93_;
  assign new_n187_ = v6 & new_n186_;
  assign \v8.25  = ~v7 & new_n187_;
  assign new_n189_ = ~v3 & new_n172_;
  assign new_n190_ = v2 & new_n189_;
  assign \v8.26  = v0 & new_n190_;
  assign new_n192_ = ~v3 & new_n141_;
  assign new_n193_ = ~v4 & new_n192_;
  assign new_n194_ = ~v5 & new_n193_;
  assign new_n195_ = v6 & new_n194_;
  assign \v8.27  = ~v7 & new_n195_;
  assign new_n197_ = v3 & new_n124_;
  assign new_n198_ = ~v4 & new_n197_;
  assign new_n199_ = ~v5 & new_n198_;
  assign new_n200_ = v6 & new_n199_;
  assign \v8.28  = v7 & new_n200_;
  assign new_n202_ = ~v6 & new_n183_;
  assign \v8.29  = v7 & new_n202_;
  assign new_n204_ = ~v5 & new_n100_;
  assign new_n205_ = v6 & new_n204_;
  assign \v8.30  = v7 & new_n205_;
  assign new_n207_ = ~v4 & v5;
  assign new_n208_ = ~new_n152_ & ~new_n207_;
  assign new_n209_ = v4 & v5;
  assign new_n210_ = ~v4 & ~v5;
  assign new_n211_ = ~new_n209_ & ~new_n210_;
  assign new_n212_ = ~v1 & v2;
  assign new_n213_ = v0 & new_n212_;
  assign new_n214_ = ~v1 & ~new_n213_;
  assign new_n215_ = ~v2 & v3;
  assign new_n216_ = v2 & ~v3;
  assign new_n217_ = ~new_n215_ & ~new_n216_;
  assign new_n218_ = ~v1 & ~new_n217_;
  assign new_n219_ = ~v0 & new_n218_;
  assign new_n220_ = new_n214_ & ~new_n219_;
  assign new_n221_ = ~new_n211_ & ~new_n220_;
  assign new_n222_ = v2 & v3;
  assign new_n223_ = ~v2 & ~v3;
  assign new_n224_ = ~new_n222_ & ~new_n223_;
  assign new_n225_ = ~v5 & ~new_n224_;
  assign new_n226_ = ~v4 & new_n225_;
  assign new_n227_ = ~v1 & new_n226_;
  assign new_n228_ = ~v0 & new_n227_;
  assign new_n229_ = ~new_n221_ & ~new_n228_;
  assign new_n230_ = new_n208_ & new_n229_;
  assign new_n231_ = ~v5 & v6;
  assign new_n232_ = ~v4 & new_n231_;
  assign new_n233_ = ~v2 & new_n232_;
  assign new_n234_ = ~v1 & new_n233_;
  assign new_n235_ = v0 & new_n234_;
  assign \v8.31  = ~new_n230_ | new_n235_;
  assign new_n237_ = ~v0 & ~new_n90_;
  assign new_n238_ = ~v1 & ~v2;
  assign new_n239_ = ~v0 & new_n238_;
  assign new_n240_ = new_n237_ & ~new_n239_;
  assign new_n241_ = new_n104_ & new_n216_;
  assign new_n242_ = new_n240_ & ~new_n241_;
  assign new_n243_ = ~new_n208_ & ~new_n242_;
  assign new_n244_ = v3 & ~v4;
  assign new_n245_ = v2 & new_n244_;
  assign new_n246_ = new_n209_ & new_n223_;
  assign new_n247_ = ~new_n245_ & ~new_n246_;
  assign new_n248_ = ~v0 & ~new_n247_;
  assign new_n249_ = v0 & ~v2;
  assign new_n250_ = ~v3 & new_n210_;
  assign new_n251_ = new_n249_ & new_n250_;
  assign new_n252_ = ~new_n248_ & ~new_n251_;
  assign new_n253_ = ~v1 & ~new_n252_;
  assign new_n254_ = ~new_n221_ & ~new_n253_;
  assign new_n255_ = ~new_n243_ & new_n254_;
  assign new_n256_ = v3 & v6;
  assign new_n257_ = v0 & new_n256_;
  assign new_n258_ = ~v3 & ~v6;
  assign new_n259_ = ~v0 & new_n258_;
  assign new_n260_ = ~new_n257_ & ~new_n259_;
  assign new_n261_ = ~v5 & ~new_n260_;
  assign new_n262_ = ~v4 & new_n261_;
  assign new_n263_ = ~v2 & new_n262_;
  assign new_n264_ = ~v1 & new_n263_;
  assign new_n265_ = new_n255_ & ~new_n264_;
  assign new_n266_ = new_n104_ & new_n223_;
  assign new_n267_ = new_n111_ & new_n210_;
  assign new_n268_ = new_n266_ & new_n267_;
  assign \v8.32  = ~new_n265_ | new_n268_;
  assign new_n270_ = v0 & ~new_n249_;
  assign new_n271_ = v2 & v4;
  assign new_n272_ = v0 & new_n271_;
  assign new_n273_ = new_n270_ & ~new_n272_;
  assign new_n274_ = v0 & v2;
  assign new_n275_ = ~v4 & ~v6;
  assign new_n276_ = new_n274_ & new_n275_;
  assign new_n277_ = new_n273_ & ~new_n276_;
  assign new_n278_ = ~v4 & new_n80_;
  assign new_n279_ = new_n274_ & new_n278_;
  assign new_n280_ = new_n277_ & ~new_n279_;
  assign new_n281_ = new_n111_ & new_n207_;
  assign new_n282_ = new_n213_ & new_n281_;
  assign new_n283_ = new_n280_ & ~new_n282_;
  assign new_n284_ = new_n97_ & new_n222_;
  assign new_n285_ = new_n267_ & new_n284_;
  assign \v8.33  = ~new_n283_ | new_n285_;
  assign new_n287_ = ~v1 & v5;
  assign new_n288_ = ~v1 & ~new_n287_;
  assign new_n289_ = v4 & ~new_n288_;
  assign new_n290_ = v1 & new_n210_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = new_n104_ & new_n152_;
  assign new_n293_ = new_n291_ & ~new_n292_;
  assign new_n294_ = v5 & v6;
  assign new_n295_ = ~new_n72_ & ~new_n294_;
  assign new_n296_ = ~v1 & ~new_n295_;
  assign new_n297_ = v1 & new_n294_;
  assign new_n298_ = ~new_n296_ & ~new_n297_;
  assign new_n299_ = ~v4 & ~new_n298_;
  assign new_n300_ = new_n293_ & ~new_n299_;
  assign new_n301_ = v5 & ~v6;
  assign new_n302_ = new_n104_ & new_n231_;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = v7 & ~new_n303_;
  assign new_n305_ = new_n81_ & new_n123_;
  assign new_n306_ = ~new_n304_ & ~new_n305_;
  assign new_n307_ = ~v4 & ~new_n306_;
  assign new_n308_ = new_n300_ & ~new_n307_;
  assign new_n309_ = ~v4 & v7;
  assign new_n310_ = ~v4 & ~new_n309_;
  assign new_n311_ = v2 & ~new_n310_;
  assign new_n312_ = v0 & new_n311_;
  assign new_n313_ = ~v0 & ~v2;
  assign new_n314_ = ~v4 & ~v7;
  assign new_n315_ = new_n313_ & new_n314_;
  assign new_n316_ = ~new_n312_ & ~new_n315_;
  assign new_n317_ = v6 & ~new_n316_;
  assign new_n318_ = v4 & ~v6;
  assign new_n319_ = v2 & new_n318_;
  assign new_n320_ = v0 & new_n319_;
  assign new_n321_ = ~new_n317_ & ~new_n320_;
  assign new_n322_ = ~v5 & ~new_n321_;
  assign new_n323_ = ~v1 & new_n322_;
  assign new_n324_ = new_n308_ & ~new_n323_;
  assign new_n325_ = ~v3 & new_n301_;
  assign new_n326_ = ~v0 & new_n212_;
  assign new_n327_ = v3 & new_n231_;
  assign new_n328_ = new_n326_ & new_n327_;
  assign new_n329_ = ~new_n325_ & ~new_n328_;
  assign new_n330_ = ~v7 & ~new_n329_;
  assign new_n331_ = ~v4 & new_n330_;
  assign \v8.34  = ~new_n324_ | new_n331_;
  assign new_n333_ = ~v1 & ~v4;
  assign new_n334_ = ~v1 & ~new_n333_;
  assign new_n335_ = new_n123_ & new_n271_;
  assign new_n336_ = new_n334_ & ~new_n335_;
  assign new_n337_ = ~v0 & v2;
  assign new_n338_ = ~new_n249_ & ~new_n337_;
  assign new_n339_ = ~v5 & ~new_n338_;
  assign new_n340_ = v4 & new_n339_;
  assign new_n341_ = ~v1 & new_n340_;
  assign new_n342_ = new_n336_ & ~new_n341_;
  assign new_n343_ = ~v3 & v5;
  assign new_n344_ = v2 & new_n343_;
  assign new_n345_ = ~new_n215_ & ~new_n344_;
  assign new_n346_ = v4 & ~new_n345_;
  assign new_n347_ = ~v1 & new_n346_;
  assign new_n348_ = ~v0 & new_n347_;
  assign \v8.35  = ~new_n342_ | new_n348_;
  assign new_n350_ = ~new_n274_ & ~new_n313_;
  assign new_n351_ = ~new_n288_ & ~new_n338_;
  assign new_n352_ = new_n350_ & ~new_n351_;
  assign new_n353_ = ~v0 & new_n271_;
  assign new_n354_ = ~v2 & ~v4;
  assign new_n355_ = v0 & new_n354_;
  assign new_n356_ = ~new_n353_ & ~new_n355_;
  assign new_n357_ = ~v5 & ~new_n356_;
  assign new_n358_ = ~v1 & new_n357_;
  assign new_n359_ = new_n352_ & ~new_n358_;
  assign new_n360_ = v3 & new_n210_;
  assign new_n361_ = new_n326_ & new_n360_;
  assign new_n362_ = new_n359_ & ~new_n361_;
  assign new_n363_ = ~v3 & ~v4;
  assign new_n364_ = new_n72_ & new_n363_;
  assign new_n365_ = new_n326_ & new_n364_;
  assign new_n366_ = new_n362_ & ~new_n365_;
  assign new_n367_ = new_n241_ & new_n267_;
  assign \v8.36  = ~new_n366_ | new_n367_;
  assign new_n369_ = v0 & ~new_n123_;
  assign new_n370_ = ~v3 & ~new_n369_;
  assign new_n371_ = v0 & ~new_n97_;
  assign new_n372_ = v4 & ~new_n371_;
  assign new_n373_ = v3 & new_n372_;
  assign new_n374_ = ~new_n370_ & ~new_n373_;
  assign new_n375_ = v1 & new_n207_;
  assign new_n376_ = ~v1 & new_n152_;
  assign new_n377_ = ~new_n375_ & ~new_n376_;
  assign new_n378_ = v0 & ~new_n377_;
  assign new_n379_ = ~v0 & new_n207_;
  assign new_n380_ = ~new_n378_ & ~new_n379_;
  assign new_n381_ = v3 & ~new_n380_;
  assign new_n382_ = new_n374_ & ~new_n381_;
  assign new_n383_ = v1 & ~v3;
  assign new_n384_ = ~v1 & new_n176_;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = v2 & ~new_n385_;
  assign new_n387_ = v0 & new_n386_;
  assign new_n388_ = new_n382_ & ~new_n387_;
  assign new_n389_ = ~new_n86_ & new_n388_;
  assign new_n390_ = v3 & new_n172_;
  assign \v8.37  = ~new_n389_ | new_n390_;
  assign new_n392_ = ~new_n161_ & ~new_n245_;
  assign new_n393_ = ~v0 & ~new_n392_;
  assign new_n394_ = new_n249_ & new_n363_;
  assign new_n395_ = ~new_n393_ & ~new_n394_;
  assign new_n396_ = ~v1 & ~new_n395_;
  assign new_n397_ = new_n220_ & ~new_n396_;
  assign new_n398_ = v0 & v3;
  assign new_n399_ = ~v0 & ~v3;
  assign new_n400_ = ~new_n398_ & ~new_n399_;
  assign new_n401_ = v5 & ~new_n400_;
  assign new_n402_ = ~v4 & new_n401_;
  assign new_n403_ = ~v2 & new_n402_;
  assign new_n404_ = ~v1 & new_n403_;
  assign new_n405_ = new_n397_ & ~new_n404_;
  assign new_n406_ = ~new_n264_ & new_n405_;
  assign \v8.38  = new_n268_ | ~new_n406_;
  assign new_n408_ = ~new_n231_ & ~new_n301_;
  assign new_n409_ = v4 & ~new_n408_;
  assign new_n410_ = new_n301_ & new_n363_;
  assign new_n411_ = ~new_n409_ & ~new_n410_;
  assign new_n412_ = ~v0 & new_n232_;
  assign new_n413_ = new_n411_ & ~new_n412_;
  assign new_n414_ = new_n295_ & new_n413_;
  assign new_n415_ = ~v6 & v7;
  assign new_n416_ = v5 & new_n415_;
  assign new_n417_ = ~new_n81_ & ~new_n416_;
  assign new_n418_ = v0 & ~new_n417_;
  assign new_n419_ = ~v0 & v5;
  assign new_n420_ = new_n415_ & new_n419_;
  assign new_n421_ = ~new_n418_ & ~new_n420_;
  assign new_n422_ = v3 & ~new_n421_;
  assign new_n423_ = v0 & ~v3;
  assign new_n424_ = new_n81_ & new_n423_;
  assign new_n425_ = ~new_n422_ & ~new_n424_;
  assign new_n426_ = ~v4 & ~new_n425_;
  assign new_n427_ = new_n414_ & ~new_n426_;
  assign new_n428_ = v1 & new_n172_;
  assign new_n429_ = v0 & new_n428_;
  assign new_n430_ = new_n427_ & ~new_n429_;
  assign new_n431_ = v2 & new_n172_;
  assign new_n432_ = ~v1 & new_n431_;
  assign new_n433_ = v0 & new_n432_;
  assign \v8.39  = ~new_n430_ | new_n433_;
  assign new_n435_ = ~new_n224_ & ~new_n237_;
  assign new_n436_ = new_n217_ & ~new_n435_;
  assign new_n437_ = ~new_n208_ & ~new_n436_;
  assign new_n438_ = ~v0 & ~new_n217_;
  assign new_n439_ = v0 & new_n222_;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = ~v0 & ~new_n399_;
  assign new_n442_ = ~v2 & ~new_n441_;
  assign new_n443_ = ~v0 & new_n222_;
  assign new_n444_ = ~new_n442_ & ~new_n443_;
  assign new_n445_ = v1 & ~new_n444_;
  assign new_n446_ = new_n440_ & ~new_n445_;
  assign new_n447_ = ~new_n211_ & ~new_n446_;
  assign new_n448_ = v0 & new_n160_;
  assign new_n449_ = new_n104_ & new_n244_;
  assign new_n450_ = ~new_n448_ & ~new_n449_;
  assign new_n451_ = v5 & ~new_n450_;
  assign new_n452_ = new_n104_ & new_n360_;
  assign new_n453_ = ~new_n451_ & ~new_n452_;
  assign new_n454_ = v2 & ~new_n453_;
  assign new_n455_ = ~v3 & new_n207_;
  assign new_n456_ = new_n239_ & new_n455_;
  assign new_n457_ = ~new_n454_ & ~new_n456_;
  assign new_n458_ = ~new_n447_ & new_n457_;
  assign new_n459_ = ~new_n437_ & new_n458_;
  assign new_n460_ = ~v2 & v6;
  assign new_n461_ = v2 & ~v6;
  assign new_n462_ = ~new_n460_ & ~new_n461_;
  assign new_n463_ = ~v1 & ~new_n462_;
  assign new_n464_ = v1 & new_n461_;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign new_n466_ = ~v3 & ~new_n465_;
  assign new_n467_ = new_n238_ & new_n256_;
  assign new_n468_ = ~new_n466_ & ~new_n467_;
  assign new_n469_ = v0 & ~new_n468_;
  assign new_n470_ = ~v2 & new_n258_;
  assign new_n471_ = new_n104_ & new_n470_;
  assign new_n472_ = ~new_n469_ & ~new_n471_;
  assign new_n473_ = ~v5 & ~new_n472_;
  assign new_n474_ = ~v4 & new_n473_;
  assign new_n475_ = new_n459_ & ~new_n474_;
  assign new_n476_ = v2 & ~v7;
  assign new_n477_ = v0 & new_n476_;
  assign new_n478_ = ~v2 & v7;
  assign new_n479_ = new_n104_ & new_n478_;
  assign new_n480_ = ~new_n477_ & ~new_n479_;
  assign new_n481_ = v6 & ~new_n480_;
  assign new_n482_ = ~v5 & new_n481_;
  assign new_n483_ = ~v4 & new_n482_;
  assign new_n484_ = ~v3 & new_n483_;
  assign \v8.40  = ~new_n475_ | new_n484_;
  assign new_n486_ = v1 & v3;
  assign new_n487_ = ~v1 & ~v3;
  assign new_n488_ = ~new_n486_ & ~new_n487_;
  assign new_n489_ = ~v1 & v3;
  assign new_n490_ = ~new_n383_ & ~new_n489_;
  assign new_n491_ = v0 & ~new_n274_;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = new_n488_ & ~new_n492_;
  assign new_n494_ = v3 & ~v5;
  assign new_n495_ = ~v2 & new_n494_;
  assign new_n496_ = ~v1 & new_n495_;
  assign new_n497_ = v0 & new_n496_;
  assign \v8.41  = ~new_n493_ | new_n497_;
  assign new_n499_ = ~v0 & ~v4;
  assign new_n500_ = new_n231_ & new_n499_;
  assign new_n501_ = ~new_n409_ & ~new_n500_;
  assign new_n502_ = new_n295_ & new_n501_;
  assign new_n503_ = ~v4 & ~new_n421_;
  assign new_n504_ = new_n502_ & ~new_n503_;
  assign new_n505_ = v1 & ~v4;
  assign new_n506_ = v0 & new_n505_;
  assign new_n507_ = new_n171_ & new_n506_;
  assign new_n508_ = new_n504_ & ~new_n507_;
  assign new_n509_ = new_n123_ & new_n216_;
  assign new_n510_ = new_n267_ & new_n509_;
  assign \v8.42  = ~new_n508_ | new_n510_;
  assign new_n512_ = ~v0 & new_n333_;
  assign new_n513_ = new_n214_ & ~new_n512_;
  assign new_n514_ = ~new_n295_ & ~new_n513_;
  assign new_n515_ = ~new_n214_ & ~new_n408_;
  assign new_n516_ = v4 & new_n515_;
  assign new_n517_ = v1 & ~v5;
  assign new_n518_ = ~new_n287_ & ~new_n517_;
  assign new_n519_ = v0 & ~new_n518_;
  assign new_n520_ = ~v0 & new_n517_;
  assign new_n521_ = ~new_n519_ & ~new_n520_;
  assign new_n522_ = ~v2 & ~new_n521_;
  assign new_n523_ = v2 & ~v5;
  assign new_n524_ = ~v0 & new_n523_;
  assign new_n525_ = ~new_n522_ & ~new_n524_;
  assign new_n526_ = v6 & ~new_n525_;
  assign new_n527_ = ~v4 & new_n526_;
  assign new_n528_ = ~new_n516_ & ~new_n527_;
  assign new_n529_ = ~new_n514_ & new_n528_;
  assign new_n530_ = ~new_n305_ & ~new_n416_;
  assign new_n531_ = new_n97_ & new_n476_;
  assign new_n532_ = ~new_n479_ & ~new_n531_;
  assign new_n533_ = v6 & ~new_n532_;
  assign new_n534_ = ~v5 & new_n533_;
  assign new_n535_ = new_n530_ & ~new_n534_;
  assign new_n536_ = ~v4 & ~new_n535_;
  assign new_n537_ = new_n529_ & ~new_n536_;
  assign new_n538_ = ~v4 & ~new_n314_;
  assign new_n539_ = ~v2 & ~new_n538_;
  assign new_n540_ = ~v1 & new_n539_;
  assign new_n541_ = ~v0 & new_n540_;
  assign new_n542_ = v2 & new_n309_;
  assign new_n543_ = new_n97_ & new_n542_;
  assign new_n544_ = ~new_n541_ & ~new_n543_;
  assign new_n545_ = v6 & ~new_n544_;
  assign new_n546_ = ~v2 & new_n318_;
  assign new_n547_ = ~v1 & new_n546_;
  assign new_n548_ = ~v0 & new_n547_;
  assign new_n549_ = ~new_n545_ & ~new_n548_;
  assign new_n550_ = ~v5 & ~new_n549_;
  assign new_n551_ = ~v2 & new_n209_;
  assign new_n552_ = ~v1 & new_n551_;
  assign new_n553_ = ~v0 & new_n552_;
  assign new_n554_ = ~new_n550_ & ~new_n553_;
  assign new_n555_ = v3 & ~new_n554_;
  assign new_n556_ = v2 & new_n160_;
  assign new_n557_ = ~v1 & new_n556_;
  assign new_n558_ = ~v0 & new_n557_;
  assign new_n559_ = ~new_n555_ & ~new_n558_;
  assign \v8.43  = ~new_n537_ | ~new_n559_;
  assign new_n561_ = v0 & v4;
  assign new_n562_ = ~new_n499_ & ~new_n561_;
  assign new_n563_ = ~v0 & v4;
  assign new_n564_ = v0 & ~v4;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = ~v1 & ~new_n212_;
  assign new_n567_ = ~v1 & new_n215_;
  assign new_n568_ = new_n566_ & ~new_n567_;
  assign new_n569_ = ~new_n565_ & ~new_n568_;
  assign new_n570_ = new_n562_ & ~new_n569_;
  assign new_n571_ = v0 & new_n238_;
  assign new_n572_ = new_n455_ & new_n571_;
  assign new_n573_ = new_n570_ & ~new_n572_;
  assign new_n574_ = new_n231_ & new_n363_;
  assign new_n575_ = new_n571_ & new_n574_;
  assign \v8.44  = ~new_n573_ | new_n575_;
  assign new_n577_ = v1 & ~v2;
  assign new_n578_ = ~new_n212_ & ~new_n577_;
  assign new_n579_ = v1 & v2;
  assign new_n580_ = ~new_n238_ & ~new_n579_;
  assign new_n581_ = v0 & ~new_n580_;
  assign new_n582_ = new_n578_ & ~new_n581_;
  assign new_n583_ = ~v2 & v4;
  assign new_n584_ = new_n104_ & new_n583_;
  assign new_n585_ = new_n582_ & ~new_n584_;
  assign new_n586_ = v5 & ~new_n580_;
  assign new_n587_ = ~v4 & new_n586_;
  assign new_n588_ = ~v0 & new_n587_;
  assign new_n589_ = new_n585_ & ~new_n588_;
  assign new_n590_ = v2 & v6;
  assign new_n591_ = v1 & new_n590_;
  assign new_n592_ = ~v2 & ~v6;
  assign new_n593_ = ~v1 & new_n592_;
  assign new_n594_ = ~new_n591_ & ~new_n593_;
  assign new_n595_ = ~v5 & ~new_n594_;
  assign new_n596_ = ~v4 & new_n595_;
  assign new_n597_ = ~v0 & new_n596_;
  assign new_n598_ = new_n589_ & ~new_n597_;
  assign new_n599_ = ~v2 & new_n82_;
  assign new_n600_ = ~v1 & new_n599_;
  assign new_n601_ = ~v0 & new_n600_;
  assign \v8.45  = ~new_n598_ | new_n601_;
  assign new_n603_ = ~v0 & ~new_n104_;
  assign new_n604_ = ~v0 & new_n579_;
  assign new_n605_ = new_n603_ & ~new_n604_;
  assign new_n606_ = new_n90_ & new_n215_;
  assign new_n607_ = new_n605_ & ~new_n606_;
  assign new_n608_ = ~v0 & new_n577_;
  assign new_n609_ = new_n455_ & new_n608_;
  assign new_n610_ = new_n607_ & ~new_n609_;
  assign new_n611_ = new_n90_ & new_n223_;
  assign new_n612_ = new_n80_ & new_n210_;
  assign new_n613_ = new_n611_ & new_n612_;
  assign \v8.46  = ~new_n610_ | new_n613_;
  assign new_n615_ = ~new_n571_ & new_n578_;
  assign new_n616_ = v0 & new_n579_;
  assign new_n617_ = ~new_n239_ & ~new_n616_;
  assign new_n618_ = v4 & ~new_n617_;
  assign new_n619_ = new_n615_ & ~new_n618_;
  assign new_n620_ = ~v0 & new_n586_;
  assign new_n621_ = new_n97_ & new_n523_;
  assign new_n622_ = ~new_n620_ & ~new_n621_;
  assign new_n623_ = ~v4 & ~new_n622_;
  assign new_n624_ = new_n619_ & ~new_n623_;
  assign new_n625_ = ~v0 & new_n595_;
  assign new_n626_ = v2 & new_n301_;
  assign new_n627_ = new_n97_ & new_n626_;
  assign new_n628_ = ~new_n625_ & ~new_n627_;
  assign new_n629_ = ~v4 & ~new_n628_;
  assign new_n630_ = new_n624_ & ~new_n629_;
  assign new_n631_ = new_n294_ & new_n363_;
  assign new_n632_ = new_n616_ & new_n631_;
  assign new_n633_ = new_n630_ & ~new_n632_;
  assign new_n634_ = ~v2 & ~v5;
  assign new_n635_ = ~v1 & new_n634_;
  assign new_n636_ = ~v0 & new_n635_;
  assign new_n637_ = v2 & new_n176_;
  assign new_n638_ = new_n97_ & new_n637_;
  assign new_n639_ = ~new_n636_ & ~new_n638_;
  assign new_n640_ = ~v7 & ~new_n639_;
  assign new_n641_ = v6 & new_n640_;
  assign new_n642_ = ~v4 & new_n641_;
  assign \v8.47  = ~new_n633_ | new_n642_;
  assign new_n644_ = new_n237_ & ~new_n326_;
  assign new_n645_ = ~new_n266_ & new_n644_;
  assign new_n646_ = ~v2 & new_n244_;
  assign new_n647_ = new_n104_ & new_n646_;
  assign new_n648_ = new_n645_ & ~new_n647_;
  assign new_n649_ = ~new_n408_ & ~new_n648_;
  assign new_n650_ = ~new_n295_ & ~new_n645_;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = new_n104_ & new_n215_;
  assign new_n653_ = new_n80_ & new_n207_;
  assign new_n654_ = new_n652_ & new_n653_;
  assign \v8.48  = ~new_n651_ | new_n654_;
  assign new_n656_ = v3 & v4;
  assign new_n657_ = v2 & new_n656_;
  assign new_n658_ = new_n104_ & new_n657_;
  assign new_n659_ = new_n240_ & ~new_n658_;
  assign new_n660_ = v2 & new_n207_;
  assign new_n661_ = ~v1 & new_n660_;
  assign new_n662_ = ~v0 & new_n661_;
  assign new_n663_ = new_n659_ & ~new_n662_;
  assign new_n664_ = v2 & new_n232_;
  assign new_n665_ = ~v1 & new_n664_;
  assign new_n666_ = ~v0 & new_n665_;
  assign \v8.49  = ~new_n663_ | new_n666_;
  assign new_n668_ = ~v2 & ~new_n583_;
  assign new_n669_ = ~v2 & new_n207_;
  assign new_n670_ = new_n668_ & ~new_n669_;
  assign new_n671_ = new_n72_ & new_n354_;
  assign new_n672_ = new_n670_ & ~new_n671_;
  assign new_n673_ = new_n81_ & new_n354_;
  assign new_n674_ = new_n672_ & ~new_n673_;
  assign new_n675_ = new_n267_ & new_n571_;
  assign new_n676_ = new_n674_ & ~new_n675_;
  assign new_n677_ = new_n97_ & new_n223_;
  assign new_n678_ = new_n267_ & new_n677_;
  assign \v8.50  = ~new_n676_ | new_n678_;
  assign new_n680_ = ~new_n90_ & ~new_n123_;
  assign new_n681_ = new_n104_ & new_n271_;
  assign new_n682_ = new_n680_ & ~new_n681_;
  assign new_n683_ = ~new_n104_ & ~new_n616_;
  assign new_n684_ = v5 & ~new_n683_;
  assign new_n685_ = ~v4 & new_n684_;
  assign new_n686_ = new_n682_ & ~new_n685_;
  assign new_n687_ = v0 & new_n486_;
  assign new_n688_ = new_n104_ & new_n160_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = new_n104_ & new_n250_;
  assign new_n691_ = new_n689_ & ~new_n690_;
  assign new_n692_ = ~v2 & ~new_n691_;
  assign new_n693_ = new_n250_ & new_n326_;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = new_n686_ & new_n694_;
  assign new_n696_ = ~v0 & new_n489_;
  assign new_n697_ = v0 & new_n383_;
  assign new_n698_ = ~new_n696_ & ~new_n697_;
  assign new_n699_ = ~new_n284_ & new_n698_;
  assign new_n700_ = v6 & ~new_n699_;
  assign new_n701_ = ~v5 & new_n700_;
  assign new_n702_ = v0 & new_n577_;
  assign new_n703_ = new_n325_ & new_n702_;
  assign new_n704_ = ~new_n701_ & ~new_n703_;
  assign new_n705_ = ~v4 & ~new_n704_;
  assign new_n706_ = new_n695_ & ~new_n705_;
  assign new_n707_ = new_n653_ & new_n677_;
  assign \v8.51  = ~new_n706_ | new_n707_;
  assign new_n709_ = ~v5 & ~new_n520_;
  assign new_n710_ = ~v4 & ~new_n709_;
  assign new_n711_ = v1 & v4;
  assign new_n712_ = ~v0 & new_n711_;
  assign new_n713_ = ~new_n710_ & ~new_n712_;
  assign new_n714_ = ~v4 & ~new_n210_;
  assign new_n715_ = v3 & ~new_n714_;
  assign new_n716_ = v0 & new_n715_;
  assign new_n717_ = new_n713_ & ~new_n716_;
  assign new_n718_ = ~v0 & ~new_n224_;
  assign new_n719_ = v0 & new_n223_;
  assign new_n720_ = ~new_n718_ & ~new_n719_;
  assign new_n721_ = v4 & ~new_n720_;
  assign new_n722_ = ~v2 & new_n250_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = ~v1 & ~new_n723_;
  assign new_n725_ = new_n717_ & ~new_n724_;
  assign new_n726_ = ~v1 & new_n216_;
  assign new_n727_ = new_n698_ & ~new_n726_;
  assign new_n728_ = v6 & ~new_n727_;
  assign new_n729_ = ~v5 & new_n728_;
  assign new_n730_ = ~v4 & new_n729_;
  assign \v8.52  = ~new_n725_ | new_n730_;
  assign new_n732_ = v4 & ~new_n224_;
  assign new_n733_ = new_n217_ & ~new_n732_;
  assign new_n734_ = ~v1 & ~new_n733_;
  assign new_n735_ = new_n160_ & new_n577_;
  assign new_n736_ = ~new_n734_ & ~new_n735_;
  assign new_n737_ = ~v1 & ~new_n224_;
  assign new_n738_ = v1 & new_n223_;
  assign new_n739_ = ~new_n737_ & ~new_n738_;
  assign new_n740_ = ~v5 & ~new_n739_;
  assign new_n741_ = v5 & ~new_n217_;
  assign new_n742_ = v1 & new_n741_;
  assign new_n743_ = ~new_n740_ & ~new_n742_;
  assign new_n744_ = ~v4 & ~new_n743_;
  assign new_n745_ = new_n736_ & ~new_n744_;
  assign new_n746_ = ~v0 & v3;
  assign new_n747_ = ~new_n448_ & ~new_n746_;
  assign new_n748_ = new_n210_ & new_n423_;
  assign new_n749_ = new_n747_ & ~new_n748_;
  assign new_n750_ = v2 & ~new_n749_;
  assign new_n751_ = new_n249_ & new_n455_;
  assign new_n752_ = ~new_n750_ & ~new_n751_;
  assign new_n753_ = v1 & ~new_n752_;
  assign new_n754_ = v3 & new_n207_;
  assign new_n755_ = new_n213_ & new_n754_;
  assign new_n756_ = ~new_n753_ & ~new_n755_;
  assign new_n757_ = new_n745_ & new_n756_;
  assign new_n758_ = ~v6 & ~new_n739_;
  assign new_n759_ = v5 & new_n758_;
  assign new_n760_ = v6 & ~new_n217_;
  assign new_n761_ = ~v5 & new_n760_;
  assign new_n762_ = v1 & new_n761_;
  assign new_n763_ = ~new_n759_ & ~new_n762_;
  assign new_n764_ = ~v0 & ~new_n763_;
  assign new_n765_ = v2 & ~new_n408_;
  assign new_n766_ = ~v2 & new_n231_;
  assign new_n767_ = ~new_n765_ & ~new_n766_;
  assign new_n768_ = v3 & ~new_n767_;
  assign new_n769_ = v1 & new_n768_;
  assign new_n770_ = new_n238_ & new_n325_;
  assign new_n771_ = ~new_n769_ & ~new_n770_;
  assign new_n772_ = v0 & ~new_n771_;
  assign new_n773_ = ~new_n764_ & ~new_n772_;
  assign new_n774_ = ~v4 & ~new_n773_;
  assign new_n775_ = new_n757_ & ~new_n774_;
  assign new_n776_ = v1 & new_n222_;
  assign new_n777_ = ~v1 & new_n223_;
  assign new_n778_ = ~new_n776_ & ~new_n777_;
  assign new_n779_ = v0 & ~new_n778_;
  assign new_n780_ = ~v0 & ~new_n739_;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = ~v7 & ~new_n781_;
  assign new_n783_ = v6 & new_n782_;
  assign new_n784_ = v5 & new_n783_;
  assign new_n785_ = ~v4 & new_n784_;
  assign \v8.53  = ~new_n775_ | new_n785_;
  assign new_n787_ = v0 & new_n333_;
  assign new_n788_ = ~v4 & ~new_n787_;
  assign new_n789_ = ~new_n217_ & ~new_n788_;
  assign new_n790_ = ~new_n284_ & ~new_n737_;
  assign new_n791_ = ~new_n160_ & ~new_n244_;
  assign new_n792_ = ~v2 & ~new_n791_;
  assign new_n793_ = v1 & new_n792_;
  assign new_n794_ = v0 & new_n793_;
  assign new_n795_ = new_n790_ & ~new_n794_;
  assign new_n796_ = ~new_n789_ & new_n795_;
  assign new_n797_ = ~v0 & ~new_n337_;
  assign new_n798_ = ~v3 & ~new_n797_;
  assign new_n799_ = ~v0 & new_n215_;
  assign new_n800_ = ~new_n798_ & ~new_n799_;
  assign new_n801_ = v1 & ~new_n800_;
  assign new_n802_ = ~new_n219_ & ~new_n801_;
  assign new_n803_ = ~v5 & ~new_n802_;
  assign new_n804_ = ~v2 & new_n343_;
  assign new_n805_ = new_n90_ & new_n804_;
  assign new_n806_ = ~new_n803_ & ~new_n805_;
  assign new_n807_ = ~v4 & ~new_n806_;
  assign new_n808_ = new_n796_ & ~new_n807_;
  assign new_n809_ = ~new_n423_ & ~new_n746_;
  assign new_n810_ = ~v0 & new_n216_;
  assign new_n811_ = new_n809_ & ~new_n810_;
  assign new_n812_ = ~v6 & ~new_n811_;
  assign new_n813_ = v5 & new_n812_;
  assign new_n814_ = v6 & ~new_n224_;
  assign new_n815_ = ~v5 & new_n814_;
  assign new_n816_ = ~v0 & new_n815_;
  assign new_n817_ = ~new_n813_ & ~new_n816_;
  assign new_n818_ = v1 & ~new_n817_;
  assign new_n819_ = ~v6 & ~new_n217_;
  assign new_n820_ = v5 & new_n819_;
  assign new_n821_ = ~v1 & new_n820_;
  assign new_n822_ = ~v0 & new_n821_;
  assign new_n823_ = ~new_n818_ & ~new_n822_;
  assign new_n824_ = ~v4 & ~new_n823_;
  assign new_n825_ = new_n808_ & ~new_n824_;
  assign new_n826_ = v1 & ~new_n811_;
  assign new_n827_ = ~new_n219_ & ~new_n826_;
  assign new_n828_ = ~v7 & ~new_n827_;
  assign new_n829_ = v6 & new_n828_;
  assign new_n830_ = v5 & new_n829_;
  assign new_n831_ = ~v4 & new_n830_;
  assign \v8.54  = ~new_n825_ | new_n831_;
  assign new_n833_ = new_n90_ & new_n207_;
  assign new_n834_ = v1 & ~new_n833_;
  assign new_n835_ = v2 & ~new_n714_;
  assign new_n836_ = ~new_n669_ & ~new_n835_;
  assign new_n837_ = v1 & ~new_n836_;
  assign new_n838_ = v0 & new_n837_;
  assign new_n839_ = new_n834_ & ~new_n838_;
  assign new_n840_ = ~new_n626_ & ~new_n766_;
  assign new_n841_ = v0 & ~new_n840_;
  assign new_n842_ = ~v0 & new_n231_;
  assign new_n843_ = ~new_n841_ & ~new_n842_;
  assign new_n844_ = ~v4 & ~new_n843_;
  assign new_n845_ = v1 & new_n844_;
  assign new_n846_ = new_n839_ & ~new_n845_;
  assign new_n847_ = ~v4 & ~\v8.0 ;
  assign new_n848_ = ~v3 & ~new_n847_;
  assign new_n849_ = ~v2 & new_n848_;
  assign new_n850_ = v1 & new_n849_;
  assign new_n851_ = v0 & new_n850_;
  assign new_n852_ = new_n846_ & ~new_n851_;
  assign new_n853_ = v2 & \v8.5 ;
  assign new_n854_ = v1 & new_n853_;
  assign new_n855_ = v0 & new_n854_;
  assign \v8.55  = ~new_n852_ | new_n855_;
  assign new_n857_ = ~v0 & ~new_n353_;
  assign new_n858_ = ~new_n239_ & new_n857_;
  assign new_n859_ = new_n212_ & new_n244_;
  assign new_n860_ = ~new_n738_ & ~new_n859_;
  assign new_n861_ = ~v0 & ~new_n860_;
  assign new_n862_ = new_n858_ & ~new_n861_;
  assign new_n863_ = ~new_n177_ & ~new_n523_;
  assign new_n864_ = v1 & ~new_n863_;
  assign new_n865_ = ~v3 & ~v5;
  assign new_n866_ = new_n212_ & new_n865_;
  assign new_n867_ = ~new_n864_ & ~new_n866_;
  assign new_n868_ = ~v4 & ~new_n867_;
  assign new_n869_ = ~v0 & new_n868_;
  assign new_n870_ = new_n862_ & ~new_n869_;
  assign new_n871_ = ~v1 & ~new_n487_;
  assign new_n872_ = ~v6 & ~new_n871_;
  assign new_n873_ = v5 & new_n872_;
  assign new_n874_ = ~v4 & new_n873_;
  assign new_n875_ = v2 & new_n874_;
  assign new_n876_ = ~v0 & new_n875_;
  assign new_n877_ = new_n870_ & ~new_n876_;
  assign new_n878_ = v2 & v5;
  assign new_n879_ = ~new_n495_ & ~new_n878_;
  assign new_n880_ = v1 & ~new_n879_;
  assign new_n881_ = new_n212_ & new_n343_;
  assign new_n882_ = ~new_n880_ & ~new_n881_;
  assign new_n883_ = ~v7 & ~new_n882_;
  assign new_n884_ = v6 & new_n883_;
  assign new_n885_ = ~v4 & new_n884_;
  assign new_n886_ = ~v0 & new_n885_;
  assign \v8.56  = ~new_n877_ | new_n886_;
  assign new_n888_ = v1 & ~new_n579_;
  assign new_n889_ = v0 & ~new_n888_;
  assign new_n890_ = ~new_n239_ & ~new_n889_;
  assign new_n891_ = ~new_n353_ & new_n890_;
  assign new_n892_ = ~v2 & ~new_n809_;
  assign new_n893_ = v1 & new_n892_;
  assign new_n894_ = v2 & new_n363_;
  assign new_n895_ = new_n104_ & new_n894_;
  assign new_n896_ = ~new_n893_ & ~new_n895_;
  assign new_n897_ = new_n891_ & new_n896_;
  assign new_n898_ = ~new_n523_ & ~new_n804_;
  assign new_n899_ = ~v0 & ~new_n898_;
  assign new_n900_ = new_n176_ & new_n249_;
  assign new_n901_ = ~new_n899_ & ~new_n900_;
  assign new_n902_ = v1 & ~new_n901_;
  assign new_n903_ = v2 & new_n494_;
  assign new_n904_ = new_n104_ & new_n903_;
  assign new_n905_ = ~new_n902_ & ~new_n904_;
  assign new_n906_ = ~v4 & ~new_n905_;
  assign new_n907_ = new_n897_ & ~new_n906_;
  assign new_n908_ = ~v1 & ~new_n489_;
  assign new_n909_ = ~v6 & ~new_n908_;
  assign new_n910_ = v5 & new_n909_;
  assign new_n911_ = ~v4 & new_n910_;
  assign new_n912_ = v2 & new_n911_;
  assign new_n913_ = ~v0 & new_n912_;
  assign new_n914_ = new_n907_ & ~new_n913_;
  assign new_n915_ = ~v2 & new_n865_;
  assign new_n916_ = ~new_n878_ & ~new_n915_;
  assign new_n917_ = ~v0 & ~new_n916_;
  assign new_n918_ = new_n249_ & new_n494_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign new_n920_ = v1 & ~new_n919_;
  assign new_n921_ = new_n104_ & new_n637_;
  assign new_n922_ = ~new_n920_ & ~new_n921_;
  assign new_n923_ = ~v7 & ~new_n922_;
  assign new_n924_ = v6 & new_n923_;
  assign new_n925_ = ~v4 & new_n924_;
  assign \v8.57  = ~new_n914_ | new_n925_;
  assign new_n927_ = ~v3 & ~new_n580_;
  assign new_n928_ = new_n123_ & new_n215_;
  assign new_n929_ = ~new_n927_ & ~new_n928_;
  assign new_n930_ = new_n578_ & new_n929_;
  assign new_n931_ = v3 & new_n618_;
  assign new_n932_ = new_n930_ & ~new_n931_;
  assign new_n933_ = v3 & new_n623_;
  assign new_n934_ = new_n932_ & ~new_n933_;
  assign new_n935_ = v3 & new_n629_;
  assign new_n936_ = new_n934_ & ~new_n935_;
  assign new_n937_ = new_n97_ & new_n878_;
  assign new_n938_ = new_n104_ & new_n634_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = ~v7 & ~new_n939_;
  assign new_n941_ = v6 & new_n940_;
  assign new_n942_ = ~v4 & new_n941_;
  assign new_n943_ = v3 & new_n942_;
  assign \v8.58  = ~new_n936_ | new_n943_;
  assign new_n945_ = ~v4 & ~new_n207_;
  assign new_n946_ = ~v0 & ~new_n945_;
  assign new_n947_ = v0 & new_n207_;
  assign new_n948_ = ~new_n946_ & ~new_n947_;
  assign new_n949_ = v0 & new_n583_;
  assign new_n950_ = new_n948_ & ~new_n949_;
  assign new_n951_ = ~new_n590_ & ~new_n592_;
  assign new_n952_ = v0 & ~new_n951_;
  assign new_n953_ = ~v0 & ~v6;
  assign new_n954_ = ~new_n952_ & ~new_n953_;
  assign new_n955_ = ~v5 & ~new_n954_;
  assign new_n956_ = ~v4 & new_n955_;
  assign new_n957_ = new_n950_ & ~new_n956_;
  assign new_n958_ = ~new_n571_ & ~new_n604_;
  assign new_n959_ = v6 & ~new_n958_;
  assign new_n960_ = ~v5 & new_n959_;
  assign new_n961_ = ~v4 & new_n960_;
  assign new_n962_ = new_n957_ & ~new_n961_;
  assign new_n963_ = ~v4 & ~new_n275_;
  assign new_n964_ = ~new_n488_ & ~new_n963_;
  assign new_n965_ = v2 & new_n964_;
  assign new_n966_ = ~v4 & v6;
  assign new_n967_ = ~v3 & new_n966_;
  assign new_n968_ = new_n577_ & new_n967_;
  assign new_n969_ = ~new_n965_ & ~new_n968_;
  assign new_n970_ = ~v5 & ~new_n969_;
  assign new_n971_ = v5 & ~new_n488_;
  assign new_n972_ = v4 & new_n971_;
  assign new_n973_ = v2 & new_n972_;
  assign new_n974_ = ~new_n970_ & ~new_n973_;
  assign new_n975_ = v0 & ~new_n974_;
  assign new_n976_ = new_n231_ & new_n244_;
  assign new_n977_ = new_n326_ & new_n976_;
  assign new_n978_ = ~new_n975_ & ~new_n977_;
  assign new_n979_ = new_n962_ & new_n978_;
  assign new_n980_ = v2 & ~new_n726_;
  assign new_n981_ = ~v0 & ~new_n980_;
  assign new_n982_ = new_n97_ & new_n215_;
  assign new_n983_ = ~new_n981_ & ~new_n982_;
  assign new_n984_ = ~v7 & ~new_n983_;
  assign new_n985_ = v6 & new_n984_;
  assign new_n986_ = ~v5 & new_n985_;
  assign new_n987_ = ~v4 & new_n986_;
  assign \v8.59  = ~new_n979_ | new_n987_;
  assign new_n989_ = ~v1 & v4;
  assign new_n990_ = ~v0 & new_n989_;
  assign new_n991_ = ~new_n506_ & ~new_n990_;
  assign new_n992_ = new_n680_ & new_n991_;
  assign new_n993_ = new_n97_ & new_n656_;
  assign new_n994_ = new_n992_ & ~new_n993_;
  assign new_n995_ = ~v4 & ~new_n217_;
  assign new_n996_ = ~v1 & new_n995_;
  assign new_n997_ = ~v0 & new_n996_;
  assign new_n998_ = new_n994_ & ~new_n997_;
  assign new_n999_ = ~new_n228_ & new_n998_;
  assign new_n1000_ = ~v6 & ~new_n224_;
  assign new_n1001_ = v5 & new_n1000_;
  assign new_n1002_ = ~v4 & new_n1001_;
  assign new_n1003_ = ~v1 & new_n1002_;
  assign new_n1004_ = ~v0 & new_n1003_;
  assign new_n1005_ = new_n999_ & ~new_n1004_;
  assign new_n1006_ = ~v7 & ~new_n224_;
  assign new_n1007_ = v6 & new_n1006_;
  assign new_n1008_ = v5 & new_n1007_;
  assign new_n1009_ = ~v4 & new_n1008_;
  assign new_n1010_ = ~v1 & new_n1009_;
  assign new_n1011_ = ~v0 & new_n1010_;
  assign \v8.60  = ~new_n1005_ | new_n1011_;
  assign new_n1013_ = new_n371_ & ~new_n571_;
  assign new_n1014_ = ~new_n509_ & new_n1013_;
  assign new_n1015_ = ~new_n755_ & new_n1014_;
  assign new_n1016_ = new_n213_ & new_n976_;
  assign \v8.61  = ~new_n1015_ | new_n1016_;
  assign new_n1018_ = new_n369_ & ~new_n687_;
  assign new_n1019_ = new_n97_ & new_n455_;
  assign new_n1020_ = new_n1018_ & ~new_n1019_;
  assign new_n1021_ = new_n232_ & new_n697_;
  assign \v8.62  = ~new_n1020_ | new_n1021_;
endmodule


