// Benchmark "x4" written by ABC on Fri Feb 25 15:12:29 2022

module x4 ( 
    a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z, a0, b0,
    c0, d0, e0, f0, g0, h0, i0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0,
    v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1,
    n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2,
    f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2,
    w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3,
    o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4,
    g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4,
    y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5  );
  input  a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y, z,
    a0, b0, c0, d0, e0, f0, g0, h0, i0, k0, l0, m0, n0, o0, p0, q0, r0, s0,
    t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1,
    l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2,
    d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2,
    v2;
  output w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3,
    n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4,
    f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4,
    x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5;
  wire new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n212_,
    new_n214_, new_n216_, new_n218_, new_n220_, new_n222_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n239_,
    new_n240_, new_n241_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n282_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n343_,
    new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_,
    new_n350_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_;
  assign new_n166_ = ~p2 & r2;
  assign new_n167_ = n2 & ~o2;
  assign new_n168_ = new_n166_ & new_n167_;
  assign new_n169_ = h0 & ~t2;
  assign new_n170_ = ~h0 & t2;
  assign new_n171_ = ~i & ~q2;
  assign new_n172_ = ~new_n170_ & ~new_n171_;
  assign new_n173_ = ~new_n169_ & new_n172_;
  assign new_n174_ = e1 & ~o2;
  assign new_n175_ = n2 & ~new_n171_;
  assign new_n176_ = new_n174_ & new_n175_;
  assign new_n177_ = new_n166_ & new_n176_;
  assign new_n178_ = new_n168_ & new_n173_;
  assign new_n179_ = e1 & new_n178_;
  assign new_n180_ = s2 & ~new_n177_;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign c3 = ~i0 & ~new_n181_;
  assign new_n183_ = ~g & ~h;
  assign new_n184_ = ~i & h0;
  assign new_n185_ = new_n183_ & new_n184_;
  assign new_n186_ = m1 & ~new_n185_;
  assign new_n187_ = f0 & v2;
  assign new_n188_ = ~k0 & ~new_n187_;
  assign new_n189_ = ~c1 & ~new_n188_;
  assign new_n190_ = ~c1 & v2;
  assign new_n191_ = g0 & ~new_n186_;
  assign new_n192_ = new_n190_ & new_n191_;
  assign d3 = new_n189_ | new_n192_;
  assign new_n194_ = ~o2 & ~p2;
  assign new_n195_ = ~q2 & ~r2;
  assign new_n196_ = new_n194_ & new_n195_;
  assign new_n197_ = n2 & new_n196_;
  assign new_n198_ = e1 & new_n197_;
  assign new_n199_ = ~l0 & ~new_n198_;
  assign e3 = ~c1 & ~new_n199_;
  assign new_n201_ = g0 & v2;
  assign new_n202_ = m0 & ~new_n201_;
  assign new_n203_ = ~i0 & ~new_n202_;
  assign new_n204_ = v2 & new_n191_;
  assign f3 = ~new_n203_ | new_n204_;
  assign new_n206_ = ~p2 & new_n195_;
  assign new_n207_ = e1 & new_n206_;
  assign new_n208_ = new_n167_ & new_n207_;
  assign new_n209_ = ~n0 & ~new_n208_;
  assign new_n210_ = ~i0 & ~c1;
  assign g3 = ~new_n209_ & new_n210_;
  assign new_n212_ = o0 & ~c1;
  assign h3 = ~i0 & new_n212_;
  assign new_n214_ = p0 & ~c1;
  assign i3 = ~i0 & new_n214_;
  assign new_n216_ = q0 & ~c1;
  assign j3 = ~i0 & new_n216_;
  assign new_n218_ = r0 & ~c1;
  assign k3 = ~i0 & new_n218_;
  assign new_n220_ = s0 & ~c1;
  assign l3 = ~i0 & new_n220_;
  assign new_n222_ = t0 & ~c1;
  assign m3 = ~i0 & new_n222_;
  assign n3 = b & ~i0;
  assign o3 = a & ~i0;
  assign p3 = ~i0 & v0;
  assign q3 = ~i0 & w0;
  assign r3 = ~i0 & x0;
  assign s3 = ~i0 & y0;
  assign t3 = ~i0 & z0;
  assign u3 = ~i0 & a1;
  assign new_n232_ = ~o2 & new_n166_;
  assign new_n233_ = ~i0 & ~new_n187_;
  assign new_n234_ = ~new_n171_ & new_n232_;
  assign new_n235_ = e1 & n2;
  assign new_n236_ = new_n234_ & new_n235_;
  assign new_n237_ = ~new_n204_ & ~new_n236_;
  assign v3 = ~new_n233_ | ~new_n237_;
  assign new_n239_ = ~g0 & ~m1;
  assign new_n240_ = i0 & ~new_n185_;
  assign new_n241_ = new_n239_ & new_n240_;
  assign w3 = v2 & new_n241_;
  assign new_n243_ = l2 & m2;
  assign new_n244_ = ~k2 & new_n243_;
  assign new_n245_ = ~d1 & ~new_n244_;
  assign new_n246_ = ~e1 & new_n245_;
  assign x3 = ~c1 & ~new_n246_;
  assign new_n248_ = o2 & new_n206_;
  assign new_n249_ = ~n2 & o2;
  assign new_n250_ = new_n207_ & new_n249_;
  assign new_n251_ = ~f1 & ~new_n250_;
  assign new_n252_ = e1 & ~n2;
  assign new_n253_ = ~o0 & new_n248_;
  assign new_n254_ = new_n252_ & new_n253_;
  assign new_n255_ = ~new_n251_ & ~new_n254_;
  assign y3 = ~c1 & new_n255_;
  assign new_n257_ = ~g1 & ~new_n250_;
  assign new_n258_ = ~p0 & new_n248_;
  assign new_n259_ = new_n252_ & new_n258_;
  assign new_n260_ = ~new_n257_ & ~new_n259_;
  assign z3 = ~c1 & new_n260_;
  assign new_n262_ = ~h1 & ~new_n250_;
  assign new_n263_ = ~q0 & new_n248_;
  assign new_n264_ = new_n252_ & new_n263_;
  assign new_n265_ = ~new_n262_ & ~new_n264_;
  assign a4 = ~c1 & new_n265_;
  assign new_n267_ = ~i1 & ~new_n250_;
  assign new_n268_ = ~r0 & new_n248_;
  assign new_n269_ = new_n252_ & new_n268_;
  assign new_n270_ = ~new_n267_ & ~new_n269_;
  assign b4 = ~c1 & new_n270_;
  assign new_n272_ = ~j1 & ~new_n250_;
  assign new_n273_ = ~s0 & new_n248_;
  assign new_n274_ = new_n252_ & new_n273_;
  assign new_n275_ = ~new_n272_ & ~new_n274_;
  assign c4 = ~c1 & new_n275_;
  assign new_n277_ = ~k1 & ~new_n250_;
  assign new_n278_ = ~t0 & new_n248_;
  assign new_n279_ = new_n252_ & new_n278_;
  assign new_n280_ = ~new_n277_ & ~new_n279_;
  assign d4 = ~c1 & new_n280_;
  assign new_n282_ = ~l1 & ~new_n198_;
  assign e4 = ~c1 & ~new_n282_;
  assign new_n284_ = ~h & ~k2;
  assign new_n285_ = ~g & new_n243_;
  assign new_n286_ = new_n284_ & new_n285_;
  assign new_n287_ = ~i0 & ~new_n201_;
  assign new_n288_ = ~m1 & ~new_n286_;
  assign f4 = new_n287_ & ~new_n288_;
  assign new_n290_ = e1 & ~o1;
  assign new_n291_ = ~h & h0;
  assign new_n292_ = ~g & new_n291_;
  assign new_n293_ = m1 & ~new_n292_;
  assign new_n294_ = v2 & new_n293_;
  assign new_n295_ = g0 & new_n294_;
  assign new_n296_ = m1 & v2;
  assign new_n297_ = ~m0 & e1;
  assign new_n298_ = h0 & new_n183_;
  assign new_n299_ = m1 & ~new_n298_;
  assign new_n300_ = g0 & new_n299_;
  assign new_n301_ = v2 & new_n300_;
  assign new_n302_ = ~new_n297_ & ~new_n301_;
  assign new_n303_ = new_n290_ & ~new_n295_;
  assign new_n304_ = ~m0 & new_n303_;
  assign new_n305_ = i & new_n296_;
  assign new_n306_ = g0 & new_n305_;
  assign new_n307_ = n1 & new_n302_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = ~new_n304_ & new_n308_;
  assign g4 = ~i0 & ~new_n309_;
  assign new_n311_ = ~h & new_n184_;
  assign new_n312_ = ~g & new_n311_;
  assign new_n313_ = ~o1 & ~new_n297_;
  assign new_n314_ = o1 & ~new_n297_;
  assign new_n315_ = p1 & ~new_n314_;
  assign new_n316_ = ~new_n313_ & ~new_n315_;
  assign new_n317_ = ~i0 & ~new_n316_;
  assign new_n318_ = g0 & ~new_n312_;
  assign new_n319_ = new_n296_ & new_n318_;
  assign h4 = ~new_n317_ | new_n319_;
  assign new_n321_ = ~i0 & new_n296_;
  assign new_n322_ = e1 & q1;
  assign new_n323_ = v2 & new_n186_;
  assign new_n324_ = g0 & new_n323_;
  assign new_n325_ = ~new_n297_ & ~new_n319_;
  assign new_n326_ = new_n322_ & ~new_n324_;
  assign new_n327_ = ~m0 & new_n326_;
  assign new_n328_ = p1 & new_n325_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~i0 & ~new_n329_;
  assign new_n331_ = k & new_n321_;
  assign new_n332_ = new_n318_ & new_n331_;
  assign i4 = new_n330_ | new_n332_;
  assign new_n334_ = e1 & r1;
  assign new_n335_ = ~new_n324_ & new_n334_;
  assign new_n336_ = ~m0 & new_n335_;
  assign new_n337_ = q1 & new_n325_;
  assign new_n338_ = ~new_n336_ & ~new_n337_;
  assign new_n339_ = ~i0 & ~new_n338_;
  assign new_n340_ = l & new_n321_;
  assign new_n341_ = new_n318_ & new_n340_;
  assign j4 = new_n339_ | new_n341_;
  assign new_n343_ = e1 & s1;
  assign new_n344_ = ~new_n324_ & new_n343_;
  assign new_n345_ = ~m0 & new_n344_;
  assign new_n346_ = r1 & new_n325_;
  assign new_n347_ = ~new_n345_ & ~new_n346_;
  assign new_n348_ = ~i0 & ~new_n347_;
  assign new_n349_ = m & new_n321_;
  assign new_n350_ = new_n318_ & new_n349_;
  assign k4 = new_n348_ | new_n350_;
  assign new_n352_ = e1 & t1;
  assign new_n353_ = ~new_n324_ & new_n352_;
  assign new_n354_ = ~m0 & new_n353_;
  assign new_n355_ = s1 & new_n325_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = ~i0 & ~new_n356_;
  assign new_n358_ = n & new_n321_;
  assign new_n359_ = new_n318_ & new_n358_;
  assign l4 = new_n357_ | new_n359_;
  assign new_n361_ = e1 & u1;
  assign new_n362_ = ~new_n324_ & new_n361_;
  assign new_n363_ = ~m0 & new_n362_;
  assign new_n364_ = t1 & new_n325_;
  assign new_n365_ = ~new_n363_ & ~new_n364_;
  assign new_n366_ = ~i0 & ~new_n365_;
  assign new_n367_ = o & new_n321_;
  assign new_n368_ = new_n318_ & new_n367_;
  assign m4 = new_n366_ | new_n368_;
  assign new_n370_ = e1 & v1;
  assign new_n371_ = ~new_n324_ & new_n370_;
  assign new_n372_ = ~m0 & new_n371_;
  assign new_n373_ = u1 & new_n325_;
  assign new_n374_ = ~new_n372_ & ~new_n373_;
  assign new_n375_ = ~i0 & ~new_n374_;
  assign new_n376_ = p & new_n321_;
  assign new_n377_ = new_n318_ & new_n376_;
  assign n4 = new_n375_ | new_n377_;
  assign new_n379_ = e1 & w1;
  assign new_n380_ = ~new_n324_ & new_n379_;
  assign new_n381_ = ~m0 & new_n380_;
  assign new_n382_ = v1 & new_n325_;
  assign new_n383_ = ~new_n381_ & ~new_n382_;
  assign new_n384_ = ~i0 & ~new_n383_;
  assign new_n385_ = q & new_n321_;
  assign new_n386_ = new_n318_ & new_n385_;
  assign o4 = new_n384_ | new_n386_;
  assign new_n388_ = e1 & x1;
  assign new_n389_ = ~new_n324_ & new_n388_;
  assign new_n390_ = ~m0 & new_n389_;
  assign new_n391_ = w1 & new_n325_;
  assign new_n392_ = ~new_n390_ & ~new_n391_;
  assign new_n393_ = ~i0 & ~new_n392_;
  assign new_n394_ = r & new_n321_;
  assign new_n395_ = new_n318_ & new_n394_;
  assign p4 = new_n393_ | new_n395_;
  assign new_n397_ = e1 & y1;
  assign new_n398_ = ~new_n324_ & new_n397_;
  assign new_n399_ = ~m0 & new_n398_;
  assign new_n400_ = x1 & new_n325_;
  assign new_n401_ = ~new_n399_ & ~new_n400_;
  assign new_n402_ = ~i0 & ~new_n401_;
  assign new_n403_ = s & new_n321_;
  assign new_n404_ = new_n318_ & new_n403_;
  assign q4 = new_n402_ | new_n404_;
  assign new_n406_ = e1 & z1;
  assign new_n407_ = ~new_n324_ & new_n406_;
  assign new_n408_ = ~m0 & new_n407_;
  assign new_n409_ = y1 & new_n325_;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = ~i0 & ~new_n410_;
  assign new_n412_ = t & new_n321_;
  assign new_n413_ = new_n318_ & new_n412_;
  assign r4 = new_n411_ | new_n413_;
  assign new_n415_ = e1 & a2;
  assign new_n416_ = ~new_n324_ & new_n415_;
  assign new_n417_ = ~m0 & new_n416_;
  assign new_n418_ = z1 & new_n325_;
  assign new_n419_ = ~new_n417_ & ~new_n418_;
  assign new_n420_ = ~i0 & ~new_n419_;
  assign new_n421_ = u & new_n321_;
  assign new_n422_ = new_n318_ & new_n421_;
  assign s4 = new_n420_ | new_n422_;
  assign new_n424_ = e1 & b2;
  assign new_n425_ = ~new_n324_ & new_n424_;
  assign new_n426_ = ~m0 & new_n425_;
  assign new_n427_ = a2 & new_n325_;
  assign new_n428_ = ~new_n426_ & ~new_n427_;
  assign new_n429_ = ~i0 & ~new_n428_;
  assign new_n430_ = v & new_n321_;
  assign new_n431_ = new_n318_ & new_n430_;
  assign t4 = new_n429_ | new_n431_;
  assign new_n433_ = e1 & c2;
  assign new_n434_ = ~new_n324_ & new_n433_;
  assign new_n435_ = ~m0 & new_n434_;
  assign new_n436_ = b2 & new_n325_;
  assign new_n437_ = ~new_n435_ & ~new_n436_;
  assign new_n438_ = ~i0 & ~new_n437_;
  assign new_n439_ = w & new_n321_;
  assign new_n440_ = new_n318_ & new_n439_;
  assign u4 = new_n438_ | new_n440_;
  assign new_n442_ = e1 & d2;
  assign new_n443_ = ~new_n324_ & new_n442_;
  assign new_n444_ = ~m0 & new_n443_;
  assign new_n445_ = c2 & new_n325_;
  assign new_n446_ = ~new_n444_ & ~new_n445_;
  assign new_n447_ = ~i0 & ~new_n446_;
  assign new_n448_ = x & new_n321_;
  assign new_n449_ = new_n318_ & new_n448_;
  assign v4 = new_n447_ | new_n449_;
  assign new_n451_ = e1 & e2;
  assign new_n452_ = ~new_n324_ & new_n451_;
  assign new_n453_ = ~m0 & new_n452_;
  assign new_n454_ = d2 & new_n325_;
  assign new_n455_ = ~new_n453_ & ~new_n454_;
  assign new_n456_ = ~i0 & ~new_n455_;
  assign new_n457_ = y & new_n321_;
  assign new_n458_ = new_n318_ & new_n457_;
  assign w4 = new_n456_ | new_n458_;
  assign new_n460_ = e1 & f2;
  assign new_n461_ = ~new_n324_ & new_n460_;
  assign new_n462_ = ~m0 & new_n461_;
  assign new_n463_ = e2 & new_n325_;
  assign new_n464_ = ~new_n462_ & ~new_n463_;
  assign new_n465_ = ~i0 & ~new_n464_;
  assign new_n466_ = z & new_n321_;
  assign new_n467_ = new_n318_ & new_n466_;
  assign x4 = new_n465_ | new_n467_;
  assign new_n469_ = e1 & g2;
  assign new_n470_ = ~new_n324_ & new_n469_;
  assign new_n471_ = ~m0 & new_n470_;
  assign new_n472_ = f2 & new_n325_;
  assign new_n473_ = ~new_n471_ & ~new_n472_;
  assign new_n474_ = ~i0 & ~new_n473_;
  assign new_n475_ = a0 & new_n321_;
  assign new_n476_ = new_n318_ & new_n475_;
  assign y4 = new_n474_ | new_n476_;
  assign new_n478_ = e1 & h2;
  assign new_n479_ = ~new_n324_ & new_n478_;
  assign new_n480_ = ~m0 & new_n479_;
  assign new_n481_ = g2 & new_n325_;
  assign new_n482_ = ~new_n480_ & ~new_n481_;
  assign new_n483_ = ~i0 & ~new_n482_;
  assign new_n484_ = b0 & new_n321_;
  assign new_n485_ = new_n318_ & new_n484_;
  assign z4 = new_n483_ | new_n485_;
  assign new_n487_ = e1 & i2;
  assign new_n488_ = ~new_n324_ & new_n487_;
  assign new_n489_ = ~m0 & new_n488_;
  assign new_n490_ = h2 & new_n325_;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = ~i0 & ~new_n491_;
  assign new_n493_ = c0 & new_n321_;
  assign new_n494_ = new_n318_ & new_n493_;
  assign a5 = new_n492_ | new_n494_;
  assign new_n496_ = e1 & j2;
  assign new_n497_ = ~new_n324_ & new_n496_;
  assign new_n498_ = ~m0 & new_n497_;
  assign new_n499_ = i2 & new_n325_;
  assign new_n500_ = ~new_n498_ & ~new_n499_;
  assign new_n501_ = ~i0 & ~new_n500_;
  assign new_n502_ = d0 & new_n321_;
  assign new_n503_ = new_n318_ & new_n502_;
  assign b5 = new_n501_ | new_n503_;
  assign new_n505_ = ~new_n312_ & new_n321_;
  assign new_n506_ = e0 & g0;
  assign new_n507_ = new_n505_ & new_n506_;
  assign new_n508_ = ~i0 & new_n325_;
  assign new_n509_ = j2 & new_n508_;
  assign c5 = new_n507_ | new_n509_;
  assign new_n511_ = b & ~u0;
  assign new_n512_ = ~u2 & ~new_n511_;
  assign new_n513_ = k2 & ~new_n512_;
  assign new_n514_ = ~c1 & ~new_n513_;
  assign new_n515_ = ~k2 & ~new_n511_;
  assign new_n516_ = ~u2 & new_n515_;
  assign d5 = new_n514_ & ~new_n516_;
  assign new_n518_ = l2 & ~m2;
  assign new_n519_ = ~k2 & ~new_n518_;
  assign new_n520_ = ~c1 & ~new_n519_;
  assign new_n521_ = ~l2 & new_n512_;
  assign new_n522_ = ~new_n513_ & ~new_n521_;
  assign new_n523_ = ~l2 & ~new_n512_;
  assign new_n524_ = ~new_n522_ & ~new_n523_;
  assign e5 = new_n520_ & ~new_n524_;
  assign new_n526_ = ~l2 & m2;
  assign new_n527_ = ~k2 & ~new_n526_;
  assign new_n528_ = ~l2 & ~m2;
  assign new_n529_ = ~c1 & ~new_n528_;
  assign new_n530_ = ~new_n527_ & new_n529_;
  assign new_n531_ = l2 & ~new_n512_;
  assign new_n532_ = ~m2 & new_n512_;
  assign new_n533_ = ~new_n531_ & ~new_n532_;
  assign new_n534_ = ~m2 & ~new_n512_;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign f5 = new_n530_ & ~new_n535_;
  assign new_n537_ = n2 & ~new_n246_;
  assign new_n538_ = ~c1 & ~new_n537_;
  assign new_n539_ = ~e1 & ~n2;
  assign new_n540_ = new_n245_ & new_n539_;
  assign g5 = new_n538_ & ~new_n540_;
  assign new_n542_ = ~e1 & ~new_n244_;
  assign new_n543_ = ~d1 & new_n542_;
  assign new_n544_ = ~n2 & ~o2;
  assign new_n545_ = ~c1 & ~new_n544_;
  assign new_n546_ = n2 & ~new_n543_;
  assign new_n547_ = ~e1 & ~o2;
  assign new_n548_ = new_n245_ & new_n547_;
  assign new_n549_ = ~new_n546_ & ~new_n548_;
  assign new_n550_ = ~o2 & ~new_n246_;
  assign new_n551_ = ~new_n549_ & ~new_n550_;
  assign h5 = new_n545_ & ~new_n551_;
  assign new_n553_ = n2 & o2;
  assign new_n554_ = ~p2 & ~new_n553_;
  assign new_n555_ = ~c1 & ~new_n554_;
  assign new_n556_ = o2 & ~new_n543_;
  assign new_n557_ = n2 & new_n556_;
  assign new_n558_ = ~e1 & ~p2;
  assign new_n559_ = new_n245_ & new_n558_;
  assign new_n560_ = ~new_n557_ & ~new_n559_;
  assign new_n561_ = ~p2 & ~new_n246_;
  assign new_n562_ = ~new_n560_ & ~new_n561_;
  assign i5 = new_n555_ & ~new_n562_;
  assign new_n564_ = p2 & q2;
  assign new_n565_ = o2 & p2;
  assign new_n566_ = n2 & new_n565_;
  assign new_n567_ = ~q2 & ~new_n566_;
  assign new_n568_ = ~c1 & ~new_n567_;
  assign new_n569_ = ~e1 & ~q2;
  assign new_n570_ = new_n245_ & new_n569_;
  assign new_n571_ = ~new_n543_ & new_n564_;
  assign new_n572_ = new_n553_ & new_n571_;
  assign new_n573_ = ~new_n570_ & ~new_n572_;
  assign j5 = new_n568_ & new_n573_;
  assign new_n575_ = q2 & r2;
  assign new_n576_ = p2 & new_n575_;
  assign new_n577_ = new_n553_ & new_n564_;
  assign new_n578_ = ~new_n246_ & new_n577_;
  assign new_n579_ = ~r2 & ~new_n578_;
  assign new_n580_ = ~new_n543_ & new_n576_;
  assign new_n581_ = new_n553_ & new_n580_;
  assign new_n582_ = ~new_n579_ & ~new_n581_;
  assign k5 = ~c1 & new_n582_;
  assign new_n584_ = ~b1 & ~new_n297_;
  assign new_n585_ = n1 & ~new_n584_;
  assign new_n586_ = b1 & ~new_n297_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign l5 = ~i0 & ~new_n587_;
  assign new_n589_ = s2 & ~t2;
  assign new_n590_ = l1 & new_n589_;
  assign new_n591_ = l1 & s2;
  assign new_n592_ = t2 & ~new_n591_;
  assign new_n593_ = ~new_n590_ & ~new_n592_;
  assign m5 = ~c1 & ~new_n593_;
  assign new_n595_ = ~i0 & ~new_n512_;
  assign new_n596_ = new_n243_ & new_n515_;
  assign n5 = new_n595_ & ~new_n596_;
  assign new_n598_ = r2 & ~new_n171_;
  assign new_n599_ = ~o2 & new_n598_;
  assign new_n600_ = ~p2 & new_n599_;
  assign new_n601_ = new_n235_ & new_n600_;
  assign new_n602_ = ~f0 & v2;
  assign new_n603_ = ~new_n601_ & ~new_n602_;
  assign o5 = new_n287_ & ~new_n603_;
  assign w2 = ~f1;
  assign x2 = ~g1;
  assign y2 = ~h1;
  assign z2 = ~i1;
  assign a3 = ~j1;
  assign b3 = ~k1;
endmodule


